

module b17_C_AntiSAT_k_256_1 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9786, n9787, n9789, n9790, n9791, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553;

  INV_X1 U11229 ( .A(n21348), .ZN(n21339) );
  OR2_X1 U11230 ( .A1(n13163), .A2(n13162), .ZN(n10292) );
  OR2_X1 U11232 ( .A1(n9851), .A2(n15485), .ZN(n15487) );
  OR2_X1 U11233 ( .A1(n15142), .A2(n15143), .ZN(n15161) );
  NOR2_X1 U11234 ( .A1(n13489), .A2(n17781), .ZN(n15398) );
  INV_X1 U11235 ( .A(n12435), .ZN(n12277) );
  INV_X1 U11236 ( .A(n9787), .ZN(n18532) );
  INV_X2 U11237 ( .A(n11790), .ZN(n20565) );
  BUF_X2 U11238 ( .A(n12907), .Z(n16946) );
  AND2_X1 U11240 ( .A1(n11455), .A2(n17691), .ZN(n13058) );
  AND2_X1 U11241 ( .A1(n9821), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11856) );
  AND2_X1 U11242 ( .A1(n13039), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12329) );
  AND2_X1 U11243 ( .A1(n9813), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11681) );
  INV_X1 U11244 ( .A(n9862), .ZN(n18473) );
  INV_X2 U11245 ( .A(n9850), .ZN(n18533) );
  INV_X2 U11246 ( .A(n18453), .ZN(n18520) );
  AND2_X1 U11247 ( .A1(n14049), .A2(n15100), .ZN(n12648) );
  OAI211_X1 U11248 ( .C1(n11514), .C2(n11501), .A(n11500), .B(n11499), .ZN(
        n11534) );
  NAND2_X1 U11250 ( .A1(n20169), .A2(n20160), .ZN(n13227) );
  NAND2_X1 U11251 ( .A1(n12688), .A2(n12732), .ZN(n13953) );
  NAND2_X1 U11252 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13228) );
  NAND2_X2 U11253 ( .A1(n20184), .A2(n20177), .ZN(n18256) );
  AND2_X1 U11254 ( .A1(n11483), .A2(n13776), .ZN(n11498) );
  CLKBUF_X2 U11256 ( .A(n11471), .Z(n13777) );
  INV_X2 U11257 ( .A(n12242), .ZN(n11482) );
  AND2_X4 U11259 ( .A1(n13885), .A2(n10368), .ZN(n10471) );
  AND2_X1 U11261 ( .A1(n10359), .A2(n10366), .ZN(n10558) );
  AND2_X1 U11262 ( .A1(n10367), .A2(n13885), .ZN(n10569) );
  AND2_X1 U11263 ( .A1(n10366), .A2(n13885), .ZN(n10539) );
  CLKBUF_X2 U11264 ( .A(n10445), .Z(n9814) );
  AND3_X2 U11265 ( .A1(n17686), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9819) );
  INV_X1 U11267 ( .A(n21553), .ZN(n9786) );
  AND2_X1 U11268 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11602), .ZN(
        n13063) );
  NOR2_X1 U11269 ( .A1(n11586), .A2(n11585), .ZN(n11835) );
  INV_X2 U11270 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17686) );
  INV_X1 U11271 ( .A(n14049), .ZN(n10532) );
  NOR2_X1 U11272 ( .A1(n10548), .A2(n10549), .ZN(n10530) );
  INV_X1 U11273 ( .A(n13067), .ZN(n12427) );
  AND2_X1 U11274 ( .A1(n11867), .A2(n11866), .ZN(n12170) );
  AOI21_X2 U11275 ( .B1(n12092), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11538), .ZN(n11540) );
  INV_X1 U11276 ( .A(n11481), .ZN(n12253) );
  AND3_X1 U11277 ( .A1(n11381), .A2(n17691), .A3(n11380), .ZN(n11384) );
  NAND2_X1 U11278 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20184), .ZN(
        n13226) );
  NAND3_X1 U11279 ( .A1(n18935), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18873) );
  INV_X1 U11280 ( .A(n15100), .ZN(n12789) );
  NOR2_X1 U11281 ( .A1(n12759), .A2(n14135), .ZN(n12747) );
  NOR2_X1 U11282 ( .A1(n14069), .A2(n14058), .ZN(n13955) );
  NAND2_X1 U11283 ( .A1(n12732), .A2(n10237), .ZN(n12764) );
  XNOR2_X1 U11284 ( .A(n10511), .B(n10512), .ZN(n14178) );
  AOI21_X2 U11285 ( .B1(n10596), .B2(n10531), .A(n10530), .ZN(n10553) );
  CLKBUF_X3 U11286 ( .A(n12092), .Z(n12129) );
  INV_X2 U11287 ( .A(n11892), .ZN(n12003) );
  BUF_X1 U11288 ( .A(n13296), .Z(n18519) );
  NAND2_X1 U11290 ( .A1(n13984), .A2(n15100), .ZN(n21543) );
  NAND2_X2 U11291 ( .A1(n14069), .A2(n17165), .ZN(n12732) );
  INV_X1 U11292 ( .A(n17165), .ZN(n13984) );
  NAND3_X1 U11293 ( .A1(n10257), .A2(n10684), .A3(n14168), .ZN(n14415) );
  INV_X1 U11294 ( .A(n16288), .ZN(n10274) );
  NAND2_X1 U11295 ( .A1(n14178), .A2(n10553), .ZN(n14030) );
  XNOR2_X1 U11296 ( .A(n13143), .B(n13144), .ZN(n16424) );
  XNOR2_X1 U11297 ( .A(n13077), .B(n13100), .ZN(n16519) );
  INV_X1 U11298 ( .A(n12290), .ZN(n10193) );
  NOR2_X1 U11299 ( .A1(n16579), .A2(n16747), .ZN(n16580) );
  NOR2_X1 U11300 ( .A1(n17967), .A2(n18893), .ZN(n17966) );
  NOR2_X1 U11301 ( .A1(n17998), .A2(n18938), .ZN(n17997) );
  INV_X1 U11302 ( .A(n18243), .ZN(n18263) );
  AND2_X1 U11303 ( .A1(n10350), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18935) );
  INV_X1 U11304 ( .A(n10237), .ZN(n14135) );
  NAND2_X1 U11305 ( .A1(n15362), .A2(n9837), .ZN(n16278) );
  INV_X1 U11306 ( .A(n17352), .ZN(n17369) );
  OR2_X1 U11307 ( .A1(n16620), .A2(n16619), .ZN(n10093) );
  NAND2_X1 U11308 ( .A1(n12918), .A2(n12917), .ZN(n16932) );
  INV_X2 U11309 ( .A(n19584), .ZN(n18624) );
  NOR2_X1 U11310 ( .A1(n17934), .A2(n17935), .ZN(n17933) );
  INV_X1 U11311 ( .A(n19071), .ZN(n19067) );
  OR2_X1 U11312 ( .A1(n13224), .A2(n13223), .ZN(n9787) );
  BUF_X2 U11313 ( .A(n11607), .Z(n9820) );
  NAND2_X2 U11314 ( .A1(n13905), .A2(n13904), .ZN(n13903) );
  AOI21_X2 U11315 ( .B1(n11253), .B2(n10872), .A(n10734), .ZN(n14888) );
  NOR2_X2 U11317 ( .A1(n13337), .A2(n19146), .ZN(n13339) );
  NAND2_X1 U11319 ( .A1(n11482), .A2(n11481), .ZN(n12240) );
  XOR2_X2 U11320 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n13531), .Z(
        n13603) );
  NOR2_X4 U11321 ( .A1(n19113), .A2(n19326), .ZN(n19018) );
  AOI22_X4 U11322 ( .A1(n19062), .A2(n19407), .B1(n19061), .B2(n19405), .ZN(
        n19113) );
  OAI21_X2 U11323 ( .B1(n10655), .B2(n14173), .A(n10253), .ZN(n14202) );
  OR2_X2 U11325 ( .A1(n13907), .A2(n11565), .ZN(n10060) );
  INV_X2 U11327 ( .A(n13259), .ZN(n13298) );
  NOR2_X2 U11328 ( .A1(n16882), .A2(n17615), .ZN(n15031) );
  OR2_X2 U11329 ( .A1(n16519), .A2(n10296), .ZN(n10293) );
  NAND2_X2 U11330 ( .A1(n11802), .A2(n11803), .ZN(n12152) );
  AND2_X2 U11331 ( .A1(n11614), .A2(n11613), .ZN(n11802) );
  CLKBUF_X3 U11332 ( .A(n11606), .Z(n13203) );
  NAND2_X1 U11333 ( .A1(n11510), .A2(n11509), .ZN(n10057) );
  NAND2_X2 U11334 ( .A1(n11367), .A2(n11366), .ZN(n11472) );
  INV_X1 U11335 ( .A(n12129), .ZN(n9789) );
  BUF_X4 U11336 ( .A(n13275), .Z(n18534) );
  XNOR2_X1 U11337 ( .A(n15424), .B(n15423), .ZN(n15434) );
  CLKBUF_X1 U11338 ( .A(n15495), .Z(n15507) );
  NAND2_X1 U11339 ( .A1(n10991), .A2(n9922), .ZN(n15495) );
  CLKBUF_X1 U11340 ( .A(n15609), .Z(n15610) );
  CLKBUF_X1 U11341 ( .A(n15367), .Z(n15634) );
  OR2_X1 U11342 ( .A1(n15150), .A2(n10797), .ZN(n10798) );
  NOR2_X1 U11343 ( .A1(n9864), .A2(n12869), .ZN(n12871) );
  NOR2_X1 U11344 ( .A1(n19369), .A2(n19038), .ZN(n19037) );
  NAND2_X2 U11345 ( .A1(n19067), .A2(n18964), .ZN(n19174) );
  CLKBUF_X1 U11346 ( .A(n14028), .Z(n16322) );
  NAND2_X1 U11347 ( .A1(n10654), .A2(n10653), .ZN(n14173) );
  OAI21_X1 U11349 ( .B1(n16326), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10615), 
        .ZN(n10616) );
  AND2_X1 U11350 ( .A1(n16823), .A2(n12259), .ZN(n17675) );
  NAND2_X2 U11351 ( .A1(n21381), .A2(n15373), .ZN(n17250) );
  BUF_X1 U11352 ( .A(n12923), .Z(n9818) );
  CLKBUF_X2 U11353 ( .A(n12815), .Z(n15194) );
  INV_X2 U11354 ( .A(n19008), .ZN(n19119) );
  OR2_X1 U11355 ( .A1(n15398), .A2(n13587), .ZN(n10011) );
  OR2_X1 U11356 ( .A1(n18706), .A2(n13332), .ZN(n13308) );
  BUF_X2 U11357 ( .A(n11546), .Z(n12074) );
  NAND2_X1 U11358 ( .A1(n12647), .A2(n13984), .ZN(n14116) );
  NOR4_X2 U11359 ( .A1(n13475), .A2(n16984), .A3(n13466), .A4(n17087), .ZN(
        n19996) );
  INV_X1 U11360 ( .A(n18732), .ZN(n19552) );
  OR2_X1 U11361 ( .A1(n12779), .A2(n12732), .ZN(n13866) );
  AND2_X1 U11362 ( .A1(n13777), .A2(n12273), .ZN(n13776) );
  NAND2_X1 U11363 ( .A1(n15373), .A2(n14049), .ZN(n10484) );
  INV_X1 U11364 ( .A(n11790), .ZN(n12273) );
  INV_X1 U11365 ( .A(n11444), .ZN(n11494) );
  NAND2_X1 U11366 ( .A1(n11418), .A2(n11417), .ZN(n11444) );
  CLKBUF_X3 U11367 ( .A(n13313), .Z(n9795) );
  CLKBUF_X3 U11368 ( .A(n13295), .Z(n9793) );
  CLKBUF_X2 U11369 ( .A(n10709), .Z(n11140) );
  CLKBUF_X2 U11370 ( .A(n10558), .Z(n11164) );
  CLKBUF_X2 U11371 ( .A(n10439), .Z(n11088) );
  CLKBUF_X2 U11372 ( .A(n10392), .Z(n11163) );
  INV_X2 U11373 ( .A(n19529), .ZN(n9790) );
  BUF_X2 U11374 ( .A(n10445), .Z(n9815) );
  CLKBUF_X2 U11375 ( .A(n10539), .Z(n11158) );
  BUF_X2 U11376 ( .A(n10445), .Z(n9816) );
  CLKBUF_X2 U11377 ( .A(n11607), .Z(n9821) );
  NAND2_X1 U11379 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20006) );
  NOR2_X4 U11380 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10366) );
  XNOR2_X1 U11381 ( .A(n10093), .B(n16623), .ZN(n16798) );
  XNOR2_X1 U11382 ( .A(n15744), .B(n15743), .ZN(n17316) );
  AND2_X1 U11383 ( .A1(n16568), .A2(n9993), .ZN(n12554) );
  AND2_X1 U11384 ( .A1(n9966), .A2(n9965), .ZN(n15744) );
  OAI21_X1 U11385 ( .B1(n12586), .B2(n17566), .A(n12569), .ZN(n12570) );
  OR2_X1 U11386 ( .A1(n12506), .A2(n17566), .ZN(n12182) );
  OR2_X1 U11387 ( .A1(n16559), .A2(n12868), .ZN(n12885) );
  NOR2_X1 U11388 ( .A1(n10241), .A2(n10240), .ZN(n10239) );
  NOR2_X1 U11389 ( .A1(n16674), .A2(n16673), .ZN(n16672) );
  NAND3_X1 U11390 ( .A1(n16412), .A2(n10292), .A3(n16421), .ZN(n16419) );
  AND2_X1 U11391 ( .A1(n16873), .A2(n17512), .ZN(n17527) );
  NAND2_X1 U11392 ( .A1(n10255), .A2(n9877), .ZN(n12629) );
  OR2_X1 U11393 ( .A1(n13145), .A2(n13144), .ZN(n10336) );
  XNOR2_X1 U11394 ( .A(n15420), .B(n15419), .ZN(n15649) );
  XNOR2_X1 U11395 ( .A(n12534), .B(n12533), .ZN(n17465) );
  XNOR2_X1 U11396 ( .A(n12523), .B(n12522), .ZN(n13218) );
  OR2_X1 U11397 ( .A1(n16405), .A2(n16404), .ZN(n12523) );
  AND2_X1 U11398 ( .A1(n9963), .A2(n9801), .ZN(n11280) );
  AOI21_X1 U11399 ( .B1(n10213), .B2(n9873), .A(n10209), .ZN(n18859) );
  OR2_X1 U11400 ( .A1(n13123), .A2(n13124), .ZN(n13125) );
  AOI21_X1 U11401 ( .B1(n9985), .B2(n16288), .A(n11276), .ZN(n11277) );
  AND2_X1 U11402 ( .A1(n9954), .A2(n10214), .ZN(n18849) );
  NAND2_X1 U11403 ( .A1(n10261), .A2(n10259), .ZN(n15343) );
  NAND2_X1 U11404 ( .A1(n10165), .A2(n10164), .ZN(n13657) );
  INV_X1 U11405 ( .A(n16379), .ZN(n10165) );
  NOR2_X1 U11406 ( .A1(n18864), .A2(n13358), .ZN(n17111) );
  NAND2_X1 U11407 ( .A1(n13360), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18863) );
  NAND2_X1 U11408 ( .A1(n9949), .A2(n11824), .ZN(n15243) );
  NAND2_X1 U11409 ( .A1(n10167), .A2(n10166), .ZN(n16379) );
  AOI21_X1 U11410 ( .B1(n12546), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12545), .ZN(n12547) );
  INV_X1 U11411 ( .A(n16393), .ZN(n10167) );
  OR2_X1 U11412 ( .A1(n12578), .A2(n12580), .ZN(n17416) );
  XNOR2_X1 U11413 ( .A(n12540), .B(n12539), .ZN(n16369) );
  OR2_X1 U11414 ( .A1(n16474), .A2(n16473), .ZN(n17414) );
  NAND2_X1 U11415 ( .A1(n10244), .A2(n10243), .ZN(n15598) );
  NOR2_X1 U11416 ( .A1(n18895), .A2(n13356), .ZN(n13357) );
  AOI21_X1 U11417 ( .B1(n10263), .B2(n10260), .A(n9884), .ZN(n10259) );
  NAND2_X1 U11418 ( .A1(n14417), .A2(n14516), .ZN(n14514) );
  NOR4_X1 U11419 ( .A1(n19219), .A2(n17742), .A3(n18925), .A4(n17741), .ZN(
        n17747) );
  NOR2_X1 U11420 ( .A1(n16503), .A2(n10198), .ZN(n16474) );
  OR2_X1 U11421 ( .A1(n16513), .A2(n16501), .ZN(n16503) );
  INV_X1 U11422 ( .A(n19174), .ZN(n19209) );
  NAND2_X1 U11423 ( .A1(n10726), .A2(n10725), .ZN(n14516) );
  OR2_X1 U11424 ( .A1(n16288), .A2(n11268), .ZN(n11269) );
  XNOR2_X1 U11425 ( .A(n11244), .B(n10730), .ZN(n11253) );
  NAND2_X1 U11426 ( .A1(n10728), .A2(n10727), .ZN(n11244) );
  OR2_X1 U11427 ( .A1(n10728), .A2(n10727), .ZN(n11243) );
  INV_X4 U11428 ( .A(n19126), .ZN(n19062) );
  AOI21_X1 U11429 ( .B1(n19007), .B2(n18900), .A(n13350), .ZN(n13351) );
  NAND2_X1 U11430 ( .A1(n10665), .A2(n10664), .ZN(n14168) );
  AND3_X1 U11431 ( .A1(n13348), .A2(n13346), .A3(n9955), .ZN(n18998) );
  XNOR2_X1 U11432 ( .A(n10708), .B(n10698), .ZN(n11231) );
  OAI22_X1 U11433 ( .A1(n11727), .A2(n11640), .B1(n11728), .B2(n11639), .ZN(
        n11641) );
  NOR2_X2 U11434 ( .A1(n19555), .A2(n17894), .ZN(n19061) );
  OAI21_X2 U11435 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19542), .A(n17894), 
        .ZN(n19212) );
  NAND2_X1 U11436 ( .A1(n11584), .A2(n11583), .ZN(n16972) );
  NAND2_X1 U11437 ( .A1(n10252), .A2(n9913), .ZN(n10708) );
  NAND2_X1 U11438 ( .A1(n19116), .A2(n17100), .ZN(n13347) );
  NAND2_X1 U11439 ( .A1(n13997), .A2(n13996), .ZN(n13995) );
  NOR2_X1 U11440 ( .A1(n14937), .A2(n14938), .ZN(n15231) );
  NAND2_X1 U11441 ( .A1(n9861), .A2(n9970), .ZN(n20865) );
  NAND2_X1 U11442 ( .A1(n10630), .A2(n10629), .ZN(n13997) );
  AND2_X1 U11443 ( .A1(n12915), .A2(n12927), .ZN(n13897) );
  NOR2_X1 U11444 ( .A1(n11578), .A2(n16918), .ZN(n11638) );
  NOR2_X1 U11445 ( .A1(n19138), .A2(n10223), .ZN(n19026) );
  NOR2_X1 U11446 ( .A1(n16902), .A2(n17624), .ZN(n16884) );
  NAND2_X1 U11447 ( .A1(n14155), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14156) );
  OR2_X1 U11448 ( .A1(n12914), .A2(n12913), .ZN(n12915) );
  OR2_X1 U11449 ( .A1(n13341), .A2(n10224), .ZN(n10223) );
  CLKBUF_X1 U11450 ( .A(n14085), .Z(n15176) );
  AOI21_X1 U11451 ( .B1(n13901), .B2(n13900), .A(n12926), .ZN(n13898) );
  NOR2_X1 U11452 ( .A1(n18448), .A2(n18081), .ZN(n18424) );
  XNOR2_X1 U11453 ( .A(n16932), .B(n12924), .ZN(n13901) );
  AOI21_X1 U11454 ( .B1(n12923), .B2(n14011), .A(n12922), .ZN(n13900) );
  NAND2_X2 U11455 ( .A1(n15733), .A2(n13998), .ZN(n15739) );
  AND2_X1 U11456 ( .A1(n10547), .A2(n10546), .ZN(n11187) );
  INV_X1 U11457 ( .A(n20004), .ZN(n15393) );
  OAI21_X1 U11458 ( .B1(n19154), .B2(n10217), .A(n10216), .ZN(n19146) );
  AND2_X2 U11459 ( .A1(n17312), .A2(n11345), .ZN(n14161) );
  CLKBUF_X1 U11460 ( .A(n19398), .Z(n19443) );
  AND2_X1 U11461 ( .A1(n13985), .A2(n13714), .ZN(n21539) );
  AND2_X1 U11462 ( .A1(n13580), .A2(n13931), .ZN(n10172) );
  OR2_X1 U11463 ( .A1(n10053), .A2(n9890), .ZN(n13985) );
  AND2_X1 U11464 ( .A1(n14977), .A2(n12693), .ZN(n14979) );
  INV_X1 U11465 ( .A(n16377), .ZN(n10166) );
  INV_X1 U11466 ( .A(n12615), .ZN(n10164) );
  NOR2_X1 U11467 ( .A1(n12295), .A2(n10179), .ZN(n10181) );
  NAND2_X1 U11468 ( .A1(n11545), .A2(n11544), .ZN(n12036) );
  NAND2_X1 U11469 ( .A1(n11533), .A2(n11532), .ZN(n11539) );
  INV_X1 U11470 ( .A(n10177), .ZN(n12294) );
  OR2_X1 U11471 ( .A1(n14151), .A2(n14150), .ZN(n14373) );
  NAND2_X1 U11472 ( .A1(n12227), .A2(n12204), .ZN(n17709) );
  AOI21_X1 U11473 ( .B1(n11516), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10345), 
        .ZN(n11519) );
  AND2_X1 U11474 ( .A1(n10513), .A2(n10507), .ZN(n10506) );
  NOR2_X1 U11475 ( .A1(n11520), .A2(n10354), .ZN(n11531) );
  XNOR2_X1 U11476 ( .A(n13327), .B(n13326), .ZN(n19183) );
  NOR2_X1 U11477 ( .A1(n11799), .A2(n11798), .ZN(n11870) );
  AND4_X1 U11478 ( .A1(n10526), .A2(n10525), .A3(n12777), .A4(n10524), .ZN(
        n10527) );
  AND2_X1 U11479 ( .A1(n13761), .A2(n13762), .ZN(n13760) );
  MUX2_X1 U11480 ( .A(n10517), .B(n10516), .S(n12662), .Z(n10528) );
  NOR2_X1 U11481 ( .A1(n10269), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10266) );
  INV_X2 U11482 ( .A(n12045), .ZN(n12524) );
  AND4_X1 U11483 ( .A1(n12650), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n21523), 
        .A4(n10522), .ZN(n10525) );
  NOR2_X1 U11484 ( .A1(n17189), .A2(n10076), .ZN(n18577) );
  NOR2_X1 U11485 ( .A1(n18712), .A2(n13509), .ZN(n13329) );
  AOI21_X1 U11486 ( .B1(n11535), .B2(P2_EBX_REG_1__SCAN_IN), .A(n10327), .ZN(
        n11505) );
  AND2_X1 U11487 ( .A1(n10490), .A2(n10519), .ZN(n11341) );
  AND2_X1 U11488 ( .A1(n10077), .A2(n17094), .ZN(n16987) );
  NAND2_X1 U11489 ( .A1(n18624), .A2(n19552), .ZN(n13466) );
  XNOR2_X1 U11490 ( .A(n13496), .B(n18716), .ZN(n13309) );
  AND2_X1 U11491 ( .A1(n10501), .A2(n11340), .ZN(n10502) );
  AND2_X1 U11492 ( .A1(n11503), .A2(n9856), .ZN(n11535) );
  AND3_X1 U11493 ( .A1(n9975), .A2(n9974), .A3(n9973), .ZN(n10500) );
  AND2_X1 U11494 ( .A1(n12208), .A2(n13777), .ZN(n11468) );
  AND2_X1 U11495 ( .A1(n11319), .A2(n11320), .ZN(n10036) );
  NAND2_X1 U11496 ( .A1(n13462), .A2(n19571), .ZN(n17087) );
  INV_X1 U11497 ( .A(n18716), .ZN(n13497) );
  AND2_X1 U11498 ( .A1(n13491), .A2(n19993), .ZN(n10077) );
  AND2_X1 U11499 ( .A1(n10489), .A2(n15373), .ZN(n10519) );
  AND3_X1 U11500 ( .A1(n13284), .A2(n10204), .A3(n13277), .ZN(n18716) );
  NAND2_X4 U11501 ( .A1(n9829), .A2(n17714), .ZN(n11789) );
  OR2_X1 U11502 ( .A1(n11687), .A2(n11686), .ZN(n11793) );
  NOR2_X1 U11503 ( .A1(n19584), .A2(n19564), .ZN(n13491) );
  INV_X1 U11504 ( .A(n13463), .ZN(n19571) );
  NOR2_X2 U11505 ( .A1(n12648), .A2(n21439), .ZN(n11338) );
  NAND2_X1 U11507 ( .A1(n11494), .A2(n12273), .ZN(n12211) );
  NOR2_X1 U11508 ( .A1(n19568), .A2(n13462), .ZN(n19993) );
  INV_X2 U11509 ( .A(n11612), .ZN(n11624) );
  INV_X1 U11510 ( .A(n10494), .ZN(n14058) );
  NOR2_X1 U11511 ( .A1(n13400), .A2(n13399), .ZN(n19564) );
  NOR2_X1 U11512 ( .A1(n13460), .A2(n13459), .ZN(n19568) );
  OR2_X1 U11513 ( .A1(n13429), .A2(n13430), .ZN(n13462) );
  NAND2_X2 U11514 ( .A1(n11430), .A2(n11429), .ZN(n11790) );
  OR2_X1 U11515 ( .A1(n10564), .A2(n10563), .ZN(n11266) );
  OR2_X2 U11516 ( .A1(n10451), .A2(n10450), .ZN(n14069) );
  AND4_X1 U11517 ( .A1(n10470), .A2(n9871), .A3(n10469), .A4(n10333), .ZN(
        n10494) );
  OR2_X2 U11518 ( .A1(n10483), .A2(n10482), .ZN(n15373) );
  OR2_X2 U11519 ( .A1(n10377), .A2(n10376), .ZN(n14049) );
  NAND2_X1 U11520 ( .A1(n11379), .A2(n11378), .ZN(n11471) );
  NAND2_X1 U11521 ( .A1(n11384), .A2(n10335), .ZN(n11394) );
  AND4_X1 U11522 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10415) );
  AND4_X1 U11523 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10435) );
  AND4_X1 U11524 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10417) );
  AND4_X1 U11525 ( .A1(n10426), .A2(n10425), .A3(n10424), .A4(n10423), .ZN(
        n10437) );
  AND4_X1 U11526 ( .A1(n10410), .A2(n10409), .A3(n10408), .A4(n10407), .ZN(
        n10416) );
  AND4_X1 U11527 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n10438) );
  AND4_X1 U11528 ( .A1(n11440), .A2(n11439), .A3(n11438), .A4(n11437), .ZN(
        n11441) );
  INV_X1 U11529 ( .A(n18486), .ZN(n18455) );
  AOI22_X1 U11530 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10381) );
  AND4_X1 U11531 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10418) );
  AND4_X1 U11532 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        n10436) );
  INV_X2 U11533 ( .A(n17881), .ZN(U215) );
  INV_X2 U11534 ( .A(n20073), .ZN(n20138) );
  NAND2_X1 U11535 ( .A1(n9997), .A2(n9996), .ZN(n18453) );
  BUF_X2 U11536 ( .A(n13296), .Z(n18498) );
  BUF_X4 U11537 ( .A(n13394), .Z(n18518) );
  BUF_X2 U11538 ( .A(n10754), .Z(n11002) );
  AND3_X1 U11539 ( .A1(n11432), .A2(n11431), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U11540 ( .A1(n9824), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9822), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11439) );
  NAND2_X2 U11541 ( .A1(n20217), .A2(n15401), .ZN(n19529) );
  INV_X2 U11542 ( .A(n9810), .ZN(n9811) );
  NAND2_X2 U11543 ( .A1(n21244), .A2(n21112), .ZN(n21163) );
  NAND2_X2 U11544 ( .A1(n9791), .A2(n17691), .ZN(n13067) );
  AND2_X2 U11545 ( .A1(n11600), .A2(n11601), .ZN(n11650) );
  INV_X1 U11546 ( .A(n17067), .ZN(n13389) );
  BUF_X4 U11547 ( .A(n13314), .Z(n9794) );
  OR2_X2 U11548 ( .A1(n11347), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17352) );
  AND2_X1 U11549 ( .A1(n10364), .A2(n10368), .ZN(n10452) );
  INV_X2 U11550 ( .A(n20195), .ZN(n20129) );
  OR2_X1 U11551 ( .A1(n13224), .A2(n13228), .ZN(n9850) );
  AND2_X1 U11552 ( .A1(n10367), .A2(n13868), .ZN(n10754) );
  INV_X2 U11553 ( .A(n17884), .ZN(n17886) );
  AND2_X2 U11554 ( .A1(n11355), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11607) );
  AND2_X2 U11555 ( .A1(n16936), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11455) );
  AND3_X2 U11556 ( .A1(n17686), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13039) );
  AND2_X1 U11557 ( .A1(n16927), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15190) );
  AND2_X2 U11558 ( .A1(n16935), .A2(n16927), .ZN(n13040) );
  NAND2_X1 U11559 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20169), .ZN(
        n13223) );
  OR2_X1 U11560 ( .A1(n20177), .A2(n13228), .ZN(n15404) );
  AND2_X2 U11561 ( .A1(n10591), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10364) );
  AND2_X1 U11562 ( .A1(n17127), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10359) );
  NAND2_X1 U11563 ( .A1(n20177), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13224) );
  NOR2_X1 U11564 ( .A1(n10620), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10367) );
  NOR2_X1 U11565 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10371) );
  NOR2_X2 U11566 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13868) );
  INV_X1 U11567 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17127) );
  INV_X1 U11568 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10591) );
  AND2_X1 U11569 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14091) );
  NOR2_X1 U11570 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U11571 ( .A1(n11511), .A2(n10057), .ZN(n11558) );
  AND2_X1 U11572 ( .A1(n11614), .A2(n11613), .ZN(n9796) );
  NAND2_X2 U11574 ( .A1(n15323), .A2(n10798), .ZN(n15335) );
  INV_X1 U11575 ( .A(n18906), .ZN(n9797) );
  NOR2_X4 U11576 ( .A1(n13227), .A2(n13226), .ZN(n13311) );
  OR2_X1 U11577 ( .A1(n11612), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12537) );
  INV_X2 U11578 ( .A(n11612), .ZN(n9829) );
  AND2_X2 U11579 ( .A1(n16936), .A2(n16927), .ZN(n9813) );
  AND2_X2 U11580 ( .A1(n16936), .A2(n16927), .ZN(n13042) );
  NAND2_X1 U11581 ( .A1(n11508), .A2(n11507), .ZN(n11511) );
  AND2_X2 U11582 ( .A1(n12847), .A2(n15199), .ZN(n12489) );
  INV_X1 U11583 ( .A(n11467), .ZN(n12272) );
  OAI22_X2 U11584 ( .A1(n17086), .A2(n19511), .B1(n17085), .B2(n19983), .ZN(
        n20036) );
  NOR2_X4 U11585 ( .A1(n20006), .A2(n13228), .ZN(n17067) );
  NAND2_X1 U11586 ( .A1(n11999), .A2(n11998), .ZN(n9798) );
  NAND2_X1 U11587 ( .A1(n11519), .A2(n11518), .ZN(n9799) );
  NAND2_X1 U11588 ( .A1(n13903), .A2(n10304), .ZN(n9800) );
  NAND2_X1 U11589 ( .A1(n13903), .A2(n10304), .ZN(n10303) );
  NAND2_X1 U11590 ( .A1(n11519), .A2(n11518), .ZN(n11550) );
  NOR2_X2 U11591 ( .A1(n18484), .A2(n18483), .ZN(n18482) );
  NOR3_X2 U11592 ( .A1(n18335), .A2(n18282), .A3(n10074), .ZN(n18331) );
  NAND4_X2 U11593 ( .A1(n12215), .A2(n20573), .A3(n13778), .A4(n12273), .ZN(
        n11502) );
  NAND2_X2 U11594 ( .A1(n11462), .A2(n11461), .ZN(n11612) );
  NOR2_X4 U11595 ( .A1(n13966), .A2(n13968), .ZN(n13969) );
  NAND2_X1 U11596 ( .A1(n18948), .A2(n13353), .ZN(n18913) );
  NAND2_X1 U11597 ( .A1(n9887), .A2(n18957), .ZN(n18896) );
  NAND2_X1 U11598 ( .A1(n11999), .A2(n11998), .ZN(n16547) );
  AOI22_X1 U11599 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11637), .B1(
        n11723), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11643) );
  NOR2_X1 U11600 ( .A1(n11586), .A2(n9970), .ZN(n10308) );
  NAND2_X1 U11601 ( .A1(n11441), .A2(n17691), .ZN(n11442) );
  NOR2_X1 U11602 ( .A1(n19211), .A2(n19201), .ZN(n19200) );
  OR2_X1 U11603 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  XNOR2_X2 U11604 ( .A(n15150), .B(n10796), .ZN(n15322) );
  NAND2_X2 U11605 ( .A1(n14887), .A2(n9909), .ZN(n15150) );
  NOR2_X4 U11606 ( .A1(n14514), .A2(n14888), .ZN(n14887) );
  NOR2_X2 U11607 ( .A1(n14415), .A2(n14416), .ZN(n14417) );
  AND2_X4 U11608 ( .A1(n13868), .A2(n10368), .ZN(n10476) );
  AND2_X1 U11609 ( .A1(n10273), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9801) );
  INV_X1 U11610 ( .A(n11263), .ZN(n9802) );
  NAND2_X1 U11611 ( .A1(n9803), .A2(n11264), .ZN(n10261) );
  NOR2_X1 U11612 ( .A1(n10262), .A2(n9802), .ZN(n9803) );
  XNOR2_X1 U11613 ( .A(n11213), .B(n11201), .ZN(n9804) );
  XNOR2_X1 U11614 ( .A(n11197), .B(n14156), .ZN(n9805) );
  NOR2_X1 U11615 ( .A1(n12633), .A2(n12789), .ZN(n9806) );
  INV_X1 U11616 ( .A(n14562), .ZN(n9807) );
  XNOR2_X1 U11617 ( .A(n11213), .B(n11201), .ZN(n14127) );
  XNOR2_X1 U11618 ( .A(n11197), .B(n14156), .ZN(n14134) );
  NOR2_X1 U11619 ( .A1(n12633), .A2(n12789), .ZN(n12773) );
  XNOR2_X1 U11620 ( .A(n10633), .B(n10632), .ZN(n11193) );
  INV_X1 U11621 ( .A(n12171), .ZN(n9808) );
  OAI21_X1 U11622 ( .B1(n11963), .B2(n10064), .A(n10062), .ZN(n9809) );
  INV_X1 U11623 ( .A(n13038), .ZN(n9810) );
  OAI21_X1 U11624 ( .B1(n11963), .B2(n10064), .A(n10062), .ZN(n16588) );
  AND3_X1 U11625 ( .A1(n11523), .A2(n11528), .A3(n11527), .ZN(n11530) );
  AND2_X1 U11626 ( .A1(n16936), .A2(n16927), .ZN(n9812) );
  NAND2_X2 U11627 ( .A1(n11476), .A2(n11474), .ZN(n12019) );
  INV_X2 U11628 ( .A(n11881), .ZN(n13570) );
  AND2_X1 U11629 ( .A1(n17714), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n21227) );
  AND2_X4 U11630 ( .A1(n10364), .A2(n10366), .ZN(n10444) );
  AND2_X1 U11631 ( .A1(n13868), .A2(n10366), .ZN(n10445) );
  NOR2_X4 U11632 ( .A1(n20416), .A2(n20417), .ZN(n15211) );
  NAND2_X1 U11633 ( .A1(n9880), .A2(n9948), .ZN(n14014) );
  NAND2_X1 U11634 ( .A1(n9947), .A2(n9948), .ZN(n20587) );
  NOR2_X4 U11635 ( .A1(n19351), .A2(n19028), .ZN(n19347) );
  INV_X2 U11636 ( .A(n9862), .ZN(n9817) );
  OR2_X1 U11637 ( .A1(n13227), .A2(n20006), .ZN(n9862) );
  NAND2_X2 U11638 ( .A1(n10313), .A2(n11907), .ZN(n17534) );
  XNOR2_X1 U11639 ( .A(n11558), .B(n11557), .ZN(n12923) );
  INV_X2 U11640 ( .A(n11716), .ZN(n11834) );
  NAND2_X2 U11642 ( .A1(n11979), .A2(n11980), .ZN(n16564) );
  NAND2_X1 U11643 ( .A1(n11444), .A2(n11790), .ZN(n12210) );
  BUF_X4 U11644 ( .A(n13040), .Z(n9822) );
  BUF_X8 U11645 ( .A(n13040), .Z(n9823) );
  NAND2_X4 U11646 ( .A1(n11443), .A2(n11442), .ZN(n11463) );
  AND2_X1 U11647 ( .A1(n11600), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9824) );
  NAND3_X2 U11648 ( .A1(n11479), .A2(n11478), .A3(n11523), .ZN(n11517) );
  NAND2_X2 U11649 ( .A1(n10308), .A2(n9818), .ZN(n11704) );
  NOR2_X4 U11650 ( .A1(n15495), .A2(n15497), .ZN(n15482) );
  NOR2_X2 U11651 ( .A1(n20573), .A2(n11481), .ZN(n12216) );
  OR2_X2 U11652 ( .A1(n16588), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11979) );
  AND2_X1 U11653 ( .A1(n10365), .A2(n10359), .ZN(n9825) );
  AND2_X1 U11654 ( .A1(n10365), .A2(n10359), .ZN(n9826) );
  AND2_X1 U11655 ( .A1(n10364), .A2(n10368), .ZN(n9827) );
  AND2_X1 U11656 ( .A1(n10364), .A2(n10368), .ZN(n9828) );
  XNOR2_X2 U11657 ( .A(n12169), .B(n12170), .ZN(n12160) );
  OR2_X1 U11658 ( .A1(n11193), .A2(n11218), .ZN(n11196) );
  INV_X4 U11659 ( .A(n11624), .ZN(n20547) );
  NOR2_X4 U11660 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16935) );
  XNOR2_X2 U11661 ( .A(n11872), .B(n15240), .ZN(n15242) );
  NAND2_X2 U11662 ( .A1(n11801), .A2(n20362), .ZN(n11872) );
  NOR2_X1 U11663 ( .A1(n11463), .A2(n17682), .ZN(n10094) );
  NAND2_X1 U11664 ( .A1(n10497), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10513) );
  AOI21_X1 U11665 ( .B1(n11534), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11506), .ZN(n11509) );
  NOR2_X1 U11666 ( .A1(n10282), .A2(n15462), .ZN(n10281) );
  INV_X1 U11667 ( .A(n15472), .ZN(n10282) );
  NAND2_X1 U11668 ( .A1(n15765), .A2(n11288), .ZN(n9965) );
  NAND2_X1 U11669 ( .A1(n12773), .A2(n9958), .ZN(n9957) );
  OR2_X1 U11670 ( .A1(n17165), .A2(n12635), .ZN(n9958) );
  INV_X1 U11671 ( .A(n19568), .ZN(n16984) );
  NAND2_X1 U11672 ( .A1(n18896), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9951) );
  NOR2_X1 U11673 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10369), .ZN(
        n10370) );
  NAND2_X1 U11674 ( .A1(n10484), .A2(n10505), .ZN(n9973) );
  NOR2_X1 U11675 ( .A1(n11502), .A2(n12240), .ZN(n11503) );
  AOI21_X1 U11676 ( .B1(n16598), .B2(n10311), .A(n9881), .ZN(n10310) );
  INV_X1 U11677 ( .A(n16605), .ZN(n10311) );
  INV_X1 U11678 ( .A(n16598), .ZN(n10312) );
  AND2_X1 U11679 ( .A1(n9856), .A2(n12206), .ZN(n11546) );
  INV_X1 U11680 ( .A(n15483), .ZN(n11109) );
  INV_X1 U11681 ( .A(n14993), .ZN(n10258) );
  INV_X1 U11682 ( .A(n15091), .ZN(n10749) );
  NOR2_X1 U11683 ( .A1(n15373), .A2(n21441), .ZN(n10659) );
  NAND2_X1 U11684 ( .A1(n10641), .A2(n10640), .ZN(n14113) );
  AND2_X1 U11685 ( .A1(n9844), .A2(n17441), .ZN(n10227) );
  NAND2_X1 U11686 ( .A1(n11624), .A2(n12898), .ZN(n13160) );
  INV_X1 U11687 ( .A(n11534), .ZN(n12042) );
  OAI21_X1 U11688 ( .B1(n17427), .B2(n11996), .A(n16576), .ZN(n12552) );
  AND2_X1 U11689 ( .A1(n10084), .A2(n12179), .ZN(n10081) );
  NAND2_X1 U11690 ( .A1(n17534), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9943) );
  NOR2_X1 U11691 ( .A1(n13227), .A2(n13224), .ZN(n13313) );
  NOR2_X1 U11692 ( .A1(n18453), .A2(n13274), .ZN(n10207) );
  NOR2_X1 U11693 ( .A1(n13225), .A2(n13224), .ZN(n13296) );
  NAND2_X1 U11694 ( .A1(n10203), .A2(n13357), .ZN(n13359) );
  INV_X1 U11695 ( .A(n13479), .ZN(n10010) );
  INV_X1 U11696 ( .A(n18794), .ZN(n13587) );
  NOR2_X1 U11697 ( .A1(n13473), .A2(n10006), .ZN(n15396) );
  NAND2_X1 U11698 ( .A1(n10007), .A2(n9874), .ZN(n10006) );
  INV_X1 U11699 ( .A(n18721), .ZN(n13496) );
  INV_X1 U11700 ( .A(n10487), .ZN(n15374) );
  OAI21_X1 U11701 ( .B1(n11174), .B2(n15746), .A(n11153), .ZN(n15462) );
  NAND2_X1 U11702 ( .A1(n12629), .A2(n16288), .ZN(n9966) );
  NAND2_X1 U11703 ( .A1(n12660), .A2(n13993), .ZN(n12795) );
  NAND2_X1 U11704 ( .A1(n10603), .A2(n10602), .ZN(n9956) );
  OR2_X1 U11705 ( .A1(n9830), .A2(n11193), .ZN(n14324) );
  NAND2_X1 U11706 ( .A1(n9917), .A2(n10351), .ZN(n10301) );
  NOR2_X1 U11707 ( .A1(n12932), .A2(n10305), .ZN(n10304) );
  INV_X1 U11708 ( .A(n12929), .ZN(n10305) );
  NAND2_X1 U11709 ( .A1(n16474), .A2(n12485), .ZN(n12540) );
  NAND2_X1 U11710 ( .A1(n12894), .A2(n20975), .ZN(n12920) );
  AND2_X1 U11711 ( .A1(n17682), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14011) );
  NAND2_X1 U11712 ( .A1(n21181), .A2(n21207), .ZN(n20971) );
  NOR2_X1 U11713 ( .A1(n20800), .A2(n21207), .ZN(n20943) );
  NAND2_X1 U11714 ( .A1(n10002), .A2(n10000), .ZN(n17191) );
  NOR2_X1 U11715 ( .A1(n17891), .A2(n10001), .ZN(n10000) );
  NAND2_X1 U11716 ( .A1(n20004), .A2(n10003), .ZN(n10002) );
  OAI221_X1 U11717 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n19119), 
        .C1(n19240), .C2(n13355), .A(n13354), .ZN(n18878) );
  INV_X1 U11718 ( .A(n20587), .ZN(n11626) );
  AND2_X2 U11719 ( .A1(n10358), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10365) );
  NAND2_X1 U11720 ( .A1(n11502), .A2(n11481), .ZN(n11469) );
  NOR2_X1 U11721 ( .A1(n12253), .A2(n17714), .ZN(n11488) );
  NAND2_X1 U11723 ( .A1(n10494), .A2(n10487), .ZN(n11189) );
  INV_X1 U11724 ( .A(n10632), .ZN(n10269) );
  NAND2_X1 U11725 ( .A1(n10500), .A2(n10485), .ZN(n12778) );
  OAI21_X1 U11726 ( .B1(n11306), .B2(n10042), .A(n10041), .ZN(n10040) );
  NAND2_X1 U11727 ( .A1(n11311), .A2(n11307), .ZN(n10041) );
  INV_X1 U11728 ( .A(n11308), .ZN(n10042) );
  INV_X1 U11729 ( .A(n11316), .ZN(n10038) );
  AND2_X1 U11730 ( .A1(n16775), .A2(n13655), .ZN(n10196) );
  INV_X1 U11731 ( .A(n11751), .ZN(n10325) );
  NAND2_X1 U11732 ( .A1(n10321), .A2(n10322), .ZN(n10320) );
  NAND2_X1 U11733 ( .A1(n10106), .A2(n10102), .ZN(n10101) );
  INV_X1 U11734 ( .A(n14784), .ZN(n10102) );
  NOR2_X1 U11735 ( .A1(n19559), .A2(n19993), .ZN(n13472) );
  NOR2_X1 U11736 ( .A1(n18703), .A2(n13308), .ZN(n13338) );
  AND2_X1 U11737 ( .A1(n16121), .A2(n9984), .ZN(n15753) );
  NAND2_X1 U11738 ( .A1(n10274), .A2(n16096), .ZN(n9984) );
  NOR2_X1 U11739 ( .A1(n15533), .A2(n15611), .ZN(n10277) );
  NOR2_X1 U11740 ( .A1(n15626), .A2(n15635), .ZN(n10284) );
  NAND2_X1 U11741 ( .A1(n15369), .A2(n15368), .ZN(n15367) );
  AND2_X1 U11742 ( .A1(n15337), .A2(n15735), .ZN(n15336) );
  NAND2_X1 U11743 ( .A1(n13975), .A2(n14166), .ZN(n10257) );
  INV_X1 U11744 ( .A(n10656), .ZN(n10872) );
  NAND2_X1 U11745 ( .A1(n16156), .A2(n9964), .ZN(n11278) );
  NOR2_X1 U11746 ( .A1(n16272), .A2(n16280), .ZN(n9964) );
  NAND2_X1 U11747 ( .A1(n15343), .A2(n11271), .ZN(n9985) );
  INV_X1 U11748 ( .A(n15574), .ZN(n10246) );
  INV_X1 U11749 ( .A(n12747), .ZN(n12768) );
  OAI21_X1 U11750 ( .B1(n10053), .B2(n10052), .A(n10494), .ZN(n10051) );
  INV_X1 U11751 ( .A(n12637), .ZN(n10052) );
  OR2_X1 U11752 ( .A1(n10575), .A2(n10574), .ZN(n11206) );
  AND2_X1 U11753 ( .A1(n11909), .A2(n9923), .ZN(n11944) );
  NAND2_X1 U11754 ( .A1(n11909), .A2(n9842), .ZN(n11935) );
  NAND2_X1 U11755 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10137) );
  NOR2_X1 U11756 ( .A1(n17511), .A2(n10149), .ZN(n10148) );
  INV_X1 U11757 ( .A(n10154), .ZN(n10153) );
  AND2_X1 U11758 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10163) );
  XNOR2_X1 U11759 ( .A(n11540), .B(n11539), .ZN(n10078) );
  AOI21_X1 U11760 ( .B1(n12092), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11549), .ZN(n12038) );
  NAND2_X1 U11761 ( .A1(n11963), .A2(n9989), .ZN(n9987) );
  NOR2_X1 U11762 ( .A1(n10312), .A2(n9992), .ZN(n10065) );
  NAND2_X1 U11763 ( .A1(n12607), .A2(n16645), .ZN(n10113) );
  NAND2_X1 U11764 ( .A1(n10115), .A2(n16645), .ZN(n10114) );
  INV_X1 U11765 ( .A(n10114), .ZN(n10110) );
  NOR2_X1 U11766 ( .A1(n12606), .A2(n10116), .ZN(n10115) );
  INV_X1 U11767 ( .A(n16655), .ZN(n10116) );
  OAI21_X1 U11768 ( .B1(n16850), .B2(n12603), .A(n16853), .ZN(n16674) );
  NOR2_X1 U11769 ( .A1(n17599), .A2(n10185), .ZN(n10184) );
  INV_X1 U11770 ( .A(n15032), .ZN(n10185) );
  NAND2_X1 U11771 ( .A1(n11895), .A2(n10314), .ZN(n10313) );
  NOR2_X1 U11772 ( .A1(n10315), .A2(n16879), .ZN(n10314) );
  INV_X1 U11773 ( .A(n10085), .ZN(n10084) );
  OAI21_X1 U11774 ( .B1(n17551), .B2(n10086), .A(n9938), .ZN(n10085) );
  INV_X1 U11775 ( .A(n17550), .ZN(n9971) );
  INV_X1 U11776 ( .A(n13964), .ZN(n10171) );
  NOR2_X1 U11777 ( .A1(n17636), .A2(n10187), .ZN(n10186) );
  INV_X1 U11778 ( .A(n17649), .ZN(n10187) );
  NAND2_X1 U11779 ( .A1(n15227), .A2(n15224), .ZN(n12161) );
  NAND2_X1 U11780 ( .A1(n10100), .A2(n10105), .ZN(n10097) );
  AND4_X1 U11781 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11783) );
  NAND2_X1 U11782 ( .A1(n11805), .A2(n11804), .ZN(n9968) );
  NOR2_X1 U11783 ( .A1(n11624), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U11784 ( .A1(n9818), .A2(n9970), .ZN(n11585) );
  NAND2_X1 U11785 ( .A1(n11423), .A2(n17691), .ZN(n11430) );
  NAND2_X1 U11786 ( .A1(n11428), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11429) );
  NOR2_X1 U11787 ( .A1(n11796), .A2(n11787), .ZN(n11788) );
  NOR2_X1 U11788 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15404), .ZN(
        n13275) );
  AND2_X1 U11789 ( .A1(n19579), .A2(n13472), .ZN(n13465) );
  INV_X1 U11790 ( .A(n19564), .ZN(n13475) );
  NOR2_X1 U11791 ( .A1(n10340), .A2(n19008), .ZN(n13345) );
  INV_X1 U11792 ( .A(n13338), .ZN(n17784) );
  INV_X1 U11793 ( .A(n19994), .ZN(n10004) );
  NOR2_X1 U11794 ( .A1(n13420), .A2(n13419), .ZN(n13463) );
  NAND2_X1 U11795 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15586), .ZN(n15566) );
  NOR2_X1 U11796 ( .A1(n10767), .A2(n21275), .ZN(n10781) );
  INV_X1 U11797 ( .A(n21315), .ZN(n10033) );
  NOR2_X1 U11798 ( .A1(n15153), .A2(n10044), .ZN(n10043) );
  NAND2_X1 U11799 ( .A1(n10045), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U11800 ( .A1(n15164), .A2(n21441), .ZN(n15117) );
  OR2_X1 U11801 ( .A1(n15736), .A2(n10505), .ZN(n15370) );
  AND2_X1 U11802 ( .A1(n21441), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15421) );
  AND2_X1 U11803 ( .A1(n10281), .A2(n11109), .ZN(n10279) );
  NAND2_X1 U11804 ( .A1(n11103), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11129) );
  NOR2_X1 U11805 ( .A1(n15521), .A2(n10276), .ZN(n10275) );
  INV_X1 U11806 ( .A(n10277), .ZN(n10276) );
  AND2_X1 U11807 ( .A1(n11064), .A2(n11063), .ZN(n15508) );
  OR2_X1 U11808 ( .A1(n16117), .A2(n11174), .ZN(n11063) );
  NAND2_X1 U11809 ( .A1(n10731), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10750) );
  AND2_X1 U11810 ( .A1(n10722), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10731) );
  INV_X1 U11811 ( .A(n9965), .ZN(n12628) );
  AND2_X1 U11812 ( .A1(n11287), .A2(n15751), .ZN(n10254) );
  NOR2_X1 U11813 ( .A1(n12795), .A2(n13856), .ZN(n14615) );
  INV_X1 U11814 ( .A(n14615), .ZN(n16220) );
  NAND2_X1 U11815 ( .A1(n10595), .A2(n10594), .ZN(n10603) );
  NAND2_X1 U11816 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  NAND2_X1 U11817 ( .A1(n14085), .A2(n21439), .ZN(n10654) );
  NAND2_X1 U11818 ( .A1(n21438), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17167) );
  NAND2_X1 U11819 ( .A1(n12515), .A2(n11986), .ZN(n17427) );
  NAND2_X1 U11820 ( .A1(n11790), .A2(n11897), .ZN(n11984) );
  NAND2_X1 U11821 ( .A1(n15194), .A2(n12890), .ZN(n10139) );
  OR2_X1 U11822 ( .A1(n16385), .A2(n9918), .ZN(n10138) );
  OR2_X1 U11823 ( .A1(n16385), .A2(n16640), .ZN(n10140) );
  NAND2_X1 U11824 ( .A1(n13078), .A2(n10297), .ZN(n10294) );
  INV_X1 U11825 ( .A(n16443), .ZN(n10297) );
  INV_X1 U11826 ( .A(n13078), .ZN(n10295) );
  OR2_X1 U11827 ( .A1(n16519), .A2(n16521), .ZN(n10298) );
  NAND2_X1 U11828 ( .A1(n14357), .A2(n10180), .ZN(n10179) );
  INV_X1 U11829 ( .A(n14361), .ZN(n10180) );
  XNOR2_X1 U11830 ( .A(n12592), .B(n12591), .ZN(n12812) );
  NAND2_X1 U11831 ( .A1(n9799), .A2(n11551), .ZN(n11556) );
  AND2_X1 U11832 ( .A1(n9848), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10290) );
  NAND2_X1 U11833 ( .A1(n16580), .A2(n9848), .ZN(n12559) );
  OR3_X1 U11834 ( .A1(n17122), .A2(n11892), .A3(n16776), .ZN(n16605) );
  NOR2_X1 U11835 ( .A1(n12612), .A2(n12611), .ZN(n16620) );
  INV_X1 U11836 ( .A(n10115), .ZN(n10112) );
  AND2_X1 U11837 ( .A1(n15031), .A2(n10184), .ZN(n17598) );
  NAND2_X1 U11838 ( .A1(n12148), .A2(n11892), .ZN(n10080) );
  INV_X1 U11839 ( .A(n10079), .ZN(n12148) );
  AOI21_X1 U11840 ( .B1(n14784), .B2(n12003), .A(n17662), .ZN(n10106) );
  NAND2_X1 U11841 ( .A1(n10079), .A2(n14784), .ZN(n10098) );
  NAND2_X1 U11842 ( .A1(n9968), .A2(n12152), .ZN(n10079) );
  XNOR2_X1 U11843 ( .A(n12294), .B(n12293), .ZN(n13741) );
  NAND2_X1 U11844 ( .A1(n13743), .A2(n9929), .ZN(n14360) );
  INV_X1 U11845 ( .A(n12295), .ZN(n10178) );
  NAND2_X1 U11846 ( .A1(n12900), .A2(n14011), .ZN(n12905) );
  INV_X1 U11847 ( .A(n20977), .ZN(n21023) );
  NAND2_X1 U11848 ( .A1(n17682), .A2(n14024), .ZN(n20977) );
  NOR2_X1 U11849 ( .A1(n17933), .A2(n18164), .ZN(n17926) );
  AND2_X1 U11850 ( .A1(n10118), .A2(n18224), .ZN(n17998) );
  NOR2_X1 U11851 ( .A1(n18668), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U11852 ( .A1(n13279), .A2(n13276), .ZN(n10208) );
  AOI21_X1 U11853 ( .B1(n9795), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(n10207), .ZN(n10206) );
  AND2_X1 U11854 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13266) );
  AOI21_X1 U11855 ( .B1(n18518), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(n9994), .ZN(n13268) );
  AOI22_X1 U11856 ( .A1(n16985), .A2(n16986), .B1(n16987), .B2(n19978), .ZN(
        n17189) );
  NAND3_X1 U11857 ( .A1(n13450), .A2(n13449), .A3(n13448), .ZN(n18732) );
  AND2_X1 U11858 ( .A1(n10348), .A2(n10123), .ZN(n10122) );
  NOR2_X1 U11859 ( .A1(n18073), .A2(n10124), .ZN(n10123) );
  NAND2_X1 U11860 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10124) );
  INV_X1 U11861 ( .A(n19138), .ZN(n10225) );
  NOR2_X1 U11862 ( .A1(n13377), .A2(n13376), .ZN(n20205) );
  NAND2_X1 U11863 ( .A1(n10201), .A2(n10202), .ZN(n10203) );
  NAND2_X1 U11864 ( .A1(n10220), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10217) );
  NAND2_X1 U11865 ( .A1(n13335), .A2(n10220), .ZN(n10216) );
  INV_X1 U11866 ( .A(n19147), .ZN(n10220) );
  OR2_X1 U11867 ( .A1(n19154), .A2(n19480), .ZN(n10219) );
  NOR2_X1 U11868 ( .A1(n19182), .A2(n13328), .ZN(n19173) );
  NOR2_X1 U11869 ( .A1(n19200), .A2(n13324), .ZN(n19191) );
  XNOR2_X1 U11870 ( .A(n18721), .B(n9952), .ZN(n19201) );
  INV_X1 U11871 ( .A(n20205), .ZN(n19555) );
  OAI21_X1 U11872 ( .B1(n15447), .B2(n21277), .A(n15441), .ZN(n10240) );
  NOR2_X1 U11873 ( .A1(n10242), .A2(n21513), .ZN(n10241) );
  INV_X1 U11874 ( .A(n15457), .ZN(n10242) );
  NAND2_X1 U11875 ( .A1(n15541), .A2(n9942), .ZN(n15456) );
  NOR2_X1 U11876 ( .A1(n21505), .A2(n21509), .ZN(n10023) );
  NOR2_X1 U11877 ( .A1(n17205), .A2(n17195), .ZN(n15541) );
  NAND2_X1 U11878 ( .A1(n9867), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n17243) );
  INV_X1 U11879 ( .A(n21308), .ZN(n21343) );
  OR3_X1 U11880 ( .A1(n15153), .A2(n17163), .A3(n15102), .ZN(n21296) );
  NAND2_X1 U11881 ( .A1(n12771), .A2(n12770), .ZN(n10243) );
  NAND2_X1 U11882 ( .A1(n12772), .A2(n10245), .ZN(n10244) );
  AND2_X1 U11883 ( .A1(n15733), .A2(n15375), .ZN(n15719) );
  INV_X1 U11884 ( .A(n15733), .ZN(n15736) );
  OR2_X1 U11885 ( .A1(n15763), .A2(n17306), .ZN(n9979) );
  XNOR2_X1 U11886 ( .A(n9981), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17322) );
  NAND2_X1 U11887 ( .A1(n9983), .A2(n9982), .ZN(n9981) );
  INV_X1 U11888 ( .A(n15755), .ZN(n9982) );
  NAND2_X1 U11889 ( .A1(n15757), .A2(n15756), .ZN(n9983) );
  INV_X1 U11890 ( .A(n14161), .ZN(n15759) );
  NAND2_X1 U11891 ( .A1(n15744), .A2(n12630), .ZN(n12631) );
  OAI21_X1 U11892 ( .B1(n17336), .B2(n10056), .A(n10055), .ZN(n17320) );
  NAND2_X1 U11893 ( .A1(n11288), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10056) );
  NOR2_X1 U11894 ( .A1(n17368), .A2(n9875), .ZN(n16256) );
  NOR2_X1 U11895 ( .A1(n12795), .A2(n12666), .ZN(n21429) );
  AND2_X1 U11896 ( .A1(n13859), .A2(n14116), .ZN(n12665) );
  NAND2_X1 U11897 ( .A1(n10271), .A2(n10270), .ZN(n10633) );
  INV_X1 U11898 ( .A(n14282), .ZN(n16328) );
  NAND2_X1 U11899 ( .A1(n15194), .A2(n10142), .ZN(n10141) );
  INV_X1 U11900 ( .A(n17403), .ZN(n10142) );
  NOR2_X1 U11901 ( .A1(n16652), .A2(n16398), .ZN(n16397) );
  NOR2_X1 U11902 ( .A1(n9914), .A2(n10301), .ZN(n10300) );
  AND2_X1 U11903 ( .A1(n20437), .A2(n13777), .ZN(n20435) );
  OAI22_X1 U11904 ( .A1(n13213), .A2(n13212), .B1(n13211), .B2(n13210), .ZN(
        n13214) );
  INV_X1 U11905 ( .A(n17591), .ZN(n17577) );
  XNOR2_X1 U11906 ( .A(n12519), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12506) );
  INV_X1 U11907 ( .A(n12502), .ZN(n10189) );
  NAND2_X1 U11908 ( .A1(n10191), .A2(n12878), .ZN(n10190) );
  INV_X1 U11909 ( .A(n13218), .ZN(n10191) );
  NAND2_X1 U11910 ( .A1(n12503), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10188) );
  INV_X1 U11911 ( .A(n17681), .ZN(n17639) );
  INV_X1 U11912 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21212) );
  OR2_X1 U11913 ( .A1(n16932), .A2(n13774), .ZN(n21207) );
  XNOR2_X1 U11914 ( .A(n13901), .B(n13900), .ZN(n21197) );
  XNOR2_X1 U11915 ( .A(n13897), .B(n13898), .ZN(n21190) );
  NAND2_X1 U11916 ( .A1(n13903), .A2(n13906), .ZN(n20800) );
  OR2_X1 U11917 ( .A1(n13904), .A2(n13905), .ZN(n13906) );
  NOR2_X1 U11918 ( .A1(n18384), .A2(n18036), .ZN(n18396) );
  NOR2_X1 U11919 ( .A1(n18606), .A2(n18738), .ZN(n18601) );
  NOR2_X1 U11920 ( .A1(n18673), .A2(n18762), .ZN(n18664) );
  NAND2_X1 U11921 ( .A1(n18724), .A2(n9998), .ZN(n18694) );
  AND2_X1 U11922 ( .A1(n18670), .A2(n9937), .ZN(n9998) );
  NOR2_X1 U11923 ( .A1(n10211), .A2(n17951), .ZN(n10210) );
  INV_X1 U11924 ( .A(n18862), .ZN(n10211) );
  NAND2_X1 U11925 ( .A1(n9953), .A2(n18850), .ZN(n10212) );
  INV_X1 U11926 ( .A(n18849), .ZN(n10213) );
  INV_X1 U11927 ( .A(n19205), .ZN(n19216) );
  INV_X1 U11928 ( .A(n19061), .ZN(n19218) );
  OAI21_X1 U11929 ( .B1(n13907), .B2(n9883), .A(n11624), .ZN(n11625) );
  NOR2_X1 U11930 ( .A1(n11618), .A2(n11617), .ZN(n11623) );
  NOR2_X1 U11931 ( .A1(n11705), .A2(n11616), .ZN(n11617) );
  AND2_X1 U11932 ( .A1(n14107), .A2(n14106), .ZN(n17139) );
  OAI22_X1 U11933 ( .A1(n11576), .A2(n11716), .B1(n20842), .B2(n11575), .ZN(
        n11577) );
  CLKBUF_X1 U11934 ( .A(n10477), .Z(n11157) );
  NAND2_X1 U11935 ( .A1(n11270), .A2(n9876), .ZN(n10262) );
  OR2_X1 U11936 ( .A1(n10675), .A2(n10674), .ZN(n11232) );
  OR2_X1 U11937 ( .A1(n10614), .A2(n10613), .ZN(n11204) );
  INV_X1 U11938 ( .A(n11341), .ZN(n10492) );
  AND2_X1 U11939 ( .A1(n11878), .A2(n11876), .ZN(n10233) );
  NOR2_X1 U11940 ( .A1(n9991), .A2(n9990), .ZN(n9989) );
  NOR2_X1 U11941 ( .A1(n11962), .A2(n9992), .ZN(n9990) );
  NAND2_X1 U11942 ( .A1(n9989), .A2(n9992), .ZN(n9988) );
  AOI21_X1 U11943 ( .B1(n10310), .B2(n10312), .A(n16754), .ZN(n10309) );
  INV_X1 U11944 ( .A(n10316), .ZN(n10315) );
  OR2_X1 U11945 ( .A1(n11865), .A2(n11864), .ZN(n11868) );
  OR2_X1 U11946 ( .A1(n11670), .A2(n11669), .ZN(n12141) );
  AND2_X1 U11947 ( .A1(n13777), .A2(n11472), .ZN(n11512) );
  NAND2_X1 U11948 ( .A1(n11492), .A2(n13681), .ZN(n11514) );
  NAND2_X1 U11949 ( .A1(n11491), .A2(n11490), .ZN(n11492) );
  NAND2_X1 U11950 ( .A1(n12272), .A2(n12253), .ZN(n11490) );
  NAND2_X1 U11951 ( .A1(n12215), .A2(n13778), .ZN(n11445) );
  INV_X1 U11952 ( .A(n11558), .ZN(n11555) );
  AND2_X1 U11953 ( .A1(n16946), .A2(n20403), .ZN(n10291) );
  NAND2_X1 U11954 ( .A1(n11455), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11352) );
  AOI22_X1 U11955 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11364) );
  NAND2_X1 U11956 ( .A1(n9861), .A2(n16946), .ZN(n11718) );
  AND2_X1 U11957 ( .A1(n21212), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11809) );
  AND2_X1 U11958 ( .A1(n12210), .A2(n12215), .ZN(n11466) );
  NAND2_X1 U11959 ( .A1(n13493), .A2(n17087), .ZN(n10007) );
  NAND2_X1 U11960 ( .A1(n9976), .A2(n10488), .ZN(n9974) );
  INV_X1 U11961 ( .A(n11189), .ZN(n9976) );
  INV_X1 U11962 ( .A(n15590), .ZN(n10247) );
  NAND2_X1 U11963 ( .A1(n11019), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11058) );
  AND2_X1 U11964 ( .A1(n15545), .A2(n10284), .ZN(n10283) );
  NOR2_X1 U11965 ( .A1(n10799), .A2(n10782), .ZN(n10863) );
  NAND2_X1 U11966 ( .A1(n15510), .A2(n10250), .ZN(n10249) );
  NOR2_X1 U11967 ( .A1(n10251), .A2(n15536), .ZN(n10250) );
  INV_X1 U11968 ( .A(n15524), .ZN(n10251) );
  INV_X1 U11969 ( .A(n10262), .ZN(n10263) );
  INV_X1 U11970 ( .A(n12764), .ZN(n12738) );
  NAND2_X1 U11971 ( .A1(n12646), .A2(n14058), .ZN(n10050) );
  OR2_X1 U11972 ( .A1(n10545), .A2(n10544), .ZN(n11205) );
  NAND2_X1 U11973 ( .A1(n10265), .A2(n10267), .ZN(n10588) );
  AOI21_X1 U11974 ( .B1(n10272), .B2(n10632), .A(n10268), .ZN(n10267) );
  INV_X1 U11975 ( .A(n11180), .ZN(n10268) );
  OR2_X1 U11976 ( .A1(n10508), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10509) );
  AND2_X1 U11977 ( .A1(n17167), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10590) );
  OR2_X1 U11978 ( .A1(n10652), .A2(n10651), .ZN(n11224) );
  INV_X1 U11979 ( .A(n9973), .ZN(n10501) );
  XNOR2_X1 U11980 ( .A(n9956), .B(n14113), .ZN(n14085) );
  INV_X1 U11981 ( .A(n9830), .ZN(n14561) );
  AND2_X1 U11982 ( .A1(n10498), .A2(n10598), .ZN(n14796) );
  OAI21_X1 U11983 ( .B1(n10040), .B2(n10039), .A(n10038), .ZN(n10037) );
  AOI21_X1 U11984 ( .B1(n10040), .B2(n10039), .A(n10036), .ZN(n10035) );
  NAND2_X1 U11985 ( .A1(n11322), .A2(n11307), .ZN(n10039) );
  AND2_X1 U11986 ( .A1(n12648), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11311) );
  NOR2_X1 U11987 ( .A1(n11656), .A2(n11655), .ZN(n12275) );
  NOR2_X1 U11988 ( .A1(n12001), .A2(n12000), .ZN(n12005) );
  INV_X1 U11989 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10228) );
  NOR2_X1 U11990 ( .A1(n11970), .A2(n10230), .ZN(n10229) );
  NOR2_X1 U11991 ( .A1(n11911), .A2(n10236), .ZN(n10235) );
  INV_X1 U11992 ( .A(n11908), .ZN(n10236) );
  NAND2_X1 U11993 ( .A1(n11900), .A2(n20286), .ZN(n20276) );
  AND2_X1 U11994 ( .A1(n11875), .A2(n10231), .ZN(n11900) );
  AND2_X1 U11995 ( .A1(n9836), .A2(n20433), .ZN(n10231) );
  NAND2_X1 U11996 ( .A1(n11875), .A2(n10233), .ZN(n11889) );
  NAND2_X1 U11997 ( .A1(n10222), .A2(n10221), .ZN(n11806) );
  NAND2_X1 U11998 ( .A1(n20565), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10221) );
  NAND2_X1 U11999 ( .A1(n12025), .A2(n11790), .ZN(n10222) );
  NAND2_X1 U12000 ( .A1(n11815), .A2(n11816), .ZN(n11814) );
  INV_X1 U12001 ( .A(n12869), .ZN(n10199) );
  INV_X1 U12002 ( .A(n16493), .ZN(n10200) );
  AOI211_X1 U12003 ( .C1(n13164), .C2(n13161), .A(n13160), .B(n16413), .ZN(
        n13162) );
  AND2_X1 U12004 ( .A1(n13100), .A2(n13099), .ZN(n13101) );
  OR2_X1 U12005 ( .A1(n16443), .A2(n16521), .ZN(n10296) );
  INV_X1 U12006 ( .A(n13069), .ZN(n13029) );
  AND2_X1 U12007 ( .A1(n9903), .A2(n10307), .ZN(n10306) );
  INV_X1 U12008 ( .A(n16462), .ZN(n10307) );
  NOR2_X1 U12009 ( .A1(n11750), .A2(n11749), .ZN(n12311) );
  NAND2_X1 U12010 ( .A1(n11494), .A2(n11790), .ZN(n11467) );
  NAND2_X1 U12011 ( .A1(n10148), .A2(n12131), .ZN(n10147) );
  NOR2_X1 U12012 ( .A1(n20309), .A2(n10155), .ZN(n10154) );
  INV_X1 U12013 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10155) );
  NAND2_X1 U12014 ( .A1(n9945), .A2(n10057), .ZN(n11554) );
  NAND2_X1 U12015 ( .A1(n9946), .A2(n11511), .ZN(n9945) );
  NAND2_X1 U12016 ( .A1(n11550), .A2(n11551), .ZN(n9946) );
  AOI22_X1 U12017 ( .A1(n11535), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11537) );
  INV_X1 U12018 ( .A(n11793), .ZN(n12289) );
  NAND2_X1 U12019 ( .A1(n10175), .A2(n16428), .ZN(n10174) );
  INV_X1 U12020 ( .A(n16446), .ZN(n10175) );
  INV_X1 U12021 ( .A(n13671), .ZN(n10195) );
  NAND2_X1 U12022 ( .A1(n10289), .A2(n12497), .ZN(n10288) );
  NAND2_X1 U12023 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10091) );
  NOR2_X1 U12024 ( .A1(n14607), .A2(n14606), .ZN(n12085) );
  INV_X1 U12025 ( .A(n12074), .ZN(n12528) );
  NAND2_X1 U12026 ( .A1(n16694), .A2(n12172), .ZN(n9972) );
  XNOR2_X1 U12027 ( .A(n12175), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17551) );
  OR2_X1 U12028 ( .A1(n12176), .A2(n11892), .ZN(n12175) );
  NAND2_X1 U12029 ( .A1(n12171), .A2(n12170), .ZN(n12176) );
  INV_X1 U12030 ( .A(n12169), .ZN(n12171) );
  NAND2_X1 U12031 ( .A1(n17590), .A2(n12150), .ZN(n12156) );
  CLKBUF_X1 U12032 ( .A(n12235), .Z(n12236) );
  INV_X1 U12033 ( .A(n12240), .ZN(n12246) );
  NOR2_X1 U12034 ( .A1(n16946), .A2(n11562), .ZN(n9947) );
  NAND2_X1 U12035 ( .A1(n11455), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11432) );
  NAND2_X1 U12036 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11431) );
  INV_X1 U12037 ( .A(n11385), .ZN(n11389) );
  NAND2_X1 U12038 ( .A1(n11455), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11386) );
  NAND2_X1 U12039 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11387) );
  AOI22_X1 U12040 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11380) );
  NAND3_X1 U12041 ( .A1(n21177), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n21023), 
        .ZN(n14018) );
  NOR2_X1 U12042 ( .A1(n20006), .A2(n13223), .ZN(n13314) );
  NAND2_X1 U12043 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20160), .ZN(
        n13225) );
  NOR2_X1 U12044 ( .A1(n13226), .A2(n13223), .ZN(n13264) );
  INV_X1 U12045 ( .A(n13223), .ZN(n9996) );
  INV_X1 U12046 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9995) );
  NOR2_X1 U12047 ( .A1(n13225), .A2(n13226), .ZN(n13295) );
  AND2_X1 U12048 ( .A1(n10348), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10126) );
  NAND2_X1 U12049 ( .A1(n18957), .A2(n18947), .ZN(n18948) );
  NAND2_X1 U12050 ( .A1(n9843), .A2(n19449), .ZN(n10224) );
  NOR2_X1 U12051 ( .A1(n19131), .A2(n19132), .ZN(n13521) );
  NAND2_X1 U12052 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19081), .ZN(
        n17739) );
  NOR2_X1 U12053 ( .A1(n13410), .A2(n13409), .ZN(n13489) );
  OR2_X1 U12054 ( .A1(n15484), .A2(n15438), .ZN(n15439) );
  NOR2_X1 U12055 ( .A1(n15444), .A2(n21495), .ZN(n10024) );
  NAND2_X1 U12056 ( .A1(n15541), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15516) );
  NAND2_X1 U12057 ( .A1(n10029), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n10028) );
  INV_X1 U12058 ( .A(n17216), .ZN(n10029) );
  AND2_X1 U12059 ( .A1(n17352), .A2(n15098), .ZN(n15099) );
  AND2_X1 U12060 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n9939), .ZN(n10034) );
  NOR2_X1 U12061 ( .A1(n21461), .A2(n15155), .ZN(n15181) );
  OR2_X1 U12062 ( .A1(n21534), .A2(n15164), .ZN(n15155) );
  INV_X1 U12063 ( .A(n12770), .ZN(n10245) );
  AND2_X1 U12064 ( .A1(n12724), .A2(n12723), .ZN(n15574) );
  NAND2_X1 U12065 ( .A1(n15362), .A2(n9899), .ZN(n15587) );
  AOI21_X1 U12066 ( .B1(n14136), .B2(n10237), .A(n12674), .ZN(n13979) );
  AND2_X1 U12067 ( .A1(n15761), .A2(n11081), .ZN(n11126) );
  INV_X1 U12068 ( .A(n15336), .ZN(n10880) );
  AND2_X1 U12069 ( .A1(n10281), .A2(n9885), .ZN(n10280) );
  NAND2_X1 U12070 ( .A1(n15753), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15756) );
  NOR2_X1 U12071 ( .A1(n15753), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15752) );
  OR2_X1 U12072 ( .A1(n15768), .A2(n11174), .ZN(n11107) );
  NOR2_X1 U12073 ( .A1(n10955), .A2(n10954), .ZN(n10956) );
  NOR2_X1 U12074 ( .A1(n10920), .A2(n10900), .ZN(n10921) );
  INV_X1 U12075 ( .A(n10919), .ZN(n10920) );
  NOR2_X1 U12076 ( .A1(n17228), .A2(n10883), .ZN(n10919) );
  NAND2_X1 U12077 ( .A1(n10832), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10882) );
  AND2_X1 U12078 ( .A1(n10817), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10832) );
  INV_X1 U12079 ( .A(n10750), .ZN(n10751) );
  AND2_X1 U12080 ( .A1(n10766), .A2(n10765), .ZN(n14993) );
  AND3_X1 U12081 ( .A1(n10748), .A2(n10747), .A3(n10746), .ZN(n15091) );
  NAND2_X1 U12082 ( .A1(n11243), .A2(n10872), .ZN(n10726) );
  CLKBUF_X1 U12083 ( .A(n14514), .Z(n14515) );
  AND2_X1 U12084 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n10699), .ZN(
        n10722) );
  NOR2_X1 U12085 ( .A1(n10680), .A2(n14629), .ZN(n10699) );
  INV_X1 U12086 ( .A(n10657), .ZN(n10658) );
  NAND2_X1 U12087 ( .A1(n10658), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10680) );
  NAND2_X1 U12088 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10657) );
  INV_X1 U12089 ( .A(n13995), .ZN(n10637) );
  AND2_X1 U12090 ( .A1(n10256), .A2(n11285), .ZN(n15765) );
  NAND2_X1 U12091 ( .A1(n16112), .A2(n15751), .ZN(n16100) );
  INV_X1 U12092 ( .A(n16121), .ZN(n16112) );
  NOR2_X1 U12093 ( .A1(n15612), .A2(n15536), .ZN(n15537) );
  NOR2_X1 U12094 ( .A1(n15612), .A2(n10248), .ZN(n15522) );
  INV_X1 U12095 ( .A(n10250), .ZN(n10248) );
  OR2_X1 U12096 ( .A1(n15620), .A2(n15614), .ZN(n15612) );
  NAND2_X1 U12097 ( .A1(n9963), .A2(n10273), .ZN(n16214) );
  OR2_X1 U12098 ( .A1(n9891), .A2(n16288), .ZN(n10273) );
  AND2_X1 U12099 ( .A1(n15630), .A2(n15549), .ZN(n15618) );
  NAND2_X1 U12100 ( .A1(n15618), .A2(n15617), .ZN(n15620) );
  AND2_X1 U12101 ( .A1(n11281), .A2(n9839), .ZN(n16137) );
  AND2_X1 U12102 ( .A1(n12731), .A2(n12730), .ZN(n16279) );
  NAND2_X1 U12103 ( .A1(n15362), .A2(n15339), .ZN(n15589) );
  NAND2_X1 U12104 ( .A1(n15124), .A2(n15123), .ZN(n10264) );
  NOR2_X1 U12105 ( .A1(n14615), .A2(n14964), .ZN(n14148) );
  NAND2_X1 U12106 ( .A1(n14127), .A2(n14126), .ZN(n9978) );
  NOR2_X1 U12107 ( .A1(n14617), .A2(n14137), .ZN(n17343) );
  NOR2_X1 U12108 ( .A1(n12795), .A2(n12791), .ZN(n16216) );
  NAND2_X1 U12109 ( .A1(n9806), .A2(n17165), .ZN(n13859) );
  NAND2_X1 U12110 ( .A1(n11196), .A2(n11195), .ZN(n14155) );
  NAND2_X1 U12111 ( .A1(n9977), .A2(n10486), .ZN(n13910) );
  INV_X1 U12112 ( .A(n10484), .ZN(n9977) );
  AND2_X2 U12113 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13885) );
  CLKBUF_X1 U12114 ( .A(n13868), .Z(n14112) );
  OR2_X1 U12115 ( .A1(n9956), .A2(n14177), .ZN(n14115) );
  NOR2_X1 U12116 ( .A1(n14703), .A2(n14561), .ZN(n14708) );
  INV_X1 U12117 ( .A(n11193), .ZN(n14562) );
  NOR2_X1 U12118 ( .A1(n14564), .A2(n14833), .ZN(n15008) );
  INV_X1 U12119 ( .A(n14637), .ZN(n14564) );
  OR2_X1 U12120 ( .A1(n9830), .A2(n14562), .ZN(n14323) );
  OAI22_X1 U12121 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14033), .B1(n14032), 
        .B2(n21545), .ZN(n14637) );
  AND2_X1 U12122 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n14637), .ZN(n14079) );
  OR2_X1 U12123 ( .A1(n16322), .A2(n14174), .ZN(n14325) );
  AOI21_X1 U12124 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n14318), .A(n14564), 
        .ZN(n14702) );
  NAND2_X1 U12125 ( .A1(n11310), .A2(n11311), .ZN(n11334) );
  NAND2_X1 U12126 ( .A1(n11333), .A2(n11332), .ZN(n12642) );
  NAND2_X1 U12127 ( .A1(n11463), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n21228) );
  AOI221_X1 U12128 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12013), 
        .C1(n17083), .C2(n12013), .A(n12012), .ZN(n12203) );
  NOR2_X1 U12129 ( .A1(n17421), .A2(n17403), .ZN(n10144) );
  NAND2_X1 U12130 ( .A1(n11989), .A2(n11990), .ZN(n12001) );
  NAND2_X1 U12131 ( .A1(n15194), .A2(n16572), .ZN(n10156) );
  NOR2_X1 U12132 ( .A1(n17447), .A2(n17434), .ZN(n10158) );
  OR2_X1 U12133 ( .A1(n17456), .A2(n15194), .ZN(n10160) );
  NOR2_X1 U12134 ( .A1(n15194), .A2(n13650), .ZN(n17118) );
  AND2_X1 U12135 ( .A1(n11926), .A2(n11924), .ZN(n20256) );
  NAND2_X1 U12136 ( .A1(n11909), .A2(n10235), .ZN(n11931) );
  NAND2_X1 U12137 ( .A1(n11909), .A2(n11908), .ZN(n20277) );
  NOR2_X1 U12138 ( .A1(n16447), .A2(n10173), .ZN(n12561) );
  OR3_X1 U12139 ( .A1(n10174), .A2(n10176), .A3(n12877), .ZN(n10173) );
  AND2_X1 U12140 ( .A1(n14351), .A2(n9932), .ZN(n10302) );
  INV_X1 U12141 ( .A(n11455), .ZN(n13041) );
  CLKBUF_X1 U12142 ( .A(n16452), .Z(n16453) );
  CLKBUF_X1 U12143 ( .A(n16454), .Z(n16455) );
  NAND2_X1 U12144 ( .A1(n9840), .A2(n13743), .ZN(n15229) );
  NAND2_X1 U12145 ( .A1(n10193), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12282) );
  AND2_X1 U12146 ( .A1(n20475), .A2(n13779), .ZN(n15216) );
  NAND2_X1 U12147 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10136) );
  NAND2_X1 U12148 ( .A1(n13643), .A2(n16391), .ZN(n16393) );
  NAND2_X1 U12149 ( .A1(n10090), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10089) );
  INV_X1 U12150 ( .A(n10091), .ZN(n10090) );
  INV_X1 U12151 ( .A(n10148), .ZN(n10146) );
  AOI21_X1 U12152 ( .B1(n16868), .B2(n16867), .A(n12602), .ZN(n17517) );
  INV_X1 U12153 ( .A(n12085), .ZN(n14609) );
  NOR2_X1 U12154 ( .A1(n9900), .A2(n10152), .ZN(n10151) );
  INV_X1 U12155 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10152) );
  AND2_X1 U12156 ( .A1(n12061), .A2(n12060), .ZN(n13964) );
  NOR2_X1 U12157 ( .A1(n16697), .A2(n10162), .ZN(n10161) );
  INV_X1 U12158 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10162) );
  AND2_X1 U12159 ( .A1(n9892), .A2(n9967), .ZN(n12164) );
  NAND2_X1 U12160 ( .A1(n10169), .A2(n12039), .ZN(n14937) );
  NOR2_X1 U12161 ( .A1(n12509), .A2(n12508), .ZN(n12510) );
  INV_X1 U12162 ( .A(n12507), .ZN(n12509) );
  NOR2_X1 U12163 ( .A1(n10352), .A2(n12543), .ZN(n12544) );
  OR3_X1 U12164 ( .A1(n12861), .A2(n11892), .A3(n12499), .ZN(n12507) );
  OR2_X1 U12165 ( .A1(n13613), .A2(n11892), .ZN(n12553) );
  INV_X1 U12166 ( .A(n12552), .ZN(n9993) );
  NOR2_X1 U12167 ( .A1(n16742), .A2(n16730), .ZN(n16718) );
  NOR3_X1 U12168 ( .A1(n16447), .A2(n10176), .A3(n16446), .ZN(n16437) );
  OR2_X1 U12169 ( .A1(n16753), .A2(n16754), .ZN(n16742) );
  OR3_X1 U12170 ( .A1(n17445), .A2(n11892), .A3(n16747), .ZN(n16576) );
  NOR2_X1 U12171 ( .A1(n16447), .A2(n16446), .ZN(n16448) );
  AND2_X1 U12172 ( .A1(n12622), .A2(n9926), .ZN(n16511) );
  AOI21_X1 U12173 ( .B1(n10065), .B2(n10063), .A(n9991), .ZN(n10062) );
  INV_X1 U12174 ( .A(n10065), .ZN(n10064) );
  INV_X1 U12175 ( .A(n11962), .ZN(n10063) );
  NOR2_X1 U12176 ( .A1(n10288), .A2(n16754), .ZN(n10286) );
  OR2_X2 U12177 ( .A1(n13667), .A2(n13668), .ZN(n16447) );
  INV_X1 U12178 ( .A(n10288), .ZN(n10285) );
  INV_X1 U12179 ( .A(n12613), .ZN(n10287) );
  NOR2_X1 U12180 ( .A1(n16644), .A2(n16799), .ZN(n16637) );
  AND2_X1 U12181 ( .A1(n12463), .A2(n12462), .ZN(n16376) );
  OR2_X1 U12182 ( .A1(n11959), .A2(n16799), .ZN(n16632) );
  INV_X1 U12183 ( .A(n10109), .ZN(n10108) );
  OAI21_X1 U12184 ( .B1(n10114), .B2(n12604), .A(n10113), .ZN(n10109) );
  OR2_X1 U12185 ( .A1(n12613), .A2(n10087), .ZN(n16644) );
  NAND2_X1 U12186 ( .A1(n10088), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10087) );
  INV_X1 U12187 ( .A(n10089), .ZN(n10088) );
  AND2_X1 U12188 ( .A1(n9904), .A2(n10183), .ZN(n10182) );
  INV_X1 U12189 ( .A(n16840), .ZN(n10183) );
  NAND2_X1 U12190 ( .A1(n12085), .A2(n10168), .ZN(n16667) );
  INV_X1 U12191 ( .A(n13626), .ZN(n10168) );
  OR2_X1 U12192 ( .A1(n12496), .A2(n12495), .ZN(n16839) );
  INV_X1 U12193 ( .A(n16839), .ZN(n16857) );
  NAND2_X1 U12194 ( .A1(n10319), .A2(n10318), .ZN(n16868) );
  NOR2_X1 U12195 ( .A1(n16899), .A2(n16684), .ZN(n10316) );
  AND2_X1 U12196 ( .A1(n12069), .A2(n12068), .ZN(n16688) );
  NAND2_X1 U12197 ( .A1(n10083), .A2(n12177), .ZN(n16893) );
  NAND2_X1 U12198 ( .A1(n17550), .A2(n17551), .ZN(n10083) );
  AND2_X2 U12199 ( .A1(n9986), .A2(n11888), .ZN(n11895) );
  OAI211_X1 U12200 ( .C1(n11884), .C2(n13569), .A(n11882), .B(n11883), .ZN(
        n9986) );
  AND2_X1 U12201 ( .A1(n12340), .A2(n12339), .ZN(n17636) );
  XNOR2_X1 U12202 ( .A(n12176), .B(n11892), .ZN(n16695) );
  NAND2_X1 U12203 ( .A1(n15234), .A2(n10172), .ZN(n13963) );
  XNOR2_X1 U12204 ( .A(n12156), .B(n12154), .ZN(n14934) );
  AOI21_X1 U12205 ( .B1(n10099), .B2(n10103), .A(n9907), .ZN(n10096) );
  NAND2_X1 U12206 ( .A1(n10079), .A2(n10097), .ZN(n10095) );
  INV_X1 U12207 ( .A(n10106), .ZN(n10103) );
  OR2_X1 U12208 ( .A1(n21190), .A2(n16968), .ZN(n20970) );
  NOR2_X1 U12209 ( .A1(n15215), .A2(n14018), .ZN(n20572) );
  NOR2_X1 U12210 ( .A1(n15214), .A2(n14018), .ZN(n20571) );
  INV_X1 U12211 ( .A(n20572), .ZN(n20579) );
  INV_X1 U12212 ( .A(n20571), .ZN(n20577) );
  INV_X1 U12213 ( .A(n20970), .ZN(n21028) );
  NAND2_X1 U12214 ( .A1(n17735), .A2(n14024), .ZN(n20574) );
  INV_X1 U12215 ( .A(n20215), .ZN(n20208) );
  NOR3_X1 U12216 ( .A1(n13587), .A2(n15394), .A3(n15393), .ZN(n19980) );
  INV_X1 U12217 ( .A(n18954), .ZN(n10119) );
  NOR2_X1 U12218 ( .A1(n18263), .A2(n18003), .ZN(n18061) );
  INV_X1 U12219 ( .A(n18061), .ZN(n18076) );
  AND2_X1 U12220 ( .A1(n9833), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10127) );
  NAND2_X1 U12221 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .ZN(n10074) );
  NOR2_X1 U12222 ( .A1(n18108), .A2(n10072), .ZN(n10071) );
  INV_X1 U12223 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n10072) );
  NOR2_X1 U12224 ( .A1(n18742), .A2(n10019), .ZN(n10018) );
  NAND2_X1 U12225 ( .A1(n18863), .A2(n19008), .ZN(n10215) );
  INV_X1 U12226 ( .A(n17910), .ZN(n17912) );
  AND2_X1 U12227 ( .A1(n18846), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17910) );
  NOR2_X1 U12228 ( .A1(n10125), .A2(n19034), .ZN(n19014) );
  NAND2_X1 U12229 ( .A1(n10126), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10125) );
  INV_X1 U12230 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19054) );
  INV_X1 U12231 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n19055) );
  NAND2_X1 U12232 ( .A1(n10117), .A2(n9838), .ZN(n18121) );
  OR2_X1 U12233 ( .A1(n19008), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13358) );
  AND2_X1 U12234 ( .A1(n15396), .A2(n10005), .ZN(n19994) );
  NAND2_X1 U12235 ( .A1(n13474), .A2(n13475), .ZN(n10005) );
  AND2_X1 U12236 ( .A1(n13461), .A2(n16986), .ZN(n10009) );
  INV_X1 U12237 ( .A(n19996), .ZN(n17781) );
  NOR2_X1 U12238 ( .A1(n19992), .A2(n19991), .ZN(n17780) );
  NAND2_X1 U12239 ( .A1(n19008), .A2(n19341), .ZN(n13346) );
  NAND2_X1 U12240 ( .A1(n13347), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9955) );
  INV_X1 U12241 ( .A(n19037), .ZN(n19028) );
  INV_X1 U12242 ( .A(n17739), .ZN(n19407) );
  NOR2_X1 U12243 ( .A1(n13463), .A2(n19559), .ZN(n17094) );
  XNOR2_X1 U12244 ( .A(n13339), .B(n13340), .ZN(n19139) );
  NOR2_X1 U12245 ( .A1(n19173), .A2(n19172), .ZN(n19171) );
  NOR2_X1 U12246 ( .A1(n19183), .A2(n19496), .ZN(n19182) );
  NAND2_X1 U12247 ( .A1(n20205), .A2(n19364), .ZN(n19511) );
  INV_X1 U12248 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20021) );
  NAND2_X1 U12249 ( .A1(n20208), .A2(n16987), .ZN(n20009) );
  INV_X1 U12250 ( .A(n13489), .ZN(n19559) );
  INV_X1 U12251 ( .A(n13462), .ZN(n19579) );
  NOR2_X1 U12252 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19550), .ZN(n19886) );
  INV_X1 U12253 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20164) );
  NAND2_X1 U12254 ( .A1(n15541), .A2(n10024), .ZN(n15506) );
  NAND2_X1 U12255 ( .A1(n10027), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n10026) );
  INV_X1 U12256 ( .A(n15443), .ZN(n10027) );
  NOR3_X1 U12257 ( .A1(n15566), .A2(n10028), .A3(n15443), .ZN(n15555) );
  NOR2_X1 U12258 ( .A1(n15566), .A2(n15443), .ZN(n17232) );
  NOR2_X1 U12259 ( .A1(n21481), .A2(n17243), .ZN(n15586) );
  NOR2_X1 U12260 ( .A1(n10032), .A2(n15442), .ZN(n10031) );
  INV_X1 U12261 ( .A(n10034), .ZN(n10032) );
  NAND2_X1 U12262 ( .A1(n10033), .A2(n10034), .ZN(n21276) );
  NOR2_X1 U12263 ( .A1(n21315), .A2(n21468), .ZN(n21298) );
  NOR2_X1 U12264 ( .A1(n21326), .A2(n15154), .ZN(n21321) );
  NAND2_X1 U12265 ( .A1(n10043), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n21326) );
  INV_X1 U12266 ( .A(n21296), .ZN(n21345) );
  INV_X1 U12267 ( .A(n21317), .ZN(n21292) );
  OR3_X1 U12268 ( .A1(n15153), .A2(n10045), .A3(n15103), .ZN(n21308) );
  AND2_X2 U12269 ( .A1(n13959), .A2(n13958), .ZN(n21381) );
  NAND2_X1 U12270 ( .A1(n21381), .A2(n15425), .ZN(n15641) );
  NAND2_X1 U12271 ( .A1(n10918), .A2(n10917), .ZN(n15627) );
  NAND2_X1 U12272 ( .A1(n15372), .A2(n15371), .ZN(n15721) );
  AND2_X1 U12273 ( .A1(n13994), .A2(n13993), .ZN(n15733) );
  OR2_X1 U12274 ( .A1(n15736), .A2(n13998), .ZN(n15732) );
  AND2_X1 U12275 ( .A1(n13925), .A2(n13924), .ZN(n21392) );
  OR2_X1 U12276 ( .A1(n15106), .A2(n15105), .ZN(n15108) );
  AND2_X1 U12277 ( .A1(n10991), .A2(n10275), .ZN(n15509) );
  NAND2_X1 U12278 ( .A1(n10991), .A2(n10990), .ZN(n15532) );
  INV_X1 U12279 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14629) );
  OR2_X1 U12280 ( .A1(n12629), .A2(n15741), .ZN(n11291) );
  NOR2_X1 U12281 ( .A1(n12807), .A2(n10054), .ZN(n17321) );
  NOR2_X1 U12282 ( .A1(n17336), .A2(n16197), .ZN(n10054) );
  NAND2_X1 U12283 ( .A1(n12800), .A2(n10046), .ZN(n17368) );
  INV_X1 U12284 ( .A(n10047), .ZN(n10046) );
  OAI21_X1 U12285 ( .B1(n16220), .B2(n17355), .A(n15351), .ZN(n10047) );
  NOR2_X1 U12286 ( .A1(n21432), .A2(n16216), .ZN(n14617) );
  AND2_X1 U12287 ( .A1(n10049), .A2(n10048), .ZN(n15351) );
  NAND2_X1 U12288 ( .A1(n16216), .A2(n14158), .ZN(n10049) );
  NAND2_X1 U12289 ( .A1(n12795), .A2(n17352), .ZN(n10048) );
  INV_X1 U12290 ( .A(n21427), .ZN(n17364) );
  INV_X1 U12291 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n14318) );
  NAND2_X1 U12292 ( .A1(n17170), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14033) );
  AOI22_X1 U12293 ( .A1(n15005), .A2(n15003), .B1(n15000), .B2(n15009), .ZN(
        n15081) );
  OR2_X1 U12294 ( .A1(n14499), .A2(n14324), .ZN(n14772) );
  OR2_X1 U12295 ( .A1(n14499), .A2(n14498), .ZN(n14748) );
  INV_X1 U12296 ( .A(n14789), .ZN(n14826) );
  OR2_X1 U12297 ( .A1(n14038), .A2(n9807), .ZN(n14865) );
  NOR2_X1 U12298 ( .A1(n14457), .A2(n14564), .ZN(n14818) );
  NOR2_X1 U12299 ( .A1(n15706), .A2(n14564), .ZN(n14810) );
  AND2_X1 U12300 ( .A1(n14708), .A2(n14562), .ZN(n14735) );
  NOR2_X1 U12301 ( .A1(n15681), .A2(n14564), .ZN(n14823) );
  NAND2_X1 U12302 ( .A1(n16328), .A2(n14283), .ZN(n14926) );
  NOR2_X1 U12303 ( .A1(n14282), .A2(n14487), .ZN(n15318) );
  INV_X1 U12304 ( .A(n15273), .ZN(n15321) );
  INV_X1 U12305 ( .A(n15315), .ZN(n15021) );
  INV_X1 U12306 ( .A(n15305), .ZN(n15078) );
  NOR2_X1 U12307 ( .A1(n15694), .A2(n14564), .ZN(n14814) );
  INV_X1 U12308 ( .A(n15298), .ZN(n15070) );
  INV_X1 U12309 ( .A(n15291), .ZN(n15063) );
  INV_X1 U12310 ( .A(n15285), .ZN(n16340) );
  INV_X1 U12311 ( .A(n14818), .ZN(n15320) );
  INV_X1 U12312 ( .A(n15280), .ZN(n16348) );
  INV_X1 U12313 ( .A(n14814), .ZN(n15302) );
  INV_X1 U12314 ( .A(n14823), .ZN(n15295) );
  INV_X2 U12315 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21441) );
  INV_X1 U12316 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n17400) );
  INV_X1 U12317 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21099) );
  AND2_X1 U12318 ( .A1(n13784), .A2(n20384), .ZN(n21239) );
  AND2_X1 U12319 ( .A1(n10145), .A2(n12816), .ZN(n17419) );
  AND3_X1 U12320 ( .A1(n10138), .A2(n15196), .A3(n10139), .ZN(n13651) );
  NAND2_X1 U12321 ( .A1(n10138), .A2(n10139), .ZN(n20246) );
  NOR2_X1 U12322 ( .A1(n12815), .A2(n16397), .ZN(n16385) );
  AND2_X1 U12323 ( .A1(n15196), .A2(n12845), .ZN(n16398) );
  INV_X1 U12324 ( .A(n20412), .ZN(n20380) );
  INV_X1 U12325 ( .A(n21086), .ZN(n20370) );
  OR2_X1 U12326 ( .A1(n12433), .A2(n12432), .ZN(n14604) );
  OR2_X1 U12327 ( .A1(n12418), .A2(n12417), .ZN(n14602) );
  OR2_X1 U12328 ( .A1(n12401), .A2(n12400), .ZN(n20420) );
  OR2_X1 U12329 ( .A1(n12385), .A2(n12384), .ZN(n20421) );
  OR2_X1 U12330 ( .A1(n12368), .A2(n12367), .ZN(n20426) );
  CLKBUF_X1 U12331 ( .A(n13969), .Z(n13970) );
  CLKBUF_X1 U12332 ( .A(n13966), .Z(n13967) );
  INV_X1 U12333 ( .A(n21197), .ZN(n16968) );
  INV_X1 U12334 ( .A(n20435), .ZN(n20428) );
  NAND2_X1 U12335 ( .A1(n12540), .A2(n12486), .ZN(n15415) );
  NOR2_X1 U12336 ( .A1(n16414), .A2(n16413), .ZN(n16416) );
  INV_X1 U12337 ( .A(n20442), .ZN(n16523) );
  CLKBUF_X1 U12338 ( .A(n16441), .Z(n16442) );
  INV_X1 U12339 ( .A(n10298), .ZN(n16520) );
  AND2_X1 U12340 ( .A1(n15216), .A2(n15214), .ZN(n20443) );
  AND2_X1 U12341 ( .A1(n15216), .A2(n15215), .ZN(n20444) );
  AND2_X1 U12342 ( .A1(n20475), .A2(n12272), .ZN(n20477) );
  NOR2_X1 U12343 ( .A1(n20492), .A2(n20477), .ZN(n20483) );
  NAND2_X1 U12344 ( .A1(n13903), .A2(n12929), .ZN(n14355) );
  INV_X1 U12345 ( .A(n20475), .ZN(n20491) );
  AND2_X1 U12346 ( .A1(n13696), .A2(n21101), .ZN(n20532) );
  INV_X1 U12347 ( .A(n20534), .ZN(n20540) );
  INV_X1 U12348 ( .A(n13920), .ZN(n13830) );
  NOR2_X1 U12349 ( .A1(n12613), .A2(n10089), .ZN(n16662) );
  INV_X1 U12350 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20287) );
  INV_X1 U12351 ( .A(n17582), .ZN(n17571) );
  INV_X1 U12352 ( .A(n17592), .ZN(n17572) );
  INV_X1 U12353 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17597) );
  NAND2_X1 U12354 ( .A1(n13682), .A2(n12130), .ZN(n17596) );
  AND2_X1 U12355 ( .A1(n17596), .A2(n13691), .ZN(n17582) );
  AND2_X1 U12356 ( .A1(n17596), .A2(n21196), .ZN(n17591) );
  INV_X1 U12357 ( .A(n17596), .ZN(n17564) );
  NOR2_X1 U12358 ( .A1(n9865), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16559) );
  NAND2_X1 U12359 ( .A1(n16607), .A2(n16606), .ZN(n11969) );
  INV_X1 U12360 ( .A(n10111), .ZN(n16648) );
  OAI21_X1 U12361 ( .B1(n16672), .B2(n10112), .A(n16656), .ZN(n10111) );
  NAND2_X1 U12362 ( .A1(n15031), .A2(n15032), .ZN(n17600) );
  NAND2_X1 U12363 ( .A1(n10098), .A2(n10106), .ZN(n17583) );
  NAND2_X1 U12364 ( .A1(n10080), .A2(n10104), .ZN(n17584) );
  NAND2_X1 U12365 ( .A1(n10079), .A2(n17588), .ZN(n17589) );
  INV_X1 U12366 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21203) );
  INV_X1 U12367 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21194) );
  NOR2_X1 U12368 ( .A1(n13742), .A2(n12295), .ZN(n14358) );
  INV_X1 U12369 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17701) );
  NAND2_X1 U12370 ( .A1(n12916), .A2(n14011), .ZN(n12918) );
  INV_X1 U12371 ( .A(n16965), .ZN(n17730) );
  INV_X1 U12372 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17083) );
  INV_X1 U12373 ( .A(n10060), .ZN(n20703) );
  OAI21_X1 U12374 ( .B1(n10060), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n10061), 
        .ZN(n20701) );
  NOR2_X1 U12375 ( .A1(n20723), .A2(n21177), .ZN(n10061) );
  NOR2_X1 U12376 ( .A1(n14378), .A2(n20931), .ZN(n20715) );
  INV_X1 U12377 ( .A(n20825), .ZN(n20828) );
  OAI21_X1 U12378 ( .B1(n20843), .B2(n20858), .A(n21023), .ZN(n20860) );
  INV_X1 U12379 ( .A(n21079), .ZN(n20999) );
  INV_X1 U12380 ( .A(n21069), .ZN(n21003) );
  OR3_X1 U12381 ( .A1(n20978), .A2(n20977), .A3(n20976), .ZN(n21011) );
  OAI21_X1 U12382 ( .B1(n20982), .B2(n20981), .A(n20980), .ZN(n21010) );
  AND2_X1 U12383 ( .A1(n20943), .A2(n20942), .ZN(n21008) );
  OAI22_X1 U12384 ( .A1(n15714), .A2(n20579), .B1(n20555), .B2(n20577), .ZN(
        n21042) );
  INV_X1 U12385 ( .A(n20996), .ZN(n21048) );
  INV_X1 U12386 ( .A(n21006), .ZN(n21066) );
  AND2_X1 U12387 ( .A1(n20943), .A2(n21028), .ZN(n21075) );
  NOR2_X1 U12388 ( .A1(n19980), .A2(n18796), .ZN(n20220) );
  INV_X1 U12389 ( .A(n20220), .ZN(n20216) );
  INV_X1 U12390 ( .A(n10011), .ZN(n17893) );
  NAND2_X2 U12391 ( .A1(n20038), .A2(n20036), .ZN(n17894) );
  AOI21_X1 U12392 ( .B1(n17934), .B2(n17935), .A(n20053), .ZN(n10135) );
  NOR2_X1 U12393 ( .A1(n17938), .A2(n10131), .ZN(n10130) );
  NAND2_X1 U12394 ( .A1(n17939), .A2(n10132), .ZN(n10131) );
  NAND2_X1 U12395 ( .A1(n18248), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n10132) );
  NOR2_X1 U12396 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18056), .ZN(n18042) );
  NOR2_X1 U12397 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18144), .ZN(n18132) );
  NOR2_X1 U12398 ( .A1(n20218), .A2(n20040), .ZN(n18243) );
  NAND4_X1 U12399 ( .A1(n19529), .A2(n20216), .A3(n20053), .A4(n20044), .ZN(
        n18273) );
  AND3_X1 U12400 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n18331), .ZN(n18319) );
  NOR2_X1 U12401 ( .A1(n18335), .A2(n10074), .ZN(n18334) );
  NOR2_X1 U12402 ( .A1(n18335), .A2(n18279), .ZN(n18340) );
  NOR2_X1 U12403 ( .A1(n18277), .A2(n18357), .ZN(n18341) );
  NOR2_X1 U12404 ( .A1(n18384), .A2(n10066), .ZN(n18369) );
  NAND2_X1 U12405 ( .A1(n19584), .A2(n10067), .ZN(n10066) );
  NOR2_X1 U12406 ( .A1(n10068), .A2(n18036), .ZN(n10067) );
  INV_X1 U12407 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U12408 ( .A1(n18482), .A2(n10069), .ZN(n18448) );
  NOR2_X1 U12409 ( .A1(n10070), .A2(n10073), .ZN(n10069) );
  INV_X1 U12410 ( .A(n10071), .ZN(n10070) );
  NAND2_X1 U12411 ( .A1(n18482), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n17074) );
  NAND2_X1 U12412 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18511), .ZN(n18483) );
  NOR2_X1 U12413 ( .A1(n18148), .A2(n18528), .ZN(n18511) );
  NAND2_X1 U12414 ( .A1(n18547), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n18528) );
  NOR2_X1 U12415 ( .A1(n18554), .A2(n10075), .ZN(n18547) );
  NAND2_X1 U12416 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .ZN(n10075) );
  NAND2_X1 U12417 ( .A1(n18565), .A2(P3_EBX_REG_5__SCAN_IN), .ZN(n18554) );
  NOR2_X1 U12418 ( .A1(n18566), .A2(n18561), .ZN(n18565) );
  NAND2_X1 U12419 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n18573), .ZN(n18566) );
  AND3_X1 U12420 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(n18577), .ZN(n18569) );
  AND2_X1 U12421 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n18569), .ZN(n18573) );
  OR3_X1 U12422 ( .A1(n19552), .A2(n20205), .A3(n20202), .ZN(n10076) );
  OAI21_X1 U12423 ( .B1(n18597), .B2(n9915), .A(n10012), .ZN(n10014) );
  NAND2_X1 U12424 ( .A1(n18646), .A2(n10013), .ZN(n10012) );
  INV_X1 U12425 ( .A(n10015), .ZN(n10013) );
  NOR2_X1 U12426 ( .A1(n18597), .A2(n10017), .ZN(n10016) );
  NAND2_X1 U12427 ( .A1(n18615), .A2(n9847), .ZN(n18606) );
  NOR2_X1 U12428 ( .A1(n18624), .A2(n18619), .ZN(n18615) );
  NAND2_X1 U12429 ( .A1(n18615), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n18614) );
  NOR2_X1 U12430 ( .A1(n18660), .A2(n10021), .ZN(n18620) );
  INV_X1 U12431 ( .A(n18625), .ZN(n10022) );
  NAND2_X1 U12432 ( .A1(n18620), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n18619) );
  NOR2_X1 U12433 ( .A1(n18624), .A2(n18660), .ZN(n18654) );
  NAND2_X1 U12434 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n18654), .ZN(n18653) );
  NAND2_X1 U12435 ( .A1(n18664), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18660) );
  OR4_X1 U12436 ( .A1(n18694), .A2(n18775), .A3(n18671), .A4(n18583), .ZN(
        n18673) );
  INV_X1 U12437 ( .A(n13499), .ZN(n18703) );
  NOR2_X1 U12438 ( .A1(n13247), .A2(n13246), .ZN(n18706) );
  NOR2_X1 U12439 ( .A1(n13257), .A2(n13256), .ZN(n18712) );
  NOR2_X1 U12440 ( .A1(n10208), .A2(n10205), .ZN(n10204) );
  NOR2_X1 U12441 ( .A1(n18669), .A2(n18668), .ZN(n18715) );
  INV_X1 U12442 ( .A(n18722), .ZN(n18717) );
  INV_X1 U12443 ( .A(n18723), .ZN(n18720) );
  NOR2_X1 U12444 ( .A1(n13267), .A2(n13266), .ZN(n13271) );
  AND2_X1 U12445 ( .A1(n9999), .A2(n20038), .ZN(n18724) );
  NAND2_X1 U12446 ( .A1(n17191), .A2(n17190), .ZN(n9999) );
  AND2_X1 U12447 ( .A1(n20015), .A2(n18724), .ZN(n18722) );
  NOR2_X1 U12448 ( .A1(n20015), .A2(n18726), .ZN(n18723) );
  NOR2_X1 U12449 ( .A1(n18796), .A2(n18730), .ZN(n18772) );
  INV_X1 U12450 ( .A(n18759), .ZN(n18789) );
  INV_X1 U12451 ( .A(n18844), .ZN(n18842) );
  NOR2_X1 U12452 ( .A1(n18973), .A2(n18972), .ZN(n13529) );
  AND2_X1 U12453 ( .A1(n19886), .A2(n19608), .ZN(n19922) );
  NOR2_X1 U12454 ( .A1(n19352), .A2(n19351), .ZN(n19350) );
  NOR2_X1 U12455 ( .A1(n19055), .A2(n19054), .ZN(n19053) );
  NAND2_X1 U12456 ( .A1(n10225), .A2(n10226), .ZN(n19118) );
  NOR2_X1 U12457 ( .A1(n13341), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10226) );
  INV_X1 U12458 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19148) );
  INV_X1 U12459 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19178) );
  INV_X1 U12460 ( .A(n10203), .ZN(n18877) );
  NAND2_X1 U12461 ( .A1(n18957), .A2(n13352), .ZN(n18907) );
  INV_X1 U12462 ( .A(n18896), .ZN(n18906) );
  OAI21_X2 U12463 ( .B1(n17780), .B2(n10008), .A(n19994), .ZN(n20014) );
  INV_X1 U12464 ( .A(n20009), .ZN(n19977) );
  NOR2_X1 U12465 ( .A1(n19533), .A2(n19291), .ZN(n19340) );
  INV_X1 U12466 ( .A(n13335), .ZN(n10218) );
  INV_X1 U12467 ( .A(n10219), .ZN(n19153) );
  NAND2_X1 U12468 ( .A1(n17090), .A2(n15397), .ZN(n19983) );
  INV_X1 U12469 ( .A(n19497), .ZN(n19525) );
  INV_X1 U12470 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20019) );
  INV_X1 U12471 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20026) );
  INV_X1 U12472 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20030) );
  INV_X1 U12473 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n20153) );
  NOR2_X1 U12475 ( .A1(n17844), .A2(n17801), .ZN(n17845) );
  OAI21_X1 U12476 ( .B1(n15598), .B2(n21296), .A(n10239), .ZN(n10238) );
  INV_X1 U12477 ( .A(n17316), .ZN(n15750) );
  NAND2_X1 U12478 ( .A1(n9980), .A2(n9872), .ZN(P1_U2971) );
  NAND2_X1 U12479 ( .A1(n17322), .A2(n17267), .ZN(n9980) );
  AND2_X1 U12480 ( .A1(n12809), .A2(n12808), .ZN(n12810) );
  AOI21_X1 U12481 ( .B1(n17412), .B2(n17411), .A(n17410), .ZN(n17413) );
  OAI21_X1 U12482 ( .B1(n13218), .B2(n17479), .A(n13217), .ZN(n13219) );
  NAND2_X1 U12483 ( .A1(n10349), .A2(n12599), .ZN(n12600) );
  INV_X1 U12484 ( .A(n12570), .ZN(n12571) );
  INV_X1 U12485 ( .A(n12548), .ZN(n12549) );
  NAND2_X1 U12486 ( .A1(n12504), .A2(n17639), .ZN(n10192) );
  INV_X1 U12487 ( .A(n12587), .ZN(n12588) );
  OAI21_X1 U12488 ( .B1(n12586), .B2(n17669), .A(n12585), .ZN(n12587) );
  OAI21_X1 U12489 ( .B1(n10134), .B2(n17933), .A(n10129), .ZN(P3_U2642) );
  AND2_X1 U12490 ( .A1(n10133), .A2(n10130), .ZN(n10129) );
  INV_X1 U12491 ( .A(n10135), .ZN(n10134) );
  OR2_X1 U12492 ( .A1(n17941), .A2(n17940), .ZN(n10133) );
  NOR3_X1 U12493 ( .A1(n18384), .A2(n18624), .A3(n18036), .ZN(n18382) );
  AND2_X1 U12494 ( .A1(n13541), .A2(n13540), .ZN(n13542) );
  OR2_X1 U12495 ( .A1(n18856), .A2(n10210), .ZN(n10209) );
  AND2_X1 U12496 ( .A1(n9813), .A2(n17691), .ZN(n11672) );
  INV_X1 U12497 ( .A(n13264), .ZN(n18486) );
  OR3_X1 U12498 ( .A1(n12826), .A2(n10137), .A3(n10136), .ZN(n9831) );
  NAND2_X1 U12499 ( .A1(n10150), .A2(n10154), .ZN(n12835) );
  AND2_X1 U12500 ( .A1(n16893), .A2(n9846), .ZN(n9832) );
  AND2_X1 U12501 ( .A1(n9841), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9833) );
  OAI21_X2 U12502 ( .B1(n12812), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12811), 
        .ZN(n15196) );
  INV_X1 U12503 ( .A(n9897), .ZN(n12481) );
  NAND2_X1 U12504 ( .A1(n11281), .A2(n16149), .ZN(n16148) );
  NAND2_X1 U12505 ( .A1(n10082), .A2(n9878), .ZN(n16579) );
  NAND2_X1 U12506 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12842) );
  NAND2_X1 U12507 ( .A1(n12843), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12841) );
  NAND2_X1 U12508 ( .A1(n10287), .A2(n10285), .ZN(n16586) );
  NAND2_X1 U12509 ( .A1(n15471), .A2(n15472), .ZN(n15461) );
  NOR2_X1 U12510 ( .A1(n9860), .A2(n11977), .ZN(n9834) );
  NAND2_X1 U12511 ( .A1(n10488), .A2(n15373), .ZN(n10505) );
  AND2_X1 U12512 ( .A1(n14887), .A2(n9906), .ZN(n14992) );
  INV_X1 U12513 ( .A(n10310), .ZN(n9991) );
  NAND2_X1 U12514 ( .A1(n10991), .A2(n10277), .ZN(n10278) );
  AND2_X1 U12515 ( .A1(n10246), .A2(n9899), .ZN(n9835) );
  AND2_X1 U12516 ( .A1(n12622), .A2(n13655), .ZN(n13653) );
  AND2_X1 U12517 ( .A1(n10233), .A2(n10232), .ZN(n9836) );
  INV_X1 U12518 ( .A(n12177), .ZN(n10086) );
  INV_X1 U12519 ( .A(n10505), .ZN(n9959) );
  AND2_X1 U12520 ( .A1(n9835), .A2(n15562), .ZN(n9837) );
  AND2_X1 U12521 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9838) );
  AND2_X1 U12522 ( .A1(n16196), .A2(n14138), .ZN(n12807) );
  INV_X1 U12523 ( .A(n12807), .ZN(n10055) );
  AND2_X1 U12524 ( .A1(n16149), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9839) );
  AND2_X1 U12525 ( .A1(n10181), .A2(n15230), .ZN(n9840) );
  INV_X1 U12526 ( .A(n10100), .ZN(n10099) );
  NAND2_X1 U12527 ( .A1(n17585), .A2(n10101), .ZN(n10100) );
  AND4_X2 U12528 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11892) );
  NAND2_X1 U12529 ( .A1(n15031), .A2(n9904), .ZN(n13624) );
  NOR3_X1 U12530 ( .A1(n12831), .A2(n10147), .A3(n16638), .ZN(n12827) );
  NOR2_X1 U12531 ( .A1(n12837), .A2(n9900), .ZN(n12836) );
  NAND2_X1 U12532 ( .A1(n15211), .A2(n9903), .ZN(n16461) );
  AND2_X1 U12533 ( .A1(n13530), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9841) );
  AND2_X1 U12534 ( .A1(n10235), .A2(n9912), .ZN(n9842) );
  INV_X1 U12535 ( .A(n13216), .ZN(n17479) );
  INV_X1 U12536 ( .A(n17479), .ZN(n20437) );
  NAND2_X1 U12537 ( .A1(n9800), .A2(n14351), .ZN(n13945) );
  NAND2_X1 U12538 ( .A1(n17650), .A2(n17649), .ZN(n17635) );
  NOR3_X1 U12539 ( .A1(n12826), .A2(n10137), .A3(n16599), .ZN(n12824) );
  NOR2_X1 U12540 ( .A1(n12826), .A2(n16625), .ZN(n12825) );
  NAND2_X1 U12541 ( .A1(n9960), .A2(n9959), .ZN(n9962) );
  INV_X1 U12542 ( .A(n17891), .ZN(n19981) );
  OAI21_X1 U12543 ( .B1(n13486), .B2(n13485), .A(n13484), .ZN(n17891) );
  AND3_X1 U12544 ( .A1(n13344), .A2(n13343), .A3(n13342), .ZN(n9843) );
  AND2_X1 U12545 ( .A1(n10229), .A2(n10228), .ZN(n9844) );
  AND2_X1 U12546 ( .A1(n18846), .A2(n9833), .ZN(n9845) );
  AND2_X1 U12547 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n9846) );
  AND2_X1 U12548 ( .A1(n10018), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n9847) );
  AND2_X1 U12549 ( .A1(n9940), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9848) );
  AND2_X1 U12550 ( .A1(n10024), .A2(n9941), .ZN(n9849) );
  NAND2_X1 U12551 ( .A1(n10552), .A2(n10553), .ZN(n10634) );
  INV_X1 U12552 ( .A(n10008), .ZN(n20003) );
  OR3_X1 U12553 ( .A1(n15394), .A2(n13587), .A3(n10009), .ZN(n10008) );
  BUF_X2 U12554 ( .A(n10800), .Z(n10689) );
  OR3_X1 U12555 ( .A1(n15612), .A2(n15498), .A3(n10249), .ZN(n9851) );
  AND2_X1 U12556 ( .A1(n12900), .A2(n11564), .ZN(n9852) );
  NAND2_X1 U12557 ( .A1(n16893), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16679) );
  AND2_X1 U12558 ( .A1(n10918), .A2(n10283), .ZN(n15546) );
  NOR2_X1 U12559 ( .A1(n12842), .A2(n17597), .ZN(n12843) );
  NOR2_X1 U12560 ( .A1(n17966), .A2(n18164), .ZN(n9853) );
  AND2_X1 U12561 ( .A1(n10163), .A2(n12843), .ZN(n9854) );
  OR2_X1 U12562 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n11985), .ZN(n9855) );
  AND2_X1 U12563 ( .A1(n10094), .A2(n11624), .ZN(n9856) );
  NOR2_X1 U12564 ( .A1(n12613), .A2(n16862), .ZN(n9857) );
  AND2_X1 U12565 ( .A1(n15541), .A2(n9849), .ZN(n9858) );
  NAND2_X1 U12566 ( .A1(n10082), .A2(n10084), .ZN(n9859) );
  AND2_X1 U12567 ( .A1(n11964), .A2(n9844), .ZN(n9860) );
  AND2_X1 U12568 ( .A1(n12900), .A2(n11566), .ZN(n9861) );
  AND2_X1 U12569 ( .A1(n10172), .A2(n10171), .ZN(n9863) );
  AND2_X1 U12570 ( .A1(n10918), .A2(n10284), .ZN(n15544) );
  OR2_X1 U12571 ( .A1(n16503), .A2(n16493), .ZN(n9864) );
  AND2_X1 U12572 ( .A1(n17517), .A2(n17514), .ZN(n16850) );
  NAND2_X1 U12573 ( .A1(n11963), .A2(n11962), .ZN(n16607) );
  AND2_X1 U12574 ( .A1(n16580), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9865) );
  NOR2_X2 U12575 ( .A1(n17790), .A2(n19216), .ZN(n19128) );
  NOR2_X1 U12576 ( .A1(n19138), .A2(n13341), .ZN(n9866) );
  INV_X1 U12577 ( .A(n11895), .ZN(n16896) );
  NAND2_X1 U12578 ( .A1(n11969), .A2(n16605), .ZN(n16597) );
  INV_X1 U12579 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19035) );
  AND2_X1 U12580 ( .A1(n10033), .A2(n10031), .ZN(n9867) );
  INV_X1 U12581 ( .A(n16606), .ZN(n9992) );
  AND2_X1 U12582 ( .A1(n16580), .A2(n10290), .ZN(n12519) );
  AND2_X1 U12583 ( .A1(n15100), .A2(n17165), .ZN(n10237) );
  NAND2_X1 U12584 ( .A1(n10121), .A2(n10126), .ZN(n13599) );
  NAND2_X1 U12585 ( .A1(n9852), .A2(n16946), .ZN(n11705) );
  NAND2_X1 U12586 ( .A1(n11555), .A2(n11556), .ZN(n11559) );
  AND2_X1 U12587 ( .A1(n11895), .A2(n10316), .ZN(n9868) );
  AND4_X1 U12588 ( .A1(n13263), .A2(n13262), .A3(n13261), .A4(n13260), .ZN(
        n9869) );
  AND2_X1 U12589 ( .A1(n16412), .A2(n10292), .ZN(n9870) );
  AND4_X1 U12590 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n9871) );
  NAND2_X1 U12591 ( .A1(n15243), .A2(n15242), .ZN(n13569) );
  NAND2_X1 U12592 ( .A1(n11895), .A2(n11894), .ZN(n16681) );
  NAND2_X1 U12593 ( .A1(n11284), .A2(n16212), .ZN(n16121) );
  NAND2_X1 U12594 ( .A1(n10143), .A2(n10141), .ZN(n17402) );
  AND2_X1 U12595 ( .A1(n9979), .A2(n15762), .ZN(n9872) );
  AND2_X1 U12596 ( .A1(n10212), .A2(n19128), .ZN(n9873) );
  INV_X2 U12597 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17691) );
  AND2_X1 U12598 ( .A1(n11560), .A2(n11556), .ZN(n12916) );
  NAND3_X1 U12599 ( .A1(n13472), .A2(n19552), .A3(n13490), .ZN(n9874) );
  AND2_X1 U12600 ( .A1(n12806), .A2(n12801), .ZN(n9875) );
  INV_X1 U12601 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18073) );
  NAND2_X1 U12602 ( .A1(n16288), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9876) );
  AND2_X1 U12603 ( .A1(n16112), .A2(n10254), .ZN(n9877) );
  AND2_X1 U12604 ( .A1(n10081), .A2(n10286), .ZN(n9878) );
  NAND2_X1 U12605 ( .A1(n10037), .A2(n10035), .ZN(n9879) );
  AND2_X1 U12606 ( .A1(n16946), .A2(n11566), .ZN(n9880) );
  NOR2_X1 U12607 ( .A1(n13665), .A2(n11974), .ZN(n9881) );
  AND2_X1 U12608 ( .A1(n9970), .A2(n11566), .ZN(n9882) );
  OR2_X1 U12609 ( .A1(n10008), .A2(n10004), .ZN(n19995) );
  INV_X1 U12610 ( .A(n19995), .ZN(n13477) );
  OR2_X1 U12611 ( .A1(n11565), .A2(n11663), .ZN(n9883) );
  NOR2_X1 U12612 ( .A1(n16503), .A2(n10197), .ZN(n12578) );
  NOR2_X1 U12613 ( .A1(n16288), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9884) );
  AND2_X1 U12614 ( .A1(n15419), .A2(n11109), .ZN(n9885) );
  AND2_X1 U12615 ( .A1(n11354), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11600) );
  INV_X1 U12616 ( .A(n10272), .ZN(n10270) );
  NOR2_X1 U12617 ( .A1(n10577), .A2(n10576), .ZN(n10272) );
  NAND2_X1 U12618 ( .A1(n10082), .A2(n10081), .ZN(n12613) );
  NAND2_X1 U12619 ( .A1(n9972), .A2(n12174), .ZN(n17550) );
  OR2_X1 U12620 ( .A1(n13760), .A2(n12286), .ZN(n9886) );
  AND2_X1 U12621 ( .A1(n13352), .A2(n18912), .ZN(n9887) );
  AND2_X1 U12622 ( .A1(n10320), .A2(n9808), .ZN(n12158) );
  OR2_X1 U12623 ( .A1(n11565), .A2(n11568), .ZN(n9888) );
  AND3_X1 U12624 ( .A1(n10189), .A2(n10190), .A3(n10188), .ZN(n9889) );
  OAI21_X1 U12625 ( .B1(n12166), .B2(n12165), .A(n12164), .ZN(n13568) );
  OR2_X1 U12626 ( .A1(n12774), .A2(n21248), .ZN(n9890) );
  AND2_X1 U12627 ( .A1(n9839), .A2(n16229), .ZN(n9891) );
  INV_X1 U12628 ( .A(n9818), .ZN(n16918) );
  NAND2_X1 U12629 ( .A1(n12163), .A2(n12162), .ZN(n9892) );
  AND2_X1 U12630 ( .A1(n9988), .A2(n10309), .ZN(n9893) );
  NAND2_X1 U12631 ( .A1(n13359), .A2(n19232), .ZN(n18864) );
  AND2_X1 U12632 ( .A1(n9863), .A2(n14006), .ZN(n9894) );
  NAND2_X1 U12633 ( .A1(n12553), .A2(n12882), .ZN(n9895) );
  AND2_X1 U12634 ( .A1(n10160), .A2(n10159), .ZN(n9896) );
  AND2_X1 U12635 ( .A1(n16577), .A2(n16566), .ZN(n11988) );
  INV_X2 U12636 ( .A(n12677), .ZN(n12755) );
  OR2_X1 U12637 ( .A1(n13777), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9897) );
  NOR2_X1 U12638 ( .A1(n12831), .A2(n10146), .ZN(n12828) );
  NAND2_X1 U12639 ( .A1(n10257), .A2(n14168), .ZN(n14169) );
  NAND2_X1 U12640 ( .A1(n14887), .A2(n10749), .ZN(n14991) );
  NAND2_X1 U12641 ( .A1(n14934), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14935) );
  NOR2_X1 U12642 ( .A1(n12831), .A2(n17511), .ZN(n12832) );
  AND2_X1 U12643 ( .A1(n15031), .A2(n10182), .ZN(n13640) );
  NOR2_X1 U12644 ( .A1(n12833), .A2(n17530), .ZN(n12834) );
  NOR2_X1 U12645 ( .A1(n12837), .A2(n20309), .ZN(n12838) );
  AND3_X1 U12646 ( .A1(n10163), .A2(n10161), .A3(n12843), .ZN(n12840) );
  INV_X1 U12647 ( .A(n10030), .ZN(n15164) );
  NAND2_X1 U12648 ( .A1(n21539), .A2(n15099), .ZN(n10030) );
  AND2_X1 U12649 ( .A1(n18615), .A2(n10018), .ZN(n9898) );
  AND2_X1 U12650 ( .A1(n15339), .A2(n10247), .ZN(n9899) );
  OR2_X1 U12651 ( .A1(n10153), .A2(n20287), .ZN(n9900) );
  INV_X1 U12652 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20975) );
  NAND2_X1 U12653 ( .A1(n18997), .A2(n19119), .ZN(n18957) );
  INV_X2 U12654 ( .A(n18646), .ZN(n18726) );
  AND2_X1 U12655 ( .A1(n18724), .A2(n18624), .ZN(n18646) );
  NAND2_X1 U12656 ( .A1(n15211), .A2(n10306), .ZN(n9901) );
  AND2_X1 U12657 ( .A1(n15362), .A2(n9835), .ZN(n9902) );
  AND2_X1 U12658 ( .A1(n15212), .A2(n17477), .ZN(n9903) );
  AND2_X1 U12659 ( .A1(n10184), .A2(n13625), .ZN(n9904) );
  NAND2_X1 U12660 ( .A1(n10264), .A2(n11270), .ZN(n15248) );
  AND2_X1 U12661 ( .A1(n15211), .A2(n15212), .ZN(n9905) );
  AND2_X1 U12662 ( .A1(n10749), .A2(n10258), .ZN(n9906) );
  AND2_X1 U12663 ( .A1(n10104), .A2(n12003), .ZN(n9907) );
  NAND2_X1 U12664 ( .A1(n10502), .A2(n11341), .ZN(n12633) );
  AND2_X1 U12665 ( .A1(n10356), .A2(n12623), .ZN(n12622) );
  AND2_X1 U12666 ( .A1(n11870), .A2(n11869), .ZN(n11875) );
  INV_X1 U12667 ( .A(n10488), .ZN(n10619) );
  OR3_X1 U12668 ( .A1(n15566), .A2(n15443), .A3(n21486), .ZN(n9908) );
  AND2_X1 U12669 ( .A1(n10295), .A2(n10298), .ZN(n16440) );
  NAND2_X1 U12670 ( .A1(n10619), .A2(n10487), .ZN(n10514) );
  AND2_X1 U12671 ( .A1(n9906), .A2(n15148), .ZN(n9909) );
  OR2_X1 U12672 ( .A1(n15612), .A2(n10249), .ZN(n9910) );
  NOR3_X1 U12673 ( .A1(n15566), .A2(n10028), .A3(n10026), .ZN(n10025) );
  NAND2_X1 U12674 ( .A1(n20565), .A2(n11914), .ZN(n9911) );
  NAND2_X1 U12675 ( .A1(n20565), .A2(n11913), .ZN(n9912) );
  NAND2_X1 U12676 ( .A1(n10677), .A2(n10676), .ZN(n9913) );
  NOR2_X1 U12677 ( .A1(n13641), .A2(n16390), .ZN(n16375) );
  INV_X1 U12678 ( .A(n10105), .ZN(n10104) );
  NAND2_X1 U12679 ( .A1(n14784), .A2(n17662), .ZN(n10105) );
  AND2_X1 U12680 ( .A1(n11893), .A2(n16908), .ZN(n16899) );
  NAND2_X1 U12681 ( .A1(n14602), .A2(n14604), .ZN(n9914) );
  BUF_X1 U12682 ( .A(n13603), .Z(n18164) );
  NAND2_X1 U12683 ( .A1(n12622), .A2(n10196), .ZN(n13670) );
  AND2_X1 U12684 ( .A1(n12727), .A2(n12726), .ZN(n15562) );
  OR2_X1 U12685 ( .A1(n10015), .A2(n10017), .ZN(n9915) );
  NAND2_X1 U12686 ( .A1(n12840), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12837) );
  OR2_X1 U12687 ( .A1(n10016), .A2(n18646), .ZN(n9916) );
  NAND2_X1 U12688 ( .A1(n11875), .A2(n9836), .ZN(n10234) );
  AND2_X1 U12689 ( .A1(n20421), .A2(n20420), .ZN(n9917) );
  NAND2_X1 U12690 ( .A1(n16613), .A2(n16612), .ZN(n13667) );
  OR2_X1 U12691 ( .A1(n20247), .A2(n16640), .ZN(n9918) );
  AND2_X1 U12692 ( .A1(n16668), .A2(n13644), .ZN(n13643) );
  AND2_X1 U12693 ( .A1(n10283), .A2(n15616), .ZN(n9919) );
  AND2_X1 U12694 ( .A1(n10186), .A2(n16903), .ZN(n9920) );
  AND2_X1 U12695 ( .A1(n10306), .A2(n13004), .ZN(n9921) );
  AND2_X1 U12696 ( .A1(n15508), .A2(n10275), .ZN(n9922) );
  AND2_X1 U12697 ( .A1(n9842), .A2(n9911), .ZN(n9923) );
  AND2_X1 U12698 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9924) );
  AND2_X1 U12699 ( .A1(n13969), .A2(n10351), .ZN(n9925) );
  NOR2_X1 U12700 ( .A1(n10301), .A2(n10299), .ZN(n14509) );
  NAND2_X1 U12701 ( .A1(n12319), .A2(n10326), .ZN(n17650) );
  AND2_X1 U12702 ( .A1(n9800), .A2(n10302), .ZN(n13930) );
  NOR2_X1 U12703 ( .A1(n17532), .A2(n17531), .ZN(n14510) );
  AND2_X1 U12704 ( .A1(n17650), .A2(n10186), .ZN(n16901) );
  INV_X1 U12705 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10149) );
  INV_X1 U12706 ( .A(n18850), .ZN(n10214) );
  NOR2_X1 U12707 ( .A1(n16687), .A2(n16688), .ZN(n14290) );
  NOR2_X1 U12708 ( .A1(n9831), .A2(n16581), .ZN(n12819) );
  NAND2_X1 U12709 ( .A1(n15229), .A2(n12316), .ZN(n13578) );
  AND2_X1 U12710 ( .A1(n10196), .A2(n10195), .ZN(n9926) );
  INV_X1 U12711 ( .A(n11965), .ZN(n10230) );
  INV_X1 U12712 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10620) );
  INV_X1 U12713 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10358) );
  BUF_X1 U12714 ( .A(n11638), .Z(n20973) );
  INV_X1 U12715 ( .A(n13969), .ZN(n10299) );
  AND2_X1 U12716 ( .A1(n18482), .A2(n10071), .ZN(n9927) );
  INV_X1 U12717 ( .A(n17447), .ZN(n10159) );
  AND2_X1 U12718 ( .A1(n10219), .A2(n10218), .ZN(n9928) );
  AND2_X1 U12719 ( .A1(n10178), .A2(n14357), .ZN(n9929) );
  AND2_X1 U12720 ( .A1(n15234), .A2(n13580), .ZN(n9930) );
  AND2_X1 U12721 ( .A1(n13743), .A2(n10181), .ZN(n9931) );
  INV_X1 U12722 ( .A(n10170), .ZN(n14005) );
  NAND2_X1 U12723 ( .A1(n15234), .A2(n9863), .ZN(n10170) );
  AND2_X1 U12724 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9932) );
  OR2_X1 U12725 ( .A1(n12826), .A2(n10137), .ZN(n9933) );
  OR2_X1 U12726 ( .A1(n12831), .A2(n10147), .ZN(n9934) );
  AND2_X1 U12727 ( .A1(n10140), .A2(n15196), .ZN(n9935) );
  AND2_X1 U12728 ( .A1(n9926), .A2(n16510), .ZN(n9936) );
  OR2_X1 U12729 ( .A1(n11703), .A2(n11702), .ZN(n12151) );
  INV_X1 U12730 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9952) );
  INV_X1 U12731 ( .A(n20206), .ZN(n10001) );
  NOR2_X1 U12732 ( .A1(n12563), .A2(n16549), .ZN(n12590) );
  NOR2_X1 U12733 ( .A1(n12817), .A2(n16558), .ZN(n12564) );
  NOR2_X1 U12734 ( .A1(n17167), .A2(n21439), .ZN(n13993) );
  NOR2_X1 U12735 ( .A1(n20049), .A2(n20047), .ZN(n20038) );
  NAND2_X1 U12736 ( .A1(n18846), .A2(n9841), .ZN(n13532) );
  INV_X1 U12737 ( .A(n10053), .ZN(n17170) );
  OAI21_X1 U12738 ( .B1(n11336), .B2(n11335), .A(n11339), .ZN(n10053) );
  NOR2_X1 U12739 ( .A1(n19034), .A2(n19035), .ZN(n18087) );
  INV_X1 U12740 ( .A(n15152), .ZN(n10045) );
  OR2_X1 U12741 ( .A1(n10523), .A2(n10504), .ZN(n13989) );
  INV_X1 U12742 ( .A(n13989), .ZN(n9960) );
  NOR2_X2 U12743 ( .A1(n13440), .A2(n13439), .ZN(n19584) );
  AND2_X1 U12744 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n9937) );
  NAND2_X1 U12745 ( .A1(n18170), .A2(n18122), .ZN(n19034) );
  NOR2_X1 U12746 ( .A1(n18121), .A2(n19148), .ZN(n18170) );
  AND2_X1 U12747 ( .A1(n9846), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9938) );
  AND2_X1 U12748 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .ZN(n9939) );
  INV_X1 U12749 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10202) );
  AND3_X1 U12750 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18193) );
  INV_X1 U12751 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10128) );
  INV_X1 U12752 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U12753 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19164) );
  INV_X1 U12754 ( .A(n19164), .ZN(n10117) );
  INV_X1 U12755 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10232) );
  AND2_X1 U12756 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9940) );
  INV_X1 U12757 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n10017) );
  INV_X1 U12758 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10020) );
  INV_X1 U12759 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n10019) );
  AND2_X1 U12760 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n9941) );
  AND2_X1 U12761 ( .A1(n9849), .A2(n10023), .ZN(n9942) );
  INV_X1 U12762 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n10073) );
  OR2_X1 U12763 ( .A1(n17394), .A2(n16334), .ZN(n17306) );
  NOR3_X2 U12764 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20050), .A3(
        n19676), .ZN(n19692) );
  NOR3_X2 U12765 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20050), .A3(
        n19767), .ZN(n19785) );
  AOI22_X2 U12766 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n20571), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n20572), .ZN(n21057) );
  NOR3_X2 U12767 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20050), .A3(
        n19607), .ZN(n19603) );
  NOR3_X4 U12768 ( .A1(n13784), .A2(n11612), .A3(n21226), .ZN(n13840) );
  AOI211_X1 U12769 ( .C1(n17929), .C2(n18225), .A(n17928), .B(n17927), .ZN(
        n17932) );
  INV_X1 U12770 ( .A(n18225), .ZN(n20053) );
  NAND3_X2 U12771 ( .A1(n10319), .A2(n10353), .A3(n10318), .ZN(n11963) );
  NAND2_X2 U12772 ( .A1(n9943), .A2(n17535), .ZN(n10319) );
  NAND2_X2 U12773 ( .A1(n9944), .A2(n11910), .ZN(n10318) );
  INV_X1 U12774 ( .A(n17534), .ZN(n9944) );
  OAI211_X2 U12775 ( .C1(n11531), .C2(n17682), .A(n11530), .B(n11529), .ZN(
        n11551) );
  NAND2_X2 U12776 ( .A1(n9948), .A2(n20403), .ZN(n11586) );
  NAND2_X2 U12777 ( .A1(n9882), .A2(n9948), .ZN(n14648) );
  INV_X2 U12778 ( .A(n12900), .ZN(n9948) );
  NAND2_X1 U12779 ( .A1(n11822), .A2(n11821), .ZN(n9949) );
  INV_X2 U12780 ( .A(n11472), .ZN(n12215) );
  NOR2_X2 U12781 ( .A1(n9950), .A2(n12210), .ZN(n11496) );
  NAND4_X1 U12782 ( .A1(n12215), .A2(n11481), .A3(n12242), .A4(n11471), .ZN(
        n9950) );
  NAND3_X1 U12783 ( .A1(n11979), .A2(n11988), .A3(n11980), .ZN(n16568) );
  NOR2_X2 U12784 ( .A1(n19139), .A2(n19456), .ZN(n19138) );
  NOR2_X1 U12785 ( .A1(n9951), .A2(n18913), .ZN(n13355) );
  NAND2_X1 U12786 ( .A1(n17192), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19211) );
  NAND3_X1 U12787 ( .A1(n13321), .A2(n13323), .A3(n13322), .ZN(n17192) );
  NAND2_X1 U12788 ( .A1(n10215), .A2(n18864), .ZN(n9954) );
  INV_X1 U12789 ( .A(n9954), .ZN(n9953) );
  INV_X2 U12790 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20177) );
  INV_X2 U12791 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20160) );
  INV_X2 U12792 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20169) );
  NAND2_X2 U12794 ( .A1(n10604), .A2(n9956), .ZN(n16326) );
  NAND3_X1 U12795 ( .A1(n9962), .A2(n14116), .A3(n9957), .ZN(n9961) );
  NAND2_X2 U12796 ( .A1(n9961), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10512) );
  NAND3_X1 U12797 ( .A1(n11277), .A2(n10274), .A3(n11278), .ZN(n9963) );
  OAI21_X1 U12798 ( .B1(n14202), .B2(n11218), .A(n11217), .ZN(n11219) );
  NAND2_X2 U12799 ( .A1(n10655), .A2(n14173), .ZN(n10253) );
  AND2_X2 U12800 ( .A1(n10616), .A2(n10617), .ZN(n10655) );
  NAND3_X1 U12801 ( .A1(n15227), .A2(n15224), .A3(n12165), .ZN(n9967) );
  NAND2_X2 U12802 ( .A1(n14935), .A2(n12157), .ZN(n15227) );
  NAND2_X2 U12803 ( .A1(n9971), .A2(n12177), .ZN(n10082) );
  NAND3_X1 U12804 ( .A1(n9968), .A2(n12152), .A3(n17587), .ZN(n17590) );
  NAND3_X1 U12805 ( .A1(n10192), .A2(n9889), .A3(n9969), .ZN(P2_U3016) );
  OR2_X1 U12806 ( .A1(n12506), .A2(n17669), .ZN(n9969) );
  INV_X2 U12807 ( .A(n16946), .ZN(n9970) );
  NAND2_X1 U12808 ( .A1(n11554), .A2(n10078), .ZN(n11543) );
  OAI22_X1 U12809 ( .A1(n13907), .A2(n9888), .B1(n14648), .B2(n11567), .ZN(
        n11569) );
  OAI22_X1 U12810 ( .A1(n10060), .A2(n11743), .B1(n20587), .B2(n11709), .ZN(
        n11710) );
  OAI22_X1 U12811 ( .A1(n10060), .A2(n13025), .B1(n14014), .B2(n14027), .ZN(
        n11828) );
  OAI21_X1 U12812 ( .B1(n10484), .B2(n10514), .A(n14069), .ZN(n9975) );
  NAND2_X1 U12813 ( .A1(n14143), .A2(n14144), .ZN(n11221) );
  XNOR2_X1 U12814 ( .A(n11219), .B(n14368), .ZN(n14144) );
  NAND2_X1 U12815 ( .A1(n9978), .A2(n11214), .ZN(n14143) );
  NAND2_X1 U12816 ( .A1(n11212), .A2(n11211), .ZN(n14126) );
  NAND2_X1 U12817 ( .A1(n10595), .A2(n14030), .ZN(n13865) );
  NAND3_X1 U12818 ( .A1(n14030), .A2(n10595), .A3(n21439), .ZN(n10547) );
  OR2_X2 U12819 ( .A1(n14178), .A2(n10553), .ZN(n10595) );
  NAND2_X1 U12820 ( .A1(n9987), .A2(n9893), .ZN(n11978) );
  NOR2_X1 U12821 ( .A1(n18453), .A2(n9995), .ZN(n9994) );
  INV_X1 U12822 ( .A(n18256), .ZN(n9997) );
  OR2_X1 U12823 ( .A1(n18794), .A2(n20205), .ZN(n10003) );
  AND2_X2 U12824 ( .A1(n10011), .A2(n10010), .ZN(n15394) );
  INV_X1 U12825 ( .A(n18597), .ZN(n18592) );
  INV_X1 U12826 ( .A(n10016), .ZN(n18591) );
  INV_X1 U12827 ( .A(n10014), .ZN(n18584) );
  NAND3_X1 U12828 ( .A1(n10022), .A2(P3_EAX_REG_17__SCAN_IN), .A3(
        P3_EAX_REG_22__SCAN_IN), .ZN(n10021) );
  INV_X1 U12829 ( .A(n10025), .ZN(n17205) );
  INV_X1 U12830 ( .A(n10043), .ZN(n21355) );
  NAND2_X1 U12831 ( .A1(n15117), .A2(n15100), .ZN(n15153) );
  INV_X1 U12832 ( .A(n11311), .ZN(n11326) );
  NAND2_X1 U12833 ( .A1(n10051), .A2(n10050), .ZN(n12659) );
  NAND2_X1 U12834 ( .A1(n16196), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17336) );
  NAND2_X2 U12835 ( .A1(n10058), .A2(n20349), .ZN(n16700) );
  NAND2_X1 U12836 ( .A1(n12160), .A2(n11892), .ZN(n10058) );
  OR2_X2 U12837 ( .A1(n12152), .A2(n10323), .ZN(n12169) );
  NAND2_X1 U12838 ( .A1(n10059), .A2(n12035), .ZN(n10169) );
  XNOR2_X2 U12839 ( .A(n10059), .B(n12035), .ZN(n12900) );
  NAND2_X1 U12840 ( .A1(n11543), .A2(n11542), .ZN(n10059) );
  NAND2_X1 U12841 ( .A1(n18369), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n18357) );
  INV_X2 U12842 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20184) );
  INV_X1 U12843 ( .A(n18331), .ZN(n18326) );
  XNOR2_X1 U12844 ( .A(n11554), .B(n10078), .ZN(n12907) );
  NOR2_X1 U12845 ( .A1(n12613), .A2(n10091), .ZN(n16822) );
  INV_X4 U12846 ( .A(n11463), .ZN(n17714) );
  NAND2_X1 U12847 ( .A1(n10095), .A2(n10096), .ZN(n14932) );
  NAND2_X1 U12848 ( .A1(n16674), .A2(n10110), .ZN(n10107) );
  NAND2_X1 U12849 ( .A1(n10107), .A2(n10108), .ZN(n16634) );
  NOR2_X1 U12850 ( .A1(n16672), .A2(n12606), .ZN(n16658) );
  NOR2_X1 U12851 ( .A1(n17979), .A2(n18164), .ZN(n17967) );
  NOR2_X2 U12852 ( .A1(n17980), .A2(n18905), .ZN(n17979) );
  INV_X1 U12853 ( .A(n10120), .ZN(n18009) );
  INV_X1 U12854 ( .A(n10118), .ZN(n18008) );
  NAND2_X1 U12855 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  OR2_X1 U12856 ( .A1(n18020), .A2(n18164), .ZN(n10120) );
  INV_X1 U12857 ( .A(n19034), .ZN(n10121) );
  NAND2_X1 U12858 ( .A1(n10122), .A2(n10121), .ZN(n19001) );
  NAND2_X1 U12859 ( .A1(n18846), .A2(n10127), .ZN(n13531) );
  INV_X1 U12860 ( .A(n10140), .ZN(n16384) );
  OR2_X1 U12861 ( .A1(n13610), .A2(n15194), .ZN(n10145) );
  AOI21_X1 U12862 ( .B1(n13610), .B2(n12816), .A(n15194), .ZN(n17404) );
  NAND2_X1 U12863 ( .A1(n13610), .A2(n10144), .ZN(n10143) );
  INV_X1 U12864 ( .A(n10145), .ZN(n17420) );
  INV_X1 U12865 ( .A(n12837), .ZN(n10150) );
  NAND2_X1 U12866 ( .A1(n10150), .A2(n10151), .ZN(n12833) );
  AOI21_X1 U12867 ( .B1(n17456), .B2(n10159), .A(n15194), .ZN(n17433) );
  NAND2_X1 U12868 ( .A1(n10157), .A2(n10156), .ZN(n17432) );
  NAND2_X1 U12869 ( .A1(n17456), .A2(n10158), .ZN(n10157) );
  INV_X1 U12870 ( .A(n10160), .ZN(n17446) );
  NAND3_X1 U12871 ( .A1(n10163), .A2(n12843), .A3(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12839) );
  NOR2_X2 U12872 ( .A1(n13657), .A2(n13656), .ZN(n16613) );
  NOR2_X2 U12873 ( .A1(n16667), .A2(n16666), .ZN(n16668) );
  NAND2_X1 U12874 ( .A1(n15234), .A2(n9894), .ZN(n16687) );
  OR3_X1 U12875 ( .A1(n16447), .A2(n10176), .A3(n10174), .ZN(n12876) );
  INV_X1 U12876 ( .A(n16435), .ZN(n10176) );
  XNOR2_X1 U12877 ( .A(n13760), .B(n12286), .ZN(n13935) );
  OAI21_X1 U12878 ( .B1(n13935), .B2(n13936), .A(n9886), .ZN(n10177) );
  NAND2_X1 U12879 ( .A1(n17650), .A2(n9920), .ZN(n16902) );
  NAND2_X2 U12880 ( .A1(n10194), .A2(n13776), .ZN(n12290) );
  NAND2_X1 U12881 ( .A1(n12622), .A2(n9936), .ZN(n16513) );
  NAND3_X1 U12882 ( .A1(n10200), .A2(n10199), .A3(n12579), .ZN(n10197) );
  NAND4_X1 U12883 ( .A1(n10200), .A2(n10199), .A3(n16472), .A4(n12579), .ZN(
        n10198) );
  INV_X1 U12884 ( .A(n13359), .ZN(n13360) );
  INV_X1 U12885 ( .A(n18878), .ZN(n10201) );
  NAND3_X1 U12886 ( .A1(n13273), .A2(n13278), .A3(n10206), .ZN(n10205) );
  XNOR2_X1 U12887 ( .A(n13334), .B(n13333), .ZN(n19154) );
  NOR2_X2 U12888 ( .A1(n11814), .A2(n11806), .ZN(n11819) );
  MUX2_X1 U12889 ( .A(n12296), .B(n11797), .S(n11789), .Z(n12025) );
  NOR2_X2 U12890 ( .A1(n18256), .A2(n13227), .ZN(n13258) );
  NAND2_X1 U12891 ( .A1(n11964), .A2(n10229), .ZN(n11975) );
  NAND2_X1 U12892 ( .A1(n11964), .A2(n11965), .ZN(n11971) );
  NAND2_X1 U12893 ( .A1(n11964), .A2(n10227), .ZN(n11985) );
  AND2_X1 U12894 ( .A1(n11875), .A2(n11878), .ZN(n11897) );
  INV_X1 U12895 ( .A(n10234), .ZN(n11899) );
  OR2_X1 U12896 ( .A1(n14135), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n12679) );
  OR2_X1 U12897 ( .A1(n14135), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n12716) );
  OR2_X1 U12898 ( .A1(n14135), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n12728) );
  OR2_X1 U12899 ( .A1(n14135), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n12734) );
  OR2_X1 U12900 ( .A1(n14135), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n12742) );
  OR2_X1 U12901 ( .A1(n14135), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n12749) );
  OR2_X1 U12902 ( .A1(n14135), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12766) );
  NOR2_X1 U12903 ( .A1(n14135), .A2(n21248), .ZN(n13958) );
  NAND2_X1 U12904 ( .A1(n13954), .A2(n10237), .ZN(n13856) );
  OR2_X1 U12905 ( .A1(n15446), .A2(n10238), .ZN(P1_U2809) );
  INV_X1 U12906 ( .A(n10253), .ZN(n10252) );
  XNOR2_X1 U12907 ( .A(n10253), .B(n9913), .ZN(n11222) );
  NOR2_X1 U12908 ( .A1(n11285), .A2(n16100), .ZN(n15764) );
  INV_X1 U12909 ( .A(n11285), .ZN(n10255) );
  NAND2_X1 U12910 ( .A1(n16121), .A2(n16096), .ZN(n10256) );
  INV_X1 U12911 ( .A(n15123), .ZN(n10260) );
  NAND2_X1 U12912 ( .A1(n10264), .A2(n10263), .ZN(n16167) );
  NAND3_X1 U12913 ( .A1(n10552), .A2(n10266), .A3(n10553), .ZN(n10265) );
  NAND3_X1 U12914 ( .A1(n10552), .A2(n10553), .A3(n21439), .ZN(n10271) );
  NAND2_X1 U12915 ( .A1(n11278), .A2(n11277), .ZN(n11281) );
  INV_X1 U12916 ( .A(n10278), .ZN(n15520) );
  AND2_X1 U12917 ( .A1(n15482), .A2(n11109), .ZN(n15471) );
  AND2_X1 U12918 ( .A1(n15482), .A2(n10279), .ZN(n15420) );
  NAND2_X1 U12919 ( .A1(n15482), .A2(n10280), .ZN(n15424) );
  NAND2_X1 U12920 ( .A1(n10918), .A2(n9919), .ZN(n15609) );
  NOR2_X1 U12921 ( .A1(n12613), .A2(n16762), .ZN(n16596) );
  INV_X1 U12922 ( .A(n16762), .ZN(n10289) );
  AND2_X1 U12923 ( .A1(n16580), .A2(n9940), .ZN(n12558) );
  NAND2_X1 U12924 ( .A1(n12900), .A2(n20403), .ZN(n11574) );
  NAND2_X1 U12925 ( .A1(n12900), .A2(n10291), .ZN(n11578) );
  NAND3_X1 U12926 ( .A1(n9796), .A2(n11803), .A3(n12151), .ZN(n10321) );
  AOI21_X2 U12927 ( .B1(n16419), .B2(n16412), .A(n16415), .ZN(n16408) );
  NOR2_X2 U12928 ( .A1(n16441), .A2(n13101), .ZN(n13123) );
  NAND2_X1 U12929 ( .A1(n10294), .A2(n10293), .ZN(n16441) );
  NAND2_X1 U12930 ( .A1(n13969), .A2(n10300), .ZN(n14603) );
  INV_X1 U12931 ( .A(n14603), .ZN(n12934) );
  NAND2_X1 U12932 ( .A1(n10303), .A2(n9924), .ZN(n13966) );
  AND2_X2 U12933 ( .A1(n15211), .A2(n9921), .ZN(n16454) );
  AND2_X4 U12934 ( .A1(n16935), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13038) );
  AND2_X2 U12935 ( .A1(n10308), .A2(n16918), .ZN(n11723) );
  NAND2_X1 U12936 ( .A1(n11988), .A2(n9895), .ZN(n10317) );
  NOR2_X2 U12937 ( .A1(n10317), .A2(n16564), .ZN(n11997) );
  AOI21_X1 U12938 ( .B1(n11997), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12552), .ZN(n11998) );
  NAND3_X1 U12939 ( .A1(n10320), .A2(n12169), .A3(n11892), .ZN(n11801) );
  NAND2_X1 U12940 ( .A1(n11752), .A2(n11751), .ZN(n10322) );
  NAND2_X1 U12941 ( .A1(n11752), .A2(n10324), .ZN(n10323) );
  NOR2_X1 U12942 ( .A1(n10325), .A2(n12306), .ZN(n10324) );
  NAND2_X1 U12943 ( .A1(n12928), .A2(n12927), .ZN(n13904) );
  OAI21_X1 U12944 ( .B1(n14028), .B2(n10656), .A(n10624), .ZN(n10625) );
  NAND2_X1 U12945 ( .A1(n11264), .A2(n11263), .ZN(n15124) );
  OR2_X1 U12946 ( .A1(n16563), .A2(n17681), .ZN(n12884) );
  NOR2_X1 U12947 ( .A1(n16098), .A2(n15754), .ZN(n11285) );
  XNOR2_X1 U12948 ( .A(n12010), .B(n12009), .ZN(n12504) );
  CLKBUF_X1 U12949 ( .A(n12900), .Z(n13907) );
  AOI21_X1 U12950 ( .B1(n12504), .B2(n17592), .A(n12140), .ZN(n12183) );
  NAND2_X1 U12951 ( .A1(n16425), .A2(n10336), .ZN(n13163) );
  NAND2_X1 U12952 ( .A1(n16424), .A2(n16426), .ZN(n16425) );
  AND2_X1 U12953 ( .A1(n15189), .A2(n12238), .ZN(n17704) );
  NAND2_X1 U12954 ( .A1(n15189), .A2(n12246), .ZN(n12234) );
  OAI22_X1 U12955 ( .A1(n11792), .A2(n11786), .B1(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n21194), .ZN(n11796) );
  OAI22_X1 U12956 ( .A1(n11704), .A2(n12378), .B1(n11728), .B2(n11580), .ZN(
        n11581) );
  AOI21_X1 U12957 ( .B1(n12235), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11485), 
        .ZN(n11486) );
  NAND2_X1 U12958 ( .A1(n12489), .A2(n11484), .ZN(n12235) );
  OR2_X1 U12959 ( .A1(n11892), .A2(n12435), .ZN(n10326) );
  AND2_X1 U12960 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10327) );
  OR2_X1 U12961 ( .A1(n10617), .A2(n10616), .ZN(n10328) );
  OR2_X1 U12962 ( .A1(n12886), .A2(n17681), .ZN(n10329) );
  AND2_X1 U12963 ( .A1(n12881), .A2(n12880), .ZN(n10330) );
  AND2_X1 U12964 ( .A1(n12627), .A2(n12626), .ZN(n10331) );
  INV_X1 U12965 ( .A(n17669), .ZN(n12521) );
  NOR2_X1 U12966 ( .A1(n12625), .A2(n10341), .ZN(n12626) );
  NOR2_X1 U12967 ( .A1(n12622), .A2(n12624), .ZN(n10332) );
  AND4_X1 U12968 ( .A1(n10468), .A2(n10467), .A3(n10466), .A4(n10465), .ZN(
        n10333) );
  INV_X1 U12969 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13344) );
  NOR2_X1 U12970 ( .A1(n14510), .A2(n17533), .ZN(n10334) );
  AND2_X1 U12971 ( .A1(n11383), .A2(n11382), .ZN(n10335) );
  NOR2_X1 U12972 ( .A1(n17240), .A2(n21292), .ZN(n10337) );
  NOR2_X1 U12973 ( .A1(n15517), .A2(n21292), .ZN(n10338) );
  OR2_X1 U12974 ( .A1(n15742), .A2(n16179), .ZN(n10339) );
  AND4_X1 U12975 ( .A1(n19385), .A2(n19369), .A3(n19078), .A4(n19351), .ZN(
        n10340) );
  INV_X1 U12976 ( .A(n14871), .ZN(n12933) );
  AND2_X1 U12977 ( .A1(n10332), .A2(n17637), .ZN(n10341) );
  INV_X1 U12978 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12591) );
  OR2_X1 U12979 ( .A1(n20398), .A2(n13684), .ZN(n10342) );
  OR2_X1 U12980 ( .A1(n11717), .A2(n11621), .ZN(n10343) );
  INV_X1 U12981 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13342) );
  INV_X1 U12982 ( .A(n16554), .ZN(n12879) );
  AND3_X1 U12983 ( .A1(n11605), .A2(n11604), .A3(n11603), .ZN(n10344) );
  OR2_X1 U12984 ( .A1(n11535), .A2(n11515), .ZN(n10345) );
  INV_X1 U12985 ( .A(n11535), .ZN(n12045) );
  NOR2_X1 U12986 ( .A1(n13225), .A2(n18256), .ZN(n13310) );
  INV_X1 U12987 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17228) );
  NAND2_X1 U12988 ( .A1(n10848), .A2(n15558), .ZN(n10346) );
  INV_X1 U12989 ( .A(n14887), .ZN(n15090) );
  INV_X2 U12990 ( .A(n18579), .ZN(n18570) );
  INV_X1 U12991 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16754) );
  OR2_X1 U12992 ( .A1(n12886), .A2(n17572), .ZN(n10347) );
  OR2_X1 U12993 ( .A1(n13682), .A2(n9829), .ZN(n17566) );
  INV_X1 U12994 ( .A(n17566), .ZN(n12599) );
  AND2_X1 U12995 ( .A1(n19053), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10348) );
  INV_X1 U12996 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13343) );
  INV_X1 U12997 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11993) );
  XOR2_X1 U12998 ( .A(n12520), .B(n12541), .Z(n10349) );
  AND2_X1 U12999 ( .A1(n18974), .A2(n13529), .ZN(n10350) );
  AND2_X1 U13000 ( .A1(n20427), .A2(n20426), .ZN(n10351) );
  AND4_X1 U13001 ( .A1(n16718), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12542), .A4(n12541), .ZN(n10352) );
  AND4_X1 U13002 ( .A1(n16622), .A2(n12604), .A3(n11947), .A4(n11946), .ZN(
        n10353) );
  AND2_X1 U13003 ( .A1(n11522), .A2(n11521), .ZN(n10354) );
  XOR2_X1 U13004 ( .A(n13747), .B(n12146), .Z(n10355) );
  AND2_X1 U13005 ( .A1(n16375), .A2(n12464), .ZN(n10356) );
  AND2_X1 U13006 ( .A1(n12893), .A2(n12892), .ZN(n10357) );
  INV_X1 U13007 ( .A(n10659), .ZN(n10969) );
  XNOR2_X1 U13008 ( .A(n10588), .B(n10586), .ZN(n10626) );
  NAND2_X1 U13009 ( .A1(n11626), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11627) );
  AND2_X1 U13010 ( .A1(n12640), .A2(n11338), .ZN(n11319) );
  AND2_X1 U13011 ( .A1(n14318), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11300) );
  AND2_X1 U13012 ( .A1(n12135), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11485) );
  AOI22_X1 U13013 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U13014 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11412) );
  NAND2_X1 U13015 ( .A1(n11295), .A2(n11294), .ZN(n11317) );
  INV_X1 U13016 ( .A(n11017), .ZN(n11018) );
  OR2_X1 U13017 ( .A1(n10719), .A2(n10718), .ZN(n11254) );
  AND2_X1 U13018 ( .A1(n10585), .A2(n10584), .ZN(n10586) );
  AND2_X1 U13019 ( .A1(n14101), .A2(n14100), .ZN(n17142) );
  AND2_X1 U13020 ( .A1(n11482), .A2(n11624), .ZN(n11475) );
  AOI22_X1 U13021 ( .A1(n9812), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11440) );
  AND2_X1 U13022 ( .A1(n19008), .A2(n19221), .ZN(n13356) );
  AOI21_X1 U13023 ( .B1(n11317), .B2(n11318), .A(n11296), .ZN(n11330) );
  AND2_X1 U13024 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n11018), .ZN(
        n11019) );
  CLKBUF_X3 U13025 ( .A(n10754), .Z(n11165) );
  INV_X1 U13026 ( .A(n14547), .ZN(n10684) );
  AND2_X1 U13027 ( .A1(n10697), .A2(n10696), .ZN(n10707) );
  OR2_X1 U13028 ( .A1(n10695), .A2(n10694), .ZN(n11245) );
  AND2_X1 U13029 ( .A1(n17469), .A2(n13100), .ZN(n13078) );
  INV_X1 U13030 ( .A(n16376), .ZN(n12464) );
  XNOR2_X1 U13031 ( .A(n12036), .B(n12038), .ZN(n12035) );
  AND4_X1 U13032 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11781) );
  INV_X1 U13033 ( .A(n16899), .ZN(n11894) );
  INV_X1 U13034 ( .A(n12160), .ZN(n12165) );
  NOR2_X1 U13035 ( .A1(n11129), .A2(n15758), .ZN(n11130) );
  NOR2_X1 U13036 ( .A1(n11058), .A2(n15526), .ZN(n11059) );
  AND2_X1 U13037 ( .A1(n10631), .A2(n16141), .ZN(n10951) );
  INV_X1 U13038 ( .A(n16286), .ZN(n11276) );
  AND2_X1 U13039 ( .A1(n15358), .A2(n15359), .ZN(n12715) );
  INV_X1 U13040 ( .A(n11218), .ZN(n11310) );
  OR2_X1 U13041 ( .A1(n10512), .A2(n10593), .ZN(n10594) );
  AOI21_X1 U13042 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12896), .A(
        n11788), .ZN(n12013) );
  AND4_X1 U13043 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12301) );
  AOI21_X1 U13044 ( .B1(n12277), .B2(n12142), .A(n12276), .ZN(n12278) );
  INV_X1 U13045 ( .A(n12555), .ZN(n11994) );
  INV_X1 U13046 ( .A(n12496), .ZN(n12179) );
  OR3_X1 U13047 ( .A1(n12176), .A2(n11892), .A3(n17643), .ZN(n12177) );
  NAND2_X1 U13048 ( .A1(n9852), .A2(n9970), .ZN(n11717) );
  INV_X1 U13049 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15955) );
  INV_X1 U13050 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18426) );
  INV_X1 U13051 ( .A(n9806), .ZN(n12774) );
  NAND2_X1 U13052 ( .A1(n13870), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11151) );
  INV_X1 U13053 ( .A(n15635), .ZN(n10917) );
  AND2_X1 U13054 ( .A1(n11102), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11103) );
  NAND2_X1 U13055 ( .A1(n11059), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11101) );
  INV_X1 U13056 ( .A(n15611), .ZN(n10990) );
  NOR2_X1 U13057 ( .A1(n10849), .A2(n17236), .ZN(n10817) );
  NAND2_X1 U13058 ( .A1(n10781), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10799) );
  INV_X1 U13059 ( .A(n10631), .ZN(n11174) );
  NAND2_X1 U13060 ( .A1(n15752), .A2(n15751), .ZN(n15757) );
  AND2_X1 U13061 ( .A1(n14145), .A2(n17343), .ZN(n14964) );
  OR2_X1 U13062 ( .A1(n14156), .A2(n11198), .ZN(n11199) );
  XNOR2_X1 U13063 ( .A(n10626), .B(n11187), .ZN(n14029) );
  INV_X1 U13064 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n17138) );
  INV_X1 U13065 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17132) );
  AND4_X1 U13066 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10469) );
  AND4_X1 U13067 ( .A1(n10456), .A2(n10455), .A3(n10454), .A4(n10453), .ZN(
        n10470) );
  NAND2_X1 U13068 ( .A1(n11944), .A2(n11943), .ZN(n11941) );
  AND2_X1 U13069 ( .A1(n14353), .A2(n12906), .ZN(n13905) );
  INV_X1 U13070 ( .A(n17672), .ZN(n12878) );
  OR2_X1 U13071 ( .A1(n13160), .A2(n12919), .ZN(n12924) );
  INV_X1 U13072 ( .A(n11717), .ZN(n20807) );
  INV_X1 U13073 ( .A(n11718), .ZN(n21017) );
  NAND2_X2 U13074 ( .A1(n20016), .A2(n20009), .ZN(n19419) );
  NOR2_X1 U13075 ( .A1(n19171), .A2(n13331), .ZN(n13334) );
  AND2_X1 U13076 ( .A1(n12737), .A2(n12736), .ZN(n15629) );
  INV_X1 U13077 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17236) );
  INV_X1 U13078 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21275) );
  INV_X1 U13079 ( .A(n11174), .ZN(n11081) );
  NOR2_X1 U13080 ( .A1(n10346), .A2(n10880), .ZN(n10881) );
  AOI21_X1 U13081 ( .B1(n11231), .B2(n10872), .A(n10706), .ZN(n14416) );
  XNOR2_X1 U13082 ( .A(n15108), .B(n15107), .ZN(n15430) );
  OR2_X1 U13083 ( .A1(n10882), .A2(n15565), .ZN(n10883) );
  NAND2_X1 U13084 ( .A1(n10863), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10849) );
  NAND2_X1 U13085 ( .A1(n10751), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10767) );
  AND2_X1 U13086 ( .A1(n16291), .A2(n11185), .ZN(n16289) );
  INV_X1 U13087 ( .A(n15010), .ZN(n15074) );
  OR2_X1 U13088 ( .A1(n14499), .A2(n14323), .ZN(n15073) );
  NAND2_X1 U13089 ( .A1(n14708), .A2(n9807), .ZN(n14864) );
  AND2_X1 U13090 ( .A1(n14281), .A2(n14280), .ZN(n14311) );
  NAND2_X1 U13091 ( .A1(n16328), .A2(n14227), .ZN(n14925) );
  OR2_X1 U13092 ( .A1(n14219), .A2(n14202), .ZN(n14282) );
  AND2_X1 U13093 ( .A1(n14643), .A2(n14642), .ZN(n14695) );
  NAND2_X1 U13094 ( .A1(n14176), .A2(n14175), .ZN(n16337) );
  NOR2_X1 U13095 ( .A1(n13663), .A2(n15194), .ZN(n17457) );
  AND2_X1 U13096 ( .A1(n11928), .A2(n11927), .ZN(n13636) );
  AND2_X1 U13097 ( .A1(n12457), .A2(n12456), .ZN(n16840) );
  AND2_X1 U13098 ( .A1(n12309), .A2(n12308), .ZN(n14361) );
  AOI21_X1 U13099 ( .B1(n20245), .B2(n17591), .A(n12891), .ZN(n12892) );
  INV_X1 U13100 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16697) );
  INV_X1 U13101 ( .A(n16375), .ZN(n16389) );
  INV_X1 U13102 ( .A(n12260), .ZN(n20324) );
  OR2_X1 U13103 ( .A1(n14012), .A2(n17730), .ZN(n14024) );
  NAND2_X1 U13104 ( .A1(n20800), .A2(n21207), .ZN(n20672) );
  INV_X1 U13105 ( .A(n21178), .ZN(n20838) );
  OR2_X1 U13106 ( .A1(n21190), .A2(n21197), .ZN(n20931) );
  INV_X1 U13107 ( .A(n20800), .ZN(n21181) );
  INV_X1 U13108 ( .A(n17924), .ZN(n17925) );
  NOR2_X1 U13109 ( .A1(n17997), .A2(n18164), .ZN(n17987) );
  NOR2_X1 U13110 ( .A1(n13603), .A2(n13602), .ZN(n18041) );
  NOR2_X1 U13111 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18178), .ZN(n18157) );
  INV_X1 U13112 ( .A(n13603), .ZN(n18224) );
  NOR2_X1 U13113 ( .A1(n13480), .A2(n13490), .ZN(n16986) );
  INV_X1 U13114 ( .A(n13281), .ZN(n13282) );
  OAI21_X1 U13115 ( .B1(n15394), .B2(n18795), .A(n17091), .ZN(n18730) );
  INV_X1 U13116 ( .A(n13538), .ZN(n13539) );
  NOR2_X1 U13117 ( .A1(n17739), .A2(n19366), .ZN(n19039) );
  INV_X1 U13118 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18138) );
  NOR2_X1 U13119 ( .A1(n13521), .A2(n19456), .ZN(n13525) );
  NAND2_X1 U13120 ( .A1(n19048), .A2(n19212), .ZN(n18964) );
  OR2_X1 U13121 ( .A1(n17742), .A2(n18857), .ZN(n17792) );
  INV_X1 U13122 ( .A(n18948), .ZN(n18992) );
  NOR2_X2 U13123 ( .A1(n17784), .A2(n17790), .ZN(n19008) );
  INV_X1 U13124 ( .A(n18698), .ZN(n17790) );
  OR2_X1 U13125 ( .A1(n19324), .A2(n19457), .ZN(n19365) );
  NAND2_X1 U13126 ( .A1(n13520), .A2(n19143), .ZN(n19132) );
  INV_X1 U13127 ( .A(n19505), .ZN(n19482) );
  AOI211_X1 U13128 ( .C1(n17090), .C2(n19982), .A(n17089), .B(n17088), .ZN(
        n17097) );
  INV_X1 U13129 ( .A(n13993), .ZN(n21248) );
  INV_X1 U13130 ( .A(n21277), .ZN(n21312) );
  NAND2_X1 U13131 ( .A1(n15129), .A2(n10030), .ZN(n21317) );
  INV_X1 U13132 ( .A(n15641), .ZN(n21376) );
  INV_X1 U13133 ( .A(n15732), .ZN(n15737) );
  INV_X1 U13134 ( .A(n14553), .ZN(n14483) );
  NAND2_X1 U13135 ( .A1(n13983), .A2(n13982), .ZN(n21419) );
  NAND2_X1 U13136 ( .A1(n10956), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U13137 ( .A1(n10921), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10955) );
  INV_X1 U13138 ( .A(n17305), .ZN(n17296) );
  AND2_X1 U13139 ( .A1(n16309), .A2(n16308), .ZN(n16311) );
  INV_X1 U13140 ( .A(n14148), .ZN(n17354) );
  NOR2_X1 U13141 ( .A1(n12795), .A2(n17128), .ZN(n21432) );
  NOR2_X1 U13142 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21523) );
  INV_X1 U13143 ( .A(n14748), .ZN(n14774) );
  INV_X1 U13144 ( .A(n14864), .ZN(n14733) );
  NOR2_X1 U13145 ( .A1(n14282), .A2(n14323), .ZN(n14597) );
  NOR2_X1 U13146 ( .A1(n14460), .A2(n14564), .ZN(n15271) );
  INV_X1 U13147 ( .A(n15269), .ZN(n15028) );
  INV_X1 U13148 ( .A(n15275), .ZN(n16360) );
  INV_X1 U13149 ( .A(n21241), .ZN(n15207) );
  OR3_X1 U13150 ( .A1(n13784), .A2(n12857), .A3(n17683), .ZN(n20396) );
  INV_X1 U13151 ( .A(n20406), .ZN(n20374) );
  INV_X1 U13152 ( .A(n20399), .ZN(n20328) );
  INV_X1 U13153 ( .A(n20402), .ZN(n20385) );
  AND2_X1 U13154 ( .A1(n21239), .A2(n12854), .ZN(n20406) );
  OR2_X1 U13155 ( .A1(n12354), .A2(n12353), .ZN(n20427) );
  INV_X1 U13156 ( .A(n13653), .ZN(n13654) );
  INV_X1 U13157 ( .A(n16543), .ZN(n20492) );
  INV_X1 U13158 ( .A(n13918), .ZN(n13845) );
  INV_X1 U13159 ( .A(n15215), .ZN(n15214) );
  AND2_X1 U13160 ( .A1(n12034), .A2(n9829), .ZN(n17592) );
  AND2_X1 U13161 ( .A1(n13965), .A2(n10170), .ZN(n17641) );
  INV_X1 U13162 ( .A(n17671), .ZN(n17637) );
  AND2_X1 U13163 ( .A1(n12233), .A2(n21241), .ZN(n12505) );
  NAND2_X1 U13164 ( .A1(n17709), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16965) );
  INV_X1 U13165 ( .A(n20645), .ZN(n20621) );
  AND2_X1 U13166 ( .A1(n21190), .A2(n16968), .ZN(n20810) );
  AND2_X1 U13167 ( .A1(n20594), .A2(n21178), .ZN(n20690) );
  NOR2_X1 U13168 ( .A1(n20672), .A2(n20931), .ZN(n20724) );
  INV_X1 U13169 ( .A(n20729), .ZN(n20744) );
  AND2_X1 U13170 ( .A1(n20800), .A2(n20407), .ZN(n20594) );
  INV_X1 U13171 ( .A(n20816), .ZN(n20830) );
  AND2_X1 U13172 ( .A1(n20943), .A2(n20810), .ZN(n20840) );
  AND2_X1 U13173 ( .A1(n21190), .A2(n21197), .ZN(n21178) );
  AND2_X1 U13174 ( .A1(n20940), .A2(n20939), .ZN(n20965) );
  AND2_X1 U13175 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12032), .ZN(n21241) );
  NAND2_X1 U13176 ( .A1(n19552), .A2(n19555), .ZN(n13479) );
  XNOR2_X1 U13177 ( .A(n17926), .B(n17925), .ZN(n17929) );
  NOR2_X1 U13178 ( .A1(n20124), .A2(n17908), .ZN(n17952) );
  INV_X1 U13179 ( .A(n18259), .ZN(n18269) );
  NOR2_X1 U13180 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18015), .ZN(n17996) );
  NOR2_X1 U13181 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18035), .ZN(n18022) );
  NOR2_X1 U13182 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18080), .ZN(n18059) );
  NOR2_X1 U13183 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18105), .ZN(n18085) );
  NOR2_X1 U13184 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18129), .ZN(n18109) );
  NOR2_X1 U13185 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18198), .ZN(n18184) );
  INV_X1 U13186 ( .A(n18260), .ZN(n18200) );
  INV_X1 U13187 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18234) );
  NOR2_X1 U13188 ( .A1(n18626), .A2(n18653), .ZN(n18641) );
  AND2_X1 U13189 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18701), .ZN(n18690) );
  NOR2_X1 U13190 ( .A1(n13283), .A2(n13282), .ZN(n13284) );
  NOR2_X1 U13191 ( .A1(n18790), .A2(n18772), .ZN(n18785) );
  NAND4_X1 U13192 ( .A1(n18732), .A2(n13491), .A3(n13463), .A4(n13465), .ZN(
        n18794) );
  NAND2_X1 U13193 ( .A1(n20038), .A2(n19981), .ZN(n18796) );
  AOI21_X1 U13194 ( .B1(n17774), .B2(n19061), .A(n13539), .ZN(n13540) );
  NAND2_X1 U13195 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19039), .ZN(
        n19352) );
  NAND2_X1 U13196 ( .A1(n13526), .A2(n19114), .ZN(n19405) );
  NOR2_X1 U13197 ( .A1(n19226), .A2(n17742), .ZN(n17794) );
  NOR3_X1 U13198 ( .A1(n17790), .A2(n19983), .A3(n19533), .ZN(n19398) );
  AOI21_X2 U13199 ( .B1(n17097), .B2(n17096), .A(n20202), .ZN(n19466) );
  INV_X1 U13200 ( .A(n19886), .ZN(n19651) );
  NOR2_X1 U13201 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20153), .ZN(
        n20178) );
  INV_X1 U13202 ( .A(n19663), .ZN(n19693) );
  INV_X1 U13203 ( .A(n19909), .ZN(n19968) );
  INV_X1 U13204 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20047) );
  NAND2_X1 U13205 ( .A1(n13555), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14552)
         );
  INV_X1 U13206 ( .A(n21331), .ZN(n21349) );
  INV_X1 U13207 ( .A(n21330), .ZN(n21273) );
  NAND2_X1 U13208 ( .A1(n10030), .A2(n15118), .ZN(n21277) );
  OR2_X1 U13209 ( .A1(n15164), .A2(n15109), .ZN(n21348) );
  INV_X1 U13210 ( .A(n17279), .ZN(n15725) );
  INV_X1 U13211 ( .A(n21392), .ZN(n21414) );
  INV_X1 U13212 ( .A(n21419), .ZN(n14553) );
  INV_X2 U13213 ( .A(n21420), .ZN(n14555) );
  NAND2_X1 U13214 ( .A1(n15759), .A2(n14162), .ZN(n17305) );
  NAND2_X2 U13215 ( .A1(n17170), .A2(n11344), .ZN(n17312) );
  AOI22_X1 U13216 ( .A1(n17316), .A2(n21429), .B1(n21427), .B2(n17315), .ZN(
        n17317) );
  INV_X1 U13217 ( .A(n21429), .ZN(n17365) );
  INV_X1 U13218 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21437) );
  OR2_X1 U13219 ( .A1(n17391), .A2(n13864), .ZN(n21526) );
  OR2_X1 U13220 ( .A1(n14499), .A2(n14487), .ZN(n14789) );
  NOR2_X1 U13221 ( .A1(n14794), .A2(n14793), .ZN(n14830) );
  INV_X1 U13222 ( .A(n14036), .ZN(n14084) );
  AOI21_X1 U13223 ( .B1(n14566), .B2(n14567), .A(n14565), .ZN(n14601) );
  INV_X1 U13224 ( .A(n15271), .ZN(n15030) );
  AOI22_X1 U13225 ( .A1(n14900), .A2(n14898), .B1(n15000), .B2(n14896), .ZN(
        n14931) );
  INV_X1 U13226 ( .A(n14810), .ZN(n15309) );
  INV_X1 U13227 ( .A(n14322), .ZN(n14414) );
  INV_X1 U13228 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21439) );
  INV_X1 U13229 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21438) );
  INV_X1 U13230 ( .A(n21520), .ZN(n21443) );
  OR2_X1 U13231 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21445), .ZN(n21549) );
  AND2_X1 U13232 ( .A1(n12865), .A2(n12864), .ZN(n12866) );
  AND2_X1 U13233 ( .A1(n13771), .A2(n21241), .ZN(n20475) );
  INV_X1 U13234 ( .A(n20468), .ZN(n20500) );
  OR2_X1 U13235 ( .A1(n20532), .A2(n20541), .ZN(n20534) );
  INV_X1 U13236 ( .A(n20532), .ZN(n20543) );
  OR2_X1 U13237 ( .A1(n13784), .A2(n9829), .ZN(n13920) );
  INV_X1 U13238 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17530) );
  INV_X1 U13239 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20309) );
  INV_X1 U13240 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20373) );
  INV_X1 U13241 ( .A(n12916), .ZN(n20403) );
  NAND2_X1 U13242 ( .A1(n12505), .A2(n21214), .ZN(n17669) );
  NAND2_X1 U13243 ( .A1(n12505), .A2(n12491), .ZN(n17671) );
  NAND2_X1 U13244 ( .A1(n12505), .A2(n21221), .ZN(n17681) );
  AOI211_X2 U13245 ( .C1(n16978), .C2(n16977), .A(n20977), .B(n16976), .ZN(
        n20585) );
  NAND2_X1 U13246 ( .A1(n20810), .A2(n20594), .ZN(n20645) );
  AOI211_X2 U13247 ( .C1(n14655), .C2(n14654), .A(n20977), .B(n14653), .ZN(
        n20666) );
  INV_X1 U13248 ( .A(n20690), .ZN(n20698) );
  INV_X1 U13249 ( .A(n20724), .ZN(n20718) );
  INV_X1 U13250 ( .A(n20715), .ZN(n20747) );
  INV_X1 U13251 ( .A(n20765), .ZN(n20762) );
  NAND2_X1 U13252 ( .A1(n21028), .A2(n20594), .ZN(n20796) );
  OR2_X1 U13253 ( .A1(n20971), .A2(n20768), .ZN(n20825) );
  INV_X1 U13254 ( .A(n20840), .ZN(n20863) );
  AND2_X1 U13255 ( .A1(n20871), .A2(n20870), .ZN(n20899) );
  NAND2_X1 U13256 ( .A1(n20943), .A2(n21178), .ZN(n20930) );
  AND2_X1 U13257 ( .A1(n20937), .A2(n20936), .ZN(n20964) );
  INV_X1 U13258 ( .A(n21042), .ZN(n20992) );
  OR2_X1 U13259 ( .A1(n20971), .A2(n20970), .ZN(n21079) );
  INV_X1 U13260 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n20204) );
  AOI211_X1 U13261 ( .C1(n17930), .C2(n18311), .A(n17919), .B(n17918), .ZN(
        n17920) );
  INV_X1 U13262 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19000) );
  INV_X1 U13263 ( .A(n18248), .ZN(n18270) );
  NAND2_X1 U13264 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18273), .ZN(n18260) );
  AND2_X1 U13265 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18690), .ZN(n18693) );
  AND2_X1 U13266 ( .A1(n18670), .A2(n18715), .ZN(n18701) );
  INV_X1 U13267 ( .A(n18785), .ZN(n18759) );
  INV_X1 U13268 ( .A(n18772), .ZN(n18792) );
  OR2_X1 U13269 ( .A1(n20039), .A2(n18796), .ZN(n18833) );
  INV_X1 U13270 ( .A(n19128), .ZN(n19101) );
  NAND2_X1 U13271 ( .A1(n19529), .A2(n19533), .ZN(n19497) );
  INV_X1 U13272 ( .A(n19466), .ZN(n19533) );
  INV_X1 U13273 ( .A(n19374), .ZN(n19536) );
  INV_X1 U13274 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20029) );
  INV_X1 U13275 ( .A(n20182), .ZN(n20185) );
  INV_X1 U13276 ( .A(n20038), .ZN(n20202) );
  INV_X1 U13277 ( .A(n20150), .ZN(n20057) );
  INV_X1 U13278 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n20071) );
  INV_X1 U13279 ( .A(n17845), .ZN(n17849) );
  NAND2_X1 U13280 ( .A1(n10347), .A2(n10357), .ZN(P2_U2994) );
  NAND2_X1 U13281 ( .A1(n10329), .A2(n10331), .ZN(P2_U3026) );
  AND2_X2 U13282 ( .A1(n10365), .A2(n13885), .ZN(n10392) );
  AND2_X4 U13283 ( .A1(n10365), .A2(n10359), .ZN(n10533) );
  AOI22_X1 U13284 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13285 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10452), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13286 ( .A1(n10558), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10539), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10361) );
  AND2_X2 U13287 ( .A1(n10367), .A2(n10364), .ZN(n10439) );
  AOI22_X1 U13288 ( .A1(n10439), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10360) );
  NAND4_X1 U13289 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10377) );
  AND2_X2 U13290 ( .A1(n10365), .A2(n13868), .ZN(n10709) );
  AOI22_X1 U13291 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10375) );
  AND2_X2 U13292 ( .A1(n10365), .A2(n10364), .ZN(n10477) );
  AOI22_X1 U13293 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13294 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10373) );
  INV_X1 U13295 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10369) );
  AND2_X2 U13296 ( .A1(n10370), .A2(n14091), .ZN(n10800) );
  AND2_X4 U13297 ( .A1(n10371), .A2(n14091), .ZN(n10534) );
  AOI22_X1 U13298 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10372) );
  NAND4_X1 U13299 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        n10376) );
  AOI22_X1 U13300 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13301 ( .A1(n9828), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10558), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13302 ( .A1(n10439), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10378) );
  NAND4_X1 U13303 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10387) );
  AOI22_X1 U13304 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U13305 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n9814), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13306 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10539), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13307 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10382) );
  NAND4_X1 U13308 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10386) );
  OR2_X2 U13309 ( .A1(n10387), .A2(n10386), .ZN(n10488) );
  AOI22_X1 U13310 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10439), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13311 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13312 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13313 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10388) );
  NAND4_X1 U13314 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10398) );
  AOI22_X1 U13315 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13316 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10558), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U13317 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10539), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13318 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10393) );
  NAND4_X1 U13319 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10397) );
  OR2_X2 U13320 ( .A1(n10398), .A2(n10397), .ZN(n10487) );
  INV_X1 U13321 ( .A(n10514), .ZN(n10486) );
  NAND2_X1 U13322 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10402) );
  NAND2_X1 U13323 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10401) );
  NAND2_X1 U13324 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10400) );
  NAND2_X1 U13325 ( .A1(n10539), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10399) );
  NAND2_X1 U13326 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10406) );
  NAND2_X1 U13327 ( .A1(n10439), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10405) );
  NAND2_X1 U13328 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13329 ( .A1(n9816), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10403) );
  NAND2_X1 U13330 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10410) );
  NAND2_X1 U13331 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10409) );
  NAND2_X1 U13332 ( .A1(n10558), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10408) );
  NAND2_X1 U13333 ( .A1(n10471), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10407) );
  NAND2_X1 U13334 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10414) );
  NAND2_X1 U13335 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10413) );
  NAND2_X1 U13336 ( .A1(n10534), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10412) );
  NAND2_X1 U13337 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10411) );
  NAND4_X4 U13338 ( .A1(n10418), .A2(n10417), .A3(n10416), .A4(n10415), .ZN(
        n17165) );
  NAND2_X1 U13339 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10422) );
  NAND2_X1 U13340 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10421) );
  NAND2_X1 U13341 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10420) );
  NAND2_X1 U13342 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10419) );
  NAND2_X1 U13343 ( .A1(n10439), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10426) );
  NAND2_X1 U13344 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10425) );
  NAND2_X1 U13345 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10424) );
  NAND2_X1 U13346 ( .A1(n10471), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10423) );
  NAND2_X1 U13347 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10430) );
  NAND2_X1 U13348 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10429) );
  NAND2_X1 U13349 ( .A1(n10558), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10428) );
  NAND2_X1 U13350 ( .A1(n10539), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10427) );
  NAND2_X1 U13351 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10434) );
  NAND2_X1 U13352 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10433) );
  NAND2_X1 U13353 ( .A1(n10534), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10432) );
  NAND2_X1 U13354 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10431) );
  NAND4_X4 U13355 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n10435), .ZN(
        n15100) );
  NAND2_X1 U13356 ( .A1(n10486), .A2(n21543), .ZN(n12651) );
  NAND2_X2 U13357 ( .A1(n10532), .A2(n10487), .ZN(n12779) );
  AOI22_X1 U13358 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10392), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13359 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10452), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13360 ( .A1(n10439), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13361 ( .A1(n10558), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10440) );
  NAND4_X1 U13362 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10451) );
  AOI22_X1 U13363 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U13364 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9816), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13365 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10539), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13366 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10446) );
  NAND4_X1 U13367 ( .A1(n10449), .A2(n10448), .A3(n10447), .A4(n10446), .ZN(
        n10450) );
  NAND2_X1 U13368 ( .A1(n12789), .A2(n17165), .ZN(n13851) );
  NAND2_X1 U13369 ( .A1(n13866), .A2(n13851), .ZN(n10518) );
  AOI21_X1 U13370 ( .B1(n14049), .B2(n12651), .A(n10518), .ZN(n10496) );
  NAND2_X1 U13371 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10456) );
  NAND2_X1 U13372 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10455) );
  NAND2_X1 U13373 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10454) );
  NAND2_X1 U13374 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10453) );
  NAND2_X1 U13375 ( .A1(n11002), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10460) );
  NAND2_X1 U13376 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10459) );
  INV_X1 U13377 ( .A(n10569), .ZN(n14090) );
  NAND2_X1 U13378 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10458) );
  NAND2_X1 U13379 ( .A1(n10471), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10457) );
  NAND2_X1 U13380 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13381 ( .A1(n10534), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10463) );
  NAND2_X1 U13382 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13383 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10461) );
  NAND2_X1 U13384 ( .A1(n10439), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10468) );
  NAND2_X1 U13385 ( .A1(n10558), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10467) );
  NAND2_X1 U13386 ( .A1(n9814), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10466) );
  NAND2_X1 U13387 ( .A1(n10539), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10465) );
  AOI22_X1 U13388 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10452), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13389 ( .A1(n10439), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10569), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13390 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10558), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13391 ( .A1(n10539), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10472) );
  NAND4_X1 U13392 ( .A1(n10475), .A2(n10474), .A3(n10473), .A4(n10472), .ZN(
        n10483) );
  AOI22_X1 U13393 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13394 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9815), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13395 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13396 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10478) );
  NAND4_X1 U13397 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10482) );
  NAND2_X1 U13398 ( .A1(n12779), .A2(n14058), .ZN(n10485) );
  NAND2_X1 U13399 ( .A1(n12778), .A2(n12789), .ZN(n10495) );
  NAND2_X1 U13400 ( .A1(n10486), .A2(n10532), .ZN(n10490) );
  NAND2_X1 U13401 ( .A1(n15374), .A2(n10488), .ZN(n10489) );
  NAND2_X1 U13402 ( .A1(n13955), .A2(n12789), .ZN(n10523) );
  INV_X1 U13403 ( .A(n10523), .ZN(n10491) );
  INV_X1 U13404 ( .A(n14069), .ZN(n10493) );
  NAND2_X1 U13405 ( .A1(n10493), .A2(n15100), .ZN(n12688) );
  NAND2_X1 U13406 ( .A1(n10494), .A2(n14069), .ZN(n12661) );
  AND2_X1 U13407 ( .A1(n15100), .A2(n14058), .ZN(n10521) );
  AOI21_X1 U13408 ( .B1(n13953), .B2(n12661), .A(n10521), .ZN(n12781) );
  NAND4_X1 U13409 ( .A1(n10496), .A2(n10495), .A3(n12783), .A4(n12781), .ZN(
        n10497) );
  NAND2_X1 U13410 ( .A1(n21523), .A2(n21439), .ZN(n11347) );
  INV_X1 U13411 ( .A(n11347), .ZN(n10639) );
  NAND2_X1 U13412 ( .A1(n14318), .A2(n17132), .ZN(n10498) );
  NAND2_X1 U13413 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10598) );
  AOI21_X1 U13414 ( .B1(n10639), .B2(n14796), .A(n10590), .ZN(n10507) );
  NOR2_X1 U13415 ( .A1(n12779), .A2(n15100), .ZN(n10499) );
  AND2_X2 U13416 ( .A1(n10500), .A2(n10499), .ZN(n12647) );
  INV_X1 U13417 ( .A(n12661), .ZN(n11340) );
  INV_X1 U13418 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n10503) );
  XNOR2_X1 U13419 ( .A(n10503), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U13420 ( .A1(n15374), .A2(n13984), .ZN(n10504) );
  NAND2_X1 U13421 ( .A1(n10506), .A2(n10512), .ZN(n10510) );
  INV_X1 U13422 ( .A(n10507), .ZN(n10508) );
  NAND2_X1 U13423 ( .A1(n10510), .A2(n10509), .ZN(n10511) );
  INV_X1 U13424 ( .A(n12778), .ZN(n10517) );
  NAND2_X1 U13425 ( .A1(n10514), .A2(n14069), .ZN(n10515) );
  NAND2_X1 U13426 ( .A1(n10515), .A2(n12732), .ZN(n10516) );
  NAND2_X1 U13427 ( .A1(n12789), .A2(n13984), .ZN(n12662) );
  INV_X1 U13428 ( .A(n10518), .ZN(n10526) );
  INV_X1 U13429 ( .A(n10519), .ZN(n10520) );
  NAND2_X1 U13430 ( .A1(n10520), .A2(n15100), .ZN(n12650) );
  INV_X1 U13431 ( .A(n10521), .ZN(n10522) );
  OR2_X1 U13432 ( .A1(n10523), .A2(n10488), .ZN(n12777) );
  NAND2_X1 U13433 ( .A1(n12651), .A2(n12648), .ZN(n10524) );
  NAND2_X1 U13434 ( .A1(n10528), .A2(n10527), .ZN(n10529) );
  AND2_X1 U13435 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10529), .ZN(
        n10531) );
  INV_X1 U13436 ( .A(n10529), .ZN(n10548) );
  INV_X1 U13437 ( .A(n17167), .ZN(n17162) );
  MUX2_X1 U13438 ( .A(n17162), .B(n11347), .S(n14318), .Z(n10549) );
  NAND2_X1 U13439 ( .A1(n10532), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10576) );
  INV_X1 U13440 ( .A(n10576), .ZN(n10583) );
  AOI22_X1 U13441 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13442 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13443 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13444 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10535) );
  NAND4_X1 U13445 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10545) );
  AOI22_X1 U13446 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13447 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9815), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13448 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13449 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10540) );
  NAND4_X1 U13450 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10544) );
  NAND2_X1 U13451 ( .A1(n10583), .A2(n11205), .ZN(n10546) );
  NAND2_X1 U13452 ( .A1(n10596), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10551) );
  AND2_X1 U13453 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  NAND2_X1 U13454 ( .A1(n10551), .A2(n10550), .ZN(n10552) );
  AOI22_X1 U13455 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13456 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13457 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13458 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10554) );
  NAND4_X1 U13459 ( .A1(n10557), .A2(n10556), .A3(n10555), .A4(n10554), .ZN(
        n10564) );
  AOI22_X1 U13460 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13461 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13462 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13463 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10559) );
  NAND4_X1 U13464 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        n10563) );
  AOI22_X1 U13465 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11140), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13466 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13467 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13468 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10565) );
  NAND4_X1 U13469 ( .A1(n10568), .A2(n10567), .A3(n10566), .A4(n10565), .ZN(
        n10575) );
  AOI22_X1 U13470 ( .A1(n10569), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13471 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9816), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13472 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13473 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10570) );
  NAND4_X1 U13474 ( .A1(n10573), .A2(n10572), .A3(n10571), .A4(n10570), .ZN(
        n10574) );
  XNOR2_X1 U13475 ( .A(n11266), .B(n11206), .ZN(n10577) );
  INV_X1 U13476 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15024) );
  INV_X1 U13477 ( .A(n11206), .ZN(n11188) );
  NAND2_X1 U13478 ( .A1(n10532), .A2(n11266), .ZN(n10578) );
  OAI211_X1 U13479 ( .C1(n11188), .C2(n15100), .A(n10578), .B(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n10579) );
  INV_X1 U13480 ( .A(n10579), .ZN(n10580) );
  OAI21_X1 U13481 ( .B1(n11326), .B2(n15024), .A(n10580), .ZN(n10632) );
  NAND2_X1 U13482 ( .A1(n10583), .A2(n11266), .ZN(n11180) );
  NAND2_X1 U13483 ( .A1(n11311), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10585) );
  INV_X1 U13484 ( .A(n11266), .ZN(n10582) );
  NOR2_X1 U13485 ( .A1(n15100), .A2(n21439), .ZN(n10581) );
  AOI22_X1 U13486 ( .A1(n10583), .A2(n10582), .B1(n10581), .B2(n11205), .ZN(
        n10584) );
  INV_X1 U13487 ( .A(n10586), .ZN(n10587) );
  NOR2_X1 U13488 ( .A1(n10588), .A2(n10587), .ZN(n10589) );
  AOI21_X1 U13489 ( .B1(n11187), .B2(n10626), .A(n10589), .ZN(n10617) );
  INV_X1 U13490 ( .A(n10590), .ZN(n10592) );
  AND2_X1 U13491 ( .A1(n10592), .A2(n10591), .ZN(n10593) );
  NAND2_X1 U13492 ( .A1(n10596), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10601) );
  INV_X1 U13493 ( .A(n10598), .ZN(n10597) );
  NAND2_X1 U13494 ( .A1(n10597), .A2(n17138), .ZN(n14488) );
  NAND2_X1 U13495 ( .A1(n10598), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10599) );
  NAND2_X1 U13496 ( .A1(n14488), .A2(n10599), .ZN(n14569) );
  AOI22_X1 U13497 ( .A1(n10639), .A2(n14569), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17167), .ZN(n10600) );
  AOI22_X1 U13498 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10392), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13499 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13500 ( .A1(n9828), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9816), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13501 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10605) );
  NAND4_X1 U13502 ( .A1(n10608), .A2(n10607), .A3(n10606), .A4(n10605), .ZN(
        n10614) );
  INV_X2 U13503 ( .A(n14090), .ZN(n11156) );
  AOI22_X1 U13504 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13505 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13506 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13507 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10609) );
  NAND4_X1 U13508 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n10613) );
  AOI22_X1 U13509 ( .A1(n11338), .A2(n11204), .B1(n11311), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10615) );
  INV_X1 U13510 ( .A(n10655), .ZN(n10618) );
  NAND2_X1 U13511 ( .A1(n10618), .A2(n10328), .ZN(n14028) );
  NAND2_X1 U13512 ( .A1(n10619), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10656) );
  NAND2_X1 U13513 ( .A1(n9959), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10662) );
  NAND2_X1 U13514 ( .A1(n10659), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10622) );
  OAI21_X1 U13515 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n10657), .ZN(n21347) );
  OAI21_X1 U13516 ( .B1(n21347), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21441), 
        .ZN(n10621) );
  OAI211_X1 U13517 ( .C1(n10662), .C2(n10358), .A(n10622), .B(n10621), .ZN(
        n10623) );
  INV_X1 U13518 ( .A(n10623), .ZN(n10624) );
  NAND2_X1 U13519 ( .A1(n15421), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14166) );
  NAND2_X1 U13520 ( .A1(n10625), .A2(n14166), .ZN(n13977) );
  INV_X1 U13521 ( .A(n13977), .ZN(n10638) );
  NAND2_X1 U13522 ( .A1(n14029), .A2(n10872), .ZN(n10630) );
  AOI22_X1 U13523 ( .A1(n10659), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21441), .ZN(n10628) );
  INV_X1 U13524 ( .A(n10662), .ZN(n10678) );
  NAND2_X1 U13525 ( .A1(n10678), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10627) );
  AND2_X1 U13526 ( .A1(n10628), .A2(n10627), .ZN(n10629) );
  NOR2_X1 U13527 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10631) );
  AOI21_X1 U13528 ( .B1(n11193), .B2(n10619), .A(n21441), .ZN(n13962) );
  AOI22_X1 U13529 ( .A1(n10659), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21441), .ZN(n10636) );
  NAND2_X1 U13530 ( .A1(n10678), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10635) );
  OAI211_X1 U13531 ( .C1(n10634), .C2(n10656), .A(n10636), .B(n10635), .ZN(
        n13960) );
  MUX2_X1 U13532 ( .A(n10631), .B(n13962), .S(n13960), .Z(n13996) );
  NAND2_X1 U13533 ( .A1(n10638), .A2(n10637), .ZN(n13975) );
  NAND2_X1 U13534 ( .A1(n10596), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10641) );
  INV_X1 U13535 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17143) );
  NOR3_X1 U13536 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17138), .A3(
        n17132), .ZN(n14701) );
  NAND2_X1 U13537 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14701), .ZN(
        n14704) );
  NAND3_X1 U13538 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14635) );
  NOR2_X1 U13539 ( .A1(n14318), .A2(n14635), .ZN(n16359) );
  AOI21_X1 U13540 ( .B1(n17143), .B2(n14704), .A(n16359), .ZN(n14795) );
  AOI22_X1 U13541 ( .A1(n10639), .A2(n14795), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17167), .ZN(n10640) );
  AOI22_X1 U13542 ( .A1(n10392), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U13543 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13544 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10644) );
  INV_X1 U13545 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13546 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10643) );
  NAND4_X1 U13547 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .ZN(
        n10652) );
  AOI22_X1 U13548 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13549 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13550 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13551 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10647) );
  NAND4_X1 U13552 ( .A1(n10650), .A2(n10649), .A3(n10648), .A4(n10647), .ZN(
        n10651) );
  AOI22_X1 U13553 ( .A1(n11338), .A2(n11224), .B1(n11311), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10653) );
  OR2_X1 U13554 ( .A1(n14202), .A2(n10656), .ZN(n10665) );
  OAI21_X1 U13555 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10658), .A(
        n10680), .ZN(n15174) );
  AOI22_X1 U13556 ( .A1(n10631), .A2(n15174), .B1(n15421), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10661) );
  INV_X1 U13557 ( .A(n10969), .ZN(n10753) );
  NAND2_X1 U13558 ( .A1(n10753), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10660) );
  OAI211_X1 U13559 ( .C1(n10662), .C2(n10369), .A(n10661), .B(n10660), .ZN(
        n10663) );
  INV_X1 U13560 ( .A(n10663), .ZN(n10664) );
  AOI22_X1 U13561 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10533), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13562 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11163), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13563 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13564 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10666) );
  NAND4_X1 U13565 ( .A1(n10669), .A2(n10668), .A3(n10667), .A4(n10666), .ZN(
        n10675) );
  AOI22_X1 U13566 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13567 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n9827), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13568 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11088), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13569 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10670) );
  NAND4_X1 U13570 ( .A1(n10673), .A2(n10672), .A3(n10671), .A4(n10670), .ZN(
        n10674) );
  NAND2_X1 U13571 ( .A1(n11338), .A2(n11232), .ZN(n10677) );
  NAND2_X1 U13572 ( .A1(n11311), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10676) );
  NAND2_X1 U13573 ( .A1(n10678), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10682) );
  AOI21_X1 U13574 ( .B1(n14629), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10679) );
  AOI21_X1 U13575 ( .B1(n10753), .B2(P1_EAX_REG_4__SCAN_IN), .A(n10679), .ZN(
        n10681) );
  AOI21_X1 U13576 ( .B1(n14629), .B2(n10680), .A(n10699), .ZN(n21340) );
  AOI22_X1 U13577 ( .A1(n10682), .A2(n10681), .B1(n10631), .B2(n21340), .ZN(
        n10683) );
  AOI21_X1 U13578 ( .B1(n11222), .B2(n10872), .A(n10683), .ZN(n14547) );
  AOI22_X1 U13579 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13580 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13581 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13582 ( .A1(n10439), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10685) );
  NAND4_X1 U13583 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        n10695) );
  AOI22_X1 U13584 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13585 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9816), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10692) );
  INV_X1 U13586 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15940) );
  AOI22_X1 U13587 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13588 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10690) );
  NAND4_X1 U13589 ( .A1(n10693), .A2(n10692), .A3(n10691), .A4(n10690), .ZN(
        n10694) );
  NAND2_X1 U13590 ( .A1(n11338), .A2(n11245), .ZN(n10697) );
  NAND2_X1 U13591 ( .A1(n11311), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10696) );
  INV_X1 U13592 ( .A(n10707), .ZN(n10698) );
  INV_X1 U13593 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n10705) );
  INV_X1 U13594 ( .A(n10722), .ZN(n10703) );
  INV_X1 U13595 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10701) );
  INV_X1 U13596 ( .A(n10699), .ZN(n10700) );
  NAND2_X1 U13597 ( .A1(n10701), .A2(n10700), .ZN(n10702) );
  NAND2_X1 U13598 ( .A1(n10703), .A2(n10702), .ZN(n21325) );
  AOI22_X1 U13599 ( .A1(n21325), .A2(n11081), .B1(n15421), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10704) );
  OAI21_X1 U13600 ( .B1(n10969), .B2(n10705), .A(n10704), .ZN(n10706) );
  AOI22_X1 U13601 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13602 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13603 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13604 ( .A1(n10439), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10710) );
  NAND4_X1 U13605 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n10719) );
  AOI22_X1 U13606 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13607 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13608 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13609 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10714) );
  NAND4_X1 U13610 ( .A1(n10717), .A2(n10716), .A3(n10715), .A4(n10714), .ZN(
        n10718) );
  NAND2_X1 U13611 ( .A1(n11338), .A2(n11254), .ZN(n10721) );
  NAND2_X1 U13612 ( .A1(n11311), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10720) );
  NAND2_X1 U13613 ( .A1(n10721), .A2(n10720), .ZN(n10727) );
  NOR2_X1 U13614 ( .A1(n10722), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10723) );
  NOR2_X1 U13615 ( .A1(n10731), .A2(n10723), .ZN(n21311) );
  INV_X1 U13616 ( .A(n15421), .ZN(n10894) );
  INV_X1 U13617 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14987) );
  OAI22_X1 U13618 ( .A1(n21311), .A2(n11174), .B1(n10894), .B2(n14987), .ZN(
        n10724) );
  AOI21_X1 U13619 ( .B1(n10753), .B2(P1_EAX_REG_6__SCAN_IN), .A(n10724), .ZN(
        n10725) );
  INV_X1 U13620 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15059) );
  NAND2_X1 U13621 ( .A1(n11338), .A2(n11266), .ZN(n10729) );
  OAI21_X1 U13622 ( .B1(n15059), .B2(n11326), .A(n10729), .ZN(n10730) );
  INV_X1 U13623 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10733) );
  OAI21_X1 U13624 ( .B1(n10731), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n10750), .ZN(n21302) );
  AOI22_X1 U13625 ( .A1(n21302), .A2(n11081), .B1(n15421), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10732) );
  OAI21_X1 U13626 ( .B1(n10969), .B2(n10733), .A(n10732), .ZN(n10734) );
  AOI22_X1 U13627 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10392), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13628 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13629 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13630 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10735) );
  NAND4_X1 U13631 ( .A1(n10738), .A2(n10737), .A3(n10736), .A4(n10735), .ZN(
        n10744) );
  AOI22_X1 U13632 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U13633 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13634 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13635 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10739) );
  NAND4_X1 U13636 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n10743) );
  OAI21_X1 U13637 ( .B1(n10744), .B2(n10743), .A(n10872), .ZN(n10748) );
  NAND2_X1 U13638 ( .A1(n10753), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10747) );
  XNOR2_X1 U13639 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n10750), .ZN(
        n21285) );
  INV_X1 U13640 ( .A(n21285), .ZN(n10745) );
  AOI22_X1 U13641 ( .A1(n15421), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n10631), .B2(n10745), .ZN(n10746) );
  XNOR2_X1 U13642 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10767), .ZN(
        n21281) );
  OAI22_X1 U13643 ( .A1(n21281), .A2(n11174), .B1(n10894), .B2(n21275), .ZN(
        n10752) );
  AOI21_X1 U13644 ( .B1(n10753), .B2(P1_EAX_REG_9__SCAN_IN), .A(n10752), .ZN(
        n10766) );
  AOI22_X1 U13645 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11140), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13646 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13647 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13648 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10755) );
  NAND4_X1 U13649 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10764) );
  AOI22_X1 U13650 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13651 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9816), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13652 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13653 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10759) );
  NAND4_X1 U13654 ( .A1(n10762), .A2(n10761), .A3(n10760), .A4(n10759), .ZN(
        n10763) );
  OAI21_X1 U13655 ( .B1(n10764), .B2(n10763), .A(n10872), .ZN(n10765) );
  INV_X1 U13656 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15167) );
  XNOR2_X1 U13657 ( .A(n15167), .B(n10781), .ZN(n17303) );
  AOI22_X1 U13658 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13659 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13660 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13661 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10768) );
  NAND4_X1 U13662 ( .A1(n10771), .A2(n10770), .A3(n10769), .A4(n10768), .ZN(
        n10777) );
  AOI22_X1 U13663 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13664 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13665 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13666 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10772) );
  NAND4_X1 U13667 ( .A1(n10775), .A2(n10774), .A3(n10773), .A4(n10772), .ZN(
        n10776) );
  OR2_X1 U13668 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  AOI22_X1 U13669 ( .A1(n10872), .A2(n10778), .B1(n15421), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10780) );
  NAND2_X1 U13670 ( .A1(n10753), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n10779) );
  OAI211_X1 U13671 ( .C1(n17303), .C2(n11174), .A(n10780), .B(n10779), .ZN(
        n15148) );
  INV_X1 U13672 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10782) );
  XNOR2_X1 U13673 ( .A(n10799), .B(n10782), .ZN(n16172) );
  NAND2_X1 U13674 ( .A1(n16172), .A2(n11081), .ZN(n10784) );
  AOI22_X1 U13675 ( .A1(n10753), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n15421), 
        .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10783) );
  NAND2_X1 U13676 ( .A1(n10784), .A2(n10783), .ZN(n10796) );
  AOI22_X1 U13677 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13678 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10439), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13679 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10786) );
  AOI22_X1 U13680 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10785) );
  NAND4_X1 U13681 ( .A1(n10788), .A2(n10787), .A3(n10786), .A4(n10785), .ZN(
        n10794) );
  AOI22_X1 U13682 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13683 ( .A1(n9816), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13684 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13685 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10789) );
  NAND4_X1 U13686 ( .A1(n10792), .A2(n10791), .A3(n10790), .A4(n10789), .ZN(
        n10793) );
  OR2_X1 U13687 ( .A1(n10794), .A2(n10793), .ZN(n10795) );
  AND2_X1 U13688 ( .A1(n10872), .A2(n10795), .ZN(n15324) );
  NAND2_X1 U13689 ( .A1(n15322), .A2(n15324), .ZN(n15323) );
  INV_X1 U13690 ( .A(n10796), .ZN(n10797) );
  XNOR2_X1 U13691 ( .A(n10882), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17278) );
  NAND2_X1 U13692 ( .A1(n17278), .A2(n11081), .ZN(n10816) );
  AOI22_X1 U13693 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10439), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13694 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9815), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13695 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13696 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11134), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10801) );
  NAND4_X1 U13697 ( .A1(n10804), .A2(n10803), .A3(n10802), .A4(n10801), .ZN(
        n10812) );
  AOI22_X1 U13698 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11140), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13699 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13700 ( .A1(n9828), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U13701 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10806) );
  AOI21_X1 U13702 ( .B1(n10534), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n10631), .ZN(n10805) );
  AND2_X1 U13703 ( .A1(n10806), .A2(n10805), .ZN(n10807) );
  NAND4_X1 U13704 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n10811) );
  INV_X1 U13705 ( .A(n13910), .ZN(n13870) );
  NAND2_X1 U13706 ( .A1(n11151), .A2(n11174), .ZN(n10950) );
  OAI21_X1 U13707 ( .B1(n10812), .B2(n10811), .A(n10950), .ZN(n10814) );
  AOI22_X1 U13708 ( .A1(n10753), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21441), .ZN(n10813) );
  NAND2_X1 U13709 ( .A1(n10814), .A2(n10813), .ZN(n10815) );
  NAND2_X1 U13710 ( .A1(n10816), .A2(n10815), .ZN(n15560) );
  INV_X1 U13711 ( .A(n15560), .ZN(n10848) );
  XNOR2_X1 U13712 ( .A(n10817), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16163) );
  AOI22_X1 U13713 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10392), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13714 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13715 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U13716 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10818) );
  NAND4_X1 U13717 ( .A1(n10821), .A2(n10820), .A3(n10819), .A4(n10818), .ZN(
        n10827) );
  AOI22_X1 U13718 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10439), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13719 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10452), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13720 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13721 ( .A1(n9816), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10822) );
  NAND4_X1 U13722 ( .A1(n10825), .A2(n10824), .A3(n10823), .A4(n10822), .ZN(
        n10826) );
  OAI21_X1 U13723 ( .B1(n10827), .B2(n10826), .A(n10872), .ZN(n10830) );
  NAND2_X1 U13724 ( .A1(n10753), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10829) );
  NAND2_X1 U13725 ( .A1(n15421), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10828) );
  NAND3_X1 U13726 ( .A1(n10830), .A2(n10829), .A3(n10828), .ZN(n10831) );
  AOI21_X1 U13727 ( .B1(n16163), .B2(n11081), .A(n10831), .ZN(n15584) );
  XOR2_X1 U13728 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n10832), .Z(
        n17283) );
  INV_X1 U13729 ( .A(n17283), .ZN(n10847) );
  AOI22_X1 U13730 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10439), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13731 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13732 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13733 ( .A1(n9828), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10833) );
  NAND4_X1 U13734 ( .A1(n10836), .A2(n10835), .A3(n10834), .A4(n10833), .ZN(
        n10842) );
  AOI22_X1 U13735 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13736 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13737 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9815), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13738 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10837) );
  NAND4_X1 U13739 ( .A1(n10840), .A2(n10839), .A3(n10838), .A4(n10837), .ZN(
        n10841) );
  OAI21_X1 U13740 ( .B1(n10842), .B2(n10841), .A(n10872), .ZN(n10845) );
  NAND2_X1 U13741 ( .A1(n10753), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10844) );
  NAND2_X1 U13742 ( .A1(n15421), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10843) );
  NAND3_X1 U13743 ( .A1(n10845), .A2(n10844), .A3(n10843), .ZN(n10846) );
  AOI21_X1 U13744 ( .B1(n10847), .B2(n11081), .A(n10846), .ZN(n15573) );
  NOR2_X1 U13745 ( .A1(n15584), .A2(n15573), .ZN(n15558) );
  XNOR2_X1 U13746 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10849), .ZN(
        n17292) );
  AOI22_X1 U13747 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13748 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13749 ( .A1(n10689), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U13750 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10850) );
  NAND4_X1 U13751 ( .A1(n10853), .A2(n10852), .A3(n10851), .A4(n10850), .ZN(
        n10859) );
  AOI22_X1 U13752 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13753 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13754 ( .A1(n9814), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13755 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10854) );
  NAND4_X1 U13756 ( .A1(n10857), .A2(n10856), .A3(n10855), .A4(n10854), .ZN(
        n10858) );
  OR2_X1 U13757 ( .A1(n10859), .A2(n10858), .ZN(n10860) );
  AOI22_X1 U13758 ( .A1(n10872), .A2(n10860), .B1(n15421), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U13759 ( .A1(n10753), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10861) );
  OAI211_X1 U13760 ( .C1(n17292), .C2(n11174), .A(n10862), .B(n10861), .ZN(
        n15337) );
  XNOR2_X1 U13761 ( .A(n10863), .B(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17245) );
  NAND2_X1 U13762 ( .A1(n17245), .A2(n11081), .ZN(n10879) );
  AOI22_X1 U13763 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11140), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13764 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13765 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10452), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13766 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10864) );
  NAND4_X1 U13767 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(
        n10874) );
  AOI22_X1 U13768 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10533), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13769 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11164), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13770 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13771 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10868) );
  NAND4_X1 U13772 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .ZN(
        n10873) );
  OAI21_X1 U13773 ( .B1(n10874), .B2(n10873), .A(n10872), .ZN(n10877) );
  NAND2_X1 U13774 ( .A1(n10753), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U13775 ( .A1(n15421), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10875) );
  AND3_X1 U13776 ( .A1(n10877), .A2(n10876), .A3(n10875), .ZN(n10878) );
  NAND2_X1 U13777 ( .A1(n10879), .A2(n10878), .ZN(n15735) );
  AND2_X2 U13778 ( .A1(n15335), .A2(n10881), .ZN(n15369) );
  INV_X1 U13779 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15565) );
  AOI21_X1 U13780 ( .B1(n17228), .B2(n10883), .A(n10919), .ZN(n17273) );
  OR2_X1 U13781 ( .A1(n17273), .A2(n11174), .ZN(n10899) );
  INV_X1 U13782 ( .A(n11151), .ZN(n11177) );
  AOI22_X1 U13783 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13784 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U13785 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U13786 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10884) );
  NAND4_X1 U13787 ( .A1(n10887), .A2(n10886), .A3(n10885), .A4(n10884), .ZN(
        n10893) );
  AOI22_X1 U13788 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13789 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9815), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13790 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U13791 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10888) );
  NAND4_X1 U13792 ( .A1(n10891), .A2(n10890), .A3(n10889), .A4(n10888), .ZN(
        n10892) );
  OR2_X1 U13793 ( .A1(n10893), .A2(n10892), .ZN(n10897) );
  INV_X1 U13794 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n10895) );
  OAI22_X1 U13795 ( .A1(n10969), .A2(n10895), .B1(n10894), .B2(n17228), .ZN(
        n10896) );
  AOI21_X1 U13796 ( .B1(n11177), .B2(n10897), .A(n10896), .ZN(n10898) );
  NAND2_X1 U13797 ( .A1(n10899), .A2(n10898), .ZN(n15368) );
  INV_X2 U13798 ( .A(n15367), .ZN(n10918) );
  INV_X1 U13799 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10900) );
  XNOR2_X1 U13800 ( .A(n10919), .B(n10900), .ZN(n17221) );
  NAND2_X1 U13801 ( .A1(n17221), .A2(n11081), .ZN(n10916) );
  AOI22_X1 U13802 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10439), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U13803 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11165), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U13804 ( .A1(n10476), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11134), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13805 ( .A1(n9816), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10901) );
  NAND4_X1 U13806 ( .A1(n10904), .A2(n10903), .A3(n10902), .A4(n10901), .ZN(
        n10912) );
  AOI22_X1 U13807 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13808 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13809 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10908) );
  NAND2_X1 U13810 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10906) );
  AOI21_X1 U13811 ( .B1(n10534), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n10631), .ZN(n10905) );
  AND2_X1 U13812 ( .A1(n10906), .A2(n10905), .ZN(n10907) );
  NAND4_X1 U13813 ( .A1(n10910), .A2(n10909), .A3(n10908), .A4(n10907), .ZN(
        n10911) );
  OAI21_X1 U13814 ( .B1(n10912), .B2(n10911), .A(n10950), .ZN(n10914) );
  AOI22_X1 U13815 ( .A1(n10753), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21441), .ZN(n10913) );
  NAND2_X1 U13816 ( .A1(n10914), .A2(n10913), .ZN(n10915) );
  NAND2_X1 U13817 ( .A1(n10916), .A2(n10915), .ZN(n15635) );
  OR2_X1 U13818 ( .A1(n10921), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10922) );
  NAND2_X1 U13819 ( .A1(n10922), .A2(n10955), .ZN(n17272) );
  AOI22_X1 U13820 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U13821 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13822 ( .A1(n9816), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U13823 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10923) );
  NAND4_X1 U13824 ( .A1(n10926), .A2(n10925), .A3(n10924), .A4(n10923), .ZN(
        n10932) );
  AOI22_X1 U13825 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U13826 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13827 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13828 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10927) );
  NAND4_X1 U13829 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n10931) );
  NOR2_X1 U13830 ( .A1(n10932), .A2(n10931), .ZN(n10933) );
  NOR2_X1 U13831 ( .A1(n11151), .A2(n10933), .ZN(n10936) );
  INV_X1 U13832 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15705) );
  NAND2_X1 U13833 ( .A1(n21441), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10934) );
  OAI211_X1 U13834 ( .C1(n10969), .C2(n15705), .A(n11174), .B(n10934), .ZN(
        n10935) );
  OAI22_X1 U13835 ( .A1(n17272), .A2(n11174), .B1(n10936), .B2(n10935), .ZN(
        n15626) );
  AOI22_X1 U13836 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11163), .B1(
        n10709), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13837 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13838 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10940) );
  NAND2_X1 U13839 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10938) );
  AOI21_X1 U13840 ( .B1(n10534), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n10631), .ZN(n10937) );
  AND2_X1 U13841 ( .A1(n10938), .A2(n10937), .ZN(n10939) );
  NAND4_X1 U13842 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10948) );
  AOI22_X1 U13843 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11088), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U13844 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10444), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U13845 ( .A1(n9816), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13846 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11134), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10943) );
  NAND4_X1 U13847 ( .A1(n10946), .A2(n10945), .A3(n10944), .A4(n10943), .ZN(
        n10947) );
  OR2_X1 U13848 ( .A1(n10948), .A2(n10947), .ZN(n10949) );
  NAND2_X1 U13849 ( .A1(n10950), .A2(n10949), .ZN(n10953) );
  AOI22_X1 U13850 ( .A1(n10753), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21441), .ZN(n10952) );
  XNOR2_X1 U13851 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n10955), .ZN(
        n16141) );
  AOI21_X1 U13852 ( .B1(n10953), .B2(n10952), .A(n10951), .ZN(n15545) );
  INV_X1 U13853 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10954) );
  OR2_X1 U13854 ( .A1(n10956), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10957) );
  NAND2_X1 U13855 ( .A1(n10957), .A2(n11017), .ZN(n17266) );
  INV_X1 U13856 ( .A(n17266), .ZN(n10973) );
  AOI22_X1 U13857 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13858 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13859 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13860 ( .A1(n9814), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10958) );
  NAND4_X1 U13861 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10967) );
  AOI22_X1 U13862 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11088), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U13863 ( .A1(n10452), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U13864 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U13865 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10962) );
  NAND4_X1 U13866 ( .A1(n10965), .A2(n10964), .A3(n10963), .A4(n10962), .ZN(
        n10966) );
  OR2_X1 U13867 ( .A1(n10967), .A2(n10966), .ZN(n10971) );
  INV_X1 U13868 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15693) );
  NAND2_X1 U13869 ( .A1(n21441), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10968) );
  OAI211_X1 U13870 ( .C1(n10969), .C2(n15693), .A(n11174), .B(n10968), .ZN(
        n10970) );
  AOI21_X1 U13871 ( .B1(n11177), .B2(n10971), .A(n10970), .ZN(n10972) );
  AOI21_X1 U13872 ( .B1(n10973), .B2(n11081), .A(n10972), .ZN(n15616) );
  INV_X2 U13873 ( .A(n15609), .ZN(n10991) );
  AOI22_X1 U13874 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U13875 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U13876 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U13877 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10974) );
  NAND4_X1 U13878 ( .A1(n10977), .A2(n10976), .A3(n10975), .A4(n10974), .ZN(
        n10983) );
  AOI22_X1 U13879 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U13880 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U13881 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U13882 ( .A1(n10800), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10978) );
  NAND4_X1 U13883 ( .A1(n10981), .A2(n10980), .A3(n10979), .A4(n10978), .ZN(
        n10982) );
  NOR2_X1 U13884 ( .A1(n10983), .A2(n10982), .ZN(n10987) );
  INV_X1 U13885 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10984) );
  AOI21_X1 U13886 ( .B1(n10984), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10985) );
  AOI21_X1 U13887 ( .B1(n10753), .B2(P1_EAX_REG_22__SCAN_IN), .A(n10985), .ZN(
        n10986) );
  OAI21_X1 U13888 ( .B1(n11151), .B2(n10987), .A(n10986), .ZN(n10989) );
  XNOR2_X1 U13889 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n11017), .ZN(
        n17257) );
  NAND2_X1 U13890 ( .A1(n10631), .A2(n17257), .ZN(n10988) );
  NAND2_X1 U13891 ( .A1(n10989), .A2(n10988), .ZN(n15611) );
  AOI22_X1 U13892 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U13893 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13894 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U13895 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10992) );
  NAND4_X1 U13896 ( .A1(n10995), .A2(n10994), .A3(n10993), .A4(n10992), .ZN(
        n11001) );
  AOI22_X1 U13897 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U13898 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U13899 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U13900 ( .A1(n10444), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10996) );
  NAND4_X1 U13901 ( .A1(n10999), .A2(n10998), .A3(n10997), .A4(n10996), .ZN(
        n11000) );
  NOR2_X1 U13902 ( .A1(n11001), .A2(n11000), .ZN(n11024) );
  AOI22_X1 U13903 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11002), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U13904 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U13905 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U13906 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11003) );
  NAND4_X1 U13907 ( .A1(n11006), .A2(n11005), .A3(n11004), .A4(n11003), .ZN(
        n11012) );
  AOI22_X1 U13908 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U13909 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U13910 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9816), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U13911 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11007) );
  NAND4_X1 U13912 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n11011) );
  NOR2_X1 U13913 ( .A1(n11012), .A2(n11011), .ZN(n11025) );
  XNOR2_X1 U13914 ( .A(n11024), .B(n11025), .ZN(n11016) );
  NAND2_X1 U13915 ( .A1(n21441), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11013) );
  NAND2_X1 U13916 ( .A1(n11174), .A2(n11013), .ZN(n11014) );
  AOI21_X1 U13917 ( .B1(n10659), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11014), .ZN(
        n11015) );
  OAI21_X1 U13918 ( .B1(n11151), .B2(n11016), .A(n11015), .ZN(n11023) );
  INV_X1 U13919 ( .A(n11019), .ZN(n11020) );
  INV_X1 U13920 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15535) );
  NAND2_X1 U13921 ( .A1(n11020), .A2(n15535), .ZN(n11021) );
  AND2_X1 U13922 ( .A1(n11058), .A2(n11021), .ZN(n15534) );
  NAND2_X1 U13923 ( .A1(n15534), .A2(n11081), .ZN(n11022) );
  NAND2_X1 U13924 ( .A1(n11023), .A2(n11022), .ZN(n15533) );
  NOR2_X1 U13925 ( .A1(n11025), .A2(n11024), .ZN(n11043) );
  AOI22_X1 U13926 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U13927 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U13928 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U13929 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11026) );
  NAND4_X1 U13930 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(
        n11035) );
  AOI22_X1 U13931 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U13932 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U13933 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U13934 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11030) );
  NAND4_X1 U13935 ( .A1(n11033), .A2(n11032), .A3(n11031), .A4(n11030), .ZN(
        n11034) );
  OR2_X1 U13936 ( .A1(n11035), .A2(n11034), .ZN(n11042) );
  XNOR2_X1 U13937 ( .A(n11043), .B(n11042), .ZN(n11039) );
  NAND2_X1 U13938 ( .A1(n21441), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11036) );
  NAND2_X1 U13939 ( .A1(n11174), .A2(n11036), .ZN(n11037) );
  AOI21_X1 U13940 ( .B1(n10659), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11037), .ZN(
        n11038) );
  OAI21_X1 U13941 ( .B1(n11039), .B2(n11151), .A(n11038), .ZN(n11041) );
  XNOR2_X1 U13942 ( .A(n11058), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15525) );
  NAND2_X1 U13943 ( .A1(n15525), .A2(n11081), .ZN(n11040) );
  NAND2_X1 U13944 ( .A1(n11041), .A2(n11040), .ZN(n15521) );
  NAND2_X1 U13945 ( .A1(n11043), .A2(n11042), .ZN(n11065) );
  AOI22_X1 U13946 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9827), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U13947 ( .A1(n10477), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U13948 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U13949 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11044) );
  NAND4_X1 U13950 ( .A1(n11047), .A2(n11046), .A3(n11045), .A4(n11044), .ZN(
        n11053) );
  AOI22_X1 U13951 ( .A1(n10533), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10439), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11051) );
  AOI22_X1 U13952 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U13953 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U13954 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11048) );
  NAND4_X1 U13955 ( .A1(n11051), .A2(n11050), .A3(n11049), .A4(n11048), .ZN(
        n11052) );
  NOR2_X1 U13956 ( .A1(n11053), .A2(n11052), .ZN(n11066) );
  XNOR2_X1 U13957 ( .A(n11065), .B(n11066), .ZN(n11057) );
  NAND2_X1 U13958 ( .A1(n21441), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11054) );
  NAND2_X1 U13959 ( .A1(n11174), .A2(n11054), .ZN(n11055) );
  AOI21_X1 U13960 ( .B1(n10659), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11055), .ZN(
        n11056) );
  OAI21_X1 U13961 ( .B1(n11057), .B2(n11151), .A(n11056), .ZN(n11064) );
  INV_X1 U13962 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15526) );
  INV_X1 U13963 ( .A(n11059), .ZN(n11061) );
  INV_X1 U13964 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11060) );
  NAND2_X1 U13965 ( .A1(n11061), .A2(n11060), .ZN(n11062) );
  NAND2_X1 U13966 ( .A1(n11101), .A2(n11062), .ZN(n16117) );
  NOR2_X1 U13967 ( .A1(n11066), .A2(n11065), .ZN(n11096) );
  AOI22_X1 U13968 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10533), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U13969 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U13970 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U13971 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11067) );
  NAND4_X1 U13972 ( .A1(n11070), .A2(n11069), .A3(n11068), .A4(n11067), .ZN(
        n11076) );
  AOI22_X1 U13973 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U13974 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9816), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U13975 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U13976 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11071) );
  NAND4_X1 U13977 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n11075) );
  OR2_X1 U13978 ( .A1(n11076), .A2(n11075), .ZN(n11095) );
  XNOR2_X1 U13979 ( .A(n11096), .B(n11095), .ZN(n11080) );
  NAND2_X1 U13980 ( .A1(n21441), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11077) );
  NAND2_X1 U13981 ( .A1(n11174), .A2(n11077), .ZN(n11078) );
  AOI21_X1 U13982 ( .B1(n10659), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11078), .ZN(
        n11079) );
  OAI21_X1 U13983 ( .B1(n11080), .B2(n11151), .A(n11079), .ZN(n11083) );
  XNOR2_X1 U13984 ( .A(n11101), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16102) );
  NAND2_X1 U13985 ( .A1(n16102), .A2(n11081), .ZN(n11082) );
  NAND2_X1 U13986 ( .A1(n11083), .A2(n11082), .ZN(n15497) );
  AOI22_X1 U13987 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10392), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U13988 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11156), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U13989 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U13990 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11084) );
  NAND4_X1 U13991 ( .A1(n11087), .A2(n11086), .A3(n11085), .A4(n11084), .ZN(
        n11094) );
  AOI22_X1 U13992 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11088), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U13993 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10533), .B1(
        n10452), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U13994 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U13995 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9815), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11089) );
  NAND4_X1 U13996 ( .A1(n11092), .A2(n11091), .A3(n11090), .A4(n11089), .ZN(
        n11093) );
  NOR2_X1 U13997 ( .A1(n11094), .A2(n11093), .ZN(n11111) );
  NAND2_X1 U13998 ( .A1(n11096), .A2(n11095), .ZN(n11110) );
  XNOR2_X1 U13999 ( .A(n11111), .B(n11110), .ZN(n11100) );
  NAND2_X1 U14000 ( .A1(n21441), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11097) );
  NAND2_X1 U14001 ( .A1(n11174), .A2(n11097), .ZN(n11098) );
  AOI21_X1 U14002 ( .B1(n10659), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11098), .ZN(
        n11099) );
  OAI21_X1 U14003 ( .B1(n11100), .B2(n11151), .A(n11099), .ZN(n11108) );
  INV_X1 U14004 ( .A(n11101), .ZN(n11102) );
  INV_X1 U14005 ( .A(n11103), .ZN(n11105) );
  INV_X1 U14006 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11104) );
  NAND2_X1 U14007 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  NAND2_X1 U14008 ( .A1(n11129), .A2(n11106), .ZN(n15768) );
  NAND2_X1 U14009 ( .A1(n11108), .A2(n11107), .ZN(n15483) );
  NOR2_X1 U14010 ( .A1(n11111), .A2(n11110), .ZN(n11148) );
  AOI22_X1 U14011 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9826), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11115) );
  AOI22_X1 U14012 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10452), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14013 ( .A1(n11164), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14014 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11112) );
  NAND4_X1 U14015 ( .A1(n11115), .A2(n11114), .A3(n11113), .A4(n11112), .ZN(
        n11121) );
  AOI22_X1 U14016 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14017 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9814), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14018 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14019 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11116) );
  NAND4_X1 U14020 ( .A1(n11119), .A2(n11118), .A3(n11117), .A4(n11116), .ZN(
        n11120) );
  OR2_X1 U14021 ( .A1(n11121), .A2(n11120), .ZN(n11147) );
  INV_X1 U14022 ( .A(n11147), .ZN(n11122) );
  XNOR2_X1 U14023 ( .A(n11148), .B(n11122), .ZN(n11123) );
  NAND2_X1 U14024 ( .A1(n11123), .A2(n11177), .ZN(n11128) );
  NAND2_X1 U14025 ( .A1(n21441), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14026 ( .A1(n11174), .A2(n11124), .ZN(n11125) );
  AOI21_X1 U14027 ( .B1(n10659), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11125), .ZN(
        n11127) );
  XNOR2_X1 U14028 ( .A(n11129), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15761) );
  AOI21_X1 U14029 ( .B1(n11128), .B2(n11127), .A(n11126), .ZN(n15472) );
  INV_X1 U14030 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15758) );
  NAND2_X1 U14031 ( .A1(n11130), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15106) );
  INV_X1 U14032 ( .A(n11130), .ZN(n11132) );
  INV_X1 U14033 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11131) );
  NAND2_X1 U14034 ( .A1(n11132), .A2(n11131), .ZN(n11133) );
  NAND2_X1 U14035 ( .A1(n15106), .A2(n11133), .ZN(n15746) );
  AOI22_X1 U14036 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11156), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14037 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11158), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11138) );
  AOI22_X1 U14038 ( .A1(n11134), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U14039 ( .A1(n9814), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11136) );
  NAND4_X1 U14040 ( .A1(n11139), .A2(n11138), .A3(n11137), .A4(n11136), .ZN(
        n11146) );
  AOI22_X1 U14041 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14042 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14043 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U14044 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11141) );
  NAND4_X1 U14045 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .ZN(
        n11145) );
  NOR2_X1 U14046 ( .A1(n11146), .A2(n11145), .ZN(n11155) );
  NAND2_X1 U14047 ( .A1(n11148), .A2(n11147), .ZN(n11154) );
  XNOR2_X1 U14048 ( .A(n11155), .B(n11154), .ZN(n11152) );
  AOI21_X1 U14049 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21441), .A(
        n10631), .ZN(n11150) );
  NAND2_X1 U14050 ( .A1(n10753), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11149) );
  OAI211_X1 U14051 ( .C1(n11152), .C2(n11151), .A(n11150), .B(n11149), .ZN(
        n11153) );
  XNOR2_X1 U14052 ( .A(n15106), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15453) );
  NOR2_X1 U14053 ( .A1(n11155), .A2(n11154), .ZN(n11173) );
  AOI22_X1 U14054 ( .A1(n11156), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14055 ( .A1(n11088), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10476), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11161) );
  AOI22_X1 U14056 ( .A1(n11157), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11134), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11160) );
  AOI22_X1 U14057 ( .A1(n11158), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10471), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11159) );
  NAND4_X1 U14058 ( .A1(n11162), .A2(n11161), .A3(n11160), .A4(n11159), .ZN(
        n11171) );
  AOI22_X1 U14059 ( .A1(n11163), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10444), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U14060 ( .A1(n9826), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11164), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11168) );
  AOI22_X1 U14061 ( .A1(n10709), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9815), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14062 ( .A1(n11165), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10534), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11166) );
  NAND4_X1 U14063 ( .A1(n11169), .A2(n11168), .A3(n11167), .A4(n11166), .ZN(
        n11170) );
  NOR2_X1 U14064 ( .A1(n11171), .A2(n11170), .ZN(n11172) );
  XNOR2_X1 U14065 ( .A(n11173), .B(n11172), .ZN(n11178) );
  INV_X1 U14066 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15105) );
  NAND2_X1 U14067 ( .A1(n10659), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11175) );
  OAI211_X1 U14068 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n15105), .A(n11175), 
        .B(n11174), .ZN(n11176) );
  AOI21_X1 U14069 ( .B1(n11178), .B2(n11177), .A(n11176), .ZN(n11179) );
  AOI21_X1 U14070 ( .B1(n11081), .B2(n15453), .A(n11179), .ZN(n15419) );
  NAND3_X1 U14071 ( .A1(n21439), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17394) );
  NAND2_X1 U14072 ( .A1(n17400), .A2(n21441), .ZN(n16334) );
  NAND2_X1 U14073 ( .A1(n17165), .A2(n10487), .ZN(n11218) );
  NOR2_X1 U14074 ( .A1(n11180), .A2(n11218), .ZN(n11181) );
  AND2_X4 U14075 ( .A1(n11244), .A2(n11181), .ZN(n16288) );
  AOI21_X1 U14076 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16288), .ZN(n15345) );
  NOR2_X1 U14077 ( .A1(n16288), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17289) );
  NAND2_X1 U14078 ( .A1(n16288), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16158) );
  OAI21_X1 U14079 ( .B1(n16288), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16158), .ZN(n17290) );
  NOR3_X1 U14080 ( .A1(n15345), .A2(n17289), .A3(n17290), .ZN(n16157) );
  OR2_X1 U14081 ( .A1(n16288), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11182) );
  NAND2_X1 U14082 ( .A1(n16157), .A2(n11182), .ZN(n16285) );
  NAND2_X1 U14083 ( .A1(n16288), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11183) );
  NAND2_X1 U14084 ( .A1(n16158), .A2(n11183), .ZN(n11275) );
  AND2_X1 U14085 ( .A1(n16288), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11184) );
  NOR2_X1 U14086 ( .A1(n11275), .A2(n11184), .ZN(n16274) );
  NAND2_X1 U14087 ( .A1(n16285), .A2(n16274), .ZN(n11186) );
  INV_X1 U14088 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16296) );
  MUX2_X1 U14089 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n16296), .S(
        n16288), .Z(n16291) );
  OR2_X1 U14090 ( .A1(n16288), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11185) );
  NAND2_X1 U14091 ( .A1(n11186), .A2(n16289), .ZN(n16272) );
  NAND2_X1 U14092 ( .A1(n11187), .A2(n11310), .ZN(n11192) );
  INV_X1 U14093 ( .A(n21543), .ZN(n11259) );
  XNOR2_X1 U14094 ( .A(n11188), .B(n11205), .ZN(n11190) );
  AOI21_X1 U14095 ( .B1(n11259), .B2(n11190), .A(n11189), .ZN(n11191) );
  NAND2_X1 U14096 ( .A1(n11192), .A2(n11191), .ZN(n11197) );
  NAND2_X1 U14097 ( .A1(n12789), .A2(n14069), .ZN(n11208) );
  OAI21_X1 U14098 ( .B1(n21543), .B2(n11206), .A(n11208), .ZN(n11194) );
  INV_X1 U14099 ( .A(n11194), .ZN(n11195) );
  NAND2_X1 U14100 ( .A1(n14134), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11200) );
  INV_X1 U14101 ( .A(n11197), .ZN(n11198) );
  NAND2_X1 U14102 ( .A1(n11200), .A2(n11199), .ZN(n11213) );
  INV_X1 U14103 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11201) );
  OR2_X1 U14104 ( .A1(n14028), .A2(n11218), .ZN(n11212) );
  INV_X1 U14105 ( .A(n11204), .ZN(n11203) );
  NAND2_X1 U14106 ( .A1(n11205), .A2(n11206), .ZN(n11202) );
  NAND2_X1 U14107 ( .A1(n11203), .A2(n11202), .ZN(n11223) );
  NAND3_X1 U14108 ( .A1(n11206), .A2(n11205), .A3(n11204), .ZN(n11207) );
  NAND2_X1 U14109 ( .A1(n11223), .A2(n11207), .ZN(n11210) );
  INV_X1 U14110 ( .A(n11208), .ZN(n11209) );
  AOI21_X1 U14111 ( .B1(n11210), .B2(n11259), .A(n11209), .ZN(n11211) );
  NAND2_X1 U14112 ( .A1(n11213), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11214) );
  INV_X1 U14113 ( .A(n11224), .ZN(n11215) );
  XNOR2_X1 U14114 ( .A(n11223), .B(n11215), .ZN(n11216) );
  NAND2_X1 U14115 ( .A1(n11216), .A2(n11259), .ZN(n11217) );
  INV_X1 U14116 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14368) );
  NAND2_X1 U14117 ( .A1(n11219), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11220) );
  NAND2_X1 U14118 ( .A1(n11221), .A2(n11220), .ZN(n14366) );
  NAND2_X1 U14119 ( .A1(n11222), .A2(n11310), .ZN(n11227) );
  NAND2_X1 U14120 ( .A1(n11224), .A2(n11223), .ZN(n11233) );
  XNOR2_X1 U14121 ( .A(n11232), .B(n11233), .ZN(n11225) );
  NAND2_X1 U14122 ( .A1(n11259), .A2(n11225), .ZN(n11226) );
  NAND2_X1 U14123 ( .A1(n11227), .A2(n11226), .ZN(n11228) );
  INV_X1 U14124 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14369) );
  XNOR2_X1 U14125 ( .A(n11228), .B(n14369), .ZN(n14367) );
  NAND2_X1 U14126 ( .A1(n14366), .A2(n14367), .ZN(n11230) );
  NAND2_X1 U14127 ( .A1(n11228), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11229) );
  NAND2_X1 U14128 ( .A1(n11230), .A2(n11229), .ZN(n14612) );
  NAND2_X1 U14129 ( .A1(n11231), .A2(n11310), .ZN(n11238) );
  INV_X1 U14130 ( .A(n11232), .ZN(n11234) );
  NOR2_X1 U14131 ( .A1(n11234), .A2(n11233), .ZN(n11246) );
  INV_X1 U14132 ( .A(n11246), .ZN(n11235) );
  XNOR2_X1 U14133 ( .A(n11245), .B(n11235), .ZN(n11236) );
  NAND2_X1 U14134 ( .A1(n11259), .A2(n11236), .ZN(n11237) );
  NAND2_X1 U14135 ( .A1(n11238), .A2(n11237), .ZN(n11240) );
  INV_X1 U14136 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11239) );
  XNOR2_X1 U14137 ( .A(n11240), .B(n11239), .ZN(n14613) );
  NAND2_X1 U14138 ( .A1(n14612), .A2(n14613), .ZN(n11242) );
  NAND2_X1 U14139 ( .A1(n11240), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11241) );
  NAND2_X1 U14140 ( .A1(n11242), .A2(n11241), .ZN(n14973) );
  NAND3_X1 U14141 ( .A1(n11244), .A2(n11243), .A3(n11310), .ZN(n11249) );
  NAND2_X1 U14142 ( .A1(n11246), .A2(n11245), .ZN(n11255) );
  XNOR2_X1 U14143 ( .A(n11254), .B(n11255), .ZN(n11247) );
  NAND2_X1 U14144 ( .A1(n11259), .A2(n11247), .ZN(n11248) );
  NAND2_X1 U14145 ( .A1(n11249), .A2(n11248), .ZN(n11250) );
  INV_X1 U14146 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14982) );
  XNOR2_X1 U14147 ( .A(n11250), .B(n14982), .ZN(n14974) );
  NAND2_X1 U14148 ( .A1(n14973), .A2(n14974), .ZN(n11252) );
  NAND2_X1 U14149 ( .A1(n11250), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11251) );
  NAND2_X1 U14150 ( .A1(n11252), .A2(n11251), .ZN(n14960) );
  NAND2_X1 U14151 ( .A1(n11253), .A2(n11310), .ZN(n11261) );
  INV_X1 U14152 ( .A(n11254), .ZN(n11256) );
  NOR2_X1 U14153 ( .A1(n11256), .A2(n11255), .ZN(n11265) );
  INV_X1 U14154 ( .A(n11265), .ZN(n11257) );
  XNOR2_X1 U14155 ( .A(n11266), .B(n11257), .ZN(n11258) );
  NAND2_X1 U14156 ( .A1(n11259), .A2(n11258), .ZN(n11260) );
  NAND2_X1 U14157 ( .A1(n11261), .A2(n11260), .ZN(n11262) );
  INV_X1 U14158 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15137) );
  XNOR2_X1 U14159 ( .A(n11262), .B(n15137), .ZN(n14961) );
  NAND2_X1 U14160 ( .A1(n14960), .A2(n14961), .ZN(n11264) );
  NAND2_X1 U14161 ( .A1(n11262), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11263) );
  NAND2_X1 U14162 ( .A1(n11266), .A2(n11265), .ZN(n11267) );
  NOR2_X1 U14163 ( .A1(n21543), .A2(n11267), .ZN(n11268) );
  INV_X1 U14164 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15138) );
  XNOR2_X1 U14165 ( .A(n11269), .B(n15138), .ZN(n15123) );
  NAND2_X1 U14166 ( .A1(n11269), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11270) );
  NOR3_X1 U14167 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11271) );
  INV_X1 U14168 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11273) );
  INV_X1 U14169 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11272) );
  INV_X1 U14170 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15356) );
  NAND3_X1 U14171 ( .A1(n11273), .A2(n11272), .A3(n15356), .ZN(n11274) );
  AND2_X1 U14172 ( .A1(n16288), .A2(n11274), .ZN(n16155) );
  NOR2_X1 U14173 ( .A1(n11275), .A2(n16155), .ZN(n16286) );
  INV_X1 U14174 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16007) );
  NAND2_X1 U14175 ( .A1(n16288), .A2(n16007), .ZN(n16138) );
  OR2_X1 U14176 ( .A1(n16288), .A2(n16007), .ZN(n11279) );
  NAND2_X1 U14177 ( .A1(n16138), .A2(n11279), .ZN(n16149) );
  INV_X1 U14178 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16253) );
  AND2_X1 U14179 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16229) );
  INV_X1 U14180 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16228) );
  NOR2_X1 U14181 ( .A1(n11280), .A2(n16288), .ZN(n16098) );
  INV_X1 U14182 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15754) );
  INV_X1 U14183 ( .A(n11280), .ZN(n11284) );
  INV_X1 U14184 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11282) );
  INV_X1 U14185 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16235) );
  NAND4_X1 U14186 ( .A1(n16007), .A2(n11282), .A3(n16253), .A4(n16235), .ZN(
        n11283) );
  OAI21_X1 U14187 ( .B1(n11281), .B2(n11283), .A(n16288), .ZN(n16212) );
  AND2_X1 U14188 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16110) );
  NAND2_X1 U14189 ( .A1(n16110), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16096) );
  NOR2_X1 U14190 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16111) );
  INV_X1 U14191 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16197) );
  AND2_X1 U14192 ( .A1(n16111), .A2(n16197), .ZN(n15751) );
  INV_X1 U14193 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16191) );
  INV_X1 U14194 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11286) );
  AND2_X1 U14195 ( .A1(n16191), .A2(n11286), .ZN(n11287) );
  INV_X1 U14196 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17319) );
  NAND2_X1 U14197 ( .A1(n16288), .A2(n17319), .ZN(n15741) );
  NAND2_X1 U14198 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17325) );
  INV_X1 U14199 ( .A(n17325), .ZN(n11288) );
  OR2_X1 U14200 ( .A1(n16288), .A2(n17319), .ZN(n15742) );
  INV_X1 U14201 ( .A(n15742), .ZN(n11289) );
  NAND2_X1 U14202 ( .A1(n12628), .A2(n11289), .ZN(n11290) );
  NAND2_X1 U14203 ( .A1(n11291), .A2(n11290), .ZN(n11292) );
  INV_X1 U14204 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16179) );
  XNOR2_X1 U14205 ( .A(n11292), .B(n16179), .ZN(n16177) );
  XNOR2_X1 U14206 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11301) );
  NAND2_X1 U14207 ( .A1(n11301), .A2(n11300), .ZN(n11304) );
  NAND2_X1 U14208 ( .A1(n17132), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11293) );
  NAND2_X1 U14209 ( .A1(n11304), .A2(n11293), .ZN(n11297) );
  XNOR2_X1 U14210 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11298) );
  NAND2_X1 U14211 ( .A1(n11297), .A2(n11298), .ZN(n11295) );
  NAND2_X1 U14212 ( .A1(n17138), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11294) );
  XNOR2_X1 U14213 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11318) );
  NOR2_X1 U14214 ( .A1(n10369), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11296) );
  NOR2_X1 U14215 ( .A1(n21437), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11331) );
  AND2_X1 U14216 ( .A1(n11330), .A2(n11331), .ZN(n11327) );
  XOR2_X1 U14217 ( .A(n11298), .B(n11297), .Z(n12640) );
  NAND2_X1 U14218 ( .A1(n13984), .A2(n10487), .ZN(n11308) );
  NAND2_X1 U14219 ( .A1(n12662), .A2(n11308), .ZN(n11320) );
  NOR2_X1 U14220 ( .A1(n10487), .A2(n21439), .ZN(n11299) );
  NOR2_X1 U14221 ( .A1(n11338), .A2(n11299), .ZN(n11306) );
  NAND2_X1 U14222 ( .A1(n11306), .A2(n17165), .ZN(n11322) );
  INV_X1 U14223 ( .A(n11300), .ZN(n11303) );
  INV_X1 U14224 ( .A(n11301), .ZN(n11302) );
  NAND2_X1 U14225 ( .A1(n11303), .A2(n11302), .ZN(n11305) );
  AND2_X1 U14226 ( .A1(n11305), .A2(n11304), .ZN(n12638) );
  INV_X1 U14227 ( .A(n12638), .ZN(n11307) );
  XNOR2_X1 U14228 ( .A(n17127), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11312) );
  INV_X1 U14229 ( .A(n11312), .ZN(n11309) );
  OAI21_X1 U14230 ( .B1(n12779), .B2(n12789), .A(n11309), .ZN(n11315) );
  INV_X1 U14231 ( .A(n11338), .ZN(n11313) );
  OAI21_X1 U14232 ( .B1(n11313), .B2(n11312), .A(n11334), .ZN(n11314) );
  OAI21_X1 U14233 ( .B1(n11320), .B2(n11315), .A(n11314), .ZN(n11316) );
  XOR2_X1 U14234 ( .A(n11318), .B(n11317), .Z(n12639) );
  OAI21_X1 U14235 ( .B1(n11320), .B2(n11319), .A(n12639), .ZN(n11321) );
  OAI21_X1 U14236 ( .B1(n11326), .B2(n12640), .A(n11321), .ZN(n11324) );
  INV_X1 U14237 ( .A(n11327), .ZN(n12644) );
  OAI22_X1 U14238 ( .A1(n11322), .A2(n12644), .B1(n12639), .B2(n11334), .ZN(
        n11323) );
  AOI21_X1 U14239 ( .B1(n9879), .B2(n11324), .A(n11323), .ZN(n11325) );
  AOI21_X1 U14240 ( .B1(n11327), .B2(n11326), .A(n11325), .ZN(n11328) );
  AOI21_X1 U14241 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21439), .A(
        n11328), .ZN(n11336) );
  NAND2_X1 U14242 ( .A1(n21437), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11329) );
  NAND2_X1 U14243 ( .A1(n11330), .A2(n11329), .ZN(n11333) );
  INV_X1 U14244 ( .A(n11331), .ZN(n11332) );
  NOR2_X1 U14245 ( .A1(n11334), .A2(n12642), .ZN(n11335) );
  INV_X1 U14246 ( .A(n12642), .ZN(n11337) );
  NAND2_X1 U14247 ( .A1(n11338), .A2(n11337), .ZN(n11339) );
  AND2_X1 U14248 ( .A1(n11341), .A2(n11340), .ZN(n11343) );
  NAND2_X1 U14249 ( .A1(n13910), .A2(n12789), .ZN(n11342) );
  NAND2_X1 U14250 ( .A1(n11343), .A2(n11342), .ZN(n12653) );
  OR2_X1 U14251 ( .A1(n12653), .A2(n12779), .ZN(n17150) );
  NOR2_X1 U14252 ( .A1(n17150), .A2(n21248), .ZN(n11344) );
  INV_X1 U14253 ( .A(n17312), .ZN(n17267) );
  NAND2_X1 U14254 ( .A1(n16177), .A2(n17267), .ZN(n11351) );
  NAND2_X1 U14255 ( .A1(n11347), .A2(n16334), .ZN(n21537) );
  NAND2_X1 U14256 ( .A1(n21537), .A2(n21439), .ZN(n11345) );
  NAND2_X1 U14257 ( .A1(n21439), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17168) );
  INV_X1 U14258 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21254) );
  NAND2_X1 U14259 ( .A1(n21254), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11346) );
  NAND2_X1 U14260 ( .A1(n17168), .A2(n11346), .ZN(n14162) );
  NAND2_X1 U14261 ( .A1(n17296), .A2(n15453), .ZN(n11348) );
  NAND2_X1 U14262 ( .A1(n17369), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16180) );
  OAI211_X1 U14263 ( .C1(n15105), .C2(n15759), .A(n11348), .B(n16180), .ZN(
        n11349) );
  INV_X1 U14264 ( .A(n11349), .ZN(n11350) );
  OAI211_X1 U14265 ( .C1(n15649), .C2(n17306), .A(n11351), .B(n11350), .ZN(
        P1_U2969) );
  AND2_X4 U14266 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16936) );
  INV_X2 U14267 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16927) );
  NAND2_X1 U14268 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11353) );
  AND2_X1 U14269 ( .A1(n11353), .A2(n11352), .ZN(n11359) );
  INV_X1 U14270 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11354) );
  AND2_X4 U14271 ( .A1(n11600), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13037) );
  AOI22_X1 U14272 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11358) );
  AND2_X4 U14273 ( .A1(n15190), .A2(n17686), .ZN(n11606) );
  AOI22_X1 U14274 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14275 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11356) );
  NAND4_X1 U14276 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11360) );
  NAND2_X1 U14277 ( .A1(n11360), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11367) );
  AOI22_X1 U14278 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14279 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14280 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11361) );
  NAND4_X1 U14281 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11365) );
  NAND2_X1 U14282 ( .A1(n11365), .A2(n17691), .ZN(n11366) );
  AOI22_X1 U14283 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11455), .B1(
        n13042), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14284 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14285 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14286 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11368) );
  NAND4_X1 U14287 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11372) );
  NAND2_X1 U14288 ( .A1(n11372), .A2(n17691), .ZN(n11379) );
  AOI22_X1 U14289 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14290 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14291 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14292 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9820), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11373) );
  NAND4_X1 U14293 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11377) );
  NAND2_X1 U14294 ( .A1(n11377), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11378) );
  AOI22_X1 U14295 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14296 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14297 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14298 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11385) );
  NAND3_X1 U14299 ( .A1(n11387), .A2(n11386), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11388) );
  NOR2_X1 U14300 ( .A1(n11389), .A2(n11388), .ZN(n11392) );
  AOI22_X1 U14301 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14302 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11390) );
  NAND3_X1 U14303 ( .A1(n11392), .A2(n11391), .A3(n11390), .ZN(n11393) );
  NAND2_X2 U14304 ( .A1(n11394), .A2(n11393), .ZN(n11481) );
  AOI22_X1 U14305 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14306 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14307 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9820), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11396) );
  NAND4_X1 U14308 ( .A1(n11398), .A2(n11397), .A3(n11396), .A4(n11395), .ZN(
        n11399) );
  NAND2_X1 U14309 ( .A1(n11399), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11406) );
  AOI22_X1 U14310 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14311 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14312 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14313 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11400) );
  NAND4_X1 U14314 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(
        n11404) );
  NAND2_X1 U14315 ( .A1(n11404), .A2(n17691), .ZN(n11405) );
  NAND2_X2 U14316 ( .A1(n11406), .A2(n11405), .ZN(n12242) );
  AOI22_X1 U14317 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14318 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14319 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14320 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11407) );
  NAND4_X1 U14321 ( .A1(n11410), .A2(n11409), .A3(n11408), .A4(n11407), .ZN(
        n11411) );
  NAND2_X1 U14322 ( .A1(n11411), .A2(n17691), .ZN(n11418) );
  AOI22_X1 U14323 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14324 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14325 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11413) );
  NAND4_X1 U14326 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(
        n11416) );
  NAND2_X1 U14327 ( .A1(n11416), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11417) );
  AOI22_X1 U14328 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14329 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14330 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U14331 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11419) );
  NAND4_X1 U14332 ( .A1(n11422), .A2(n11421), .A3(n11420), .A4(n11419), .ZN(
        n11423) );
  AOI22_X1 U14333 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14334 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14335 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14336 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11424) );
  NAND4_X1 U14337 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(
        n11428) );
  AOI22_X1 U14338 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9822), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14339 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14340 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U14341 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n11443) );
  AOI22_X1 U14342 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14343 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11607), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11437) );
  NOR2_X1 U14344 ( .A1(n11496), .A2(n17714), .ZN(n11449) );
  OAI21_X1 U14345 ( .B1(n12215), .B2(n20573), .A(n11445), .ZN(n11447) );
  AND2_X1 U14346 ( .A1(n12210), .A2(n11482), .ZN(n11446) );
  OAI211_X1 U14347 ( .C1(n12272), .C2(n11481), .A(n11447), .B(n11446), .ZN(
        n11448) );
  NAND2_X1 U14348 ( .A1(n11449), .A2(n11448), .ZN(n12250) );
  AOI22_X1 U14349 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11450) );
  AND2_X1 U14350 ( .A1(n11450), .A2(n17691), .ZN(n11454) );
  AOI22_X1 U14351 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9820), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14352 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14353 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11451) );
  NAND4_X1 U14354 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(
        n11462) );
  AOI22_X1 U14355 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11455), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14356 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9820), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11456) );
  AND3_X1 U14357 ( .A1(n11457), .A2(n11456), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14358 ( .A1(n11606), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13038), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14359 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11458) );
  NAND3_X1 U14360 ( .A1(n11460), .A2(n11459), .A3(n11458), .ZN(n11461) );
  AND2_X1 U14361 ( .A1(n11467), .A2(n11612), .ZN(n12245) );
  INV_X2 U14362 ( .A(n11471), .ZN(n20573) );
  NAND2_X1 U14363 ( .A1(n12245), .A2(n11502), .ZN(n11521) );
  NAND2_X1 U14364 ( .A1(n11521), .A2(n11463), .ZN(n11464) );
  NAND2_X1 U14365 ( .A1(n12250), .A2(n11464), .ZN(n11520) );
  NAND2_X1 U14366 ( .A1(n11520), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11479) );
  NAND2_X1 U14368 ( .A1(n11466), .A2(n12211), .ZN(n12221) );
  NAND2_X1 U14369 ( .A1(n11467), .A2(n11472), .ZN(n12208) );
  NAND2_X1 U14370 ( .A1(n12221), .A2(n11468), .ZN(n12251) );
  NAND2_X1 U14371 ( .A1(n12251), .A2(n12253), .ZN(n11470) );
  NAND2_X1 U14372 ( .A1(n11470), .A2(n11469), .ZN(n11522) );
  NAND2_X1 U14373 ( .A1(n11522), .A2(n9856), .ZN(n11478) );
  NOR2_X1 U14374 ( .A1(n12242), .A2(n11472), .ZN(n11473) );
  AND2_X2 U14375 ( .A1(n12216), .A2(n11473), .ZN(n11476) );
  INV_X1 U14376 ( .A(n12210), .ZN(n11474) );
  NAND2_X1 U14377 ( .A1(n12019), .A2(n11475), .ZN(n11477) );
  INV_X1 U14378 ( .A(n12211), .ZN(n11489) );
  NAND2_X2 U14379 ( .A1(n11476), .A2(n11489), .ZN(n11493) );
  AND2_X2 U14380 ( .A1(n11477), .A2(n11493), .ZN(n12487) );
  NAND2_X1 U14381 ( .A1(n12487), .A2(n21227), .ZN(n11523) );
  NAND2_X1 U14382 ( .A1(n11517), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11487) );
  INV_X1 U14383 ( .A(n11493), .ZN(n11480) );
  NAND2_X1 U14384 ( .A1(n11480), .A2(n17714), .ZN(n12847) );
  NAND2_X1 U14385 ( .A1(n11496), .A2(n11463), .ZN(n15199) );
  NOR2_X1 U14386 ( .A1(n11624), .A2(n12240), .ZN(n11483) );
  NAND3_X1 U14387 ( .A1(n11498), .A2(n11463), .A3(n13778), .ZN(n11484) );
  NOR2_X1 U14388 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12135) );
  AND2_X2 U14389 ( .A1(n11487), .A2(n11486), .ZN(n11510) );
  INV_X1 U14390 ( .A(n11510), .ZN(n11508) );
  NAND2_X1 U14391 ( .A1(n11489), .A2(n11488), .ZN(n11491) );
  NAND2_X1 U14392 ( .A1(n11612), .A2(n11463), .ZN(n12239) );
  NAND2_X2 U14393 ( .A1(n11789), .A2(n12239), .ZN(n13681) );
  NAND3_X1 U14394 ( .A1(n12246), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11512), 
        .ZN(n11501) );
  INV_X1 U14395 ( .A(n11493), .ZN(n12206) );
  NAND3_X1 U14396 ( .A1(n12206), .A2(n11612), .A3(n21227), .ZN(n11500) );
  NOR2_X1 U14397 ( .A1(n21228), .A2(n11494), .ZN(n11497) );
  NOR2_X1 U14398 ( .A1(n21228), .A2(n11624), .ZN(n11495) );
  NAND2_X1 U14399 ( .A1(n11546), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11504) );
  NAND2_X1 U14400 ( .A1(n11505), .A2(n11504), .ZN(n11506) );
  INV_X1 U14401 ( .A(n11509), .ZN(n11507) );
  INV_X1 U14402 ( .A(n11512), .ZN(n11513) );
  NOR2_X2 U14403 ( .A1(n11514), .A2(n11513), .ZN(n15189) );
  INV_X1 U14404 ( .A(n12234), .ZN(n11516) );
  INV_X1 U14405 ( .A(n12135), .ZN(n11525) );
  NOR2_X1 U14406 ( .A1(n11525), .A2(n21212), .ZN(n11515) );
  NAND2_X1 U14407 ( .A1(n11517), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11518) );
  NAND2_X1 U14408 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14409 ( .A1(n11525), .A2(n11524), .ZN(n11526) );
  AOI21_X1 U14410 ( .B1(n11535), .B2(P2_EBX_REG_0__SCAN_IN), .A(n11526), .ZN(
        n11528) );
  NAND2_X1 U14411 ( .A1(n11546), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11527) );
  NAND2_X1 U14412 ( .A1(n11534), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11529) );
  NAND2_X1 U14413 ( .A1(n11517), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11533) );
  AOI21_X1 U14414 ( .B1(n17682), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11532) );
  INV_X2 U14415 ( .A(n12042), .ZN(n12092) );
  NAND2_X1 U14416 ( .A1(n11546), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11536) );
  NAND2_X1 U14417 ( .A1(n11537), .A2(n11536), .ZN(n11538) );
  INV_X1 U14418 ( .A(n11539), .ZN(n11541) );
  NAND2_X1 U14419 ( .A1(n11541), .A2(n11540), .ZN(n11542) );
  NAND2_X1 U14420 ( .A1(n11517), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11545) );
  NAND2_X1 U14421 ( .A1(n12135), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11544) );
  AOI22_X1 U14422 ( .A1(n11535), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11548) );
  NAND2_X1 U14423 ( .A1(n12074), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U14424 ( .A1(n11548), .A2(n11547), .ZN(n11549) );
  INV_X1 U14425 ( .A(n9799), .ZN(n11553) );
  INV_X1 U14426 ( .A(n11551), .ZN(n11552) );
  NAND2_X1 U14427 ( .A1(n11553), .A2(n11552), .ZN(n11560) );
  INV_X1 U14428 ( .A(n11556), .ZN(n11557) );
  NAND2_X1 U14429 ( .A1(n20973), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11573) );
  AND2_X1 U14430 ( .A1(n11558), .A2(n12916), .ZN(n11564) );
  INV_X1 U14431 ( .A(n11560), .ZN(n11561) );
  NOR2_X1 U14432 ( .A1(n11559), .A2(n11561), .ZN(n11566) );
  AOI22_X1 U14433 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20807), .B1(
        n21017), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11572) );
  INV_X1 U14434 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12982) );
  INV_X1 U14435 ( .A(n11564), .ZN(n11562) );
  INV_X1 U14436 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11563) );
  OAI22_X1 U14437 ( .A1(n12982), .A2(n14014), .B1(n20587), .B2(n11563), .ZN(
        n11570) );
  INV_X1 U14438 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U14439 ( .A1(n16946), .A2(n11564), .ZN(n11565) );
  INV_X1 U14440 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11567) );
  NOR2_X1 U14441 ( .A1(n11570), .A2(n11569), .ZN(n11571) );
  AND3_X1 U14442 ( .A1(n11573), .A2(n11572), .A3(n11571), .ZN(n11595) );
  INV_X1 U14443 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11576) );
  OR2_X1 U14444 ( .A1(n16946), .A2(n9818), .ZN(n11582) );
  OR2_X2 U14445 ( .A1(n11582), .A2(n11574), .ZN(n11716) );
  OR2_X2 U14446 ( .A1(n11585), .A2(n11574), .ZN(n20842) );
  INV_X1 U14447 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11575) );
  AOI21_X1 U14448 ( .B1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n11723), .A(
        n11577), .ZN(n11594) );
  INV_X1 U14449 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12378) );
  INV_X1 U14450 ( .A(n11578), .ZN(n11579) );
  NAND2_X1 U14451 ( .A1(n11579), .A2(n16918), .ZN(n11728) );
  INV_X1 U14452 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11580) );
  INV_X1 U14453 ( .A(n11581), .ZN(n11593) );
  INV_X1 U14454 ( .A(n11586), .ZN(n11584) );
  INV_X1 U14455 ( .A(n11582), .ZN(n11583) );
  INV_X1 U14456 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12899) );
  NAND2_X1 U14457 ( .A1(n11835), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11587) );
  OAI21_X1 U14458 ( .B1(n16972), .B2(n12899), .A(n11587), .ZN(n11591) );
  INV_X1 U14459 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11589) );
  INV_X1 U14460 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11588) );
  OAI22_X1 U14461 ( .A1(n11589), .A2(n11705), .B1(n20865), .B2(n11588), .ZN(
        n11590) );
  NOR2_X1 U14462 ( .A1(n11591), .A2(n11590), .ZN(n11592) );
  NAND4_X1 U14463 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11614) );
  AND2_X2 U14464 ( .A1(n13203), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11736) );
  AND2_X2 U14465 ( .A1(n13038), .A2(n17691), .ZN(n11767) );
  AOI22_X1 U14466 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11736), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11599) );
  AND2_X2 U14467 ( .A1(n13037), .A2(n17691), .ZN(n13018) );
  AND2_X2 U14468 ( .A1(n9823), .A2(n17691), .ZN(n12322) );
  AOI22_X1 U14469 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12322), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11598) );
  AND2_X2 U14470 ( .A1(n9823), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12321) );
  AND2_X2 U14471 ( .A1(n9811), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11753) );
  AOI22_X1 U14472 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n12321), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14473 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11596) );
  NAND4_X1 U14474 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n11611) );
  NAND2_X1 U14475 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13043) );
  INV_X1 U14476 ( .A(n13043), .ZN(n11601) );
  NAND3_X1 U14477 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12011) );
  INV_X1 U14478 ( .A(n12011), .ZN(n11602) );
  AOI22_X1 U14479 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n13063), .ZN(n11605) );
  NAND2_X1 U14480 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11604) );
  AND2_X2 U14481 ( .A1(n9819), .A2(n17691), .ZN(n13069) );
  NAND2_X1 U14482 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11603) );
  AND2_X2 U14483 ( .A1(n13203), .A2(n17691), .ZN(n11855) );
  AOI22_X1 U14484 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .B2(n11856), .ZN(n11609) );
  AOI22_X1 U14485 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12329), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11608) );
  NAND3_X1 U14486 ( .A1(n10344), .A2(n11609), .A3(n11608), .ZN(n11610) );
  NOR2_X1 U14487 ( .A1(n11611), .A2(n11610), .ZN(n12296) );
  NAND2_X1 U14488 ( .A1(n12296), .A2(n20547), .ZN(n11613) );
  INV_X1 U14489 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11615) );
  NOR2_X1 U14490 ( .A1(n20865), .A2(n11615), .ZN(n11618) );
  INV_X1 U14491 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11616) );
  INV_X1 U14492 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12954) );
  INV_X1 U14493 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11619) );
  OAI22_X1 U14494 ( .A1(n14014), .A2(n12954), .B1(n11619), .B2(n14648), .ZN(
        n11620) );
  INV_X1 U14495 ( .A(n11620), .ZN(n11622) );
  INV_X1 U14496 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11621) );
  NAND3_X1 U14497 ( .A1(n11623), .A2(n11622), .A3(n10343), .ZN(n11631) );
  INV_X1 U14498 ( .A(n11625), .ZN(n11629) );
  NAND2_X1 U14499 ( .A1(n11834), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11628) );
  INV_X1 U14500 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15963) );
  NAND3_X1 U14501 ( .A1(n11629), .A2(n11628), .A3(n11627), .ZN(n11630) );
  NOR2_X1 U14502 ( .A1(n11631), .A2(n11630), .ZN(n11645) );
  INV_X1 U14503 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12919) );
  INV_X1 U14504 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11632) );
  OAI22_X1 U14505 ( .A1(n16972), .A2(n12919), .B1(n11718), .B2(n11632), .ZN(
        n11636) );
  INV_X1 U14506 ( .A(n11835), .ZN(n20617) );
  INV_X1 U14507 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11634) );
  INV_X1 U14508 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11633) );
  OAI22_X1 U14509 ( .A1(n20617), .A2(n11634), .B1(n20842), .B2(n11633), .ZN(
        n11635) );
  NOR2_X1 U14510 ( .A1(n11636), .A2(n11635), .ZN(n11644) );
  INV_X1 U14511 ( .A(n11704), .ZN(n11637) );
  INV_X1 U14512 ( .A(n11638), .ZN(n11727) );
  INV_X1 U14513 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11640) );
  INV_X1 U14514 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11639) );
  INV_X1 U14515 ( .A(n11641), .ZN(n11642) );
  NAND4_X1 U14516 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11689) );
  AOI22_X1 U14517 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14518 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11672), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14519 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14520 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11646) );
  NAND4_X1 U14521 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n11656) );
  AOI22_X1 U14522 ( .A1(n12322), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11650), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14523 ( .A1(n11767), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13069), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14524 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13063), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14525 ( .A1(n11753), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11651) );
  NAND4_X1 U14526 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11655) );
  AOI22_X1 U14527 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14528 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14529 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14530 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11657) );
  NAND4_X1 U14531 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n11670) );
  AOI22_X1 U14532 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n11856), .ZN(n11668) );
  INV_X1 U14533 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11663) );
  NAND2_X1 U14534 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11662) );
  NAND2_X1 U14535 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11661) );
  OAI211_X1 U14536 ( .C1(n13067), .C2(n11663), .A(n11662), .B(n11661), .ZN(
        n11664) );
  INV_X1 U14537 ( .A(n11664), .ZN(n11667) );
  AOI22_X1 U14538 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14539 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11665) );
  NAND4_X1 U14540 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11669) );
  INV_X1 U14541 ( .A(n12141), .ZN(n12285) );
  NOR2_X1 U14542 ( .A1(n12275), .A2(n12285), .ZN(n11671) );
  NAND2_X1 U14543 ( .A1(n20547), .A2(n11671), .ZN(n12145) );
  AOI22_X1 U14544 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14545 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12322), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14546 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14547 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11673) );
  NAND4_X1 U14548 ( .A1(n11676), .A2(n11675), .A3(n11674), .A4(n11673), .ZN(
        n11687) );
  AOI22_X1 U14549 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n11856), .ZN(n11685) );
  INV_X1 U14550 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11679) );
  NAND2_X1 U14551 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11678) );
  NAND2_X1 U14552 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11677) );
  OAI211_X1 U14553 ( .C1(n13029), .C2(n11679), .A(n11678), .B(n11677), .ZN(
        n11680) );
  INV_X1 U14554 ( .A(n11680), .ZN(n11684) );
  AOI22_X1 U14555 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12329), .B1(
        n12427), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11683) );
  NAND2_X1 U14556 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11682) );
  NAND4_X1 U14557 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11686) );
  NAND2_X1 U14558 ( .A1(n12145), .A2(n12289), .ZN(n11688) );
  AND2_X2 U14559 ( .A1(n11689), .A2(n11688), .ZN(n11803) );
  AOI22_X1 U14560 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11855), .B1(
        n12322), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14561 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14562 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12321), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14563 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11690) );
  NAND4_X1 U14564 ( .A1(n11693), .A2(n11692), .A3(n11691), .A4(n11690), .ZN(
        n11703) );
  AOI22_X1 U14565 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__4__SCAN_IN), .B2(n12427), .ZN(n11701) );
  INV_X1 U14566 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U14567 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11695) );
  NAND2_X1 U14568 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11694) );
  OAI211_X1 U14569 ( .C1(n13029), .C2(n11696), .A(n11695), .B(n11694), .ZN(
        n11697) );
  INV_X1 U14570 ( .A(n11697), .ZN(n11700) );
  AOI22_X1 U14571 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12329), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11699) );
  NAND2_X1 U14572 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11698) );
  NAND4_X1 U14573 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n11698), .ZN(
        n11702) );
  INV_X1 U14574 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12411) );
  INV_X1 U14575 ( .A(n11705), .ZN(n11706) );
  INV_X1 U14576 ( .A(n20865), .ZN(n20873) );
  AOI22_X1 U14577 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n11706), .B1(
        n20873), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11713) );
  INV_X1 U14578 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11708) );
  INV_X1 U14579 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11707) );
  OAI22_X1 U14580 ( .A1(n11708), .A2(n14014), .B1(n14648), .B2(n11707), .ZN(
        n11711) );
  INV_X1 U14581 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11743) );
  INV_X1 U14582 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11709) );
  NOR2_X1 U14583 ( .A1(n11711), .A2(n11710), .ZN(n11712) );
  OAI211_X1 U14584 ( .C1(n12411), .C2(n11704), .A(n11713), .B(n11712), .ZN(
        n11714) );
  INV_X1 U14585 ( .A(n11714), .ZN(n11735) );
  INV_X1 U14586 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13946) );
  INV_X1 U14587 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11715) );
  OAI22_X1 U14588 ( .A1(n16972), .A2(n13946), .B1(n11716), .B2(n11715), .ZN(
        n11722) );
  INV_X1 U14589 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11720) );
  INV_X1 U14590 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11719) );
  OAI22_X1 U14591 ( .A1(n11720), .A2(n11717), .B1(n11718), .B2(n11719), .ZN(
        n11721) );
  NOR2_X1 U14592 ( .A1(n11722), .A2(n11721), .ZN(n11734) );
  INV_X1 U14593 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11725) );
  INV_X1 U14594 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11724) );
  OAI22_X1 U14595 ( .A1(n20617), .A2(n11725), .B1(n20842), .B2(n11724), .ZN(
        n11726) );
  AOI21_X1 U14596 ( .B1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B2(n11723), .A(
        n11726), .ZN(n11733) );
  INV_X1 U14597 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11730) );
  INV_X1 U14598 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11729) );
  OAI22_X1 U14599 ( .A1(n11730), .A2(n11727), .B1(n11728), .B2(n11729), .ZN(
        n11731) );
  INV_X1 U14600 ( .A(n11731), .ZN(n11732) );
  NAND4_X1 U14601 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n11752) );
  AOI22_X1 U14602 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14603 ( .A1(n12322), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14604 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14605 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11737) );
  NAND4_X1 U14606 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n11750) );
  AOI22_X1 U14607 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11748) );
  NAND2_X1 U14608 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U14609 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11741) );
  OAI211_X1 U14610 ( .C1(n13067), .C2(n11743), .A(n11742), .B(n11741), .ZN(
        n11744) );
  INV_X1 U14611 ( .A(n11744), .ZN(n11747) );
  AOI22_X1 U14612 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11746) );
  NAND2_X1 U14613 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11745) );
  NAND4_X1 U14614 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n11749) );
  NAND2_X1 U14615 ( .A1(n12311), .A2(n20547), .ZN(n11751) );
  NAND2_X1 U14616 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11759) );
  INV_X1 U14617 ( .A(n11753), .ZN(n11755) );
  INV_X1 U14618 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11754) );
  OR2_X1 U14619 ( .A1(n11755), .A2(n11754), .ZN(n11758) );
  NAND2_X1 U14620 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11757) );
  NAND2_X1 U14621 ( .A1(n13058), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11756) );
  INV_X1 U14622 ( .A(n11855), .ZN(n13026) );
  INV_X1 U14623 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n20665) );
  INV_X1 U14624 ( .A(n12329), .ZN(n13028) );
  INV_X1 U14625 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11760) );
  OAI22_X1 U14626 ( .A1(n13026), .A2(n20665), .B1(n13028), .B2(n11760), .ZN(
        n11764) );
  INV_X1 U14627 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11762) );
  INV_X1 U14628 ( .A(n11856), .ZN(n13024) );
  INV_X1 U14629 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11761) );
  OAI22_X1 U14630 ( .A1(n11762), .A2(n13029), .B1(n13024), .B2(n11761), .ZN(
        n11763) );
  NOR2_X1 U14631 ( .A1(n11764), .A2(n11763), .ZN(n11782) );
  NAND2_X1 U14632 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11775) );
  INV_X1 U14633 ( .A(n12321), .ZN(n11766) );
  INV_X1 U14634 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11765) );
  OR2_X1 U14635 ( .A1(n11766), .A2(n11765), .ZN(n11774) );
  INV_X1 U14636 ( .A(n11767), .ZN(n11769) );
  INV_X1 U14637 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11768) );
  OR2_X1 U14638 ( .A1(n11769), .A2(n11768), .ZN(n11773) );
  INV_X1 U14639 ( .A(n12322), .ZN(n11771) );
  INV_X1 U14640 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11770) );
  OR2_X1 U14641 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  INV_X1 U14642 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14643 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n13063), .ZN(n11777) );
  NAND2_X1 U14644 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11776) );
  OAI211_X1 U14645 ( .C1(n13067), .C2(n11778), .A(n11777), .B(n11776), .ZN(
        n11779) );
  INV_X1 U14646 ( .A(n11779), .ZN(n11780) );
  XNOR2_X1 U14647 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12021) );
  NAND2_X1 U14648 ( .A1(n12021), .A2(n11809), .ZN(n11785) );
  NAND2_X1 U14649 ( .A1(n21203), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11784) );
  NAND2_X1 U14650 ( .A1(n11785), .A2(n11784), .ZN(n11792) );
  NOR2_X1 U14651 ( .A1(n17686), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11786) );
  MUX2_X1 U14652 ( .A(n12896), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11795) );
  INV_X1 U14653 ( .A(n11795), .ZN(n11787) );
  NAND3_X1 U14654 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12013), .A3(
        n17083), .ZN(n12197) );
  INV_X1 U14655 ( .A(n11789), .ZN(n12184) );
  MUX2_X1 U14656 ( .A(n12197), .B(n12151), .S(n12184), .Z(n12027) );
  INV_X1 U14657 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12041) );
  MUX2_X1 U14658 ( .A(n12027), .B(n12041), .S(n20565), .Z(n11820) );
  XNOR2_X1 U14659 ( .A(n17686), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11791) );
  XNOR2_X1 U14660 ( .A(n11792), .B(n11791), .ZN(n12187) );
  MUX2_X1 U14661 ( .A(n11793), .B(n12187), .S(n11789), .Z(n12022) );
  INV_X1 U14662 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14878) );
  MUX2_X1 U14663 ( .A(n12022), .B(n14878), .S(n20565), .Z(n11815) );
  NOR2_X1 U14664 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11794) );
  MUX2_X1 U14665 ( .A(n12141), .B(n11794), .S(n20565), .Z(n11816) );
  XNOR2_X1 U14666 ( .A(n11796), .B(n11795), .ZN(n12196) );
  INV_X1 U14667 ( .A(n12196), .ZN(n11797) );
  NAND2_X1 U14668 ( .A1(n11820), .A2(n11819), .ZN(n11799) );
  MUX2_X1 U14669 ( .A(n12311), .B(P2_EBX_REG_5__SCAN_IN), .S(n20565), .Z(
        n11798) );
  AND2_X1 U14670 ( .A1(n11799), .A2(n11798), .ZN(n11800) );
  OR2_X1 U14671 ( .A1(n11800), .A2(n11870), .ZN(n20362) );
  INV_X1 U14672 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15240) );
  INV_X1 U14673 ( .A(n9796), .ZN(n11805) );
  INV_X1 U14674 ( .A(n11803), .ZN(n11804) );
  INV_X1 U14675 ( .A(n11819), .ZN(n11808) );
  NAND2_X1 U14676 ( .A1(n11814), .A2(n11806), .ZN(n11807) );
  NAND2_X1 U14677 ( .A1(n11808), .A2(n11807), .ZN(n14784) );
  INV_X1 U14678 ( .A(n11809), .ZN(n12014) );
  NAND2_X1 U14679 ( .A1(n16927), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U14680 ( .A1(n12014), .A2(n11810), .ZN(n12191) );
  MUX2_X1 U14681 ( .A(n12275), .B(n12191), .S(n11789), .Z(n12024) );
  INV_X1 U14682 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n20397) );
  MUX2_X1 U14683 ( .A(n12024), .B(n20397), .S(n20565), .Z(n20398) );
  INV_X1 U14684 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13684) );
  INV_X1 U14685 ( .A(n11816), .ZN(n11812) );
  NAND3_X1 U14686 ( .A1(n20565), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U14687 ( .A1(n11812), .A2(n11811), .ZN(n16709) );
  NOR2_X1 U14688 ( .A1(n10342), .A2(n16709), .ZN(n11813) );
  NAND2_X1 U14689 ( .A1(n10342), .A2(n16709), .ZN(n16708) );
  OAI21_X1 U14690 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11813), .A(
        n16708), .ZN(n13706) );
  OAI21_X1 U14691 ( .B1(n11816), .B2(n11815), .A(n11814), .ZN(n11817) );
  INV_X1 U14692 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13747) );
  XNOR2_X1 U14693 ( .A(n11817), .B(n13747), .ZN(n13705) );
  OR2_X1 U14694 ( .A1(n13706), .A2(n13705), .ZN(n13708) );
  INV_X1 U14695 ( .A(n11817), .ZN(n14880) );
  NAND2_X1 U14696 ( .A1(n14880), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11818) );
  AND2_X1 U14697 ( .A1(n13708), .A2(n11818), .ZN(n17585) );
  INV_X1 U14698 ( .A(n14932), .ZN(n11822) );
  XNOR2_X1 U14699 ( .A(n11820), .B(n11819), .ZN(n20381) );
  INV_X1 U14700 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15942) );
  XNOR2_X1 U14701 ( .A(n20381), .B(n15942), .ZN(n14933) );
  INV_X1 U14702 ( .A(n14933), .ZN(n11821) );
  INV_X1 U14703 ( .A(n20381), .ZN(n11823) );
  NAND2_X1 U14704 ( .A1(n11823), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11824) );
  INV_X1 U14705 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11826) );
  INV_X1 U14706 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11825) );
  OAI22_X1 U14707 ( .A1(n11826), .A2(n20587), .B1(n14648), .B2(n11825), .ZN(
        n11830) );
  INV_X1 U14708 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13023) );
  INV_X1 U14709 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11827) );
  OAI22_X1 U14710 ( .A1(n13023), .A2(n11718), .B1(n20865), .B2(n11827), .ZN(
        n11829) );
  INV_X1 U14711 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14027) );
  INV_X1 U14712 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13025) );
  OR3_X2 U14713 ( .A1(n11830), .A2(n11829), .A3(n11828), .ZN(n11833) );
  INV_X1 U14714 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11831) );
  NOR2_X1 U14715 ( .A1(n11728), .A2(n11831), .ZN(n11832) );
  NOR2_X1 U14716 ( .A1(n11833), .A2(n11832), .ZN(n11850) );
  INV_X1 U14717 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U14718 ( .A1(n11834), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11837) );
  NAND2_X1 U14719 ( .A1(n11835), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11836) );
  OAI211_X1 U14720 ( .C1(n11704), .C2(n13030), .A(n11837), .B(n11836), .ZN(
        n11838) );
  INV_X1 U14721 ( .A(n11838), .ZN(n11849) );
  INV_X1 U14722 ( .A(n11723), .ZN(n11840) );
  INV_X1 U14723 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11839) );
  INV_X1 U14724 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13027) );
  OAI22_X1 U14725 ( .A1(n11840), .A2(n11839), .B1(n11727), .B2(n13027), .ZN(
        n11841) );
  INV_X1 U14726 ( .A(n11841), .ZN(n11848) );
  INV_X1 U14727 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16981) );
  INV_X1 U14728 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11842) );
  OAI22_X1 U14729 ( .A1(n16972), .A2(n16981), .B1(n20842), .B2(n11842), .ZN(
        n11846) );
  INV_X1 U14730 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11844) );
  INV_X1 U14731 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11843) );
  OAI22_X1 U14732 ( .A1(n11844), .A2(n11705), .B1(n11717), .B2(n11843), .ZN(
        n11845) );
  NOR2_X1 U14733 ( .A1(n11846), .A2(n11845), .ZN(n11847) );
  NAND4_X1 U14734 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11867) );
  AOI22_X1 U14735 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14736 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14737 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14738 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11851) );
  NAND4_X1 U14739 ( .A1(n11854), .A2(n11853), .A3(n11852), .A4(n11851), .ZN(
        n11865) );
  AOI22_X1 U14740 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n11856), .ZN(n11863) );
  NAND2_X1 U14741 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11858) );
  NAND2_X1 U14742 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11857) );
  OAI211_X1 U14743 ( .C1(n13067), .C2(n13025), .A(n11858), .B(n11857), .ZN(
        n11859) );
  INV_X1 U14744 ( .A(n11859), .ZN(n11862) );
  AOI22_X1 U14745 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11861) );
  NAND2_X1 U14746 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11860) );
  NAND4_X1 U14747 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(
        n11864) );
  INV_X1 U14748 ( .A(n11868), .ZN(n12315) );
  NAND2_X1 U14749 ( .A1(n12315), .A2(n20547), .ZN(n11866) );
  INV_X1 U14750 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n20348) );
  MUX2_X1 U14751 ( .A(n11868), .B(n20348), .S(n20565), .Z(n11869) );
  NOR2_X1 U14752 ( .A1(n11870), .A2(n11869), .ZN(n11871) );
  OR2_X1 U14753 ( .A1(n11875), .A2(n11871), .ZN(n20349) );
  NOR2_X1 U14754 ( .A1(n16700), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11884) );
  AND2_X2 U14755 ( .A1(n11872), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11881) );
  INV_X1 U14756 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13571) );
  NAND2_X1 U14757 ( .A1(n13570), .A2(n13571), .ZN(n11873) );
  NAND2_X1 U14758 ( .A1(n11873), .A2(n16700), .ZN(n11883) );
  INV_X1 U14759 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11874) );
  MUX2_X1 U14760 ( .A(n12003), .B(n11874), .S(n20565), .Z(n11878) );
  NAND2_X1 U14761 ( .A1(n20565), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11876) );
  OR2_X1 U14762 ( .A1(n11897), .A2(n11876), .ZN(n11877) );
  NAND2_X1 U14763 ( .A1(n11889), .A2(n11877), .ZN(n20323) );
  NOR2_X1 U14764 ( .A1(n20323), .A2(n11892), .ZN(n11885) );
  NAND2_X1 U14765 ( .A1(n11885), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17557) );
  INV_X1 U14766 ( .A(n11878), .ZN(n11879) );
  XNOR2_X1 U14767 ( .A(n11875), .B(n11879), .ZN(n11887) );
  NAND2_X1 U14768 ( .A1(n11887), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17553) );
  NAND2_X1 U14769 ( .A1(n17557), .A2(n17553), .ZN(n11880) );
  AOI21_X1 U14770 ( .B1(n11881), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11880), .ZN(n11882) );
  INV_X1 U14771 ( .A(n11885), .ZN(n11886) );
  INV_X1 U14772 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17643) );
  NAND2_X1 U14773 ( .A1(n11886), .A2(n17643), .ZN(n17556) );
  INV_X1 U14774 ( .A(n11887), .ZN(n20341) );
  INV_X1 U14775 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17657) );
  NAND2_X1 U14776 ( .A1(n20341), .A2(n17657), .ZN(n17552) );
  AND2_X1 U14777 ( .A1(n17556), .A2(n17552), .ZN(n11888) );
  NAND2_X1 U14778 ( .A1(n20565), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11890) );
  MUX2_X1 U14779 ( .A(n20565), .B(n11890), .S(n11889), .Z(n11891) );
  NAND2_X1 U14780 ( .A1(n10234), .A2(n11891), .ZN(n20310) );
  OR2_X1 U14781 ( .A1(n20310), .A2(n11892), .ZN(n11893) );
  INV_X1 U14782 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16908) );
  NAND2_X1 U14783 ( .A1(n20565), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11896) );
  MUX2_X1 U14784 ( .A(n11896), .B(P2_EBX_REG_10__SCAN_IN), .S(n11899), .Z(
        n11898) );
  AND2_X1 U14785 ( .A1(n11898), .A2(n11984), .ZN(n20300) );
  AOI21_X1 U14786 ( .B1(n20300), .B2(n12003), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16684) );
  INV_X1 U14787 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n20433) );
  INV_X1 U14788 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n20286) );
  NAND2_X2 U14789 ( .A1(n20276), .A2(n11984), .ZN(n11909) );
  INV_X1 U14790 ( .A(n11900), .ZN(n11901) );
  AND3_X1 U14791 ( .A1(n20565), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n11901), .ZN(
        n11902) );
  OR2_X1 U14792 ( .A1(n11909), .A2(n11902), .ZN(n20288) );
  INV_X1 U14793 ( .A(n20288), .ZN(n11903) );
  AOI21_X1 U14794 ( .B1(n11903), .B2(n12003), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16879) );
  INV_X1 U14795 ( .A(n20300), .ZN(n11904) );
  INV_X1 U14796 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16680) );
  OR3_X1 U14797 ( .A1(n11904), .A2(n11892), .A3(n16680), .ZN(n16682) );
  NAND2_X1 U14798 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11905) );
  OR2_X1 U14799 ( .A1(n20310), .A2(n11905), .ZN(n16897) );
  NAND2_X1 U14800 ( .A1(n16682), .A2(n16897), .ZN(n16877) );
  NAND2_X1 U14801 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11906) );
  NOR2_X1 U14802 ( .A1(n20288), .A2(n11906), .ZN(n16878) );
  NOR2_X1 U14803 ( .A1(n16877), .A2(n16878), .ZN(n11907) );
  NAND2_X1 U14804 ( .A1(n20565), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11908) );
  NAND2_X1 U14805 ( .A1(n20277), .A2(n12003), .ZN(n17535) );
  INV_X1 U14806 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11910) );
  AND2_X1 U14807 ( .A1(n20565), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11911) );
  INV_X1 U14808 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11912) );
  INV_X1 U14809 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n20266) );
  NAND2_X1 U14810 ( .A1(n11912), .A2(n20266), .ZN(n11913) );
  INV_X1 U14811 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11920) );
  INV_X1 U14812 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n16468) );
  NAND2_X1 U14813 ( .A1(n11920), .A2(n16468), .ZN(n11914) );
  NAND2_X1 U14814 ( .A1(n20565), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11943) );
  AND2_X1 U14815 ( .A1(n20565), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11915) );
  OR2_X2 U14816 ( .A1(n11941), .A2(n11915), .ZN(n11940) );
  NOR2_X2 U14817 ( .A1(n11940), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11918) );
  INV_X1 U14818 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11916) );
  NAND2_X1 U14819 ( .A1(n11918), .A2(n11916), .ZN(n11966) );
  NAND2_X1 U14820 ( .A1(n11966), .A2(n11984), .ZN(n11964) );
  NAND2_X1 U14821 ( .A1(n20565), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11917) );
  NOR2_X1 U14822 ( .A1(n11918), .A2(n11917), .ZN(n11919) );
  OR2_X1 U14823 ( .A1(n11964), .A2(n11919), .ZN(n13652) );
  INV_X1 U14824 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16787) );
  OAI21_X1 U14825 ( .B1(n13652), .B2(n11892), .A(n16787), .ZN(n16622) );
  INV_X1 U14826 ( .A(n11935), .ZN(n11921) );
  NAND2_X1 U14827 ( .A1(n11921), .A2(n11920), .ZN(n11926) );
  AND2_X1 U14828 ( .A1(n20565), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11923) );
  INV_X1 U14829 ( .A(n11984), .ZN(n11922) );
  AOI21_X1 U14830 ( .B1(n11935), .B2(n11923), .A(n11922), .ZN(n11924) );
  NAND2_X1 U14831 ( .A1(n20256), .A2(n12003), .ZN(n11925) );
  XNOR2_X1 U14832 ( .A(n11925), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12604) );
  INV_X1 U14833 ( .A(n11944), .ZN(n11928) );
  NAND3_X1 U14834 ( .A1(n11926), .A2(P2_EBX_REG_17__SCAN_IN), .A3(n20565), 
        .ZN(n11927) );
  NAND2_X1 U14835 ( .A1(n13636), .A2(n12003), .ZN(n11929) );
  INV_X1 U14836 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16834) );
  NAND2_X1 U14837 ( .A1(n11929), .A2(n16834), .ZN(n16656) );
  NAND2_X1 U14838 ( .A1(n20565), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11930) );
  MUX2_X1 U14839 ( .A(n20565), .B(n11930), .S(n11931), .Z(n11932) );
  OR2_X1 U14840 ( .A1(n11931), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11934) );
  AND2_X1 U14841 ( .A1(n11932), .A2(n11934), .ZN(n20268) );
  NAND2_X1 U14842 ( .A1(n20268), .A2(n12003), .ZN(n11955) );
  INV_X1 U14843 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17601) );
  NAND2_X1 U14844 ( .A1(n11955), .A2(n17601), .ZN(n17514) );
  AND2_X1 U14845 ( .A1(n20565), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11933) );
  NAND2_X1 U14846 ( .A1(n11934), .A2(n11933), .ZN(n11936) );
  AND2_X1 U14847 ( .A1(n11936), .A2(n11935), .ZN(n13622) );
  NAND2_X1 U14848 ( .A1(n13622), .A2(n12003), .ZN(n11937) );
  INV_X1 U14849 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16862) );
  NAND2_X1 U14850 ( .A1(n11937), .A2(n16862), .ZN(n16853) );
  NAND2_X1 U14851 ( .A1(n20565), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11938) );
  XNOR2_X1 U14852 ( .A(n20277), .B(n11938), .ZN(n15033) );
  NAND2_X1 U14853 ( .A1(n15033), .A2(n12003), .ZN(n11954) );
  INV_X1 U14854 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11953) );
  NAND2_X1 U14855 ( .A1(n11954), .A2(n11953), .ZN(n16866) );
  AND4_X1 U14856 ( .A1(n16656), .A2(n17514), .A3(n16853), .A4(n16866), .ZN(
        n11947) );
  NAND2_X1 U14857 ( .A1(n20565), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11939) );
  XNOR2_X1 U14858 ( .A(n11940), .B(n11939), .ZN(n20244) );
  AOI21_X1 U14859 ( .B1(n20244), .B2(n12003), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16619) );
  NAND2_X1 U14860 ( .A1(n20565), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11942) );
  XNOR2_X1 U14861 ( .A(n11941), .B(n11942), .ZN(n16382) );
  NAND2_X1 U14862 ( .A1(n16382), .A2(n12003), .ZN(n11959) );
  INV_X1 U14863 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16799) );
  NAND2_X1 U14864 ( .A1(n11959), .A2(n16799), .ZN(n16631) );
  OR2_X1 U14865 ( .A1(n11944), .A2(n11943), .ZN(n11945) );
  NAND2_X1 U14866 ( .A1(n11941), .A2(n11945), .ZN(n11949) );
  INV_X1 U14867 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16814) );
  OAI21_X1 U14868 ( .B1(n11949), .B2(n11892), .A(n16814), .ZN(n16646) );
  NAND2_X1 U14869 ( .A1(n16631), .A2(n16646), .ZN(n12608) );
  NOR2_X1 U14870 ( .A1(n16619), .A2(n12608), .ZN(n11946) );
  NAND2_X1 U14871 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11948) );
  OR2_X1 U14872 ( .A1(n13652), .A2(n11948), .ZN(n16621) );
  INV_X1 U14873 ( .A(n11949), .ZN(n16401) );
  AND2_X1 U14874 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U14875 ( .A1(n16401), .A2(n11950), .ZN(n16645) );
  AND2_X1 U14876 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11951) );
  NAND2_X1 U14877 ( .A1(n13636), .A2(n11951), .ZN(n16655) );
  AND2_X1 U14878 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11952) );
  NAND2_X1 U14879 ( .A1(n20256), .A2(n11952), .ZN(n12605) );
  OR2_X1 U14880 ( .A1(n11954), .A2(n11953), .ZN(n16867) );
  NAND4_X1 U14881 ( .A1(n16645), .A2(n16655), .A3(n12605), .A4(n16867), .ZN(
        n11958) );
  INV_X1 U14882 ( .A(n11955), .ZN(n11956) );
  NAND2_X1 U14883 ( .A1(n11956), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17515) );
  AND2_X1 U14884 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11957) );
  NAND2_X1 U14885 ( .A1(n13622), .A2(n11957), .ZN(n16852) );
  NAND2_X1 U14886 ( .A1(n17515), .A2(n16852), .ZN(n12603) );
  NOR2_X1 U14887 ( .A1(n11958), .A2(n12603), .ZN(n11961) );
  AND2_X1 U14888 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11960) );
  NAND2_X1 U14889 ( .A1(n20244), .A2(n11960), .ZN(n12609) );
  AND4_X1 U14890 ( .A1(n16621), .A2(n11961), .A3(n16632), .A4(n12609), .ZN(
        n11962) );
  NAND2_X1 U14891 ( .A1(n20565), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11965) );
  NAND2_X1 U14892 ( .A1(n11966), .A2(n10230), .ZN(n11967) );
  NAND2_X1 U14893 ( .A1(n11971), .A2(n11967), .ZN(n17122) );
  OR2_X1 U14894 ( .A1(n17122), .A2(n11892), .ZN(n11968) );
  INV_X1 U14895 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16776) );
  NAND2_X1 U14896 ( .A1(n11968), .A2(n16776), .ZN(n16606) );
  AND2_X1 U14897 ( .A1(n20565), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11970) );
  NAND2_X1 U14898 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  NAND2_X1 U14899 ( .A1(n11975), .A2(n11972), .ZN(n13665) );
  OR2_X1 U14900 ( .A1(n13665), .A2(n11892), .ZN(n11973) );
  XNOR2_X1 U14901 ( .A(n11973), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16598) );
  NAND2_X1 U14902 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11974) );
  NAND3_X1 U14903 ( .A1(n11975), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n20565), 
        .ZN(n11976) );
  NAND2_X1 U14904 ( .A1(n11976), .A2(n11984), .ZN(n11977) );
  NAND2_X1 U14905 ( .A1(n9834), .A2(n12003), .ZN(n16589) );
  NAND2_X1 U14906 ( .A1(n11978), .A2(n16589), .ZN(n11980) );
  NAND2_X1 U14907 ( .A1(n20565), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11981) );
  MUX2_X1 U14908 ( .A(n11981), .B(P2_EBX_REG_25__SCAN_IN), .S(n9860), .Z(
        n11982) );
  NAND2_X1 U14909 ( .A1(n11982), .A2(n11984), .ZN(n17445) );
  OR2_X1 U14910 ( .A1(n17445), .A2(n11892), .ZN(n11983) );
  INV_X1 U14911 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16747) );
  NAND2_X1 U14912 ( .A1(n11983), .A2(n16747), .ZN(n16577) );
  INV_X1 U14913 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n17441) );
  NAND2_X1 U14914 ( .A1(n11984), .A2(n9855), .ZN(n11989) );
  INV_X1 U14915 ( .A(n11989), .ZN(n12515) );
  NAND3_X1 U14916 ( .A1(n20565), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n11985), 
        .ZN(n11986) );
  OR2_X1 U14917 ( .A1(n17427), .A2(n11892), .ZN(n11987) );
  XNOR2_X1 U14918 ( .A(n11987), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16566) );
  NAND2_X1 U14919 ( .A1(n20565), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11990) );
  INV_X1 U14920 ( .A(n11990), .ZN(n11991) );
  NAND2_X1 U14921 ( .A1(n11991), .A2(n9855), .ZN(n11992) );
  NAND2_X1 U14922 ( .A1(n12001), .A2(n11992), .ZN(n13613) );
  INV_X1 U14923 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12882) );
  NAND2_X1 U14924 ( .A1(n11993), .A2(n12882), .ZN(n11995) );
  AND2_X1 U14925 ( .A1(n20565), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12000) );
  XOR2_X1 U14926 ( .A(n12000), .B(n12001), .Z(n17415) );
  NAND2_X1 U14927 ( .A1(n17415), .A2(n12003), .ZN(n12555) );
  OAI21_X1 U14928 ( .B1(n11997), .B2(n11995), .A(n11994), .ZN(n11999) );
  NAND2_X1 U14929 ( .A1(n12003), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11996) );
  NAND2_X1 U14930 ( .A1(n20565), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12004) );
  XNOR2_X1 U14931 ( .A(n12005), .B(n12004), .ZN(n12002) );
  INV_X1 U14932 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16717) );
  OAI21_X1 U14933 ( .B1(n12002), .B2(n11892), .A(n16717), .ZN(n16546) );
  NAND2_X1 U14934 ( .A1(n16547), .A2(n16546), .ZN(n12512) );
  INV_X1 U14935 ( .A(n12002), .ZN(n17407) );
  NAND3_X1 U14936 ( .A1(n17407), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12003), .ZN(n16545) );
  NAND2_X1 U14937 ( .A1(n12512), .A2(n16545), .ZN(n12010) );
  NAND2_X1 U14938 ( .A1(n12005), .A2(n12004), .ZN(n12513) );
  NAND2_X1 U14939 ( .A1(n20565), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12006) );
  XNOR2_X1 U14940 ( .A(n12513), .B(n12006), .ZN(n12007) );
  AOI21_X1 U14941 ( .B1(n12007), .B2(n12003), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12511) );
  INV_X1 U14942 ( .A(n12511), .ZN(n12008) );
  INV_X1 U14943 ( .A(n12007), .ZN(n12861) );
  INV_X1 U14944 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12499) );
  NAND2_X1 U14945 ( .A1(n12008), .A2(n12507), .ZN(n12009) );
  NAND2_X1 U14946 ( .A1(n17083), .A2(n12011), .ZN(n17712) );
  INV_X1 U14947 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13683) );
  OAI21_X1 U14948 ( .B1(n17712), .B2(n11650), .A(n13683), .ZN(n21204) );
  NOR2_X1 U14949 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17701), .ZN(
        n12012) );
  XNOR2_X1 U14950 ( .A(n12021), .B(n12014), .ZN(n12188) );
  AND4_X1 U14951 ( .A1(n12197), .A2(n12187), .A3(n12196), .A4(n12188), .ZN(
        n12015) );
  OR2_X1 U14952 ( .A1(n12203), .A2(n12015), .ZN(n17706) );
  INV_X1 U14953 ( .A(n12191), .ZN(n12016) );
  AND4_X1 U14954 ( .A1(n12197), .A2(n12016), .A3(n12187), .A4(n12196), .ZN(
        n12017) );
  NOR2_X1 U14955 ( .A1(n17706), .A2(n12017), .ZN(n12018) );
  MUX2_X1 U14956 ( .A(n21204), .B(n12018), .S(n12040), .Z(n17725) );
  INV_X1 U14957 ( .A(n12019), .ZN(n17715) );
  NAND3_X1 U14958 ( .A1(n17725), .A2(n17715), .A3(n11624), .ZN(n12031) );
  INV_X1 U14959 ( .A(n12203), .ZN(n21217) );
  AND2_X1 U14960 ( .A1(n17714), .A2(n20547), .ZN(n12213) );
  INV_X1 U14961 ( .A(n12213), .ZN(n12020) );
  NOR2_X1 U14962 ( .A1(n12019), .A2(n12020), .ZN(n21214) );
  INV_X1 U14963 ( .A(n12021), .ZN(n12190) );
  INV_X1 U14964 ( .A(n12022), .ZN(n12023) );
  OAI21_X1 U14965 ( .B1(n12024), .B2(n12190), .A(n12023), .ZN(n12029) );
  INV_X1 U14966 ( .A(n12025), .ZN(n12026) );
  NAND2_X1 U14967 ( .A1(n12027), .A2(n12026), .ZN(n12200) );
  INV_X1 U14968 ( .A(n12200), .ZN(n12028) );
  NAND2_X1 U14969 ( .A1(n12029), .A2(n12028), .ZN(n21216) );
  NAND3_X1 U14970 ( .A1(n21217), .A2(n21214), .A3(n21216), .ZN(n12030) );
  NAND2_X1 U14971 ( .A1(n12031), .A2(n12030), .ZN(n12205) );
  NAND2_X1 U14972 ( .A1(n12040), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12852) );
  INV_X1 U14973 ( .A(n12852), .ZN(n12032) );
  NOR2_X1 U14974 ( .A1(n11463), .A2(n15207), .ZN(n12033) );
  NAND2_X1 U14975 ( .A1(n12205), .A2(n12033), .ZN(n13682) );
  INV_X1 U14976 ( .A(n13682), .ZN(n12034) );
  INV_X1 U14977 ( .A(n12036), .ZN(n12037) );
  NAND2_X1 U14978 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  INV_X1 U14979 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n12040) );
  INV_X1 U14980 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20379) );
  OAI22_X1 U14981 ( .A1(n12045), .A2(n12041), .B1(n12040), .B2(n20379), .ZN(
        n12044) );
  NOR2_X1 U14982 ( .A1(n9789), .A2(n15942), .ZN(n12043) );
  AOI211_X1 U14983 ( .C1(n12074), .C2(P2_REIP_REG_4__SCAN_IN), .A(n12044), .B(
        n12043), .ZN(n14938) );
  NAND2_X1 U14984 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12049) );
  AOI22_X1 U14985 ( .A1(n12524), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12047) );
  NAND2_X1 U14986 ( .A1(n12074), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12046) );
  AND2_X1 U14987 ( .A1(n12047), .A2(n12046), .ZN(n12048) );
  NAND2_X1 U14988 ( .A1(n12049), .A2(n12048), .ZN(n15232) );
  AND2_X2 U14989 ( .A1(n15231), .A2(n15232), .ZN(n15234) );
  NAND2_X1 U14990 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12053) );
  AOI22_X1 U14991 ( .A1(n12524), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12051) );
  NAND2_X1 U14992 ( .A1(n12074), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12050) );
  AND2_X1 U14993 ( .A1(n12051), .A2(n12050), .ZN(n12052) );
  NAND2_X1 U14994 ( .A1(n12053), .A2(n12052), .ZN(n13580) );
  NAND2_X1 U14995 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12057) );
  AOI22_X1 U14996 ( .A1(n12524), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12055) );
  NAND2_X1 U14997 ( .A1(n12074), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12054) );
  AND2_X1 U14998 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  NAND2_X1 U14999 ( .A1(n12057), .A2(n12056), .ZN(n13931) );
  NAND2_X1 U15000 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12061) );
  AOI22_X1 U15001 ( .A1(n12524), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12059) );
  NAND2_X1 U15002 ( .A1(n12074), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12058) );
  AND2_X1 U15003 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  NAND2_X1 U15004 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12065) );
  AOI22_X1 U15005 ( .A1(n12524), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12063) );
  NAND2_X1 U15006 ( .A1(n12074), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12062) );
  AND2_X1 U15007 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  NAND2_X1 U15008 ( .A1(n12065), .A2(n12064), .ZN(n14006) );
  NAND2_X1 U15009 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12069) );
  AOI22_X1 U15010 ( .A1(n12524), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12067) );
  NAND2_X1 U15011 ( .A1(n12074), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12066) );
  AND2_X1 U15012 ( .A1(n12067), .A2(n12066), .ZN(n12068) );
  NAND2_X1 U15013 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12073) );
  AOI22_X1 U15014 ( .A1(n12524), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12071) );
  NAND2_X1 U15015 ( .A1(n12074), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12070) );
  AND2_X1 U15016 ( .A1(n12071), .A2(n12070), .ZN(n12072) );
  NAND2_X1 U15017 ( .A1(n12073), .A2(n12072), .ZN(n14291) );
  NAND2_X1 U15018 ( .A1(n14290), .A2(n14291), .ZN(n17532) );
  INV_X1 U15019 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12077) );
  NAND2_X1 U15020 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12076) );
  NAND2_X1 U15021 ( .A1(n12524), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12075) );
  OAI211_X1 U15022 ( .C1(n12528), .C2(n12077), .A(n12076), .B(n12075), .ZN(
        n12078) );
  AOI21_X1 U15023 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12078), .ZN(n17531) );
  INV_X1 U15024 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15036) );
  NAND2_X1 U15025 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12080) );
  AOI22_X1 U15026 ( .A1(n12524), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n12079) );
  OAI211_X1 U15027 ( .C1(n12528), .C2(n15036), .A(n12080), .B(n12079), .ZN(
        n14511) );
  NAND2_X1 U15028 ( .A1(n14510), .A2(n14511), .ZN(n14607) );
  INV_X1 U15029 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12083) );
  NAND2_X1 U15030 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12082) );
  NAND2_X1 U15031 ( .A1(n12524), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12081) );
  OAI211_X1 U15032 ( .C1(n12528), .C2(n12083), .A(n12082), .B(n12081), .ZN(
        n12084) );
  AOI21_X1 U15033 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n12084), .ZN(n14606) );
  INV_X1 U15034 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n12438) );
  NAND2_X1 U15035 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12087) );
  NAND2_X1 U15036 ( .A1(n12524), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12086) );
  OAI211_X1 U15037 ( .C1(n12528), .C2(n12438), .A(n12087), .B(n12086), .ZN(
        n12088) );
  AOI21_X1 U15038 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12088), .ZN(n13626) );
  INV_X1 U15039 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n12455) );
  NAND2_X1 U15040 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12090) );
  NAND2_X1 U15041 ( .A1(n12524), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12089) );
  OAI211_X1 U15042 ( .C1(n12528), .C2(n12455), .A(n12090), .B(n12089), .ZN(
        n12091) );
  AOI21_X1 U15043 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12091), .ZN(n16666) );
  INV_X1 U15044 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n21137) );
  NAND2_X1 U15045 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12094) );
  AOI22_X1 U15046 ( .A1(n12524), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12093) );
  OAI211_X1 U15047 ( .C1(n12528), .C2(n21137), .A(n12094), .B(n12093), .ZN(
        n13644) );
  INV_X1 U15048 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n21139) );
  NAND2_X1 U15049 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12096) );
  AOI22_X1 U15050 ( .A1(n12524), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12095) );
  OAI211_X1 U15051 ( .C1(n12528), .C2(n21139), .A(n12096), .B(n12095), .ZN(
        n16391) );
  INV_X1 U15052 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n21141) );
  NAND2_X1 U15053 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U15054 ( .A1(n12524), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12097) );
  OAI211_X1 U15055 ( .C1(n12528), .C2(n21141), .A(n12098), .B(n12097), .ZN(
        n12099) );
  AOI21_X1 U15056 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12099), .ZN(n16377) );
  INV_X1 U15057 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n21143) );
  NAND2_X1 U15058 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12101) );
  NAND2_X1 U15059 ( .A1(n12524), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12100) );
  OAI211_X1 U15060 ( .C1(n12528), .C2(n21143), .A(n12101), .B(n12100), .ZN(
        n12102) );
  AOI21_X1 U15061 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12102), .ZN(n12615) );
  INV_X1 U15062 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n21145) );
  NAND2_X1 U15063 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12104) );
  NAND2_X1 U15064 ( .A1(n12524), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12103) );
  OAI211_X1 U15065 ( .C1(n12528), .C2(n21145), .A(n12104), .B(n12103), .ZN(
        n12105) );
  AOI21_X1 U15066 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12105), .ZN(n13656) );
  INV_X1 U15067 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n17121) );
  NAND2_X1 U15068 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12107) );
  AOI22_X1 U15069 ( .A1(n12524), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12106) );
  OAI211_X1 U15070 ( .C1(n12528), .C2(n17121), .A(n12107), .B(n12106), .ZN(
        n16612) );
  INV_X1 U15071 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n21148) );
  NAND2_X1 U15072 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12109) );
  NAND2_X1 U15073 ( .A1(n12524), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12108) );
  OAI211_X1 U15074 ( .C1(n12528), .C2(n21148), .A(n12109), .B(n12108), .ZN(
        n12110) );
  AOI21_X1 U15075 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12110), .ZN(n13668) );
  INV_X1 U15076 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n12471) );
  NAND2_X1 U15077 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12112) );
  NAND2_X1 U15078 ( .A1(n12524), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12111) );
  OAI211_X1 U15079 ( .C1(n12528), .C2(n12471), .A(n12112), .B(n12111), .ZN(
        n12113) );
  AOI21_X1 U15080 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12113), .ZN(n16446) );
  INV_X1 U15081 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n21151) );
  NAND2_X1 U15082 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12115) );
  AOI22_X1 U15083 ( .A1(n12524), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12114) );
  OAI211_X1 U15084 ( .C1(n12528), .C2(n21151), .A(n12115), .B(n12114), .ZN(
        n16435) );
  INV_X1 U15085 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n21153) );
  NAND2_X1 U15086 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12117) );
  AOI22_X1 U15087 ( .A1(n12524), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12116) );
  OAI211_X1 U15088 ( .C1(n12528), .C2(n21153), .A(n12117), .B(n12116), .ZN(
        n16428) );
  INV_X1 U15089 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n21156) );
  NAND2_X1 U15090 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12119) );
  NAND2_X1 U15091 ( .A1(n12524), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12118) );
  OAI211_X1 U15092 ( .C1(n12528), .C2(n21156), .A(n12119), .B(n12118), .ZN(
        n12120) );
  AOI21_X1 U15093 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12120), .ZN(n12877) );
  INV_X1 U15094 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n21157) );
  NAND2_X1 U15095 ( .A1(n12129), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12122) );
  AOI22_X1 U15096 ( .A1(n12524), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12121) );
  OAI211_X1 U15097 ( .C1(n12528), .C2(n21157), .A(n12122), .B(n12121), .ZN(
        n12560) );
  NAND2_X1 U15098 ( .A1(n12561), .A2(n12560), .ZN(n16405) );
  INV_X1 U15099 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n21159) );
  NAND2_X1 U15100 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12124) );
  NAND2_X1 U15101 ( .A1(n12524), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12123) );
  OAI211_X1 U15102 ( .C1(n12528), .C2(n21159), .A(n12124), .B(n12123), .ZN(
        n12125) );
  AOI21_X1 U15103 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12125), .ZN(n16404) );
  INV_X1 U15104 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12860) );
  NAND2_X1 U15105 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12127) );
  NAND2_X1 U15106 ( .A1(n12524), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12126) );
  OAI211_X1 U15107 ( .C1(n12528), .C2(n12860), .A(n12127), .B(n12126), .ZN(
        n12128) );
  AOI21_X1 U15108 ( .B1(n12129), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12128), .ZN(n12522) );
  NOR2_X2 U15109 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n21177) );
  NOR2_X1 U15110 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n21082) );
  OR2_X1 U15111 ( .A1(n21177), .A2(n21082), .ZN(n21195) );
  NAND2_X1 U15112 ( .A1(n21195), .A2(n17682), .ZN(n12130) );
  AND2_X1 U15113 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n21196) );
  NAND2_X1 U15114 ( .A1(n12834), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12831) );
  INV_X1 U15115 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17511) );
  AND2_X1 U15116 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12131) );
  INV_X1 U15117 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16638) );
  NAND2_X1 U15118 ( .A1(n12827), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12826) );
  INV_X1 U15119 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16625) );
  INV_X1 U15120 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16599) );
  INV_X1 U15121 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16581) );
  INV_X1 U15122 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U15123 ( .A1(n12819), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12817) );
  INV_X1 U15124 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16558) );
  NAND2_X1 U15125 ( .A1(n12564), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12563) );
  INV_X1 U15126 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16549) );
  INV_X1 U15127 ( .A(n12590), .ZN(n12814) );
  INV_X1 U15128 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12136) );
  XNOR2_X1 U15129 ( .A(n12814), .B(n12136), .ZN(n16367) );
  INV_X1 U15130 ( .A(n16367), .ZN(n12138) );
  INV_X1 U15131 ( .A(n14011), .ZN(n12134) );
  INV_X1 U15132 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n12132) );
  NAND2_X1 U15133 ( .A1(n12132), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12133) );
  NAND2_X1 U15134 ( .A1(n12134), .A2(n12133), .ZN(n13691) );
  AND2_X1 U15135 ( .A1(n21177), .A2(n12135), .ZN(n12260) );
  INV_X2 U15136 ( .A(n20324), .ZN(n20376) );
  NAND2_X1 U15137 ( .A1(n20376), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12501) );
  OAI21_X1 U15138 ( .B1(n17596), .B2(n12136), .A(n12501), .ZN(n12137) );
  AOI21_X1 U15139 ( .B1(n12138), .B2(n17582), .A(n12137), .ZN(n12139) );
  OAI21_X1 U15140 ( .B1(n13218), .B2(n17577), .A(n12139), .ZN(n12140) );
  OR2_X1 U15141 ( .A1(n12275), .A2(n11624), .ZN(n13687) );
  NAND2_X1 U15142 ( .A1(n13687), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13686) );
  INV_X1 U15143 ( .A(n12275), .ZN(n12142) );
  XNOR2_X1 U15144 ( .A(n12142), .B(n12141), .ZN(n12143) );
  NOR2_X1 U15145 ( .A1(n13686), .A2(n12143), .ZN(n12144) );
  INV_X1 U15146 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16713) );
  XNOR2_X1 U15147 ( .A(n13686), .B(n12143), .ZN(n16712) );
  NOR2_X1 U15148 ( .A1(n16713), .A2(n16712), .ZN(n16711) );
  NOR2_X1 U15149 ( .A1(n12144), .A2(n16711), .ZN(n12146) );
  XNOR2_X1 U15150 ( .A(n12145), .B(n12289), .ZN(n13704) );
  NAND2_X1 U15151 ( .A1(n10355), .A2(n13704), .ZN(n13703) );
  OR2_X1 U15152 ( .A1(n12146), .A2(n13747), .ZN(n12147) );
  NAND2_X1 U15153 ( .A1(n13703), .A2(n12147), .ZN(n12149) );
  INV_X1 U15154 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17662) );
  XNOR2_X1 U15155 ( .A(n12149), .B(n17662), .ZN(n17587) );
  NAND2_X1 U15156 ( .A1(n12149), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12150) );
  INV_X1 U15157 ( .A(n12151), .ZN(n12306) );
  NAND2_X1 U15158 ( .A1(n12152), .A2(n12306), .ZN(n12153) );
  NAND2_X1 U15159 ( .A1(n10321), .A2(n12153), .ZN(n12154) );
  INV_X1 U15160 ( .A(n12154), .ZN(n12155) );
  NAND2_X1 U15161 ( .A1(n12156), .A2(n12155), .ZN(n12157) );
  INV_X1 U15162 ( .A(n12158), .ZN(n12159) );
  NAND2_X1 U15163 ( .A1(n12159), .A2(n15240), .ZN(n15224) );
  NAND2_X1 U15164 ( .A1(n12158), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15225) );
  NAND2_X1 U15165 ( .A1(n12161), .A2(n15225), .ZN(n12166) );
  INV_X1 U15166 ( .A(n15225), .ZN(n12163) );
  INV_X1 U15167 ( .A(n12170), .ZN(n12162) );
  NAND2_X1 U15168 ( .A1(n13568), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12168) );
  NAND2_X1 U15169 ( .A1(n12166), .A2(n12160), .ZN(n12167) );
  NAND2_X1 U15170 ( .A1(n12168), .A2(n12167), .ZN(n16694) );
  NAND2_X1 U15171 ( .A1(n16695), .A2(n17657), .ZN(n12172) );
  INV_X1 U15172 ( .A(n16695), .ZN(n12173) );
  NAND2_X1 U15173 ( .A1(n12173), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12174) );
  INV_X1 U15174 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16886) );
  NAND2_X1 U15175 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17614) );
  INV_X1 U15176 ( .A(n17614), .ZN(n12178) );
  NAND2_X1 U15177 ( .A1(n12178), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12496) );
  AND3_X1 U15178 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16813) );
  AND3_X1 U15179 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n16813), .ZN(n12181) );
  AND2_X1 U15180 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12180) );
  NAND2_X1 U15181 ( .A1(n12181), .A2(n12180), .ZN(n16762) );
  AND2_X1 U15182 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12497) );
  NAND2_X1 U15183 ( .A1(n12183), .A2(n12182), .ZN(P2_U2984) );
  NOR2_X1 U15184 ( .A1(n21227), .A2(n20547), .ZN(n12185) );
  MUX2_X1 U15185 ( .A(n12185), .B(n12184), .S(n12187), .Z(n12186) );
  INV_X1 U15186 ( .A(n12186), .ZN(n12195) );
  NAND2_X1 U15187 ( .A1(n20547), .A2(n12191), .ZN(n12189) );
  AOI22_X1 U15188 ( .A1(n12189), .A2(n12188), .B1(n20547), .B2(n12187), .ZN(
        n12193) );
  NOR2_X1 U15189 ( .A1(n12191), .A2(n12190), .ZN(n12192) );
  OAI22_X1 U15190 ( .A1(n12193), .A2(n17714), .B1(n12192), .B2(n11789), .ZN(
        n12194) );
  NAND2_X1 U15191 ( .A1(n12195), .A2(n12194), .ZN(n12199) );
  AND2_X1 U15192 ( .A1(n12197), .A2(n12196), .ZN(n12198) );
  AOI22_X1 U15193 ( .A1(n12200), .A2(n11789), .B1(n12199), .B2(n12198), .ZN(
        n12201) );
  OR2_X1 U15194 ( .A1(n12201), .A2(n12203), .ZN(n12202) );
  MUX2_X1 U15195 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12202), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12227) );
  NAND2_X1 U15196 ( .A1(n12203), .A2(n21227), .ZN(n12204) );
  NAND2_X1 U15197 ( .A1(n17709), .A2(n11624), .ZN(n13695) );
  INV_X1 U15198 ( .A(n13695), .ZN(n15201) );
  NAND2_X1 U15199 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n21236) );
  INV_X1 U15200 ( .A(n21236), .ZN(n21226) );
  NAND2_X1 U15201 ( .A1(n21099), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21245) );
  INV_X2 U15202 ( .A(n21245), .ZN(n21244) );
  NAND2_X2 U15203 ( .A1(n21244), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n21161) );
  NOR2_X1 U15204 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n21095) );
  INV_X1 U15205 ( .A(n21095), .ZN(n21106) );
  NAND3_X1 U15206 ( .A1(n21099), .A2(n21161), .A3(n21106), .ZN(n21229) );
  NOR2_X1 U15207 ( .A1(n21226), .A2(n21229), .ZN(n15197) );
  NAND3_X1 U15208 ( .A1(n15201), .A2(n15197), .A3(n12242), .ZN(n12232) );
  INV_X1 U15209 ( .A(n12205), .ZN(n12231) );
  NAND2_X1 U15210 ( .A1(n11480), .A2(n15197), .ZN(n12207) );
  OR2_X1 U15211 ( .A1(n17706), .A2(n12207), .ZN(n12223) );
  INV_X1 U15212 ( .A(n15199), .ZN(n12849) );
  NAND2_X1 U15213 ( .A1(n12208), .A2(n11482), .ZN(n12209) );
  NAND2_X1 U15214 ( .A1(n15199), .A2(n12209), .ZN(n12220) );
  NAND2_X1 U15215 ( .A1(n12211), .A2(n12210), .ZN(n12212) );
  NAND2_X1 U15216 ( .A1(n12212), .A2(n13777), .ZN(n12214) );
  NAND2_X1 U15217 ( .A1(n12214), .A2(n12213), .ZN(n12252) );
  OAI21_X1 U15218 ( .B1(n11624), .B2(n12215), .A(n11463), .ZN(n12217) );
  NAND2_X1 U15219 ( .A1(n12217), .A2(n12216), .ZN(n12218) );
  NAND2_X1 U15220 ( .A1(n12218), .A2(n11482), .ZN(n12219) );
  AND4_X1 U15221 ( .A1(n12221), .A2(n12220), .A3(n12252), .A4(n12219), .ZN(
        n12222) );
  NAND2_X1 U15222 ( .A1(n12223), .A2(n12222), .ZN(n15202) );
  MUX2_X1 U15223 ( .A(n11480), .B(n12242), .S(n20547), .Z(n12224) );
  NAND2_X1 U15224 ( .A1(n12224), .A2(n21236), .ZN(n12225) );
  NOR2_X1 U15225 ( .A1(n17706), .A2(n12225), .ZN(n12226) );
  NOR2_X1 U15226 ( .A1(n15202), .A2(n12226), .ZN(n12230) );
  AOI21_X1 U15227 ( .B1(n12227), .B2(n11463), .A(n12215), .ZN(n12228) );
  NAND2_X1 U15228 ( .A1(n13695), .A2(n12228), .ZN(n12229) );
  NAND4_X1 U15229 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12233) );
  NOR2_X1 U15230 ( .A1(n12019), .A2(n11789), .ZN(n21221) );
  NAND2_X1 U15231 ( .A1(n12236), .A2(n20547), .ZN(n12237) );
  NAND2_X1 U15232 ( .A1(n12234), .A2(n12237), .ZN(n12531) );
  NAND2_X1 U15233 ( .A1(n12505), .A2(n12531), .ZN(n17672) );
  AND3_X1 U15234 ( .A1(n11790), .A2(n20547), .A3(n11482), .ZN(n12238) );
  NAND2_X1 U15235 ( .A1(n12505), .A2(n17704), .ZN(n16823) );
  NOR2_X1 U15236 ( .A1(n12240), .A2(n12239), .ZN(n12241) );
  INV_X1 U15237 ( .A(n11502), .ZN(n12257) );
  NAND2_X1 U15238 ( .A1(n12241), .A2(n12257), .ZN(n13770) );
  NAND2_X1 U15239 ( .A1(n17714), .A2(n12242), .ZN(n12243) );
  OAI211_X1 U15240 ( .C1(n12215), .C2(n13681), .A(n13770), .B(n12243), .ZN(
        n12244) );
  INV_X1 U15241 ( .A(n12244), .ZN(n12249) );
  OAI21_X1 U15242 ( .B1(n12245), .B2(n12257), .A(n13681), .ZN(n12247) );
  NAND2_X1 U15243 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  AND3_X1 U15244 ( .A1(n12250), .A2(n12249), .A3(n12248), .ZN(n12256) );
  NAND2_X1 U15245 ( .A1(n12251), .A2(n9829), .ZN(n15187) );
  NAND2_X1 U15246 ( .A1(n15187), .A2(n12252), .ZN(n12254) );
  NAND2_X1 U15247 ( .A1(n12254), .A2(n12253), .ZN(n12255) );
  NAND2_X1 U15248 ( .A1(n12256), .A2(n12255), .ZN(n16964) );
  OR2_X1 U15249 ( .A1(n16964), .A2(n12257), .ZN(n12258) );
  NAND2_X1 U15250 ( .A1(n12505), .A2(n12258), .ZN(n12259) );
  INV_X1 U15251 ( .A(n17675), .ZN(n16922) );
  NAND2_X1 U15252 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15228) );
  NOR2_X1 U15253 ( .A1(n13571), .A2(n15228), .ZN(n17634) );
  NAND2_X1 U15254 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17634), .ZN(
        n13575) );
  NOR2_X1 U15255 ( .A1(n17657), .A2(n13575), .ZN(n17644) );
  NAND2_X1 U15256 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17644), .ZN(
        n12493) );
  NAND2_X1 U15257 ( .A1(n16922), .A2(n12493), .ZN(n12264) );
  INV_X1 U15258 ( .A(n12259), .ZN(n16825) );
  NAND3_X1 U15259 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U15260 ( .A1(n16825), .A2(n13749), .ZN(n12262) );
  INV_X1 U15261 ( .A(n12505), .ZN(n12261) );
  INV_X1 U15262 ( .A(n12260), .ZN(n20347) );
  NAND2_X1 U15263 ( .A1(n12261), .A2(n20347), .ZN(n17670) );
  AND2_X1 U15264 ( .A1(n12262), .A2(n17670), .ZN(n13574) );
  INV_X1 U15265 ( .A(n16823), .ZN(n13752) );
  NAND2_X1 U15266 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16921) );
  NAND2_X1 U15267 ( .A1(n13747), .A2(n16921), .ZN(n13748) );
  INV_X1 U15268 ( .A(n13748), .ZN(n12492) );
  NAND2_X1 U15269 ( .A1(n13752), .A2(n12492), .ZN(n12263) );
  AND3_X1 U15270 ( .A1(n12264), .A2(n13574), .A3(n12263), .ZN(n16909) );
  NAND2_X1 U15271 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12494) );
  OAI21_X1 U15272 ( .B1(n16908), .B2(n12494), .A(n16922), .ZN(n12265) );
  NAND2_X1 U15273 ( .A1(n16909), .A2(n12265), .ZN(n17616) );
  NOR2_X1 U15274 ( .A1(n17675), .A2(n12179), .ZN(n12266) );
  OR2_X1 U15275 ( .A1(n17616), .A2(n12266), .ZN(n16861) );
  NOR2_X1 U15276 ( .A1(n17675), .A2(n10289), .ZN(n12267) );
  OR2_X1 U15277 ( .A1(n16861), .A2(n12267), .ZN(n16792) );
  OAI21_X1 U15278 ( .B1(n17675), .B2(n12497), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12268) );
  NOR2_X1 U15279 ( .A1(n16792), .A2(n12268), .ZN(n16752) );
  NAND2_X1 U15280 ( .A1(n17675), .A2(n17670), .ZN(n14944) );
  INV_X1 U15281 ( .A(n14944), .ZN(n12269) );
  OR2_X1 U15282 ( .A1(n16752), .A2(n12269), .ZN(n16746) );
  INV_X1 U15283 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16729) );
  OR2_X1 U15284 ( .A1(n16747), .A2(n16729), .ZN(n16730) );
  NAND2_X1 U15285 ( .A1(n14944), .A2(n16730), .ZN(n12270) );
  NAND2_X1 U15286 ( .A1(n16746), .A2(n12270), .ZN(n12875) );
  AND3_X1 U15287 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12542) );
  NOR2_X1 U15288 ( .A1(n17675), .A2(n12542), .ZN(n12271) );
  NOR2_X1 U15289 ( .A1(n12875), .A2(n12271), .ZN(n12535) );
  INV_X1 U15290 ( .A(n12535), .ZN(n12503) );
  NAND2_X1 U15291 ( .A1(n12482), .A2(n12272), .ZN(n12287) );
  NOR2_X1 U15292 ( .A1(n12273), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12274) );
  OAI22_X1 U15294 ( .A1(n13777), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n21212), 
        .B2(n20975), .ZN(n12276) );
  NAND2_X1 U15295 ( .A1(n12287), .A2(n12278), .ZN(n13761) );
  INV_X1 U15296 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n20395) );
  NAND2_X1 U15297 ( .A1(n20573), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12279) );
  OAI211_X1 U15298 ( .C1(n20547), .C2(n13684), .A(n12279), .B(n20975), .ZN(
        n12280) );
  INV_X1 U15299 ( .A(n12280), .ZN(n12281) );
  NAND2_X1 U15300 ( .A1(n12282), .A2(n12281), .ZN(n13762) );
  INV_X1 U15301 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n20539) );
  INV_X1 U15302 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n21114) );
  OAI222_X1 U15303 ( .A1(n12537), .A2(n16713), .B1(n9897), .B2(n20539), .C1(
        n12290), .C2(n21114), .ZN(n12286) );
  NOR3_X1 U15304 ( .A1(n12272), .A2(n20573), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12283) );
  AOI21_X1 U15305 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_3__SCAN_IN), .A(n12283), .ZN(n12284) );
  OAI21_X1 U15306 ( .B1(n12285), .B2(n12435), .A(n12284), .ZN(n13936) );
  NAND2_X1 U15307 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12288) );
  OAI211_X1 U15308 ( .C1(n12435), .C2(n12289), .A(n12288), .B(n12287), .ZN(
        n12293) );
  INV_X1 U15309 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n21116) );
  OR2_X1 U15310 ( .A1(n12290), .A2(n21116), .ZN(n12292) );
  INV_X2 U15311 ( .A(n12537), .ZN(n12482) );
  AOI22_X1 U15312 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12291) );
  NAND2_X1 U15313 ( .A1(n12292), .A2(n12291), .ZN(n13740) );
  NOR2_X1 U15314 ( .A1(n13741), .A2(n13740), .ZN(n13742) );
  NOR2_X1 U15315 ( .A1(n12294), .A2(n12293), .ZN(n12295) );
  OR2_X1 U15316 ( .A1(n12290), .A2(n21118), .ZN(n12302) );
  OR2_X1 U15317 ( .A1(n12435), .A2(n12296), .ZN(n12300) );
  NAND2_X1 U15318 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12299) );
  NAND2_X1 U15319 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12298) );
  NAND2_X1 U15320 ( .A1(n12481), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12297) );
  NAND2_X1 U15321 ( .A1(n12302), .A2(n12301), .ZN(n14357) );
  INV_X1 U15322 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12303) );
  OR2_X1 U15323 ( .A1(n12290), .A2(n12303), .ZN(n12309) );
  NAND2_X1 U15324 ( .A1(n12481), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n12305) );
  NAND2_X1 U15325 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12304) );
  OAI211_X1 U15326 ( .C1(n12435), .C2(n12306), .A(n12305), .B(n12304), .ZN(
        n12307) );
  INV_X1 U15327 ( .A(n12307), .ZN(n12308) );
  INV_X1 U15328 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15235) );
  OAI22_X1 U15329 ( .A1(n12290), .A2(n15235), .B1(n12537), .B2(n15240), .ZN(
        n12310) );
  INV_X1 U15330 ( .A(n12310), .ZN(n12314) );
  INV_X1 U15331 ( .A(n12311), .ZN(n12312) );
  AOI22_X1 U15332 ( .A1(n12277), .A2(n12312), .B1(n12481), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n12313) );
  NAND2_X1 U15333 ( .A1(n12314), .A2(n12313), .ZN(n15230) );
  OR2_X1 U15334 ( .A1(n12435), .A2(n12315), .ZN(n12316) );
  INV_X1 U15335 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n21121) );
  OR2_X1 U15336 ( .A1(n12290), .A2(n21121), .ZN(n12318) );
  AOI22_X1 U15337 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U15338 ( .A1(n12318), .A2(n12317), .ZN(n13579) );
  NAND2_X1 U15339 ( .A1(n13578), .A2(n13579), .ZN(n12319) );
  INV_X1 U15340 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20525) );
  INV_X1 U15341 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n21123) );
  OAI222_X1 U15342 ( .A1(n17657), .A2(n12537), .B1(n9897), .B2(n20525), .C1(
        n12290), .C2(n21123), .ZN(n17649) );
  INV_X1 U15343 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12320) );
  OR2_X1 U15344 ( .A1(n12290), .A2(n12320), .ZN(n12340) );
  AOI22_X1 U15345 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15346 ( .A1(n12322), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15347 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U15348 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12323) );
  NAND4_X1 U15349 ( .A1(n12326), .A2(n12325), .A3(n12324), .A4(n12323), .ZN(
        n12335) );
  AOI22_X1 U15350 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15351 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13063), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U15352 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12327) );
  AND2_X1 U15353 ( .A1(n12328), .A2(n12327), .ZN(n12332) );
  AOI22_X1 U15354 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12331) );
  NAND2_X1 U15355 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12330) );
  NAND4_X1 U15356 ( .A1(n12333), .A2(n12332), .A3(n12331), .A4(n12330), .ZN(
        n12334) );
  NOR2_X1 U15357 ( .A1(n12335), .A2(n12334), .ZN(n13968) );
  NAND2_X1 U15358 ( .A1(n12481), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n12337) );
  NAND2_X1 U15359 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12336) );
  OAI211_X1 U15360 ( .C1(n12435), .C2(n13968), .A(n12337), .B(n12336), .ZN(
        n12338) );
  INV_X1 U15361 ( .A(n12338), .ZN(n12339) );
  AOI22_X1 U15362 ( .A1(n10193), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n12482), 
        .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15363 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15364 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15365 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15366 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12341) );
  NAND4_X1 U15367 ( .A1(n12344), .A2(n12343), .A3(n12342), .A4(n12341), .ZN(
        n12354) );
  AOI22_X1 U15368 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n11856), .ZN(n12352) );
  INV_X1 U15369 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12347) );
  NAND2_X1 U15370 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12346) );
  NAND2_X1 U15371 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12345) );
  OAI211_X1 U15372 ( .C1(n13067), .C2(n12347), .A(n12346), .B(n12345), .ZN(
        n12348) );
  INV_X1 U15373 ( .A(n12348), .ZN(n12351) );
  AOI22_X1 U15374 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12350) );
  NAND2_X1 U15375 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12349) );
  NAND4_X1 U15376 ( .A1(n12352), .A2(n12351), .A3(n12350), .A4(n12349), .ZN(
        n12353) );
  AOI22_X1 U15377 ( .A1(n12277), .A2(n20427), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n12481), .ZN(n12355) );
  NAND2_X1 U15378 ( .A1(n12356), .A2(n12355), .ZN(n16903) );
  AOI22_X1 U15379 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n11736), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15380 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12322), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15381 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15382 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11681), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12357) );
  NAND4_X1 U15383 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n12357), .ZN(
        n12368) );
  AOI22_X1 U15384 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15385 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n13063), .ZN(n12362) );
  NAND2_X1 U15386 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12361) );
  AND2_X1 U15387 ( .A1(n12362), .A2(n12361), .ZN(n12365) );
  AOI22_X1 U15388 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12364) );
  NAND2_X1 U15389 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12363) );
  NAND4_X1 U15390 ( .A1(n12366), .A2(n12365), .A3(n12364), .A4(n12363), .ZN(
        n12367) );
  INV_X1 U15391 ( .A(n20426), .ZN(n12370) );
  AOI22_X1 U15392 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12369) );
  OAI21_X1 U15393 ( .B1(n12370), .B2(n12435), .A(n12369), .ZN(n12371) );
  AOI21_X1 U15394 ( .B1(n10193), .B2(P2_REIP_REG_10__SCAN_IN), .A(n12371), 
        .ZN(n17624) );
  AOI22_X1 U15395 ( .A1(n10193), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n12482), .ZN(n12387) );
  AOI22_X1 U15396 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15397 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15398 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12373) );
  AOI22_X1 U15399 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12372) );
  NAND4_X1 U15400 ( .A1(n12375), .A2(n12374), .A3(n12373), .A4(n12372), .ZN(
        n12385) );
  INV_X1 U15401 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15997) );
  AOI22_X1 U15402 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12383) );
  NAND2_X1 U15403 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12377) );
  NAND2_X1 U15404 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12376) );
  OAI211_X1 U15405 ( .C1(n13067), .C2(n12378), .A(n12377), .B(n12376), .ZN(
        n12379) );
  INV_X1 U15406 ( .A(n12379), .ZN(n12382) );
  AOI22_X1 U15407 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12381) );
  NAND2_X1 U15408 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12380) );
  NAND4_X1 U15409 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n12380), .ZN(
        n12384) );
  AOI22_X1 U15410 ( .A1(n12277), .A2(n20421), .B1(P2_EAX_REG_11__SCAN_IN), 
        .B2(n12481), .ZN(n12386) );
  NAND2_X1 U15411 ( .A1(n12387), .A2(n12386), .ZN(n16883) );
  NAND2_X1 U15412 ( .A1(n16884), .A2(n16883), .ZN(n16882) );
  AOI22_X1 U15413 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11855), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12391) );
  AOI22_X1 U15414 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11767), .B1(
        n12322), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12390) );
  AOI22_X1 U15415 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15416 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11681), .B1(
        n11672), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12388) );
  NAND4_X1 U15417 ( .A1(n12391), .A2(n12390), .A3(n12389), .A4(n12388), .ZN(
        n12401) );
  AOI22_X1 U15418 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__4__SCAN_IN), .B2(n11856), .ZN(n12399) );
  INV_X1 U15419 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12394) );
  NAND2_X1 U15420 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12393) );
  NAND2_X1 U15421 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12392) );
  OAI211_X1 U15422 ( .C1(n13067), .C2(n12394), .A(n12393), .B(n12392), .ZN(
        n12395) );
  INV_X1 U15423 ( .A(n12395), .ZN(n12398) );
  AOI22_X1 U15424 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12397) );
  NAND2_X1 U15425 ( .A1(n13058), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12396) );
  NAND4_X1 U15426 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12400) );
  INV_X1 U15427 ( .A(n20420), .ZN(n12403) );
  AOI22_X1 U15428 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12402) );
  OAI21_X1 U15429 ( .B1(n12403), .B2(n12435), .A(n12402), .ZN(n12404) );
  AOI21_X1 U15430 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n10193), .A(n12404), 
        .ZN(n17615) );
  AOI22_X1 U15431 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15432 ( .A1(n12321), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12322), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15433 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15434 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12405) );
  NAND4_X1 U15435 ( .A1(n12408), .A2(n12407), .A3(n12406), .A4(n12405), .ZN(
        n12418) );
  AOI22_X1 U15436 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12416) );
  NAND2_X1 U15437 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12410) );
  NAND2_X1 U15438 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12409) );
  OAI211_X1 U15439 ( .C1(n13067), .C2(n12411), .A(n12410), .B(n12409), .ZN(
        n12412) );
  INV_X1 U15440 ( .A(n12412), .ZN(n12415) );
  AOI22_X1 U15441 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12414) );
  NAND2_X1 U15442 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12413) );
  NAND4_X1 U15443 ( .A1(n12416), .A2(n12415), .A3(n12414), .A4(n12413), .ZN(
        n12417) );
  AOI22_X1 U15444 ( .A1(n10193), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n12277), 
        .B2(n14602), .ZN(n12420) );
  AOI22_X1 U15445 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U15446 ( .A1(n12420), .A2(n12419), .ZN(n15032) );
  AOI22_X1 U15447 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11855), .B1(
        n12322), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U15448 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11767), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U15449 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15450 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n13058), .B1(
        n11672), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12421) );
  NAND4_X1 U15451 ( .A1(n12424), .A2(n12423), .A3(n12422), .A4(n12421), .ZN(
        n12433) );
  AOI22_X1 U15452 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n11856), .ZN(n12431) );
  AOI22_X1 U15453 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n13063), .ZN(n12426) );
  NAND2_X1 U15454 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12425) );
  AND2_X1 U15455 ( .A1(n12426), .A2(n12425), .ZN(n12430) );
  AOI22_X1 U15456 ( .A1(n12427), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12429) );
  NAND2_X1 U15457 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12428) );
  NAND4_X1 U15458 ( .A1(n12431), .A2(n12430), .A3(n12429), .A4(n12428), .ZN(
        n12432) );
  INV_X1 U15459 ( .A(n14604), .ZN(n12436) );
  AOI22_X1 U15460 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12434) );
  OAI21_X1 U15461 ( .B1(n12436), .B2(n12435), .A(n12434), .ZN(n12437) );
  AOI21_X1 U15462 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n10193), .A(n12437), 
        .ZN(n17599) );
  INV_X1 U15463 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13921) );
  OAI22_X1 U15464 ( .A1(n12290), .A2(n12438), .B1(n9897), .B2(n13921), .ZN(
        n12439) );
  INV_X1 U15465 ( .A(n12439), .ZN(n12454) );
  AOI22_X1 U15466 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U15467 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U15468 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U15469 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12440) );
  NAND4_X1 U15470 ( .A1(n12443), .A2(n12442), .A3(n12441), .A4(n12440), .ZN(
        n12452) );
  AOI22_X1 U15471 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n11856), .ZN(n12450) );
  INV_X1 U15472 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15872) );
  NAND2_X1 U15473 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12445) );
  NAND2_X1 U15474 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12444) );
  OAI211_X1 U15475 ( .C1(n13067), .C2(n15872), .A(n12445), .B(n12444), .ZN(
        n12446) );
  INV_X1 U15476 ( .A(n12446), .ZN(n12449) );
  AOI22_X1 U15477 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12448) );
  NAND2_X1 U15478 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12447) );
  NAND4_X1 U15479 ( .A1(n12450), .A2(n12449), .A3(n12448), .A4(n12447), .ZN(
        n12451) );
  NOR2_X1 U15480 ( .A1(n12452), .A2(n12451), .ZN(n14871) );
  AOI22_X1 U15481 ( .A1(n12277), .A2(n12933), .B1(n12482), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12453) );
  NAND2_X1 U15482 ( .A1(n12454), .A2(n12453), .ZN(n13625) );
  OR2_X1 U15483 ( .A1(n12290), .A2(n12455), .ZN(n12457) );
  AOI22_X1 U15484 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n12456) );
  OR2_X1 U15485 ( .A1(n12290), .A2(n21137), .ZN(n12459) );
  AOI22_X1 U15486 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12458) );
  NAND2_X1 U15487 ( .A1(n12459), .A2(n12458), .ZN(n13642) );
  NAND2_X1 U15488 ( .A1(n13640), .A2(n13642), .ZN(n13641) );
  OR2_X1 U15489 ( .A1(n12290), .A2(n21139), .ZN(n12461) );
  AOI22_X1 U15490 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12460) );
  AND2_X1 U15491 ( .A1(n12461), .A2(n12460), .ZN(n16390) );
  OR2_X1 U15492 ( .A1(n12290), .A2(n21141), .ZN(n12463) );
  AOI22_X1 U15493 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12462) );
  OR2_X1 U15494 ( .A1(n12290), .A2(n21143), .ZN(n12466) );
  AOI22_X1 U15495 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12465) );
  NAND2_X1 U15496 ( .A1(n12466), .A2(n12465), .ZN(n12623) );
  INV_X1 U15497 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13700) );
  OAI222_X1 U15498 ( .A1(n12290), .A2(n21145), .B1(n9897), .B2(n13700), .C1(
        n16787), .C2(n12537), .ZN(n13655) );
  OR2_X1 U15499 ( .A1(n12290), .A2(n17121), .ZN(n12468) );
  AOI22_X1 U15500 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12467) );
  NAND2_X1 U15501 ( .A1(n12468), .A2(n12467), .ZN(n16775) );
  INV_X1 U15502 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12469) );
  INV_X1 U15503 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16522) );
  OAI22_X1 U15504 ( .A1(n12537), .A2(n12469), .B1(n9897), .B2(n16522), .ZN(
        n12470) );
  AOI21_X1 U15505 ( .B1(n10193), .B2(P2_REIP_REG_23__SCAN_IN), .A(n12470), 
        .ZN(n13671) );
  OR2_X1 U15506 ( .A1(n12290), .A2(n12471), .ZN(n12473) );
  AOI22_X1 U15507 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12472) );
  NAND2_X1 U15508 ( .A1(n12473), .A2(n12472), .ZN(n16510) );
  INV_X1 U15509 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n16504) );
  OAI22_X1 U15510 ( .A1(n12537), .A2(n16747), .B1(n9897), .B2(n16504), .ZN(
        n12474) );
  AOI21_X1 U15511 ( .B1(n10193), .B2(P2_REIP_REG_25__SCAN_IN), .A(n12474), 
        .ZN(n16501) );
  INV_X1 U15512 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n16495) );
  OAI22_X1 U15513 ( .A1(n12537), .A2(n16729), .B1(n9897), .B2(n16495), .ZN(
        n12475) );
  AOI21_X1 U15514 ( .B1(n10193), .B2(P2_REIP_REG_26__SCAN_IN), .A(n12475), 
        .ZN(n16493) );
  INV_X1 U15515 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n16487) );
  OAI22_X1 U15516 ( .A1(n12537), .A2(n12882), .B1(n9897), .B2(n16487), .ZN(
        n12476) );
  AOI21_X1 U15517 ( .B1(n10193), .B2(P2_REIP_REG_27__SCAN_IN), .A(n12476), 
        .ZN(n12869) );
  OR2_X1 U15518 ( .A1(n12290), .A2(n21157), .ZN(n12478) );
  AOI22_X1 U15519 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12477) );
  NAND2_X1 U15520 ( .A1(n12478), .A2(n12477), .ZN(n12579) );
  OR2_X1 U15521 ( .A1(n12290), .A2(n21159), .ZN(n12480) );
  AOI22_X1 U15522 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U15523 ( .A1(n12480), .A2(n12479), .ZN(n16472) );
  OR2_X1 U15524 ( .A1(n12290), .A2(n12860), .ZN(n12484) );
  AOI22_X1 U15525 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n12481), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n12483) );
  NAND2_X1 U15526 ( .A1(n12484), .A2(n12483), .ZN(n12485) );
  OR2_X1 U15527 ( .A1(n16474), .A2(n12485), .ZN(n12486) );
  INV_X1 U15528 ( .A(n12487), .ZN(n12488) );
  AND2_X1 U15529 ( .A1(n12488), .A2(n15189), .ZN(n17708) );
  NOR2_X1 U15530 ( .A1(n12489), .A2(n20547), .ZN(n12490) );
  OR2_X1 U15531 ( .A1(n17708), .A2(n12490), .ZN(n12491) );
  AOI211_X1 U15532 ( .C1(n16823), .C2(n13749), .A(n12492), .B(n17675), .ZN(
        n17663) );
  INV_X1 U15533 ( .A(n17663), .ZN(n13572) );
  NOR2_X1 U15534 ( .A1(n12493), .A2(n13572), .ZN(n16905) );
  NAND2_X1 U15535 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16905), .ZN(
        n17625) );
  NOR2_X2 U15536 ( .A1(n12494), .A2(n17625), .ZN(n17619) );
  INV_X1 U15537 ( .A(n17619), .ZN(n12495) );
  INV_X1 U15538 ( .A(n12497), .ZN(n16763) );
  NOR2_X1 U15539 ( .A1(n16762), .A2(n16763), .ZN(n12498) );
  NAND2_X1 U15540 ( .A1(n16857), .A2(n12498), .ZN(n16753) );
  NAND3_X1 U15541 ( .A1(n16718), .A2(n12499), .A3(n12542), .ZN(n12500) );
  OAI211_X1 U15542 ( .C1(n15415), .C2(n17671), .A(n12501), .B(n12500), .ZN(
        n12502) );
  INV_X1 U15543 ( .A(n16545), .ZN(n12508) );
  OAI21_X2 U15544 ( .B1(n12512), .B2(n12511), .A(n12510), .ZN(n12518) );
  NOR2_X1 U15545 ( .A1(n12513), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12514) );
  MUX2_X1 U15546 ( .A(n12515), .B(n12514), .S(n20565), .Z(n16372) );
  NAND2_X1 U15547 ( .A1(n16372), .A2(n12003), .ZN(n12516) );
  INV_X1 U15548 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12541) );
  XNOR2_X1 U15549 ( .A(n12516), .B(n12541), .ZN(n12517) );
  XNOR2_X1 U15550 ( .A(n12518), .B(n12517), .ZN(n12598) );
  NAND2_X1 U15551 ( .A1(n12598), .A2(n17639), .ZN(n12551) );
  NAND2_X1 U15552 ( .A1(n12519), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12520) );
  NAND2_X1 U15553 ( .A1(n10349), .A2(n12521), .ZN(n12550) );
  NOR2_X2 U15554 ( .A1(n12523), .A2(n12522), .ZN(n12534) );
  NAND2_X1 U15555 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12811) );
  INV_X1 U15556 ( .A(n12811), .ZN(n12530) );
  INV_X1 U15557 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U15558 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12526) );
  NAND2_X1 U15559 ( .A1(n12524), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12525) );
  OAI211_X1 U15560 ( .C1(n12528), .C2(n12527), .A(n12526), .B(n12525), .ZN(
        n12529) );
  AOI21_X1 U15561 ( .B1(n12531), .B2(n12530), .A(n12529), .ZN(n12532) );
  INV_X1 U15562 ( .A(n12532), .ZN(n12533) );
  OAI21_X1 U15563 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17675), .A(
        n12535), .ZN(n12546) );
  INV_X1 U15564 ( .A(P2_EAX_REG_31__SCAN_IN), .ZN(n12536) );
  OAI22_X1 U15565 ( .A1(n12537), .A2(n12541), .B1(n9897), .B2(n12536), .ZN(
        n12538) );
  AOI21_X1 U15566 ( .B1(n10193), .B2(P2_REIP_REG_31__SCAN_IN), .A(n12538), 
        .ZN(n12539) );
  NAND2_X1 U15567 ( .A1(n20376), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12593) );
  INV_X1 U15568 ( .A(n12593), .ZN(n12543) );
  OAI21_X1 U15569 ( .B1(n16369), .B2(n17671), .A(n12544), .ZN(n12545) );
  OAI21_X1 U15570 ( .B1(n17465), .B2(n17672), .A(n12547), .ZN(n12548) );
  NAND3_X1 U15571 ( .A1(n12551), .A2(n12550), .A3(n12549), .ZN(P2_U3015) );
  XNOR2_X1 U15572 ( .A(n12554), .B(n12553), .ZN(n12883) );
  OAI22_X1 U15573 ( .A1(n12883), .A2(n12882), .B1(n12554), .B2(n12553), .ZN(
        n12557) );
  XOR2_X1 U15574 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n12555), .Z(
        n12556) );
  XNOR2_X1 U15575 ( .A(n12557), .B(n12556), .ZN(n12573) );
  NAND2_X1 U15576 ( .A1(n12573), .A2(n17592), .ZN(n12572) );
  OAI21_X1 U15577 ( .B1(n12558), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12559), .ZN(n12586) );
  OR2_X1 U15578 ( .A1(n12561), .A2(n12560), .ZN(n12562) );
  NAND2_X1 U15579 ( .A1(n16405), .A2(n12562), .ZN(n17417) );
  INV_X1 U15580 ( .A(n17417), .ZN(n12568) );
  OR2_X1 U15581 ( .A1(n12564), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12565) );
  NAND2_X1 U15582 ( .A1(n12563), .A2(n12565), .ZN(n12816) );
  NAND2_X1 U15583 ( .A1(n20376), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12581) );
  NAND2_X1 U15584 ( .A1(n17564), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12566) );
  OAI211_X1 U15585 ( .C1(n17571), .C2(n12816), .A(n12581), .B(n12566), .ZN(
        n12567) );
  AOI21_X1 U15586 ( .B1(n12568), .B2(n17591), .A(n12567), .ZN(n12569) );
  NAND2_X1 U15587 ( .A1(n12572), .A2(n12571), .ZN(P2_U2986) );
  NAND2_X1 U15588 ( .A1(n12573), .A2(n17639), .ZN(n12589) );
  INV_X1 U15589 ( .A(n12875), .ZN(n12576) );
  NAND2_X1 U15590 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U15591 ( .A1(n16718), .A2(n12574), .ZN(n12575) );
  NAND2_X1 U15592 ( .A1(n12576), .A2(n12575), .ZN(n16722) );
  INV_X1 U15593 ( .A(n16718), .ZN(n12577) );
  OAI21_X1 U15594 ( .B1(n12577), .B2(n12882), .A(n11993), .ZN(n12584) );
  NOR2_X1 U15595 ( .A1(n12871), .A2(n12579), .ZN(n12580) );
  OAI21_X1 U15596 ( .B1(n17671), .B2(n17416), .A(n12581), .ZN(n12583) );
  NOR2_X1 U15597 ( .A1(n17417), .A2(n17672), .ZN(n12582) );
  AOI211_X1 U15598 ( .C1(n16722), .C2(n12584), .A(n12583), .B(n12582), .ZN(
        n12585) );
  NAND2_X1 U15599 ( .A1(n12589), .A2(n12588), .ZN(P2_U3018) );
  NAND2_X1 U15600 ( .A1(n12590), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12592) );
  INV_X1 U15601 ( .A(n12812), .ZN(n12595) );
  OAI21_X1 U15602 ( .B1(n17596), .B2(n12591), .A(n12593), .ZN(n12594) );
  AOI21_X1 U15603 ( .B1(n17582), .B2(n12595), .A(n12594), .ZN(n12596) );
  OAI21_X1 U15604 ( .B1(n17465), .B2(n17577), .A(n12596), .ZN(n12597) );
  AOI21_X1 U15605 ( .B1(n12598), .B2(n17592), .A(n12597), .ZN(n12601) );
  NAND2_X1 U15606 ( .A1(n12601), .A2(n12600), .ZN(P2_U2983) );
  INV_X1 U15607 ( .A(n16866), .ZN(n12602) );
  INV_X1 U15608 ( .A(n12604), .ZN(n16673) );
  INV_X1 U15609 ( .A(n12605), .ZN(n12606) );
  INV_X1 U15610 ( .A(n16656), .ZN(n12607) );
  AOI21_X2 U15611 ( .B1(n16634), .B2(n16632), .A(n12608), .ZN(n12612) );
  INV_X1 U15612 ( .A(n16619), .ZN(n12610) );
  NAND2_X1 U15613 ( .A1(n12610), .A2(n12609), .ZN(n12611) );
  AOI21_X1 U15614 ( .B1(n12612), .B2(n12611), .A(n16620), .ZN(n12886) );
  XNOR2_X1 U15615 ( .A(n16637), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12887) );
  OR2_X1 U15616 ( .A1(n12887), .A2(n17669), .ZN(n12627) );
  NAND2_X1 U15617 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16813), .ZN(
        n12616) );
  AOI21_X1 U15618 ( .B1(n16922), .B2(n12616), .A(n16861), .ZN(n16812) );
  INV_X1 U15619 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12621) );
  INV_X1 U15620 ( .A(n13657), .ZN(n12614) );
  AOI21_X1 U15621 ( .B1(n12615), .B2(n16379), .A(n12614), .ZN(n20245) );
  NOR2_X1 U15622 ( .A1(n20324), .A2(n21143), .ZN(n12888) );
  NOR2_X1 U15623 ( .A1(n16839), .A2(n12616), .ZN(n16800) );
  INV_X1 U15624 ( .A(n16800), .ZN(n12618) );
  NAND2_X1 U15625 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16785) );
  OAI21_X1 U15626 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n16785), .ZN(n12617) );
  NOR2_X1 U15627 ( .A1(n12618), .A2(n12617), .ZN(n12619) );
  AOI211_X1 U15628 ( .C1(n20245), .C2(n12878), .A(n12888), .B(n12619), .ZN(
        n12620) );
  OAI21_X1 U15629 ( .B1(n16812), .B2(n12621), .A(n12620), .ZN(n12625) );
  NOR2_X1 U15630 ( .A1(n10356), .A2(n12623), .ZN(n12624) );
  NOR2_X1 U15631 ( .A1(n15741), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12630) );
  OAI21_X1 U15632 ( .B1(n15744), .B2(n10339), .A(n12631), .ZN(n12632) );
  XNOR2_X1 U15633 ( .A(n12632), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15433) );
  INV_X1 U15634 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12634) );
  NAND2_X1 U15635 ( .A1(n12635), .A2(n12634), .ZN(n17186) );
  NAND2_X1 U15636 ( .A1(n13984), .A2(n17186), .ZN(n15101) );
  NAND2_X1 U15637 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21452) );
  NAND2_X1 U15638 ( .A1(n15101), .A2(n21452), .ZN(n12636) );
  OAI211_X1 U15639 ( .C1(n12633), .C2(n12636), .A(n15100), .B(n10505), .ZN(
        n12637) );
  NAND3_X1 U15640 ( .A1(n12640), .A2(n12639), .A3(n12638), .ZN(n12641) );
  NAND2_X1 U15641 ( .A1(n12642), .A2(n12641), .ZN(n12643) );
  NAND2_X1 U15642 ( .A1(n12644), .A2(n12643), .ZN(n13722) );
  INV_X1 U15643 ( .A(n21452), .ZN(n21541) );
  AOI21_X1 U15644 ( .B1(n17165), .B2(n17186), .A(n21541), .ZN(n12645) );
  NAND2_X1 U15645 ( .A1(n13722), .A2(n12645), .ZN(n12646) );
  NAND2_X1 U15646 ( .A1(n13870), .A2(n17165), .ZN(n12656) );
  INV_X1 U15647 ( .A(n12647), .ZN(n12655) );
  INV_X1 U15648 ( .A(n12648), .ZN(n12649) );
  NAND3_X1 U15649 ( .A1(n12650), .A2(n10514), .A3(n12649), .ZN(n12652) );
  AND2_X1 U15650 ( .A1(n12652), .A2(n12651), .ZN(n12782) );
  OR2_X1 U15651 ( .A1(n12653), .A2(n12782), .ZN(n12654) );
  NAND2_X1 U15652 ( .A1(n12655), .A2(n12654), .ZN(n13853) );
  OAI21_X1 U15653 ( .B1(n17170), .B2(n12656), .A(n13853), .ZN(n12657) );
  INV_X1 U15654 ( .A(n12657), .ZN(n12658) );
  NAND2_X1 U15655 ( .A1(n12659), .A2(n12658), .ZN(n12660) );
  NOR2_X1 U15656 ( .A1(n13910), .A2(n12661), .ZN(n13954) );
  INV_X1 U15657 ( .A(n12662), .ZN(n15116) );
  NAND2_X1 U15658 ( .A1(n13954), .A2(n15116), .ZN(n13858) );
  OAI211_X1 U15659 ( .C1(n10532), .C2(n9962), .A(n17150), .B(n13858), .ZN(
        n12663) );
  INV_X1 U15660 ( .A(n12663), .ZN(n12664) );
  AND2_X1 U15661 ( .A1(n12665), .A2(n12664), .ZN(n12666) );
  NAND2_X1 U15662 ( .A1(n13953), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U15663 ( .A1(n14135), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12667) );
  NAND2_X1 U15664 ( .A1(n12668), .A2(n12667), .ZN(n15452) );
  INV_X1 U15665 ( .A(n12732), .ZN(n13715) );
  MUX2_X1 U15666 ( .A(n12764), .B(n12732), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n12670) );
  OR2_X1 U15667 ( .A1(n13953), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12669) );
  NAND2_X1 U15668 ( .A1(n12670), .A2(n12669), .ZN(n12674) );
  INV_X1 U15669 ( .A(n12688), .ZN(n12677) );
  INV_X1 U15670 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12671) );
  OR2_X1 U15671 ( .A1(n12755), .A2(n12671), .ZN(n12673) );
  NAND2_X1 U15672 ( .A1(n13715), .A2(n12671), .ZN(n12672) );
  NAND2_X1 U15673 ( .A1(n12673), .A2(n12672), .ZN(n13951) );
  XNOR2_X1 U15674 ( .A(n12674), .B(n13951), .ZN(n14136) );
  MUX2_X1 U15675 ( .A(n12764), .B(n12759), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12676) );
  OR2_X1 U15676 ( .A1(n13953), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12675) );
  AND2_X1 U15677 ( .A1(n12676), .A2(n12675), .ZN(n13978) );
  NAND2_X1 U15678 ( .A1(n13979), .A2(n13978), .ZN(n14151) );
  INV_X1 U15679 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12678) );
  NAND2_X1 U15680 ( .A1(n12747), .A2(n12678), .ZN(n12682) );
  NAND2_X1 U15681 ( .A1(n12755), .A2(n14368), .ZN(n12680) );
  NAND3_X1 U15682 ( .A1(n12680), .A2(n12759), .A3(n12679), .ZN(n12681) );
  AND2_X1 U15683 ( .A1(n12682), .A2(n12681), .ZN(n14150) );
  NAND2_X1 U15684 ( .A1(n12759), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12683) );
  OAI211_X1 U15685 ( .C1(n14135), .C2(P1_EBX_REG_4__SCAN_IN), .A(n12755), .B(
        n12683), .ZN(n12684) );
  OAI21_X1 U15686 ( .B1(n12764), .B2(P1_EBX_REG_4__SCAN_IN), .A(n12684), .ZN(
        n14372) );
  NOR2_X2 U15687 ( .A1(n14373), .A2(n14372), .ZN(n14977) );
  INV_X1 U15688 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21369) );
  NAND2_X1 U15689 ( .A1(n12738), .A2(n21369), .ZN(n12687) );
  NAND2_X1 U15690 ( .A1(n12759), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12685) );
  OAI211_X1 U15691 ( .C1(n14135), .C2(P1_EBX_REG_6__SCAN_IN), .A(n12755), .B(
        n12685), .ZN(n12686) );
  AND2_X1 U15692 ( .A1(n12687), .A2(n12686), .ZN(n14975) );
  OR2_X1 U15693 ( .A1(n12768), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n12692) );
  NAND2_X1 U15694 ( .A1(n12732), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12689) );
  NAND2_X1 U15695 ( .A1(n12755), .A2(n12689), .ZN(n12690) );
  OAI21_X1 U15696 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n14135), .A(n12690), .ZN(
        n12691) );
  NAND2_X1 U15697 ( .A1(n12692), .A2(n12691), .ZN(n14976) );
  AND2_X1 U15698 ( .A1(n14975), .A2(n14976), .ZN(n12693) );
  OR2_X1 U15699 ( .A1(n12768), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n12697) );
  NAND2_X1 U15700 ( .A1(n12759), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12694) );
  NAND2_X1 U15701 ( .A1(n12755), .A2(n12694), .ZN(n12695) );
  OAI21_X1 U15702 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n14135), .A(n12695), .ZN(
        n12696) );
  NAND2_X1 U15703 ( .A1(n12697), .A2(n12696), .ZN(n14889) );
  NAND2_X1 U15704 ( .A1(n14979), .A2(n14889), .ZN(n15142) );
  NAND2_X1 U15705 ( .A1(n12759), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12698) );
  OAI211_X1 U15706 ( .C1(n14135), .C2(P1_EBX_REG_8__SCAN_IN), .A(n12755), .B(
        n12698), .ZN(n12699) );
  OAI21_X1 U15707 ( .B1(n12764), .B2(P1_EBX_REG_8__SCAN_IN), .A(n12699), .ZN(
        n15143) );
  MUX2_X1 U15708 ( .A(n12764), .B(n12759), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12701) );
  OR2_X1 U15709 ( .A1(n13953), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12700) );
  NAND2_X1 U15710 ( .A1(n12701), .A2(n12700), .ZN(n15159) );
  INV_X1 U15711 ( .A(n15159), .ZN(n12706) );
  OR2_X1 U15712 ( .A1(n12768), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n12705) );
  NAND2_X1 U15713 ( .A1(n12732), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12702) );
  NAND2_X1 U15714 ( .A1(n12755), .A2(n12702), .ZN(n12703) );
  OAI21_X1 U15715 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n14135), .A(n12703), .ZN(
        n12704) );
  NAND2_X1 U15716 ( .A1(n12705), .A2(n12704), .ZN(n15094) );
  NAND2_X1 U15717 ( .A1(n12706), .A2(n15094), .ZN(n12707) );
  NOR2_X2 U15718 ( .A1(n15161), .A2(n12707), .ZN(n15360) );
  INV_X1 U15719 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n17256) );
  NAND2_X1 U15720 ( .A1(n12738), .A2(n17256), .ZN(n12710) );
  NAND2_X1 U15721 ( .A1(n12759), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12708) );
  OAI211_X1 U15722 ( .C1(n14135), .C2(P1_EBX_REG_12__SCAN_IN), .A(n12755), .B(
        n12708), .ZN(n12709) );
  AND2_X1 U15723 ( .A1(n12710), .A2(n12709), .ZN(n15358) );
  OR2_X1 U15724 ( .A1(n12768), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n12714) );
  NAND2_X1 U15725 ( .A1(n12759), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12711) );
  NAND2_X1 U15726 ( .A1(n12755), .A2(n12711), .ZN(n12712) );
  OAI21_X1 U15727 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(n14135), .A(n12712), .ZN(
        n12713) );
  NAND2_X1 U15728 ( .A1(n12714), .A2(n12713), .ZN(n15359) );
  AND2_X2 U15729 ( .A1(n15360), .A2(n12715), .ZN(n15362) );
  INV_X1 U15730 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n17237) );
  NAND2_X1 U15731 ( .A1(n12747), .A2(n17237), .ZN(n12719) );
  INV_X1 U15732 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U15733 ( .A1(n12755), .A2(n12799), .ZN(n12717) );
  NAND3_X1 U15734 ( .A1(n12717), .A2(n12759), .A3(n12716), .ZN(n12718) );
  NAND2_X1 U15735 ( .A1(n12719), .A2(n12718), .ZN(n15339) );
  MUX2_X1 U15736 ( .A(n12764), .B(n12759), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12720) );
  OAI21_X1 U15737 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n13953), .A(
        n12720), .ZN(n15590) );
  OR2_X1 U15738 ( .A1(n12768), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n12724) );
  NAND2_X1 U15739 ( .A1(n12759), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12721) );
  NAND2_X1 U15740 ( .A1(n12755), .A2(n12721), .ZN(n12722) );
  OAI21_X1 U15741 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(n14135), .A(n12722), .ZN(
        n12723) );
  INV_X1 U15742 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15640) );
  NAND2_X1 U15743 ( .A1(n12738), .A2(n15640), .ZN(n12727) );
  NAND2_X1 U15744 ( .A1(n12759), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12725) );
  OAI211_X1 U15745 ( .C1(n14135), .C2(P1_EBX_REG_16__SCAN_IN), .A(n12755), .B(
        n12725), .ZN(n12726) );
  INV_X1 U15746 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n17253) );
  NAND2_X1 U15747 ( .A1(n12747), .A2(n17253), .ZN(n12731) );
  NAND2_X1 U15748 ( .A1(n12755), .A2(n16280), .ZN(n12729) );
  NAND3_X1 U15749 ( .A1(n12729), .A2(n12759), .A3(n12728), .ZN(n12730) );
  MUX2_X1 U15750 ( .A(n12764), .B(n12732), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12733) );
  OAI21_X1 U15751 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n13953), .A(
        n12733), .ZN(n15636) );
  OR3_X2 U15752 ( .A1(n16278), .A2(n16279), .A3(n15636), .ZN(n15637) );
  INV_X1 U15753 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n17212) );
  NAND2_X1 U15754 ( .A1(n12747), .A2(n17212), .ZN(n12737) );
  NAND2_X1 U15755 ( .A1(n12755), .A2(n16253), .ZN(n12735) );
  NAND3_X1 U15756 ( .A1(n12735), .A2(n12759), .A3(n12734), .ZN(n12736) );
  NOR2_X2 U15757 ( .A1(n15637), .A2(n15629), .ZN(n15630) );
  INV_X1 U15758 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15623) );
  NAND2_X1 U15759 ( .A1(n12738), .A2(n15623), .ZN(n12741) );
  NAND2_X1 U15760 ( .A1(n12759), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12739) );
  OAI211_X1 U15761 ( .C1(n14135), .C2(P1_EBX_REG_20__SCAN_IN), .A(n12755), .B(
        n12739), .ZN(n12740) );
  AND2_X1 U15762 ( .A1(n12741), .A2(n12740), .ZN(n15549) );
  INV_X1 U15763 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n17200) );
  NAND2_X1 U15764 ( .A1(n12747), .A2(n17200), .ZN(n12745) );
  NAND2_X1 U15765 ( .A1(n12755), .A2(n16235), .ZN(n12743) );
  NAND3_X1 U15766 ( .A1(n12743), .A2(n12759), .A3(n12742), .ZN(n12744) );
  NAND2_X1 U15767 ( .A1(n12745), .A2(n12744), .ZN(n15617) );
  MUX2_X1 U15768 ( .A(n12764), .B(n12759), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12746) );
  OAI21_X1 U15769 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n13953), .A(
        n12746), .ZN(n15614) );
  INV_X1 U15770 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n12748) );
  NAND2_X1 U15771 ( .A1(n12747), .A2(n12748), .ZN(n12752) );
  INV_X1 U15772 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16207) );
  NAND2_X1 U15773 ( .A1(n12755), .A2(n16207), .ZN(n12750) );
  NAND3_X1 U15774 ( .A1(n12750), .A2(n12759), .A3(n12749), .ZN(n12751) );
  AND2_X1 U15775 ( .A1(n12752), .A2(n12751), .ZN(n15536) );
  MUX2_X1 U15776 ( .A(n12764), .B(n12759), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12754) );
  OR2_X1 U15777 ( .A1(n13953), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12753) );
  AND2_X1 U15778 ( .A1(n12754), .A2(n12753), .ZN(n15524) );
  OR2_X1 U15779 ( .A1(n12768), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n12758) );
  NAND2_X1 U15780 ( .A1(n12755), .A2(n16197), .ZN(n12756) );
  OAI211_X1 U15781 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n14135), .A(n12756), .B(
        n12759), .ZN(n12757) );
  NAND2_X1 U15782 ( .A1(n12758), .A2(n12757), .ZN(n15510) );
  MUX2_X1 U15783 ( .A(n12764), .B(n12759), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12760) );
  OAI21_X1 U15784 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n13953), .A(
        n12760), .ZN(n15498) );
  OR2_X1 U15785 ( .A1(n12768), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n12763) );
  NAND2_X1 U15786 ( .A1(n12755), .A2(n16191), .ZN(n12761) );
  OAI211_X1 U15787 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n14135), .A(n12761), .B(
        n12759), .ZN(n12762) );
  AND2_X1 U15788 ( .A1(n12763), .A2(n12762), .ZN(n15485) );
  MUX2_X1 U15789 ( .A(n12764), .B(n12759), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12765) );
  OAI21_X1 U15790 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n13953), .A(
        n12765), .ZN(n15473) );
  NOR2_X2 U15791 ( .A1(n15487), .A2(n15473), .ZN(n15474) );
  OR2_X1 U15792 ( .A1(n13953), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12767) );
  INV_X1 U15793 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15601) );
  NAND2_X1 U15794 ( .A1(n12767), .A2(n12766), .ZN(n15449) );
  OAI22_X1 U15795 ( .A1(n15449), .A2(n13715), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12768), .ZN(n15465) );
  NAND2_X1 U15796 ( .A1(n15474), .A2(n15465), .ZN(n15464) );
  MUX2_X1 U15797 ( .A(n15452), .B(n13715), .S(n15464), .Z(n12772) );
  INV_X1 U15798 ( .A(n15464), .ZN(n15450) );
  NAND2_X1 U15799 ( .A1(n15450), .A2(n15452), .ZN(n12771) );
  AND2_X1 U15800 ( .A1(n14135), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12769) );
  AOI21_X1 U15801 ( .B1(n13953), .B2(P1_EBX_REG_31__SCAN_IN), .A(n12769), .ZN(
        n12770) );
  INV_X1 U15802 ( .A(n15598), .ZN(n12793) );
  OAI22_X1 U15803 ( .A1(n12774), .A2(n17165), .B1(n14049), .B2(n9962), .ZN(
        n12775) );
  INV_X1 U15804 ( .A(n12775), .ZN(n12776) );
  NOR2_X2 U15805 ( .A1(n12795), .A2(n12776), .ZN(n21427) );
  INV_X1 U15806 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21513) );
  NOR2_X1 U15807 ( .A1(n17352), .A2(n21513), .ZN(n15428) );
  AOI21_X1 U15808 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14149) );
  NOR2_X1 U15809 ( .A1(n14369), .A2(n14368), .ZN(n14618) );
  NAND2_X1 U15810 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14618), .ZN(
        n12796) );
  NOR2_X1 U15811 ( .A1(n14149), .A2(n12796), .ZN(n14614) );
  INV_X1 U15812 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13876) );
  NOR2_X1 U15813 ( .A1(n13876), .A2(n11201), .ZN(n14145) );
  NAND2_X1 U15814 ( .A1(n12647), .A2(n17165), .ZN(n17128) );
  INV_X1 U15815 ( .A(n13866), .ZN(n12790) );
  INV_X1 U15816 ( .A(n12777), .ZN(n12788) );
  NAND2_X1 U15817 ( .A1(n12778), .A2(n15116), .ZN(n12787) );
  INV_X1 U15818 ( .A(n13851), .ZN(n15104) );
  NAND2_X1 U15819 ( .A1(n15104), .A2(n12779), .ZN(n12780) );
  AND2_X1 U15820 ( .A1(n12781), .A2(n12780), .ZN(n12786) );
  INV_X1 U15821 ( .A(n12782), .ZN(n12785) );
  OR2_X1 U15822 ( .A1(n12783), .A2(n13984), .ZN(n12784) );
  NAND4_X1 U15823 ( .A1(n12787), .A2(n12786), .A3(n12785), .A4(n12784), .ZN(
        n13883) );
  AOI211_X1 U15824 ( .C1(n12790), .C2(n12789), .A(n12788), .B(n13883), .ZN(
        n12791) );
  NOR2_X1 U15825 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21432), .ZN(
        n14137) );
  NAND2_X1 U15826 ( .A1(n14614), .A2(n17354), .ZN(n14981) );
  NOR3_X1 U15827 ( .A1(n15138), .A2(n15137), .A3(n14982), .ZN(n15386) );
  NAND3_X1 U15828 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n15386), .ZN(n15355) );
  NOR2_X1 U15829 ( .A1(n11273), .A2(n15355), .ZN(n12794) );
  NAND2_X1 U15830 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n12794), .ZN(
        n12798) );
  INV_X1 U15831 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16280) );
  NAND2_X1 U15832 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16300) );
  NOR2_X1 U15833 ( .A1(n16280), .A2(n16300), .ZN(n16267) );
  NAND3_X1 U15834 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n16267), .ZN(n12801) );
  NOR2_X1 U15835 ( .A1(n12799), .A2(n12801), .ZN(n16227) );
  NAND3_X1 U15836 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n16227), .ZN(n16222) );
  NOR2_X1 U15837 ( .A1(n12798), .A2(n16222), .ZN(n12802) );
  NAND3_X1 U15838 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n12802), .ZN(n16204) );
  NOR2_X1 U15839 ( .A1(n14981), .A2(n16204), .ZN(n17349) );
  NAND3_X1 U15840 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17349), .ZN(n17335) );
  NOR2_X1 U15841 ( .A1(n16197), .A2(n17335), .ZN(n17338) );
  NAND2_X1 U15842 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17338), .ZN(
        n16187) );
  NOR2_X1 U15843 ( .A1(n17325), .A2(n16187), .ZN(n17313) );
  NAND2_X1 U15844 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17313), .ZN(
        n16178) );
  NOR3_X1 U15845 ( .A1(n16178), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16179), .ZN(n12792) );
  AOI211_X1 U15846 ( .C1(n12793), .C2(n21427), .A(n15428), .B(n12792), .ZN(
        n12809) );
  OR2_X1 U15847 ( .A1(n14615), .A2(n16216), .ZN(n21430) );
  OR2_X1 U15848 ( .A1(n21432), .A2(n21430), .ZN(n12806) );
  INV_X1 U15849 ( .A(n12806), .ZN(n14138) );
  NAND2_X1 U15850 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12805) );
  INV_X1 U15851 ( .A(n14617), .ZN(n15349) );
  NOR2_X1 U15852 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n16220), .ZN(
        n12804) );
  NAND2_X1 U15853 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12803) );
  AND2_X1 U15854 ( .A1(n12794), .A2(n14614), .ZN(n15353) );
  NAND2_X1 U15855 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15353), .ZN(
        n16219) );
  NOR2_X1 U15856 ( .A1(n12799), .A2(n16219), .ZN(n17355) );
  INV_X1 U15857 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14158) );
  INV_X1 U15858 ( .A(n12796), .ZN(n12797) );
  NAND2_X1 U15859 ( .A1(n14145), .A2(n12797), .ZN(n15350) );
  NOR2_X1 U15860 ( .A1(n15350), .A2(n12798), .ZN(n16221) );
  INV_X1 U15861 ( .A(n16221), .ZN(n16218) );
  OAI21_X1 U15862 ( .B1(n12799), .B2(n16218), .A(n15349), .ZN(n12800) );
  NAND2_X1 U15863 ( .A1(n14138), .A2(n15351), .ZN(n16262) );
  INV_X1 U15864 ( .A(n16262), .ZN(n16263) );
  AOI21_X1 U15865 ( .B1(n16256), .B2(n12802), .A(n16263), .ZN(n16239) );
  AOI21_X1 U15866 ( .B1(n12806), .B2(n12803), .A(n16239), .ZN(n16208) );
  OAI21_X1 U15867 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16220), .A(
        n16208), .ZN(n17341) );
  AOI211_X1 U15868 ( .C1(n12805), .C2(n15349), .A(n12804), .B(n17341), .ZN(
        n16196) );
  OAI211_X1 U15869 ( .C1(n14138), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17320), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16184) );
  NAND3_X1 U15870 ( .A1(n16184), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n10055), .ZN(n12808) );
  OAI21_X1 U15871 ( .B1(n15433), .B2(n17365), .A(n12810), .ZN(P1_U3000) );
  INV_X2 U15872 ( .A(n15196), .ZN(n12815) );
  NAND2_X1 U15873 ( .A1(n12563), .A2(n16549), .ZN(n12813) );
  AND2_X1 U15874 ( .A1(n12814), .A2(n12813), .ZN(n17403) );
  INV_X1 U15875 ( .A(n12816), .ZN(n17421) );
  AND2_X1 U15876 ( .A1(n12817), .A2(n16558), .ZN(n12818) );
  NOR2_X1 U15877 ( .A1(n12564), .A2(n12818), .ZN(n16555) );
  INV_X1 U15878 ( .A(n12819), .ZN(n12823) );
  NAND2_X1 U15879 ( .A1(n12823), .A2(n12820), .ZN(n12821) );
  NAND2_X1 U15880 ( .A1(n12817), .A2(n12821), .ZN(n16572) );
  INV_X1 U15881 ( .A(n16572), .ZN(n17434) );
  NAND2_X1 U15882 ( .A1(n9831), .A2(n16581), .ZN(n12822) );
  AND2_X1 U15883 ( .A1(n12823), .A2(n12822), .ZN(n17447) );
  OAI21_X1 U15884 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12824), .A(
        n9831), .ZN(n16591) );
  INV_X1 U15885 ( .A(n16591), .ZN(n17458) );
  OAI21_X1 U15886 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12825), .A(
        n9933), .ZN(n16611) );
  INV_X1 U15887 ( .A(n16611), .ZN(n17119) );
  AOI21_X1 U15888 ( .B1(n16625), .B2(n12826), .A(n12825), .ZN(n16627) );
  OAI21_X1 U15889 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12827), .A(
        n12826), .ZN(n12890) );
  INV_X1 U15890 ( .A(n12890), .ZN(n20247) );
  NAND2_X1 U15891 ( .A1(n12828), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12829) );
  INV_X1 U15892 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16649) );
  NAND2_X1 U15893 ( .A1(n12829), .A2(n16649), .ZN(n12830) );
  AND2_X1 U15894 ( .A1(n12830), .A2(n9934), .ZN(n16652) );
  XNOR2_X1 U15895 ( .A(n12828), .B(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16661) );
  INV_X1 U15896 ( .A(n16661), .ZN(n13635) );
  AOI21_X1 U15897 ( .B1(n17511), .B2(n12831), .A(n12832), .ZN(n17501) );
  AOI21_X1 U15898 ( .B1(n17530), .B2(n12833), .A(n12834), .ZN(n17524) );
  AOI21_X1 U15899 ( .B1(n20287), .B2(n12835), .A(n12836), .ZN(n20293) );
  AOI21_X1 U15900 ( .B1(n20309), .B2(n12837), .A(n12838), .ZN(n20315) );
  AOI21_X1 U15901 ( .B1(n16697), .B2(n12839), .A(n12840), .ZN(n20337) );
  AOI21_X1 U15902 ( .B1(n20373), .B2(n12841), .A(n9854), .ZN(n20366) );
  AOI21_X1 U15903 ( .B1(n17597), .B2(n12842), .A(n12843), .ZN(n17581) );
  OAI22_X1 U15904 ( .A1(n17682), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n15195) );
  INV_X1 U15905 ( .A(n15195), .ZN(n20409) );
  AOI22_X1 U15906 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16713), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17682), .ZN(n14950) );
  NOR2_X1 U15907 ( .A1(n20409), .A2(n14950), .ZN(n14949) );
  OAI21_X1 U15908 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n12842), .ZN(n14874) );
  NAND2_X1 U15909 ( .A1(n14949), .A2(n14874), .ZN(n14778) );
  NOR2_X1 U15910 ( .A1(n17581), .A2(n14778), .ZN(n20387) );
  OAI21_X1 U15911 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12843), .A(
        n12841), .ZN(n20386) );
  NAND2_X1 U15912 ( .A1(n20387), .A2(n20386), .ZN(n20364) );
  NOR2_X1 U15913 ( .A1(n20366), .A2(n20364), .ZN(n20352) );
  OAI21_X1 U15914 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9854), .A(
        n12839), .ZN(n20353) );
  NAND2_X1 U15915 ( .A1(n20352), .A2(n20353), .ZN(n20336) );
  NOR2_X1 U15916 ( .A1(n20337), .A2(n20336), .ZN(n20320) );
  OAI21_X1 U15917 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12840), .A(
        n12837), .ZN(n20321) );
  NAND2_X1 U15918 ( .A1(n20320), .A2(n20321), .ZN(n20313) );
  NOR2_X1 U15919 ( .A1(n20315), .A2(n20313), .ZN(n20303) );
  OAI21_X1 U15920 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12838), .A(
        n12835), .ZN(n20304) );
  NAND2_X1 U15921 ( .A1(n20303), .A2(n20304), .ZN(n20291) );
  NOR2_X1 U15922 ( .A1(n20293), .A2(n20291), .ZN(n20273) );
  OAI21_X1 U15923 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12836), .A(
        n12833), .ZN(n20274) );
  NAND2_X1 U15924 ( .A1(n20273), .A2(n20274), .ZN(n15042) );
  NOR2_X1 U15925 ( .A1(n17524), .A2(n15042), .ZN(n15041) );
  OAI21_X1 U15926 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12834), .A(
        n12831), .ZN(n20263) );
  NAND2_X1 U15927 ( .A1(n15041), .A2(n20263), .ZN(n13619) );
  NOR2_X1 U15928 ( .A1(n17501), .A2(n13619), .ZN(n20253) );
  INV_X1 U15929 ( .A(n12832), .ZN(n12844) );
  AOI21_X1 U15930 ( .B1(n10149), .B2(n12844), .A(n12828), .ZN(n20255) );
  INV_X1 U15931 ( .A(n20255), .ZN(n16671) );
  NAND2_X1 U15932 ( .A1(n20253), .A2(n16671), .ZN(n13634) );
  NOR2_X1 U15933 ( .A1(n13635), .A2(n13634), .ZN(n13633) );
  INV_X1 U15934 ( .A(n13633), .ZN(n12845) );
  AOI21_X1 U15935 ( .B1(n16638), .B2(n9934), .A(n12827), .ZN(n16640) );
  NOR2_X1 U15936 ( .A1(n16627), .A2(n13651), .ZN(n13650) );
  NOR2_X1 U15937 ( .A1(n17119), .A2(n17118), .ZN(n17117) );
  NOR2_X1 U15938 ( .A1(n15194), .A2(n17117), .ZN(n13664) );
  AOI21_X1 U15939 ( .B1(n16599), .B2(n9933), .A(n12824), .ZN(n16601) );
  NOR2_X1 U15940 ( .A1(n13664), .A2(n16601), .ZN(n13663) );
  NOR2_X1 U15941 ( .A1(n17458), .A2(n17457), .ZN(n17456) );
  NOR2_X1 U15942 ( .A1(n15194), .A2(n17432), .ZN(n13611) );
  NOR2_X1 U15943 ( .A1(n16555), .A2(n13611), .ZN(n13610) );
  NOR2_X1 U15944 ( .A1(n12815), .A2(n17402), .ZN(n12846) );
  XNOR2_X1 U15945 ( .A(n12846), .B(n12138), .ZN(n12867) );
  INV_X1 U15946 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n21225) );
  NAND4_X1 U15947 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21225), .A3(n17682), 
        .A4(n12132), .ZN(n21086) );
  NOR2_X1 U15948 ( .A1(n17706), .A2(n15207), .ZN(n12850) );
  INV_X1 U15949 ( .A(n12847), .ZN(n12848) );
  NAND2_X1 U15950 ( .A1(n12850), .A2(n12848), .ZN(n13784) );
  NAND2_X1 U15951 ( .A1(n12850), .A2(n12849), .ZN(n20384) );
  NAND2_X1 U15952 ( .A1(n12132), .A2(n21236), .ZN(n12858) );
  OR3_X1 U15953 ( .A1(n21239), .A2(n11789), .A3(n12858), .ZN(n20402) );
  NAND2_X1 U15954 ( .A1(n12132), .A2(n15197), .ZN(n12856) );
  OR2_X2 U15955 ( .A1(n13920), .A2(n12856), .ZN(n20401) );
  OAI22_X1 U15956 ( .A1(n13218), .A2(n20402), .B1(n20401), .B2(n15415), .ZN(
        n12851) );
  INV_X1 U15957 ( .A(n12851), .ZN(n12865) );
  NAND2_X1 U15958 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n21225), .ZN(n14020) );
  NOR2_X1 U15959 ( .A1(n12852), .A2(n14020), .ZN(n17685) );
  OR2_X1 U15960 ( .A1(n17685), .A2(n20376), .ZN(n12853) );
  NOR2_X1 U15961 ( .A1(n20370), .A2(n12853), .ZN(n12854) );
  NOR2_X2 U15962 ( .A1(n20406), .A2(n20975), .ZN(n20412) );
  AOI21_X1 U15963 ( .B1(n12132), .B2(n21236), .A(P2_EBX_REG_31__SCAN_IN), .ZN(
        n12855) );
  NOR2_X1 U15964 ( .A1(n20547), .A2(n12855), .ZN(n12857) );
  INV_X1 U15965 ( .A(n12856), .ZN(n17683) );
  INV_X1 U15966 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12862) );
  NAND2_X1 U15967 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12858), .ZN(n12859) );
  OR3_X1 U15968 ( .A1(n21239), .A2(n11789), .A3(n12859), .ZN(n20399) );
  OAI222_X1 U15969 ( .A1(n20396), .A2(n12862), .B1(n20399), .B2(n12861), .C1(
        n12860), .C2(n20374), .ZN(n12863) );
  AOI21_X1 U15970 ( .B1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20412), .A(
        n12863), .ZN(n12864) );
  OAI21_X1 U15971 ( .B1(n12867), .B2(n21086), .A(n12866), .ZN(P2_U2825) );
  OR2_X1 U15972 ( .A1(n12558), .A2(n17669), .ZN(n12868) );
  AND2_X1 U15973 ( .A1(n9864), .A2(n12869), .ZN(n12870) );
  NOR2_X1 U15974 ( .A1(n12871), .A2(n12870), .ZN(n16489) );
  INV_X1 U15975 ( .A(n16489), .ZN(n13614) );
  NAND2_X1 U15976 ( .A1(n20376), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n16556) );
  INV_X1 U15977 ( .A(n16556), .ZN(n12872) );
  AOI21_X1 U15978 ( .B1(n16718), .B2(n12882), .A(n12872), .ZN(n12873) );
  OAI21_X1 U15979 ( .B1(n17671), .B2(n13614), .A(n12873), .ZN(n12874) );
  AOI21_X1 U15980 ( .B1(n12875), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12874), .ZN(n12881) );
  XNOR2_X1 U15981 ( .A(n12876), .B(n12877), .ZN(n16554) );
  NAND2_X1 U15982 ( .A1(n12879), .A2(n12878), .ZN(n12880) );
  XNOR2_X1 U15983 ( .A(n12883), .B(n12882), .ZN(n16563) );
  NAND3_X1 U15984 ( .A1(n12885), .A2(n10330), .A3(n12884), .ZN(P2_U3019) );
  OR2_X1 U15985 ( .A1(n12887), .A2(n17566), .ZN(n12893) );
  AOI21_X1 U15986 ( .B1(n17564), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12888), .ZN(n12889) );
  OAI21_X1 U15987 ( .B1(n17571), .B2(n12890), .A(n12889), .ZN(n12891) );
  NAND2_X1 U15988 ( .A1(n13778), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U15989 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20972) );
  INV_X1 U15990 ( .A(n20972), .ZN(n21015) );
  AND2_X1 U15991 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21015), .ZN(
        n12895) );
  NAND2_X1 U15992 ( .A1(n12895), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21019) );
  INV_X1 U15993 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12896) );
  INV_X1 U15994 ( .A(n12895), .ZN(n12908) );
  NAND2_X1 U15995 ( .A1(n12896), .A2(n12908), .ZN(n12897) );
  AND3_X1 U15996 ( .A1(n21019), .A2(n21177), .A3(n12897), .ZN(n20900) );
  AOI21_X1 U15997 ( .B1(n12920), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n20900), .ZN(n12903) );
  INV_X1 U15998 ( .A(n12903), .ZN(n12930) );
  NOR2_X1 U15999 ( .A1(n13778), .A2(n17682), .ZN(n12898) );
  NOR2_X1 U16000 ( .A1(n13160), .A2(n12899), .ZN(n12901) );
  NAND2_X1 U16001 ( .A1(n12930), .A2(n12901), .ZN(n14353) );
  INV_X1 U16002 ( .A(n12901), .ZN(n12902) );
  AND2_X1 U16003 ( .A1(n12903), .A2(n12902), .ZN(n12904) );
  NAND2_X1 U16004 ( .A1(n12905), .A2(n12904), .ZN(n12906) );
  NAND2_X1 U16005 ( .A1(n12907), .A2(n14011), .ZN(n12911) );
  NAND2_X1 U16006 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n14649) );
  NAND2_X1 U16007 ( .A1(n14649), .A2(n21194), .ZN(n12909) );
  AND2_X1 U16008 ( .A1(n12909), .A2(n12908), .ZN(n20669) );
  AOI22_X1 U16009 ( .A1(n12920), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21177), .B2(n20669), .ZN(n12910) );
  NAND2_X1 U16010 ( .A1(n12911), .A2(n12910), .ZN(n12914) );
  INV_X1 U16011 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12912) );
  NOR2_X1 U16012 ( .A1(n13160), .A2(n12912), .ZN(n12913) );
  NAND2_X1 U16013 ( .A1(n12914), .A2(n12913), .ZN(n12927) );
  AOI22_X1 U16014 ( .A1(n12920), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n21177), .B2(n21212), .ZN(n12917) );
  NAND2_X1 U16015 ( .A1(n12920), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12921) );
  NAND2_X1 U16016 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21203), .ZN(
        n20797) );
  NAND2_X1 U16017 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21212), .ZN(
        n20833) );
  NAND2_X1 U16018 ( .A1(n20797), .A2(n20833), .ZN(n20667) );
  NAND2_X1 U16019 ( .A1(n21177), .A2(n20667), .ZN(n20836) );
  NAND2_X1 U16020 ( .A1(n12921), .A2(n20836), .ZN(n12922) );
  INV_X1 U16021 ( .A(n12924), .ZN(n12925) );
  NOR2_X1 U16022 ( .A1(n16932), .A2(n12925), .ZN(n12926) );
  NAND2_X1 U16023 ( .A1(n13897), .A2(n13898), .ZN(n12928) );
  NAND2_X1 U16024 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13778), .ZN(
        n12929) );
  AND2_X1 U16025 ( .A1(n12930), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12932) );
  INV_X1 U16026 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12931) );
  NOR2_X1 U16027 ( .A1(n13160), .A2(n12931), .ZN(n14351) );
  NAND2_X1 U16028 ( .A1(n12934), .A2(n12933), .ZN(n20416) );
  AOI22_X1 U16029 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U16030 ( .A1(n12321), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12322), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U16031 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U16032 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12935) );
  NAND4_X1 U16033 ( .A1(n12938), .A2(n12937), .A3(n12936), .A4(n12935), .ZN(
        n12947) );
  AOI22_X1 U16034 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12945) );
  INV_X1 U16035 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n20750) );
  NAND2_X1 U16036 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12940) );
  NAND2_X1 U16037 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12939) );
  OAI211_X1 U16038 ( .C1(n13067), .C2(n20750), .A(n12940), .B(n12939), .ZN(
        n12941) );
  INV_X1 U16039 ( .A(n12941), .ZN(n12944) );
  AOI22_X1 U16040 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12943) );
  NAND2_X1 U16041 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12942) );
  NAND4_X1 U16042 ( .A1(n12945), .A2(n12944), .A3(n12943), .A4(n12942), .ZN(
        n12946) );
  NOR2_X1 U16043 ( .A1(n12947), .A2(n12946), .ZN(n20417) );
  AOI22_X1 U16044 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U16045 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U16046 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U16047 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12948) );
  NAND4_X1 U16048 ( .A1(n12951), .A2(n12950), .A3(n12949), .A4(n12948), .ZN(
        n12961) );
  AOI22_X1 U16049 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n11856), .ZN(n12959) );
  NAND2_X1 U16050 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12953) );
  NAND2_X1 U16051 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12952) );
  OAI211_X1 U16052 ( .C1(n13067), .C2(n12954), .A(n12953), .B(n12952), .ZN(
        n12955) );
  INV_X1 U16053 ( .A(n12955), .ZN(n12958) );
  AOI22_X1 U16054 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12957) );
  NAND2_X1 U16055 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12956) );
  NAND4_X1 U16056 ( .A1(n12959), .A2(n12958), .A3(n12957), .A4(n12956), .ZN(
        n12960) );
  OR2_X1 U16057 ( .A1(n12961), .A2(n12960), .ZN(n15212) );
  AOI22_X1 U16058 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U16059 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U16060 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16061 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12962) );
  NAND4_X1 U16062 ( .A1(n12965), .A2(n12964), .A3(n12963), .A4(n12962), .ZN(
        n12975) );
  AOI22_X1 U16063 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n11856), .ZN(n12973) );
  INV_X1 U16064 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12968) );
  NAND2_X1 U16065 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12967) );
  NAND2_X1 U16066 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12966) );
  OAI211_X1 U16067 ( .C1(n13067), .C2(n12968), .A(n12967), .B(n12966), .ZN(
        n12969) );
  INV_X1 U16068 ( .A(n12969), .ZN(n12972) );
  AOI22_X1 U16069 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12971) );
  NAND2_X1 U16070 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12970) );
  NAND4_X1 U16071 ( .A1(n12973), .A2(n12972), .A3(n12971), .A4(n12970), .ZN(
        n12974) );
  OR2_X1 U16072 ( .A1(n12975), .A2(n12974), .ZN(n17477) );
  AOI22_X1 U16073 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12979) );
  AOI22_X1 U16074 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12978) );
  AOI22_X1 U16075 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12977) );
  AOI22_X1 U16076 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12976) );
  NAND4_X1 U16077 ( .A1(n12979), .A2(n12978), .A3(n12977), .A4(n12976), .ZN(
        n12989) );
  AOI22_X1 U16078 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n11856), .ZN(n12987) );
  NAND2_X1 U16079 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12981) );
  NAND2_X1 U16080 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12980) );
  OAI211_X1 U16081 ( .C1(n13067), .C2(n12982), .A(n12981), .B(n12980), .ZN(
        n12983) );
  INV_X1 U16082 ( .A(n12983), .ZN(n12986) );
  AOI22_X1 U16083 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12985) );
  NAND2_X1 U16084 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12984) );
  NAND4_X1 U16085 ( .A1(n12987), .A2(n12986), .A3(n12985), .A4(n12984), .ZN(
        n12988) );
  NOR2_X1 U16086 ( .A1(n12989), .A2(n12988), .ZN(n16462) );
  AOI22_X1 U16087 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16088 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16089 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16090 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12990) );
  NAND4_X1 U16091 ( .A1(n12993), .A2(n12992), .A3(n12991), .A4(n12990), .ZN(
        n13003) );
  AOI22_X1 U16092 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n11856), .ZN(n13001) );
  INV_X1 U16093 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U16094 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12995) );
  NAND2_X1 U16095 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12994) );
  OAI211_X1 U16096 ( .C1(n13067), .C2(n12996), .A(n12995), .B(n12994), .ZN(
        n12997) );
  INV_X1 U16097 ( .A(n12997), .ZN(n13000) );
  AOI22_X1 U16098 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16099 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12998) );
  NAND4_X1 U16100 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        n13002) );
  NOR2_X1 U16101 ( .A1(n13003), .A2(n13002), .ZN(n17474) );
  INV_X1 U16102 ( .A(n17474), .ZN(n13004) );
  AOI22_X1 U16103 ( .A1(n11736), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U16104 ( .A1(n12321), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12322), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U16105 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U16106 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13005) );
  NAND4_X1 U16107 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13017) );
  AOI22_X1 U16108 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13015) );
  NAND2_X1 U16109 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13010) );
  NAND2_X1 U16110 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13009) );
  OAI211_X1 U16111 ( .C1(n13067), .C2(n11708), .A(n13010), .B(n13009), .ZN(
        n13011) );
  INV_X1 U16112 ( .A(n13011), .ZN(n13014) );
  AOI22_X1 U16113 ( .A1(n13069), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U16114 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13012) );
  NAND4_X1 U16115 ( .A1(n13015), .A2(n13014), .A3(n13013), .A4(n13012), .ZN(
        n13016) );
  OR2_X1 U16116 ( .A1(n13017), .A2(n13016), .ZN(n16456) );
  NAND2_X1 U16117 ( .A1(n16454), .A2(n16456), .ZN(n16452) );
  AOI22_X1 U16118 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11736), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U16119 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12322), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16120 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11767), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U16121 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13019) );
  NAND4_X1 U16122 ( .A1(n13022), .A2(n13021), .A3(n13020), .A4(n13019), .ZN(
        n13036) );
  OAI22_X1 U16123 ( .A1(n13026), .A2(n13025), .B1(n13024), .B2(n13023), .ZN(
        n13035) );
  OAI22_X1 U16124 ( .A1(n13030), .A2(n13029), .B1(n13028), .B2(n13027), .ZN(
        n13034) );
  NAND2_X1 U16125 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n13032) );
  AOI22_X1 U16126 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n13063), .ZN(n13031) );
  OAI211_X1 U16127 ( .C1(n13067), .C2(n14027), .A(n13032), .B(n13031), .ZN(
        n13033) );
  NOR4_X1 U16128 ( .A1(n13036), .A2(n13035), .A3(n13034), .A4(n13033), .ZN(
        n17470) );
  NOR2_X2 U16129 ( .A1(n16452), .A2(n17470), .ZN(n13077) );
  AOI22_X1 U16130 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U16131 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9819), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13048) );
  INV_X1 U16132 ( .A(n13041), .ZN(n16939) );
  AOI22_X1 U16133 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13047) );
  NAND2_X1 U16134 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13045) );
  NAND2_X1 U16135 ( .A1(n9791), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13044) );
  OAI21_X1 U16136 ( .B1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n13043), .ZN(n13206) );
  AND3_X1 U16137 ( .A1(n13045), .A2(n13044), .A3(n13206), .ZN(n13046) );
  NAND4_X1 U16138 ( .A1(n13049), .A2(n13048), .A3(n13047), .A4(n13046), .ZN(
        n13057) );
  AOI22_X1 U16139 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16140 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9819), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16141 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13053) );
  NAND2_X1 U16142 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13051) );
  NAND2_X1 U16143 ( .A1(n9791), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13050) );
  INV_X1 U16144 ( .A(n13206), .ZN(n13185) );
  AND3_X1 U16145 ( .A1(n13051), .A2(n13050), .A3(n13185), .ZN(n13052) );
  NAND4_X1 U16146 ( .A1(n13055), .A2(n13054), .A3(n13053), .A4(n13052), .ZN(
        n13056) );
  NAND2_X1 U16147 ( .A1(n13057), .A2(n13056), .ZN(n13098) );
  NOR2_X1 U16148 ( .A1(n20547), .A2(n13098), .ZN(n13076) );
  AOI22_X1 U16149 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n11736), .B1(
        n12321), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U16150 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11767), .B1(
        n12322), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U16151 ( .A1(n13018), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11753), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U16152 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11672), .B1(
        n13058), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13059) );
  NAND4_X1 U16153 ( .A1(n13062), .A2(n13061), .A3(n13060), .A4(n13059), .ZN(
        n13075) );
  AOI22_X1 U16154 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n11856), .ZN(n13073) );
  INV_X1 U16155 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13066) );
  NAND2_X1 U16156 ( .A1(n11650), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13065) );
  NAND2_X1 U16157 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13064) );
  OAI211_X1 U16158 ( .C1(n13067), .C2(n13066), .A(n13065), .B(n13064), .ZN(
        n13068) );
  INV_X1 U16159 ( .A(n13068), .ZN(n13072) );
  AOI22_X1 U16160 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13069), .B1(
        n12329), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13071) );
  NAND2_X1 U16161 ( .A1(n11681), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13070) );
  NAND4_X1 U16162 ( .A1(n13073), .A2(n13072), .A3(n13071), .A4(n13070), .ZN(
        n13074) );
  NOR2_X1 U16163 ( .A1(n13075), .A2(n13074), .ZN(n13093) );
  XNOR2_X1 U16164 ( .A(n13076), .B(n13093), .ZN(n13100) );
  INV_X1 U16165 ( .A(n13098), .ZN(n13094) );
  NAND2_X1 U16166 ( .A1(n20547), .A2(n13094), .ZN(n16521) );
  AOI22_X1 U16168 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U16169 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11607), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U16170 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13082) );
  NAND2_X1 U16171 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13080) );
  NAND2_X1 U16172 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13079) );
  AND3_X1 U16173 ( .A1(n13080), .A2(n13079), .A3(n13206), .ZN(n13081) );
  NAND4_X1 U16174 ( .A1(n13084), .A2(n13083), .A3(n13082), .A4(n13081), .ZN(
        n13092) );
  AOI22_X1 U16175 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16176 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U16177 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13088) );
  NAND2_X1 U16178 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13086) );
  NAND2_X1 U16179 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13085) );
  AND3_X1 U16180 ( .A1(n13086), .A2(n13085), .A3(n13185), .ZN(n13087) );
  NAND4_X1 U16181 ( .A1(n13090), .A2(n13089), .A3(n13088), .A4(n13087), .ZN(
        n13091) );
  NAND2_X1 U16182 ( .A1(n13092), .A2(n13091), .ZN(n13102) );
  INV_X1 U16183 ( .A(n13093), .ZN(n13095) );
  NAND2_X1 U16184 ( .A1(n13095), .A2(n13094), .ZN(n13103) );
  XOR2_X1 U16185 ( .A(n13102), .B(n13103), .Z(n13096) );
  INV_X1 U16186 ( .A(n13160), .ZN(n13118) );
  NAND2_X1 U16187 ( .A1(n13096), .A2(n13118), .ZN(n16443) );
  INV_X1 U16188 ( .A(n13102), .ZN(n13097) );
  NAND2_X1 U16189 ( .A1(n20547), .A2(n13097), .ZN(n16445) );
  NOR2_X1 U16190 ( .A1(n16445), .A2(n13098), .ZN(n13099) );
  NOR2_X1 U16191 ( .A1(n13103), .A2(n13102), .ZN(n13119) );
  AOI22_X1 U16192 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U16193 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9820), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13108) );
  AOI22_X1 U16194 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13107) );
  NAND2_X1 U16195 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13105) );
  NAND2_X1 U16196 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13104) );
  AND3_X1 U16197 ( .A1(n13105), .A2(n13104), .A3(n13206), .ZN(n13106) );
  NAND4_X1 U16198 ( .A1(n13109), .A2(n13108), .A3(n13107), .A4(n13106), .ZN(
        n13117) );
  AOI22_X1 U16199 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U16200 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16201 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13113) );
  NAND2_X1 U16202 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13111) );
  NAND2_X1 U16203 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13110) );
  AND3_X1 U16204 ( .A1(n13111), .A2(n13110), .A3(n13185), .ZN(n13112) );
  NAND4_X1 U16205 ( .A1(n13115), .A2(n13114), .A3(n13113), .A4(n13112), .ZN(
        n13116) );
  AND2_X1 U16206 ( .A1(n13117), .A2(n13116), .ZN(n13121) );
  NAND2_X1 U16207 ( .A1(n13119), .A2(n13121), .ZN(n13140) );
  OAI211_X1 U16208 ( .C1(n13119), .C2(n13121), .A(n13140), .B(n13118), .ZN(
        n13124) );
  INV_X1 U16209 ( .A(n13124), .ZN(n13120) );
  XNOR2_X1 U16210 ( .A(n13123), .B(n13120), .ZN(n16432) );
  INV_X1 U16211 ( .A(n13121), .ZN(n13122) );
  NOR2_X1 U16212 ( .A1(n11624), .A2(n13122), .ZN(n16434) );
  NAND2_X1 U16213 ( .A1(n16432), .A2(n16434), .ZN(n16433) );
  AOI22_X1 U16214 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16215 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U16216 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U16217 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13127) );
  NAND2_X1 U16218 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13126) );
  AND3_X1 U16219 ( .A1(n13127), .A2(n13126), .A3(n13206), .ZN(n13128) );
  NAND4_X1 U16220 ( .A1(n13131), .A2(n13130), .A3(n13129), .A4(n13128), .ZN(
        n13139) );
  AOI22_X1 U16221 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16222 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9821), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U16223 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13135) );
  NAND2_X1 U16224 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13133) );
  NAND2_X1 U16225 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13132) );
  AND3_X1 U16226 ( .A1(n13133), .A2(n13132), .A3(n13185), .ZN(n13134) );
  NAND4_X1 U16227 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        n13138) );
  NAND2_X1 U16228 ( .A1(n13139), .A2(n13138), .ZN(n13142) );
  AOI21_X1 U16229 ( .B1(n13140), .B2(n13142), .A(n13160), .ZN(n13141) );
  OR2_X1 U16230 ( .A1(n13140), .A2(n13142), .ZN(n13161) );
  NAND2_X1 U16231 ( .A1(n13141), .A2(n13161), .ZN(n13144) );
  NOR2_X1 U16232 ( .A1(n11624), .A2(n13142), .ZN(n16426) );
  INV_X1 U16233 ( .A(n13143), .ZN(n13145) );
  AOI22_X1 U16234 ( .A1(n9824), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9811), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13151) );
  AOI22_X1 U16235 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9819), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U16236 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U16237 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13147) );
  NAND2_X1 U16238 ( .A1(n9791), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13146) );
  AND3_X1 U16239 ( .A1(n13147), .A2(n13146), .A3(n13206), .ZN(n13148) );
  NAND4_X1 U16240 ( .A1(n13151), .A2(n13150), .A3(n13149), .A4(n13148), .ZN(
        n13159) );
  AOI22_X1 U16241 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16242 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13156) );
  INV_X1 U16243 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20957) );
  AOI22_X1 U16244 ( .A1(n9811), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9812), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13155) );
  INV_X1 U16245 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20887) );
  NAND2_X1 U16246 ( .A1(n16939), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13153) );
  NAND2_X1 U16247 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13152) );
  AND3_X1 U16248 ( .A1(n13153), .A2(n13152), .A3(n13185), .ZN(n13154) );
  NAND4_X1 U16249 ( .A1(n13157), .A2(n13156), .A3(n13155), .A4(n13154), .ZN(
        n13158) );
  NAND2_X1 U16250 ( .A1(n13159), .A2(n13158), .ZN(n13164) );
  NOR2_X1 U16251 ( .A1(n13161), .A2(n13164), .ZN(n16413) );
  NAND2_X1 U16252 ( .A1(n13163), .A2(n13162), .ZN(n16412) );
  NOR2_X1 U16253 ( .A1(n9829), .A2(n13164), .ZN(n16421) );
  AOI22_X1 U16254 ( .A1(n9824), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n9811), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13170) );
  AOI22_X1 U16255 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9820), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13169) );
  AOI22_X1 U16256 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13168) );
  NAND2_X1 U16257 ( .A1(n9812), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13166) );
  NAND2_X1 U16258 ( .A1(n9819), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13165) );
  AND3_X1 U16259 ( .A1(n13166), .A2(n13165), .A3(n13206), .ZN(n13167) );
  NAND4_X1 U16260 ( .A1(n13170), .A2(n13169), .A3(n13168), .A4(n13167), .ZN(
        n13178) );
  AOI22_X1 U16261 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13176) );
  AOI22_X1 U16262 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11607), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16263 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13174) );
  NAND2_X1 U16264 ( .A1(n13042), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13172) );
  NAND2_X1 U16265 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13171) );
  AND3_X1 U16266 ( .A1(n13172), .A2(n13171), .A3(n13185), .ZN(n13173) );
  NAND4_X1 U16267 ( .A1(n13176), .A2(n13175), .A3(n13174), .A4(n13173), .ZN(
        n13177) );
  NAND2_X1 U16268 ( .A1(n13178), .A2(n13177), .ZN(n16415) );
  AOI22_X1 U16269 ( .A1(n13037), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9811), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13184) );
  AOI22_X1 U16270 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9819), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13183) );
  AOI22_X1 U16271 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U16272 ( .A1(n9812), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13180) );
  NAND2_X1 U16273 ( .A1(n9821), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13179) );
  AND3_X1 U16274 ( .A1(n13180), .A2(n13179), .A3(n13206), .ZN(n13181) );
  NAND4_X1 U16275 ( .A1(n13184), .A2(n13183), .A3(n13182), .A4(n13181), .ZN(
        n13193) );
  AOI22_X1 U16276 ( .A1(n9824), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9811), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U16277 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9819), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U16278 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16939), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13189) );
  NAND2_X1 U16279 ( .A1(n9813), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13187) );
  NAND2_X1 U16280 ( .A1(n9791), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n13186) );
  AND3_X1 U16281 ( .A1(n13187), .A2(n13186), .A3(n13185), .ZN(n13188) );
  NAND4_X1 U16282 ( .A1(n13191), .A2(n13190), .A3(n13189), .A4(n13188), .ZN(
        n13192) );
  NAND2_X1 U16283 ( .A1(n13193), .A2(n13192), .ZN(n13196) );
  NOR2_X1 U16284 ( .A1(n20547), .A2(n16415), .ZN(n13194) );
  NAND2_X1 U16285 ( .A1(n16413), .A2(n13194), .ZN(n13195) );
  NOR2_X1 U16286 ( .A1(n13195), .A2(n13196), .ZN(n13197) );
  AOI21_X1 U16287 ( .B1(n13196), .B2(n13195), .A(n13197), .ZN(n16407) );
  NAND2_X1 U16288 ( .A1(n16408), .A2(n16407), .ZN(n16409) );
  INV_X1 U16289 ( .A(n13197), .ZN(n13198) );
  NAND2_X1 U16290 ( .A1(n16409), .A2(n13198), .ZN(n13215) );
  AOI22_X1 U16291 ( .A1(n9824), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9811), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13200) );
  AOI22_X1 U16292 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9791), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13199) );
  NAND2_X1 U16293 ( .A1(n13200), .A2(n13199), .ZN(n13213) );
  INV_X1 U16294 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n20898) );
  AOI22_X1 U16295 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9812), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13202) );
  AOI21_X1 U16296 ( .B1(n9819), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n13206), .ZN(n13201) );
  OAI211_X1 U16297 ( .C1(n13041), .C2(n20898), .A(n13202), .B(n13201), .ZN(
        n13212) );
  AOI22_X1 U16298 ( .A1(n9824), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9811), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U16299 ( .A1(n13203), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9819), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U16300 ( .A1(n13205), .A2(n13204), .ZN(n13211) );
  AOI22_X1 U16301 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13042), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13209) );
  NAND2_X1 U16302 ( .A1(n9791), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13208) );
  NAND2_X1 U16303 ( .A1(n16939), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n13207) );
  NAND4_X1 U16304 ( .A1(n13209), .A2(n13208), .A3(n13207), .A4(n13206), .ZN(
        n13210) );
  XNOR2_X1 U16305 ( .A(n13215), .B(n13214), .ZN(n15417) );
  INV_X1 U16306 ( .A(n17709), .ZN(n17705) );
  NAND2_X1 U16307 ( .A1(n17705), .A2(n17708), .ZN(n15203) );
  OR2_X1 U16308 ( .A1(n16964), .A2(n11502), .ZN(n16952) );
  AOI21_X2 U16309 ( .B1(n15203), .B2(n16952), .A(n15207), .ZN(n13216) );
  NAND2_X1 U16310 ( .A1(n15417), .A2(n20435), .ZN(n13221) );
  NAND2_X1 U16311 ( .A1(n17479), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13217) );
  INV_X1 U16312 ( .A(n13219), .ZN(n13220) );
  NAND2_X1 U16313 ( .A1(n13221), .A2(n13220), .ZN(P2_U2857) );
  INV_X1 U16314 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U16315 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13237) );
  AOI22_X1 U16316 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13236) );
  NOR2_X2 U16317 ( .A1(n18256), .A2(n13228), .ZN(n13259) );
  INV_X4 U16318 ( .A(n13298), .ZN(n18539) );
  INV_X1 U16319 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18454) );
  AOI22_X1 U16320 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13222) );
  OAI21_X1 U16321 ( .B1(n18454), .B2(n9787), .A(n13222), .ZN(n13234) );
  AOI22_X1 U16322 ( .A1(n18473), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13232) );
  AOI22_X1 U16323 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n9794), .B1(
        n18472), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13231) );
  AOI22_X1 U16324 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13230) );
  AOI22_X1 U16325 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13229) );
  NAND4_X1 U16326 ( .A1(n13232), .A2(n13231), .A3(n13230), .A4(n13229), .ZN(
        n13233) );
  AOI211_X1 U16327 ( .C1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .C2(n18539), .A(
        n13234), .B(n13233), .ZN(n13235) );
  NAND3_X1 U16328 ( .A1(n13237), .A2(n13236), .A3(n13235), .ZN(n13499) );
  INV_X2 U16329 ( .A(n9787), .ZN(n17066) );
  AOI22_X1 U16330 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13241) );
  AOI22_X1 U16331 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13240) );
  AOI22_X1 U16332 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U16333 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18534), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13238) );
  NAND4_X1 U16334 ( .A1(n13241), .A2(n13240), .A3(n13239), .A4(n13238), .ZN(
        n13247) );
  AOI22_X1 U16335 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U16336 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16337 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n9795), .B1(n9817), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U16338 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13242) );
  NAND4_X1 U16339 ( .A1(n13245), .A2(n13244), .A3(n13243), .A4(n13242), .ZN(
        n13246) );
  AOI22_X1 U16340 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13251) );
  AOI22_X1 U16341 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U16342 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13249) );
  AOI22_X1 U16343 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13248) );
  NAND4_X1 U16344 ( .A1(n13251), .A2(n13250), .A3(n13249), .A4(n13248), .ZN(
        n13257) );
  AOI22_X1 U16345 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13255) );
  AOI22_X1 U16346 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13254) );
  INV_X1 U16347 ( .A(n13258), .ZN(n17029) );
  INV_X2 U16348 ( .A(n17029), .ZN(n18503) );
  AOI22_X1 U16349 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18503), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13253) );
  AOI22_X1 U16350 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n9794), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13252) );
  NAND4_X1 U16351 ( .A1(n13255), .A2(n13254), .A3(n13253), .A4(n13252), .ZN(
        n13256) );
  AOI22_X1 U16352 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13263) );
  AOI22_X1 U16353 ( .A1(n13296), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13310), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U16354 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13258), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13261) );
  AOI22_X1 U16355 ( .A1(n13259), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13260) );
  AOI22_X1 U16356 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13272) );
  AOI22_X1 U16357 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13295), .B1(
        n13264), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13265) );
  INV_X1 U16358 ( .A(n13265), .ZN(n13267) );
  INV_X1 U16359 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17030) );
  OAI21_X1 U16360 ( .B1(n17030), .B2(n9862), .A(n13268), .ZN(n13269) );
  INV_X1 U16361 ( .A(n13269), .ZN(n13270) );
  NAND4_X1 U16362 ( .A1(n9869), .A2(n13272), .A3(n13271), .A4(n13270), .ZN(
        n18721) );
  INV_X1 U16363 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U16364 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13273) );
  AOI22_X1 U16365 ( .A1(n13310), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18473), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13279) );
  AOI22_X1 U16366 ( .A1(n13296), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U16367 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U16368 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13276) );
  AOI22_X1 U16369 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13280) );
  INV_X1 U16370 ( .A(n13280), .ZN(n13283) );
  AOI22_X1 U16371 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13281) );
  NAND2_X1 U16372 ( .A1(n18721), .A2(n13497), .ZN(n13509) );
  AOI22_X1 U16373 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18503), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13294) );
  AOI22_X1 U16374 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n17066), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U16375 ( .A1(n13259), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13285) );
  OAI21_X1 U16376 ( .B1(n15955), .B2(n9862), .A(n13285), .ZN(n13291) );
  AOI22_X1 U16377 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13289) );
  AOI22_X1 U16378 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9794), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13288) );
  AOI22_X1 U16379 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U16380 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18534), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13286) );
  NAND4_X1 U16381 ( .A1(n13289), .A2(n13288), .A3(n13287), .A4(n13286), .ZN(
        n13290) );
  AOI211_X1 U16382 ( .C1(n18519), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n13291), .B(n13290), .ZN(n13292) );
  NAND3_X1 U16383 ( .A1(n13294), .A2(n13293), .A3(n13292), .ZN(n13498) );
  NAND2_X1 U16384 ( .A1(n13329), .A2(n13498), .ZN(n13332) );
  AOI22_X1 U16385 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13307) );
  AOI22_X1 U16386 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13306) );
  INV_X1 U16387 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15976) );
  AOI22_X1 U16388 ( .A1(n18520), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13297) );
  OAI21_X1 U16389 ( .B1(n15976), .B2(n13298), .A(n13297), .ZN(n13304) );
  AOI22_X1 U16390 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U16391 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9794), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U16392 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U16393 ( .A1(n18534), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13299) );
  NAND4_X1 U16394 ( .A1(n13302), .A2(n13301), .A3(n13300), .A4(n13299), .ZN(
        n13303) );
  AOI211_X1 U16395 ( .C1(n9817), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n13304), .B(n13303), .ZN(n13305) );
  NAND3_X1 U16396 ( .A1(n13307), .A2(n13306), .A3(n13305), .ZN(n18698) );
  INV_X1 U16397 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19240) );
  XOR2_X1 U16398 ( .A(n13308), .B(n13499), .Z(n13336) );
  INV_X1 U16399 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19468) );
  NOR2_X1 U16400 ( .A1(n13336), .A2(n19468), .ZN(n13337) );
  INV_X1 U16401 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19507) );
  NOR2_X1 U16402 ( .A1(n19507), .A2(n13309), .ZN(n13325) );
  XNOR2_X1 U16403 ( .A(n19507), .B(n13309), .ZN(n19190) );
  AOI22_X1 U16404 ( .A1(n18519), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U16405 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13322) );
  AOI22_X1 U16406 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13312) );
  OAI21_X1 U16407 ( .B1(n13389), .B2(n18426), .A(n13312), .ZN(n13320) );
  AOI22_X1 U16408 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U16409 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U16410 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9794), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U16411 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13315) );
  NAND4_X1 U16412 ( .A1(n13318), .A2(n13317), .A3(n13316), .A4(n13315), .ZN(
        n13319) );
  AOI211_X1 U16413 ( .C1(n18472), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n13320), .B(n13319), .ZN(n13321) );
  AND2_X1 U16414 ( .A1(n13496), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13324) );
  NOR2_X1 U16415 ( .A1(n19190), .A2(n19191), .ZN(n19189) );
  NOR2_X2 U16416 ( .A1(n13325), .A2(n19189), .ZN(n13327) );
  XNOR2_X1 U16417 ( .A(n13509), .B(n18712), .ZN(n13326) );
  NOR2_X1 U16418 ( .A1(n13327), .A2(n13326), .ZN(n13328) );
  INV_X1 U16419 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19496) );
  INV_X1 U16420 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19488) );
  INV_X1 U16421 ( .A(n13498), .ZN(n18709) );
  XOR2_X1 U16422 ( .A(n18709), .B(n13329), .Z(n13330) );
  XNOR2_X1 U16423 ( .A(n19488), .B(n13330), .ZN(n19172) );
  NOR2_X1 U16424 ( .A1(n19488), .A2(n13330), .ZN(n13331) );
  XNOR2_X1 U16425 ( .A(n13332), .B(n18706), .ZN(n13333) );
  NOR2_X1 U16426 ( .A1(n13334), .A2(n13333), .ZN(n13335) );
  INV_X1 U16427 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n19480) );
  XNOR2_X1 U16428 ( .A(n13336), .B(n19468), .ZN(n19147) );
  OAI21_X1 U16429 ( .B1(n13338), .B2(n18698), .A(n19119), .ZN(n13340) );
  NOR2_X1 U16430 ( .A1(n13339), .A2(n13340), .ZN(n13341) );
  INV_X1 U16431 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19456) );
  INV_X1 U16432 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n19449) );
  NOR2_X1 U16433 ( .A1(n19008), .A2(n19026), .ZN(n19057) );
  INV_X1 U16434 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n19385) );
  INV_X1 U16435 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n19369) );
  INV_X1 U16436 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19078) );
  INV_X1 U16437 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19351) );
  NOR2_X1 U16438 ( .A1(n19057), .A2(n13345), .ZN(n13348) );
  NOR2_X2 U16439 ( .A1(n9866), .A2(n19449), .ZN(n19116) );
  NOR2_X1 U16440 ( .A1(n13343), .A2(n13342), .ZN(n19412) );
  NAND2_X1 U16441 ( .A1(n19412), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19392) );
  NOR2_X1 U16442 ( .A1(n19392), .A2(n19078), .ZN(n19361) );
  NAND2_X1 U16443 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19361), .ZN(
        n19366) );
  INV_X1 U16444 ( .A(n19366), .ZN(n19363) );
  NAND2_X1 U16445 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19363), .ZN(
        n19349) );
  NOR2_X1 U16446 ( .A1(n19351), .A2(n19349), .ZN(n17100) );
  INV_X1 U16447 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n19341) );
  INV_X1 U16448 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19333) );
  NAND2_X1 U16449 ( .A1(n18998), .A2(n19333), .ZN(n18997) );
  NAND2_X1 U16450 ( .A1(n13348), .A2(n13347), .ZN(n19007) );
  NAND2_X1 U16451 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19318) );
  INV_X1 U16452 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18983) );
  INV_X1 U16453 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18961) );
  NOR2_X1 U16454 ( .A1(n18983), .A2(n18961), .ZN(n19280) );
  NAND3_X1 U16455 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n19280), .ZN(n18929) );
  NOR2_X1 U16456 ( .A1(n19318), .A2(n18929), .ZN(n18926) );
  NAND2_X1 U16457 ( .A1(n18926), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17099) );
  INV_X1 U16458 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18924) );
  NOR2_X1 U16459 ( .A1(n17099), .A2(n18924), .ZN(n18900) );
  NOR2_X1 U16460 ( .A1(n19008), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18991) );
  NAND2_X1 U16461 ( .A1(n18991), .A2(n18983), .ZN(n13349) );
  NOR2_X1 U16462 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13349), .ZN(
        n18949) );
  INV_X1 U16463 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n19296) );
  NAND2_X1 U16464 ( .A1(n18949), .A2(n19296), .ZN(n18928) );
  NOR3_X1 U16465 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n18928), .ZN(n13350) );
  INV_X1 U16466 ( .A(n13351), .ZN(n13352) );
  INV_X1 U16467 ( .A(n19318), .ZN(n18959) );
  NAND2_X1 U16468 ( .A1(n18959), .A2(n19007), .ZN(n18947) );
  INV_X1 U16469 ( .A(n18929), .ZN(n17783) );
  NAND2_X1 U16470 ( .A1(n17783), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17098) );
  INV_X1 U16471 ( .A(n17098), .ZN(n13353) );
  NAND2_X1 U16472 ( .A1(n19119), .A2(n18896), .ZN(n13354) );
  NOR2_X1 U16473 ( .A1(n13355), .A2(n19119), .ZN(n18895) );
  NAND2_X1 U16474 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19221) );
  INV_X1 U16475 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17758) );
  NAND2_X1 U16476 ( .A1(n17111), .A2(n17758), .ZN(n17176) );
  NAND2_X1 U16477 ( .A1(n19119), .A2(n17176), .ZN(n13363) );
  NAND2_X1 U16478 ( .A1(n19008), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13361) );
  NOR2_X2 U16479 ( .A1(n18863), .A2(n13361), .ZN(n17112) );
  NAND2_X1 U16480 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17112), .ZN(
        n17177) );
  AOI22_X1 U16481 ( .A1(n13363), .A2(n17751), .B1(n17177), .B2(n19008), .ZN(
        n13362) );
  INV_X1 U16482 ( .A(n13362), .ZN(n13367) );
  INV_X1 U16483 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20165) );
  AOI22_X1 U16484 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n19008), .B1(
        n19119), .B2(n20165), .ZN(n13366) );
  OAI211_X1 U16485 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17751), .A(
        n17177), .B(n13363), .ZN(n13365) );
  NOR2_X1 U16486 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n20165), .ZN(
        n17773) );
  NOR2_X1 U16487 ( .A1(n13366), .A2(n17773), .ZN(n13364) );
  AOI22_X2 U16488 ( .A1(n13367), .A2(n13366), .B1(n13365), .B2(n13364), .ZN(
        n17775) );
  AOI22_X1 U16489 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13371) );
  AOI22_X1 U16490 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18518), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13370) );
  AOI22_X1 U16491 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18472), .B1(
        n18503), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13369) );
  AOI22_X1 U16492 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13368) );
  NAND4_X1 U16493 ( .A1(n13371), .A2(n13370), .A3(n13369), .A4(n13368), .ZN(
        n13377) );
  AOI22_X1 U16494 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13375) );
  AOI22_X1 U16495 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U16496 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18473), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U16497 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13372) );
  NAND4_X1 U16498 ( .A1(n13375), .A2(n13374), .A3(n13373), .A4(n13372), .ZN(
        n13376) );
  NAND2_X1 U16499 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20164), .ZN(n20049) );
  AOI22_X1 U16500 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n20021), .B2(n20177), .ZN(
        n13482) );
  AOI22_X1 U16501 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20169), .B1(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20026), .ZN(n13387) );
  NAND2_X1 U16502 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20019), .ZN(
        n13483) );
  NAND2_X1 U16503 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20021), .ZN(
        n13378) );
  AOI22_X1 U16504 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20177), .B1(
        n13483), .B2(n13378), .ZN(n13386) );
  NAND2_X1 U16505 ( .A1(n13387), .A2(n13386), .ZN(n13379) );
  OAI21_X1 U16506 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20169), .A(
        n13379), .ZN(n13380) );
  OAI22_X1 U16507 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20030), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13380), .ZN(n13384) );
  NOR2_X1 U16508 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20030), .ZN(
        n13381) );
  NAND2_X1 U16509 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13380), .ZN(
        n13382) );
  AOI22_X1 U16510 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13384), .B1(
        n13381), .B2(n13382), .ZN(n13388) );
  OAI211_X1 U16511 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20019), .A(
        n13388), .B(n13483), .ZN(n13487) );
  INV_X1 U16512 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19987) );
  AND2_X1 U16513 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13382), .ZN(
        n13383) );
  OAI22_X1 U16514 ( .A1(n19987), .A2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n13384), .B2(n13383), .ZN(n13385) );
  INV_X1 U16515 ( .A(n13385), .ZN(n13484) );
  XOR2_X1 U16516 ( .A(n13387), .B(n13386), .Z(n13481) );
  NAND2_X1 U16517 ( .A1(n13388), .A2(n13481), .ZN(n13485) );
  OAI211_X1 U16518 ( .C1(n13482), .C2(n13487), .A(n13484), .B(n13485), .ZN(
        n17086) );
  AOI22_X1 U16519 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13393) );
  AOI22_X1 U16520 ( .A1(n18520), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13392) );
  AOI22_X1 U16521 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13391) );
  AOI22_X1 U16522 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13390) );
  NAND4_X1 U16523 ( .A1(n13393), .A2(n13392), .A3(n13391), .A4(n13390), .ZN(
        n13400) );
  AOI22_X1 U16524 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18472), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U16525 ( .A1(n18519), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13397) );
  AOI22_X1 U16526 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18539), .B1(
        n18473), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U16527 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13395) );
  NAND4_X1 U16528 ( .A1(n13398), .A2(n13397), .A3(n13396), .A4(n13395), .ZN(
        n13399) );
  AOI22_X1 U16529 ( .A1(n18473), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13404) );
  AOI22_X1 U16530 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U16531 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U16532 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13401) );
  NAND4_X1 U16533 ( .A1(n13404), .A2(n13403), .A3(n13402), .A4(n13401), .ZN(
        n13410) );
  AOI22_X1 U16534 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13408) );
  AOI22_X1 U16535 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13311), .B1(
        n18519), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U16536 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13406) );
  AOI22_X1 U16537 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n17066), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13405) );
  NAND4_X1 U16538 ( .A1(n13408), .A2(n13407), .A3(n13406), .A4(n13405), .ZN(
        n13409) );
  NAND2_X1 U16539 ( .A1(n19564), .A2(n13489), .ZN(n13480) );
  AOI22_X1 U16540 ( .A1(n18519), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9794), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13414) );
  AOI22_X1 U16541 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U16542 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U16543 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n13311), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13411) );
  NAND4_X1 U16544 ( .A1(n13414), .A2(n13413), .A3(n13412), .A4(n13411), .ZN(
        n13420) );
  AOI22_X1 U16545 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U16546 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n17067), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U16547 ( .A1(n18520), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U16548 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13415) );
  NAND4_X1 U16549 ( .A1(n13418), .A2(n13417), .A3(n13416), .A4(n13415), .ZN(
        n13419) );
  AOI22_X1 U16550 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U16551 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9794), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13423) );
  AOI22_X1 U16552 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18539), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13422) );
  AOI22_X1 U16553 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13421) );
  NAND4_X1 U16554 ( .A1(n13424), .A2(n13423), .A3(n13422), .A4(n13421), .ZN(
        n13430) );
  AOI22_X1 U16555 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18533), .B1(
        n18472), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U16556 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18455), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13427) );
  AOI22_X1 U16557 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U16558 ( .A1(n18519), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13425) );
  NAND4_X1 U16559 ( .A1(n13428), .A2(n13427), .A3(n13426), .A4(n13425), .ZN(
        n13429) );
  NAND2_X1 U16560 ( .A1(n13463), .A2(n13462), .ZN(n13490) );
  AOI22_X1 U16561 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U16562 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n18539), .ZN(n13433) );
  AOI22_X1 U16563 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17067), .ZN(n13432) );
  AOI22_X1 U16564 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18534), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n18473), .ZN(n13431) );
  NAND4_X1 U16565 ( .A1(n13434), .A2(n13433), .A3(n13432), .A4(n13431), .ZN(
        n13440) );
  AOI22_X1 U16566 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18533), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n18518), .ZN(n13438) );
  AOI22_X1 U16567 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13311), .B1(
        n18472), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13437) );
  AOI22_X1 U16568 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17066), .ZN(n13436) );
  INV_X2 U16569 ( .A(n18486), .ZN(n18513) );
  AOI22_X1 U16570 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9793), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13435) );
  NAND4_X1 U16571 ( .A1(n13438), .A2(n13437), .A3(n13436), .A4(n13435), .ZN(
        n13439) );
  AOI22_X1 U16572 ( .A1(n18473), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13450) );
  AOI22_X1 U16573 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18472), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13449) );
  AOI22_X1 U16574 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13441) );
  OAI21_X1 U16575 ( .B1(n17029), .B2(n18426), .A(n13441), .ZN(n13447) );
  AOI22_X1 U16576 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13445) );
  AOI22_X1 U16577 ( .A1(n18519), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13444) );
  AOI22_X1 U16578 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13443) );
  AOI22_X1 U16579 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13275), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13442) );
  NAND4_X1 U16580 ( .A1(n13445), .A2(n13444), .A3(n13443), .A4(n13442), .ZN(
        n13446) );
  AOI211_X1 U16581 ( .C1(n9793), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n13447), .B(n13446), .ZN(n13448) );
  NOR2_X1 U16582 ( .A1(n19555), .A2(n13466), .ZN(n13461) );
  AOI22_X1 U16583 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n17067), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U16584 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9794), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13453) );
  AOI22_X1 U16585 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13452) );
  AOI22_X1 U16586 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18472), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13451) );
  NAND4_X1 U16587 ( .A1(n13454), .A2(n13453), .A3(n13452), .A4(n13451), .ZN(
        n13460) );
  AOI22_X1 U16588 ( .A1(n18473), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13458) );
  AOI22_X1 U16589 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18455), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U16590 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U16591 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n9795), .B1(
        n18519), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13455) );
  NAND4_X1 U16592 ( .A1(n13458), .A2(n13457), .A3(n13456), .A4(n13455), .ZN(
        n13459) );
  NOR2_X1 U16593 ( .A1(n13463), .A2(n13462), .ZN(n20015) );
  INV_X1 U16594 ( .A(n20015), .ZN(n13468) );
  NAND2_X1 U16595 ( .A1(n18732), .A2(n20205), .ZN(n13478) );
  AOI21_X1 U16596 ( .B1(n18624), .B2(n13468), .A(n13478), .ZN(n13464) );
  INV_X1 U16597 ( .A(n13464), .ZN(n15395) );
  OAI21_X1 U16598 ( .B1(n17094), .B2(n13465), .A(n15395), .ZN(n13474) );
  NAND2_X1 U16599 ( .A1(n13479), .A2(n13489), .ZN(n13493) );
  NAND2_X1 U16600 ( .A1(n18624), .A2(n17087), .ZN(n13470) );
  NAND2_X1 U16601 ( .A1(n19564), .A2(n13466), .ZN(n13467) );
  OAI21_X1 U16602 ( .B1(n13468), .B2(n16984), .A(n13467), .ZN(n13469) );
  AOI21_X1 U16603 ( .B1(n16984), .B2(n13470), .A(n13469), .ZN(n13471) );
  INV_X1 U16604 ( .A(n13471), .ZN(n13473) );
  INV_X1 U16605 ( .A(n17781), .ZN(n13476) );
  NAND2_X2 U16606 ( .A1(n13477), .A2(n13476), .ZN(n20004) );
  NOR2_X4 U16607 ( .A1(n15393), .A2(n10008), .ZN(n20016) );
  NAND2_X1 U16608 ( .A1(n13479), .A2(n13478), .ZN(n20215) );
  INV_X1 U16609 ( .A(n13480), .ZN(n19992) );
  NOR2_X1 U16610 ( .A1(n20205), .A2(n13491), .ZN(n19991) );
  NOR2_X4 U16611 ( .A1(n19419), .A2(n20014), .ZN(n19364) );
  INV_X1 U16612 ( .A(n13481), .ZN(n13488) );
  XNOR2_X1 U16613 ( .A(n13483), .B(n13482), .ZN(n13486) );
  OAI21_X1 U16614 ( .B1(n13488), .B2(n13487), .A(n19981), .ZN(n17085) );
  NAND2_X1 U16615 ( .A1(n13489), .A2(n19555), .ZN(n17092) );
  NOR2_X1 U16616 ( .A1(n19579), .A2(n17092), .ZN(n17090) );
  OAI211_X1 U16617 ( .C1(n19568), .C2(n20015), .A(n13491), .B(n13490), .ZN(
        n13492) );
  NOR2_X1 U16618 ( .A1(n13493), .A2(n13492), .ZN(n15397) );
  NOR2_X4 U16619 ( .A1(n20205), .A2(n17894), .ZN(n19205) );
  NAND2_X1 U16620 ( .A1(n17775), .A2(n19128), .ZN(n13543) );
  NAND2_X1 U16621 ( .A1(n9866), .A2(n19119), .ZN(n19081) );
  INV_X1 U16622 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18912) );
  NOR2_X1 U16623 ( .A1(n18924), .A2(n18912), .ZN(n19244) );
  NAND3_X1 U16624 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n19244), .ZN(n19219) );
  NOR2_X1 U16625 ( .A1(n17099), .A2(n19219), .ZN(n17104) );
  NAND2_X1 U16626 ( .A1(n19350), .A2(n17104), .ZN(n19226) );
  NAND2_X1 U16627 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17742) );
  NOR3_X1 U16628 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17751), .A3(
        n17758), .ZN(n13495) );
  NOR2_X1 U16629 ( .A1(n17742), .A2(n17758), .ZN(n13527) );
  INV_X1 U16630 ( .A(n13527), .ZN(n17181) );
  NOR2_X1 U16631 ( .A1(n19226), .A2(n17181), .ZN(n17109) );
  AOI21_X1 U16632 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17109), .A(
        n20165), .ZN(n13494) );
  AOI21_X1 U16633 ( .B1(n17794), .B2(n13495), .A(n13494), .ZN(n17778) );
  NAND2_X2 U16634 ( .A1(n17790), .A2(n19205), .ZN(n19126) );
  OR2_X1 U16635 ( .A1(n17778), .A2(n19126), .ZN(n13541) );
  INV_X1 U16636 ( .A(n13495), .ZN(n17768) );
  INV_X1 U16637 ( .A(n17192), .ZN(n13511) );
  NOR2_X1 U16638 ( .A1(n13496), .A2(n13511), .ZN(n13512) );
  NOR2_X1 U16639 ( .A1(n13512), .A2(n13497), .ZN(n13507) );
  NOR2_X1 U16640 ( .A1(n18712), .A2(n13507), .ZN(n13504) );
  NAND2_X1 U16641 ( .A1(n13504), .A2(n13498), .ZN(n13502) );
  NOR2_X1 U16642 ( .A1(n18706), .A2(n13502), .ZN(n13501) );
  NAND2_X1 U16643 ( .A1(n13501), .A2(n13499), .ZN(n13500) );
  NOR2_X1 U16644 ( .A1(n17790), .A2(n13500), .ZN(n13522) );
  XNOR2_X1 U16645 ( .A(n18698), .B(n13500), .ZN(n19131) );
  XNOR2_X1 U16646 ( .A(n18703), .B(n13501), .ZN(n13518) );
  XOR2_X1 U16647 ( .A(n18706), .B(n13502), .Z(n13503) );
  NAND2_X1 U16648 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13503), .ZN(
        n13517) );
  XNOR2_X1 U16649 ( .A(n19480), .B(n13503), .ZN(n19157) );
  XNOR2_X1 U16650 ( .A(n18709), .B(n13504), .ZN(n13505) );
  NAND2_X1 U16651 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13505), .ZN(
        n13516) );
  XNOR2_X1 U16652 ( .A(n19488), .B(n13505), .ZN(n19168) );
  XOR2_X1 U16653 ( .A(n18712), .B(n13507), .Z(n13506) );
  NAND2_X1 U16654 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13506), .ZN(
        n13515) );
  XNOR2_X1 U16655 ( .A(n19496), .B(n13506), .ZN(n19181) );
  INV_X1 U16656 ( .A(n13507), .ZN(n13508) );
  OAI21_X1 U16657 ( .B1(n13511), .B2(n13509), .A(n13508), .ZN(n13510) );
  NAND2_X1 U16658 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13510), .ZN(
        n13514) );
  XOR2_X1 U16659 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13510), .Z(
        n19194) );
  NOR2_X1 U16660 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18721), .ZN(
        n13513) );
  INV_X1 U16661 ( .A(n19201), .ZN(n19203) );
  INV_X1 U16662 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20181) );
  NAND2_X1 U16663 ( .A1(n13511), .A2(n20181), .ZN(n19210) );
  NOR2_X1 U16664 ( .A1(n19203), .A2(n19210), .ZN(n19202) );
  NOR3_X1 U16665 ( .A1(n13513), .A2(n13512), .A3(n19202), .ZN(n19193) );
  NAND2_X1 U16666 ( .A1(n19194), .A2(n19193), .ZN(n19192) );
  NAND2_X1 U16667 ( .A1(n13514), .A2(n19192), .ZN(n19180) );
  NAND2_X1 U16668 ( .A1(n19181), .A2(n19180), .ZN(n19179) );
  NAND2_X1 U16669 ( .A1(n13515), .A2(n19179), .ZN(n19167) );
  NAND2_X1 U16670 ( .A1(n19168), .A2(n19167), .ZN(n19166) );
  NAND2_X1 U16671 ( .A1(n13516), .A2(n19166), .ZN(n19156) );
  NAND2_X1 U16672 ( .A1(n19157), .A2(n19156), .ZN(n19155) );
  NAND2_X1 U16673 ( .A1(n13517), .A2(n19155), .ZN(n13519) );
  NAND2_X1 U16674 ( .A1(n13518), .A2(n13519), .ZN(n13520) );
  XOR2_X1 U16675 ( .A(n13519), .B(n13518), .Z(n19144) );
  NAND2_X1 U16676 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19144), .ZN(
        n19143) );
  NAND2_X1 U16677 ( .A1(n13522), .A2(n13525), .ZN(n13526) );
  INV_X1 U16678 ( .A(n13522), .ZN(n13524) );
  NAND2_X1 U16679 ( .A1(n19131), .A2(n19132), .ZN(n19130) );
  NAND2_X1 U16680 ( .A1(n13525), .A2(n13524), .ZN(n13523) );
  OAI211_X1 U16681 ( .C1(n13525), .C2(n13524), .A(n19130), .B(n13523), .ZN(
        n19115) );
  NAND2_X1 U16682 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19115), .ZN(
        n19114) );
  NAND2_X1 U16683 ( .A1(n19363), .A2(n19405), .ZN(n19038) );
  NAND2_X1 U16684 ( .A1(n17104), .A2(n19347), .ZN(n18857) );
  INV_X1 U16685 ( .A(n18857), .ZN(n19224) );
  NAND2_X1 U16686 ( .A1(n13527), .A2(n19224), .ZN(n17756) );
  OAI21_X1 U16687 ( .B1(n17751), .B2(n17756), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13528) );
  OAI21_X1 U16688 ( .B1(n17768), .B2(n17792), .A(n13528), .ZN(n17774) );
  AOI21_X1 U16689 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n20201)
         );
  INV_X1 U16690 ( .A(n20201), .ZN(n19542) );
  NOR3_X4 U16691 ( .A1(n19163), .A2(P3_STATEBS16_REG_SCAN_IN), .A3(n20164), 
        .ZN(n19071) );
  INV_X1 U16692 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18888) );
  NAND3_X1 U16693 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19092) );
  NOR2_X1 U16694 ( .A1(n19092), .A2(n18138), .ZN(n18122) );
  NOR2_X2 U16695 ( .A1(n19001), .A2(n19000), .ZN(n18974) );
  INV_X1 U16696 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18973) );
  INV_X1 U16697 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18972) );
  NOR2_X4 U16698 ( .A1(n18888), .A2(n18873), .ZN(n18887) );
  AND4_X2 U16699 ( .A1(n18887), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18846) );
  NAND2_X1 U16700 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18852) );
  INV_X1 U16701 ( .A(n18852), .ZN(n13530) );
  INV_X1 U16702 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17936) );
  INV_X1 U16703 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20135) );
  NAND2_X1 U16704 ( .A1(n20164), .A2(n20153), .ZN(n20154) );
  NOR2_X1 U16705 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n20154), .ZN(n20217) );
  INV_X1 U16706 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n15401) );
  NOR2_X1 U16707 ( .A1(n20135), .A2(n19529), .ZN(n17771) );
  NAND3_X1 U16708 ( .A1(n18846), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17753) );
  NOR2_X1 U16709 ( .A1(n17936), .A2(n17753), .ZN(n13533) );
  INV_X1 U16710 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19208) );
  NOR2_X1 U16711 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20047), .ZN(n19048) );
  NAND2_X1 U16712 ( .A1(n20164), .A2(n20047), .ZN(n20056) );
  NAND2_X1 U16713 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19538) );
  AOI21_X1 U16714 ( .B1(n20056), .B2(n19538), .A(n20178), .ZN(n19550) );
  NOR3_X1 U16715 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n20204), .ZN(n19608) );
  INV_X2 U16716 ( .A(n19922), .ZN(n19652) );
  OAI21_X2 U16717 ( .B1(n19208), .B2(n18964), .A(n19652), .ZN(n19052) );
  NAND2_X1 U16718 ( .A1(n13533), .A2(n19052), .ZN(n17745) );
  INV_X1 U16719 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17922) );
  XOR2_X1 U16720 ( .A(n17922), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n13536) );
  NOR2_X1 U16721 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18964), .ZN(
        n17762) );
  INV_X1 U16722 ( .A(n13532), .ZN(n13535) );
  INV_X1 U16723 ( .A(n19048), .ZN(n19011) );
  OR2_X1 U16724 ( .A1(n19652), .A2(n13533), .ZN(n13534) );
  OAI211_X1 U16725 ( .C1(n13535), .C2(n19011), .A(n19212), .B(n13534), .ZN(
        n17755) );
  NOR2_X1 U16726 ( .A1(n17762), .A2(n17755), .ZN(n17744) );
  OAI22_X1 U16727 ( .A1(n17745), .A2(n13536), .B1(n17744), .B2(n17922), .ZN(
        n13537) );
  AOI211_X1 U16728 ( .C1(n19071), .C2(n18224), .A(n17771), .B(n13537), .ZN(
        n13538) );
  NAND2_X1 U16729 ( .A1(n13543), .A2(n13542), .ZN(P3_U2799) );
  INV_X1 U16730 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n21213) );
  NOR2_X1 U16731 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n21213), .ZN(n13545) );
  NOR4_X1 U16732 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13544) );
  INV_X1 U16733 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n21166) );
  NAND4_X1 U16734 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13545), .A3(n13544), .A4(
        n21166), .ZN(n13567) );
  NOR2_X1 U16735 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13567), .ZN(n17875)
         );
  NOR4_X1 U16736 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13549) );
  NOR4_X1 U16737 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n13548) );
  NOR4_X1 U16738 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13547) );
  NOR4_X1 U16739 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_10__SCAN_IN), .ZN(n13546) );
  AND4_X1 U16740 ( .A1(n13549), .A2(n13548), .A3(n13547), .A4(n13546), .ZN(
        n13554) );
  NOR4_X1 U16741 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_6__SCAN_IN), .ZN(n13552) );
  NOR4_X1 U16742 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n13551) );
  NOR4_X1 U16743 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13550) );
  INV_X1 U16744 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21464) );
  AND4_X1 U16745 ( .A1(n13552), .A2(n13551), .A3(n13550), .A4(n21464), .ZN(
        n13553) );
  NAND2_X1 U16746 ( .A1(n13554), .A2(n13553), .ZN(n13555) );
  INV_X2 U16747 ( .A(n14552), .ZN(n15371) );
  INV_X1 U16748 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21536) );
  NOR3_X1 U16749 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21536), .ZN(n13557) );
  NOR4_X1 U16750 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13556) );
  NAND4_X1 U16751 ( .A1(n15371), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13557), .A4(
        n13556), .ZN(U214) );
  NOR4_X1 U16752 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13561) );
  NOR4_X1 U16753 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13560) );
  NOR4_X1 U16754 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13559) );
  NOR4_X1 U16755 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13558) );
  NAND4_X1 U16756 ( .A1(n13561), .A2(n13560), .A3(n13559), .A4(n13558), .ZN(
        n13566) );
  NOR4_X1 U16757 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13564) );
  NOR4_X1 U16758 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13563) );
  NOR4_X1 U16759 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13562) );
  INV_X1 U16760 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n21117) );
  NAND4_X1 U16761 ( .A1(n13564), .A2(n13563), .A3(n13562), .A4(n21117), .ZN(
        n13565) );
  OAI21_X2 U16762 ( .B1(n13566), .B2(n13565), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n15215) );
  NOR2_X1 U16763 ( .A1(n15215), .A2(n13567), .ZN(n17801) );
  NAND2_X1 U16764 ( .A1(n17801), .A2(U214), .ZN(U212) );
  XNOR2_X1 U16765 ( .A(n13568), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17567) );
  NOR2_X1 U16766 ( .A1(n17567), .A2(n17669), .ZN(n13586) );
  NAND2_X1 U16767 ( .A1(n13569), .A2(n13570), .ZN(n16703) );
  XNOR2_X1 U16768 ( .A(n16700), .B(n13571), .ZN(n16702) );
  XNOR2_X1 U16769 ( .A(n16703), .B(n16702), .ZN(n17565) );
  NOR2_X1 U16770 ( .A1(n17565), .A2(n17681), .ZN(n13585) );
  NOR2_X1 U16771 ( .A1(n17662), .A2(n13572), .ZN(n17633) );
  INV_X1 U16772 ( .A(n17633), .ZN(n13573) );
  NOR2_X1 U16773 ( .A1(n15228), .A2(n13573), .ZN(n13577) );
  OAI21_X1 U16774 ( .B1(n17675), .B2(n13748), .A(n13574), .ZN(n17664) );
  OAI21_X1 U16775 ( .B1(n13575), .B2(n17664), .A(n14944), .ZN(n17656) );
  INV_X1 U16776 ( .A(n17656), .ZN(n13576) );
  MUX2_X1 U16777 ( .A(n13577), .B(n13576), .S(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n13584) );
  XNOR2_X1 U16778 ( .A(n13578), .B(n13579), .ZN(n20474) );
  NOR2_X1 U16779 ( .A1(n15234), .A2(n13580), .ZN(n13581) );
  NOR2_X1 U16780 ( .A1(n9930), .A2(n13581), .ZN(n20355) );
  AOI22_X1 U16781 ( .A1(n12878), .A2(n20355), .B1(n20376), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n13582) );
  OAI21_X1 U16782 ( .B1(n20474), .B2(n17671), .A(n13582), .ZN(n13583) );
  OR4_X1 U16783 ( .A1(n13586), .A2(n13585), .A3(n13584), .A4(n13583), .ZN(
        P2_U3040) );
  NOR3_X1 U16784 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18239) );
  NAND2_X1 U16785 ( .A1(n18239), .A2(n18234), .ZN(n18233) );
  NOR2_X1 U16786 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18233), .ZN(n18211) );
  INV_X1 U16787 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18204) );
  NAND2_X1 U16788 ( .A1(n18211), .A2(n18204), .ZN(n18198) );
  INV_X1 U16789 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18549) );
  NAND2_X1 U16790 ( .A1(n18184), .A2(n18549), .ZN(n18178) );
  INV_X1 U16791 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18148) );
  NAND2_X1 U16792 ( .A1(n18157), .A2(n18148), .ZN(n18144) );
  INV_X1 U16793 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n18484) );
  NAND2_X1 U16794 ( .A1(n18132), .A2(n18484), .ZN(n18129) );
  INV_X1 U16795 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n18108) );
  NAND2_X1 U16796 ( .A1(n18109), .A2(n18108), .ZN(n18105) );
  INV_X1 U16797 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n18081) );
  NAND2_X1 U16798 ( .A1(n18085), .A2(n18081), .ZN(n18080) );
  INV_X1 U16799 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n18398) );
  NAND2_X1 U16800 ( .A1(n18059), .A2(n18398), .ZN(n18056) );
  INV_X1 U16801 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n18036) );
  NAND2_X1 U16802 ( .A1(n18042), .A2(n18036), .ZN(n18035) );
  INV_X1 U16803 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18368) );
  NAND2_X1 U16804 ( .A1(n18022), .A2(n18368), .ZN(n18015) );
  INV_X1 U16805 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n18278) );
  NAND2_X1 U16806 ( .A1(n17996), .A2(n18278), .ZN(n17992) );
  NOR2_X1 U16807 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17992), .ZN(n17965) );
  INV_X1 U16808 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n18281) );
  NAND2_X1 U16809 ( .A1(n17965), .A2(n18281), .ZN(n13589) );
  NOR2_X1 U16810 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n13589), .ZN(n17960) );
  NAND2_X1 U16811 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n20206) );
  NAND2_X1 U16812 ( .A1(n20220), .A2(n18732), .ZN(n20218) );
  NAND2_X1 U16813 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19555), .ZN(n13588) );
  AOI211_X4 U16814 ( .C1(n20204), .C2(n20206), .A(n20218), .B(n13588), .ZN(
        n18259) );
  AOI211_X1 U16815 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n13589), .A(n17960), .B(
        n18269), .ZN(n13609) );
  INV_X1 U16816 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20124) );
  NAND2_X1 U16817 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n20071), .ZN(n20195) );
  INV_X1 U16818 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n20074) );
  NOR2_X1 U16819 ( .A1(n20195), .A2(n20074), .ZN(n20073) );
  NOR2_X1 U16820 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n20058) );
  NOR3_X1 U16821 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n20073), .A3(n20058), 
        .ZN(n17091) );
  INV_X1 U16822 ( .A(n17091), .ZN(n20203) );
  AOI211_X1 U16823 ( .C1(n20205), .C2(n20203), .A(n10001), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n13604) );
  INV_X1 U16824 ( .A(n13604), .ZN(n20040) );
  INV_X1 U16825 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20118) );
  INV_X1 U16826 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20098) );
  INV_X1 U16827 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20095) );
  INV_X1 U16828 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20086) );
  INV_X1 U16829 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20082) );
  INV_X1 U16830 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20078) );
  NAND2_X1 U16831 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n18242) );
  NOR2_X1 U16832 ( .A1(n20078), .A2(n18242), .ZN(n18218) );
  NAND2_X1 U16833 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18218), .ZN(n18203) );
  NOR2_X1 U16834 ( .A1(n20082), .A2(n18203), .ZN(n18177) );
  NAND2_X1 U16835 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18177), .ZN(n18174) );
  NOR2_X1 U16836 ( .A1(n20086), .A2(n18174), .ZN(n18159) );
  NAND2_X1 U16837 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18159), .ZN(n18158) );
  NAND2_X1 U16838 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n18133) );
  NOR3_X1 U16839 ( .A1(n20095), .A2(n18158), .A3(n18133), .ZN(n18112) );
  NAND2_X1 U16840 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18112), .ZN(n18096) );
  NOR2_X1 U16841 ( .A1(n20098), .A2(n18096), .ZN(n18086) );
  NAND2_X1 U16842 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n18086), .ZN(n18003) );
  INV_X1 U16843 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20114) );
  INV_X1 U16844 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20110) );
  INV_X1 U16845 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20108) );
  NAND3_X1 U16846 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(P3_REIP_REG_17__SCAN_IN), 
        .A3(P3_REIP_REG_16__SCAN_IN), .ZN(n18031) );
  NOR3_X1 U16847 ( .A1(n20110), .A2(n20108), .A3(n18031), .ZN(n18019) );
  NAND2_X1 U16848 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18019), .ZN(n18004) );
  NOR2_X1 U16849 ( .A1(n20114), .A2(n18004), .ZN(n18002) );
  NAND2_X1 U16850 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n18002), .ZN(n17989) );
  NOR3_X1 U16851 ( .A1(n20118), .A2(n18003), .A3(n17989), .ZN(n17976) );
  NAND2_X1 U16852 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17976), .ZN(n13590) );
  NOR2_X1 U16853 ( .A1(n18263), .A2(n13590), .ZN(n17972) );
  NAND2_X1 U16854 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17972), .ZN(n17908) );
  NAND3_X1 U16855 ( .A1(n15401), .A2(n20047), .A3(n20204), .ZN(n20055) );
  NOR2_X1 U16856 ( .A1(n20164), .A2(n20055), .ZN(n18225) );
  INV_X1 U16857 ( .A(n20049), .ZN(n19213) );
  NOR2_X2 U16858 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n20153), .ZN(n20050) );
  NAND2_X1 U16859 ( .A1(n19213), .A2(n20050), .ZN(n20044) );
  NAND2_X1 U16860 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n18273), .ZN(n17970) );
  OR2_X1 U16861 ( .A1(n13590), .A2(n17970), .ZN(n13591) );
  NAND2_X1 U16862 ( .A1(n18263), .A2(n18273), .ZN(n18271) );
  OAI21_X1 U16863 ( .B1(n20124), .B2(n13591), .A(n18271), .ZN(n17914) );
  AOI21_X1 U16864 ( .B1(n20124), .B2(n17908), .A(n17914), .ZN(n13608) );
  INV_X1 U16865 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13605) );
  NAND2_X1 U16866 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18936) );
  NAND2_X1 U16867 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18935), .ZN(
        n13597) );
  NOR2_X1 U16868 ( .A1(n18936), .A2(n13597), .ZN(n13595) );
  NAND2_X1 U16869 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18889) );
  NOR2_X1 U16870 ( .A1(n18888), .A2(n18889), .ZN(n18874) );
  NAND2_X1 U16871 ( .A1(n13595), .A2(n18874), .ZN(n18848) );
  AOI21_X1 U16872 ( .B1(n13605), .B2(n18848), .A(n17910), .ZN(n18881) );
  INV_X1 U16873 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18891) );
  NAND3_X1 U16874 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18887), .A3(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13593) );
  INV_X1 U16875 ( .A(n18848), .ZN(n13592) );
  AOI21_X1 U16876 ( .B1(n18891), .B2(n13593), .A(n13592), .ZN(n18893) );
  NAND2_X1 U16877 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18887), .ZN(
        n13594) );
  XNOR2_X1 U16878 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n13594), .ZN(
        n18905) );
  INV_X1 U16879 ( .A(n13595), .ZN(n18885) );
  AOI22_X1 U16880 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18887), .B1(
        n18888), .B2(n18885), .ZN(n18916) );
  INV_X1 U16881 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18940) );
  INV_X1 U16882 ( .A(n13597), .ZN(n13598) );
  NAND2_X1 U16883 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13598), .ZN(
        n13596) );
  AOI21_X1 U16884 ( .B1(n18940), .B2(n13596), .A(n13595), .ZN(n18938) );
  INV_X1 U16885 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18945) );
  AOI22_X1 U16886 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13598), .B1(
        n13597), .B2(n18945), .ZN(n18954) );
  INV_X1 U16887 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18933) );
  NAND2_X1 U16888 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10350), .ZN(
        n18931) );
  AOI21_X1 U16889 ( .B1(n18933), .B2(n18931), .A(n13598), .ZN(n18965) );
  NOR2_X1 U16890 ( .A1(n19208), .A2(n13599), .ZN(n19012) );
  NAND2_X1 U16891 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19012), .ZN(
        n18072) );
  INV_X1 U16892 ( .A(n18072), .ZN(n18066) );
  NAND2_X1 U16893 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18066), .ZN(
        n18065) );
  NOR2_X1 U16894 ( .A1(n19000), .A2(n18065), .ZN(n18976) );
  NAND2_X1 U16895 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18976), .ZN(
        n13601) );
  INV_X1 U16896 ( .A(n18931), .ZN(n13600) );
  AOI21_X1 U16897 ( .B1(n18972), .B2(n13601), .A(n13600), .ZN(n18977) );
  XOR2_X1 U16898 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B(n18976), .Z(
        n18985) );
  NOR2_X1 U16899 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19208), .ZN(
        n18252) );
  AND2_X1 U16900 ( .A1(n18974), .A2(n18252), .ZN(n13602) );
  NOR2_X1 U16901 ( .A1(n18985), .A2(n18041), .ZN(n18040) );
  NOR2_X1 U16902 ( .A1(n18040), .A2(n18164), .ZN(n18029) );
  NOR2_X1 U16903 ( .A1(n18977), .A2(n18029), .ZN(n18028) );
  NOR2_X1 U16904 ( .A1(n18028), .A2(n18164), .ZN(n18021) );
  NOR2_X1 U16905 ( .A1(n18965), .A2(n18021), .ZN(n18020) );
  NOR2_X1 U16906 ( .A1(n18916), .A2(n17987), .ZN(n17986) );
  NOR2_X1 U16907 ( .A1(n17986), .A2(n18164), .ZN(n17980) );
  NOR2_X1 U16908 ( .A1(n18881), .A2(n9853), .ZN(n17913) );
  AOI211_X1 U16909 ( .C1(n18881), .C2(n9853), .A(n17913), .B(n20053), .ZN(
        n13607) );
  AOI211_X4 U16910 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n19555), .A(n13604), .B(
        n20218), .ZN(n18248) );
  INV_X1 U16911 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n18282) );
  OAI22_X1 U16912 ( .A1(n13605), .A2(n18260), .B1(n18270), .B2(n18282), .ZN(
        n13606) );
  OR4_X1 U16913 ( .A1(n13609), .A2(n13608), .A3(n13607), .A4(n13606), .ZN(
        P3_U2645) );
  AOI211_X1 U16914 ( .C1(n16555), .C2(n13611), .A(n13610), .B(n21086), .ZN(
        n13618) );
  INV_X1 U16915 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n13612) );
  OAI22_X1 U16916 ( .A1(n13613), .A2(n20399), .B1(n13612), .B2(n20396), .ZN(
        n13617) );
  OAI22_X1 U16917 ( .A1(n16558), .A2(n20380), .B1(n21156), .B2(n20374), .ZN(
        n13616) );
  OAI22_X1 U16918 ( .A1(n16554), .A2(n20402), .B1(n20401), .B2(n13614), .ZN(
        n13615) );
  OR4_X1 U16919 ( .A1(n13618), .A2(n13617), .A3(n13616), .A4(n13615), .ZN(
        P2_U2828) );
  NOR2_X1 U16920 ( .A1(n21086), .A2(n12815), .ZN(n20410) );
  INV_X1 U16921 ( .A(n20410), .ZN(n13632) );
  AOI211_X1 U16922 ( .C1(n17501), .C2(n13619), .A(n20253), .B(n13632), .ZN(
        n13631) );
  INV_X1 U16923 ( .A(n17501), .ZN(n13621) );
  NAND2_X1 U16924 ( .A1(n20370), .A2(n12815), .ZN(n14951) );
  INV_X1 U16925 ( .A(n20396), .ZN(n20359) );
  AOI22_X1 U16926 ( .A1(n20406), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_EBX_REG_15__SCAN_IN), .B2(n20359), .ZN(n13620) );
  OAI211_X1 U16927 ( .C1(n13621), .C2(n14951), .A(n13620), .B(n20347), .ZN(
        n13630) );
  INV_X1 U16928 ( .A(n13622), .ZN(n13623) );
  OAI22_X1 U16929 ( .A1(n13623), .A2(n20399), .B1(n17511), .B2(n20380), .ZN(
        n13629) );
  OAI21_X1 U16930 ( .B1(n17598), .B2(n13625), .A(n13624), .ZN(n20451) );
  NAND2_X1 U16931 ( .A1(n14609), .A2(n13626), .ZN(n13627) );
  NAND2_X1 U16932 ( .A1(n16667), .A2(n13627), .ZN(n17507) );
  OAI22_X1 U16933 ( .A1(n20451), .A2(n20401), .B1(n20402), .B2(n17507), .ZN(
        n13628) );
  OR4_X1 U16934 ( .A1(n13631), .A2(n13630), .A3(n13629), .A4(n13628), .ZN(
        P2_U2840) );
  AOI211_X1 U16935 ( .C1(n13635), .C2(n13634), .A(n13633), .B(n13632), .ZN(
        n13649) );
  NAND2_X1 U16936 ( .A1(n13636), .A2(n20328), .ZN(n13638) );
  AOI21_X1 U16937 ( .B1(n20359), .B2(P2_EBX_REG_17__SCAN_IN), .A(n20376), .ZN(
        n13637) );
  OAI211_X1 U16938 ( .C1(n20374), .C2(n21137), .A(n13638), .B(n13637), .ZN(
        n13648) );
  INV_X1 U16939 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13639) );
  OAI22_X1 U16940 ( .A1(n13639), .A2(n20380), .B1(n16661), .B2(n14951), .ZN(
        n13647) );
  OAI21_X1 U16941 ( .B1(n13640), .B2(n13642), .A(n13641), .ZN(n16832) );
  NOR2_X1 U16942 ( .A1(n16668), .A2(n13644), .ZN(n13645) );
  OR2_X1 U16943 ( .A1(n13643), .A2(n13645), .ZN(n16659) );
  OAI22_X1 U16944 ( .A1(n16832), .A2(n20401), .B1(n20402), .B2(n16659), .ZN(
        n13646) );
  OR4_X1 U16945 ( .A1(n13649), .A2(n13648), .A3(n13647), .A4(n13646), .ZN(
        P2_U2838) );
  AOI211_X1 U16946 ( .C1(n16627), .C2(n13651), .A(n13650), .B(n21086), .ZN(
        n13662) );
  OAI22_X1 U16947 ( .A1(n13652), .A2(n20399), .B1(n21145), .B2(n20374), .ZN(
        n13661) );
  OAI22_X1 U16948 ( .A1(n20396), .A2(n11916), .B1(n16625), .B2(n20380), .ZN(
        n13660) );
  OAI21_X1 U16949 ( .B1(n12622), .B2(n13655), .A(n13654), .ZN(n16794) );
  AND2_X1 U16950 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  OR2_X1 U16951 ( .A1(n13658), .A2(n16613), .ZN(n16790) );
  OAI22_X1 U16952 ( .A1(n16794), .A2(n20401), .B1(n20402), .B2(n16790), .ZN(
        n13659) );
  OR4_X1 U16953 ( .A1(n13662), .A2(n13661), .A3(n13660), .A4(n13659), .ZN(
        P2_U2834) );
  AOI211_X1 U16954 ( .C1(n16601), .C2(n13664), .A(n13663), .B(n21086), .ZN(
        n13676) );
  OAI22_X1 U16955 ( .A1(n13665), .A2(n20399), .B1(n21148), .B2(n20374), .ZN(
        n13675) );
  INV_X1 U16956 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n13666) );
  OAI22_X1 U16957 ( .A1(n20396), .A2(n13666), .B1(n16599), .B2(n20380), .ZN(
        n13674) );
  NAND2_X1 U16958 ( .A1(n13667), .A2(n13668), .ZN(n13669) );
  NAND2_X1 U16959 ( .A1(n16447), .A2(n13669), .ZN(n17468) );
  AND2_X1 U16960 ( .A1(n13670), .A2(n13671), .ZN(n13672) );
  OR2_X1 U16961 ( .A1(n13672), .A2(n16511), .ZN(n16766) );
  OAI22_X1 U16962 ( .A1(n17468), .A2(n20402), .B1(n20401), .B2(n16766), .ZN(
        n13673) );
  OR4_X1 U16963 ( .A1(n13676), .A2(n13675), .A3(n13674), .A4(n13673), .ZN(
        P2_U2832) );
  AND2_X1 U16964 ( .A1(n21177), .A2(n12040), .ZN(n13678) );
  INV_X1 U16965 ( .A(n13784), .ZN(n13783) );
  AOI211_X1 U16966 ( .C1(P2_MEMORYFETCH_REG_SCAN_IN), .C2(n20384), .A(n13678), 
        .B(n13783), .ZN(n13677) );
  INV_X1 U16967 ( .A(n13677), .ZN(P2_U2814) );
  INV_X1 U16968 ( .A(n13681), .ZN(n13680) );
  OAI21_X1 U16969 ( .B1(n13678), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n21239), 
        .ZN(n13679) );
  OAI21_X1 U16970 ( .B1(n13680), .B2(n21239), .A(n13679), .ZN(P2_U3612) );
  AND2_X1 U16971 ( .A1(n13681), .A2(n21236), .ZN(n13767) );
  NOR4_X1 U16972 ( .A1(n17706), .A2(n12489), .A3(n13767), .A4(n15197), .ZN(
        n17713) );
  NOR2_X1 U16973 ( .A1(n17713), .A2(n15207), .ZN(n21223) );
  OAI21_X1 U16974 ( .B1(n13683), .B2(n21223), .A(n13682), .ZN(P2_U2819) );
  NAND2_X1 U16975 ( .A1(n20398), .A2(n13684), .ZN(n13685) );
  NAND2_X1 U16976 ( .A1(n10342), .A2(n13685), .ZN(n17680) );
  INV_X1 U16977 ( .A(n17680), .ZN(n13690) );
  NAND2_X1 U16978 ( .A1(n20376), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n17678) );
  INV_X1 U16979 ( .A(n17678), .ZN(n13689) );
  OAI21_X1 U16980 ( .B1(n13687), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13686), .ZN(n17668) );
  NOR2_X1 U16981 ( .A1(n17566), .A2(n17668), .ZN(n13688) );
  AOI211_X1 U16982 ( .C1(n17592), .C2(n13690), .A(n13689), .B(n13688), .ZN(
        n13693) );
  OAI21_X1 U16983 ( .B1(n17564), .B2(n13691), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13692) );
  OAI211_X1 U16984 ( .C1(n17577), .C2(n20403), .A(n13693), .B(n13692), .ZN(
        P2_U3014) );
  OR2_X1 U16985 ( .A1(n15199), .A2(n15207), .ZN(n13694) );
  OAI21_X1 U16986 ( .B1(n13695), .B2(n13694), .A(n13920), .ZN(n13696) );
  INV_X1 U16987 ( .A(n21229), .ZN(n21101) );
  NAND2_X1 U16988 ( .A1(n20532), .A2(n21227), .ZN(n20502) );
  INV_X1 U16989 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n16475) );
  NAND2_X1 U16990 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n21205) );
  OR2_X1 U16991 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n21205), .ZN(n20507) );
  INV_X1 U16992 ( .A(P2_UWORD_REG_13__SCAN_IN), .ZN(n13697) );
  INV_X2 U16993 ( .A(n20507), .ZN(n20541) );
  INV_X1 U16994 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n17879) );
  OAI222_X1 U16995 ( .A1(n20502), .A2(n16475), .B1(n20507), .B2(n13697), .C1(
        n20534), .C2(n17879), .ZN(P2_U2922) );
  INV_X1 U16996 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13698) );
  INV_X1 U16997 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n15898) );
  INV_X1 U16998 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n17880) );
  OAI222_X1 U16999 ( .A1(n20502), .A2(n13698), .B1(n20507), .B2(n15898), .C1(
        n20534), .C2(n17880), .ZN(P2_U2921) );
  INV_X1 U17000 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n17871) );
  INV_X1 U17001 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13699) );
  OAI222_X1 U17002 ( .A1(n20502), .A2(n13700), .B1(n20534), .B2(n17871), .C1(
        n13699), .C2(n20507), .ZN(P2_U2930) );
  INV_X1 U17003 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13702) );
  INV_X1 U17004 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n17869) );
  INV_X1 U17005 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13701) );
  OAI222_X1 U17006 ( .A1(n20502), .A2(n13702), .B1(n20534), .B2(n17869), .C1(
        n13701), .C2(n20507), .ZN(P2_U2932) );
  INV_X1 U17007 ( .A(n14874), .ZN(n13711) );
  OAI21_X1 U17008 ( .B1(n10355), .B2(n13704), .A(n13703), .ZN(n13755) );
  INV_X1 U17009 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14877) );
  OAI22_X1 U17010 ( .A1(n13755), .A2(n17566), .B1(n17596), .B2(n14877), .ZN(
        n13710) );
  NAND2_X1 U17011 ( .A1(n13706), .A2(n13705), .ZN(n13707) );
  NAND2_X1 U17012 ( .A1(n13708), .A2(n13707), .ZN(n13745) );
  NAND2_X1 U17013 ( .A1(n20376), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13746) );
  OAI21_X1 U17014 ( .B1(n13745), .B2(n17572), .A(n13746), .ZN(n13709) );
  AOI211_X1 U17015 ( .C1(n17582), .C2(n13711), .A(n13710), .B(n13709), .ZN(
        n13712) );
  OAI21_X1 U17016 ( .B1(n9970), .B2(n17577), .A(n13712), .ZN(P2_U3012) );
  NAND3_X1 U17017 ( .A1(n12647), .A2(n13993), .A3(n13722), .ZN(n13714) );
  INV_X1 U17018 ( .A(n13714), .ZN(n13713) );
  INV_X1 U17019 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21551) );
  INV_X2 U17020 ( .A(n16334), .ZN(n16320) );
  NAND2_X1 U17021 ( .A1(n16320), .A2(n21438), .ZN(n15165) );
  OAI211_X1 U17022 ( .C1(n13713), .C2(n21551), .A(n13985), .B(n15165), .ZN(
        P1_U2801) );
  NOR2_X1 U17023 ( .A1(n15116), .A2(n13715), .ZN(n13718) );
  INV_X1 U17024 ( .A(n15165), .ZN(n13716) );
  OAI21_X1 U17025 ( .B1(n13716), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n21539), 
        .ZN(n13717) );
  OAI21_X1 U17026 ( .B1(n21539), .B2(n13718), .A(n13717), .ZN(P1_U3487) );
  NAND2_X1 U17027 ( .A1(n12647), .A2(n13722), .ZN(n13719) );
  NAND2_X1 U17028 ( .A1(n12774), .A2(n13719), .ZN(n13720) );
  OAI21_X1 U17029 ( .B1(n17170), .B2(n15116), .A(n13720), .ZN(n21249) );
  AND2_X1 U17030 ( .A1(n13851), .A2(n21543), .ZN(n13886) );
  INV_X1 U17031 ( .A(n17186), .ZN(n13924) );
  OR2_X1 U17032 ( .A1(n13886), .A2(n13924), .ZN(n13721) );
  AND2_X1 U17033 ( .A1(n13721), .A2(n21452), .ZN(n21542) );
  NOR2_X1 U17034 ( .A1(n21249), .A2(n21542), .ZN(n17153) );
  NOR2_X1 U17035 ( .A1(n17153), .A2(n21248), .ZN(n21256) );
  INV_X1 U17036 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13728) );
  AND3_X1 U17037 ( .A1(n12774), .A2(n17150), .A3(n13858), .ZN(n13726) );
  INV_X1 U17038 ( .A(n13722), .ZN(n13860) );
  NAND2_X1 U17039 ( .A1(n12647), .A2(n13860), .ZN(n13725) );
  INV_X1 U17040 ( .A(n13856), .ZN(n13723) );
  NAND2_X1 U17041 ( .A1(n17170), .A2(n13723), .ZN(n13724) );
  OAI211_X1 U17042 ( .C1(n17170), .C2(n13726), .A(n13725), .B(n13724), .ZN(
        n17152) );
  NAND2_X1 U17043 ( .A1(n21256), .A2(n17152), .ZN(n13727) );
  OAI21_X1 U17044 ( .B1(n21256), .B2(n13728), .A(n13727), .ZN(P1_U3484) );
  INV_X1 U17045 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17046 ( .A1(n20541), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13729) );
  OAI21_X1 U17047 ( .B1(n13844), .B2(n20502), .A(n13729), .ZN(P2_U2927) );
  AOI22_X1 U17048 ( .A1(n20541), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13730) );
  OAI21_X1 U17049 ( .B1(n16504), .B2(n20502), .A(n13730), .ZN(P2_U2926) );
  INV_X1 U17050 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n16481) );
  AOI22_X1 U17051 ( .A1(n20541), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13731) );
  OAI21_X1 U17052 ( .B1(n16481), .B2(n20502), .A(n13731), .ZN(P2_U2923) );
  INV_X1 U17053 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13733) );
  AOI22_X1 U17054 ( .A1(n20541), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13732) );
  OAI21_X1 U17055 ( .B1(n13733), .B2(n20502), .A(n13732), .ZN(P2_U2934) );
  AOI22_X1 U17056 ( .A1(n20541), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13734) );
  OAI21_X1 U17057 ( .B1(n16495), .B2(n20502), .A(n13734), .ZN(P2_U2925) );
  AOI22_X1 U17058 ( .A1(n20541), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13735) );
  OAI21_X1 U17059 ( .B1(n16487), .B2(n20502), .A(n13735), .ZN(P2_U2924) );
  INV_X1 U17060 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13834) );
  AOI22_X1 U17061 ( .A1(n20541), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13736) );
  OAI21_X1 U17062 ( .B1(n13834), .B2(n20502), .A(n13736), .ZN(P2_U2935) );
  INV_X1 U17063 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13738) );
  AOI22_X1 U17064 ( .A1(n20541), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13737) );
  OAI21_X1 U17065 ( .B1(n13738), .B2(n20502), .A(n13737), .ZN(P2_U2933) );
  AOI22_X1 U17066 ( .A1(n20541), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13739) );
  OAI21_X1 U17067 ( .B1(n16522), .B2(n20502), .A(n13739), .ZN(P2_U2928) );
  NAND2_X1 U17068 ( .A1(n13741), .A2(n13740), .ZN(n13744) );
  INV_X1 U17069 ( .A(n13742), .ZN(n13743) );
  AND2_X1 U17070 ( .A1(n13744), .A2(n13743), .ZN(n14882) );
  INV_X1 U17071 ( .A(n13745), .ZN(n13758) );
  OAI21_X1 U17072 ( .B1(n17670), .B2(n13747), .A(n13746), .ZN(n13757) );
  NAND2_X1 U17073 ( .A1(n13749), .A2(n13748), .ZN(n13751) );
  INV_X1 U17074 ( .A(n13751), .ZN(n13750) );
  AOI22_X1 U17075 ( .A1(n16946), .A2(n12878), .B1(n16825), .B2(n13750), .ZN(
        n13754) );
  NAND2_X1 U17076 ( .A1(n13752), .A2(n13751), .ZN(n13753) );
  OAI211_X1 U17077 ( .C1(n17669), .C2(n13755), .A(n13754), .B(n13753), .ZN(
        n13756) );
  AOI211_X1 U17078 ( .C1(n17639), .C2(n13758), .A(n13757), .B(n13756), .ZN(
        n13759) );
  OAI21_X1 U17079 ( .B1(n14882), .B2(n17671), .A(n13759), .ZN(P2_U3044) );
  INV_X1 U17080 ( .A(n13760), .ZN(n13766) );
  INV_X1 U17081 ( .A(n13761), .ZN(n13764) );
  INV_X1 U17082 ( .A(n13762), .ZN(n13763) );
  NAND2_X1 U17083 ( .A1(n13764), .A2(n13763), .ZN(n13765) );
  NAND2_X1 U17084 ( .A1(n13766), .A2(n13765), .ZN(n20400) );
  INV_X1 U17085 ( .A(n12489), .ZN(n17707) );
  NAND2_X1 U17086 ( .A1(n17707), .A2(n13767), .ZN(n13768) );
  NOR2_X1 U17087 ( .A1(n17706), .A2(n13768), .ZN(n13769) );
  AOI21_X1 U17088 ( .B1(n17709), .B2(n17704), .A(n13769), .ZN(n15205) );
  NAND2_X1 U17089 ( .A1(n15205), .A2(n13770), .ZN(n13771) );
  NAND2_X1 U17090 ( .A1(n20475), .A2(n20573), .ZN(n16543) );
  INV_X1 U17091 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20546) );
  AND2_X1 U17092 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20975), .ZN(n13772) );
  OAI211_X1 U17093 ( .C1(n20547), .C2(n20546), .A(n11494), .B(n13772), .ZN(
        n13773) );
  INV_X1 U17094 ( .A(n13773), .ZN(n13774) );
  INV_X1 U17095 ( .A(n20477), .ZN(n20496) );
  NOR2_X1 U17096 ( .A1(n21207), .A2(n20400), .ZN(n20495) );
  AOI211_X1 U17097 ( .C1(n21207), .C2(n20400), .A(n20496), .B(n20495), .ZN(
        n13775) );
  AOI21_X1 U17098 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n20491), .A(n13775), .ZN(
        n13782) );
  AND2_X1 U17099 ( .A1(n20475), .A2(n13776), .ZN(n20442) );
  AND2_X1 U17100 ( .A1(n13778), .A2(n13777), .ZN(n13779) );
  INV_X1 U17101 ( .A(n15216), .ZN(n13780) );
  NAND2_X1 U17102 ( .A1(n16523), .A2(n13780), .ZN(n20468) );
  INV_X1 U17103 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n17850) );
  INV_X1 U17104 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19547) );
  AOI22_X1 U17105 ( .A1(n15214), .A2(n17850), .B1(n19547), .B2(n15215), .ZN(
        n20441) );
  NAND2_X1 U17106 ( .A1(n20468), .A2(n20441), .ZN(n13781) );
  OAI211_X1 U17107 ( .C1(n20400), .C2(n16543), .A(n13782), .B(n13781), .ZN(
        P2_U2919) );
  OAI21_X1 U17108 ( .B1(n20547), .B2(n21236), .A(n13783), .ZN(n13827) );
  INV_X1 U17109 ( .A(n13827), .ZN(n13918) );
  AOI22_X1 U17110 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13786) );
  AOI22_X1 U17111 ( .A1(n15214), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15215), .ZN(n20576) );
  INV_X1 U17112 ( .A(n20576), .ZN(n13785) );
  NAND2_X1 U17113 ( .A1(n13840), .A2(n13785), .ZN(n13828) );
  NAND2_X1 U17114 ( .A1(n13786), .A2(n13828), .ZN(P2_U2959) );
  AOI22_X1 U17115 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13787) );
  AOI22_X1 U17116 ( .A1(n15214), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15215), .ZN(n20566) );
  INV_X1 U17117 ( .A(n20566), .ZN(n16529) );
  NAND2_X1 U17118 ( .A1(n13840), .A2(n16529), .ZN(n13802) );
  NAND2_X1 U17119 ( .A1(n13787), .A2(n13802), .ZN(P2_U2957) );
  AOI22_X1 U17120 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U17121 ( .A1(n15214), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15215), .ZN(n20548) );
  INV_X1 U17122 ( .A(n20548), .ZN(n15217) );
  NAND2_X1 U17123 ( .A1(n13840), .A2(n15217), .ZN(n13795) );
  NAND2_X1 U17124 ( .A1(n13788), .A2(n13795), .ZN(P2_U2953) );
  AOI22_X1 U17125 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13789) );
  INV_X1 U17126 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17843) );
  INV_X1 U17127 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19560) );
  AOI22_X1 U17128 ( .A1(n15214), .A2(n17843), .B1(n19560), .B2(n15215), .ZN(
        n20553) );
  NAND2_X1 U17129 ( .A1(n13840), .A2(n20553), .ZN(n13797) );
  NAND2_X1 U17130 ( .A1(n13789), .A2(n13797), .ZN(P2_U2954) );
  AOI22_X1 U17131 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13790) );
  AOI22_X1 U17132 ( .A1(n15214), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15215), .ZN(n20558) );
  INV_X1 U17133 ( .A(n20558), .ZN(n16536) );
  NAND2_X1 U17134 ( .A1(n13840), .A2(n16536), .ZN(n13799) );
  NAND2_X1 U17135 ( .A1(n13790), .A2(n13799), .ZN(P2_U2955) );
  AOI22_X1 U17136 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13827), .B1(n13830), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13791) );
  INV_X1 U17137 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n17837) );
  INV_X1 U17138 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n19577) );
  AOI22_X1 U17139 ( .A1(n15214), .A2(n17837), .B1(n19577), .B2(n15215), .ZN(
        n17484) );
  NAND2_X1 U17140 ( .A1(n13840), .A2(n17484), .ZN(n13793) );
  NAND2_X1 U17141 ( .A1(n13791), .A2(n13793), .ZN(P2_U2973) );
  AOI22_X1 U17142 ( .A1(P2_UWORD_REG_14__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n13792) );
  AOI22_X1 U17143 ( .A1(n15214), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n15215), .ZN(n20453) );
  INV_X1 U17144 ( .A(n20453), .ZN(n15412) );
  NAND2_X1 U17145 ( .A1(n13840), .A2(n15412), .ZN(n13825) );
  NAND2_X1 U17146 ( .A1(n13792), .A2(n13825), .ZN(P2_U2966) );
  AOI22_X1 U17147 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13794) );
  NAND2_X1 U17148 ( .A1(n13794), .A2(n13793), .ZN(P2_U2958) );
  AOI22_X1 U17149 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n13827), .B1(n13830), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13796) );
  NAND2_X1 U17150 ( .A1(n13796), .A2(n13795), .ZN(P2_U2968) );
  AOI22_X1 U17151 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n13827), .B1(n13830), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13798) );
  NAND2_X1 U17152 ( .A1(n13798), .A2(n13797), .ZN(P2_U2969) );
  AOI22_X1 U17153 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n13827), .B1(n13830), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13800) );
  NAND2_X1 U17154 ( .A1(n13800), .A2(n13799), .ZN(P2_U2970) );
  AOI22_X1 U17155 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n13827), .B1(n13830), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13801) );
  OAI22_X1 U17156 ( .A1(n15215), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n15214), .ZN(n20561) );
  INV_X1 U17157 ( .A(n20561), .ZN(n17491) );
  NAND2_X1 U17158 ( .A1(n13840), .A2(n17491), .ZN(n13817) );
  NAND2_X1 U17159 ( .A1(n13801), .A2(n13817), .ZN(P2_U2971) );
  AOI22_X1 U17160 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n13827), .B1(n13830), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13803) );
  NAND2_X1 U17161 ( .A1(n13803), .A2(n13802), .ZN(P2_U2972) );
  AOI22_X1 U17162 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13807) );
  INV_X1 U17163 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n13804) );
  NOR2_X1 U17164 ( .A1(n15214), .A2(n13804), .ZN(n13805) );
  AOI21_X1 U17165 ( .B1(BUF1_REG_9__SCAN_IN), .B2(n15214), .A(n13805), .ZN(
        n20466) );
  INV_X1 U17166 ( .A(n20466), .ZN(n13806) );
  NAND2_X1 U17167 ( .A1(n13840), .A2(n13806), .ZN(n13815) );
  NAND2_X1 U17168 ( .A1(n13807), .A2(n13815), .ZN(P2_U2961) );
  AOI22_X1 U17169 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13810) );
  NOR2_X1 U17170 ( .A1(n15214), .A2(n18838), .ZN(n13808) );
  AOI21_X1 U17171 ( .B1(BUF1_REG_13__SCAN_IN), .B2(n15214), .A(n13808), .ZN(
        n20456) );
  INV_X1 U17172 ( .A(n20456), .ZN(n13809) );
  NAND2_X1 U17173 ( .A1(n13840), .A2(n13809), .ZN(n13823) );
  NAND2_X1 U17174 ( .A1(n13810), .A2(n13823), .ZN(P2_U2965) );
  AOI22_X1 U17175 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n13814) );
  INV_X1 U17176 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n13811) );
  NOR2_X1 U17177 ( .A1(n15214), .A2(n13811), .ZN(n13812) );
  AOI21_X1 U17178 ( .B1(BUF1_REG_11__SCAN_IN), .B2(n15214), .A(n13812), .ZN(
        n20461) );
  INV_X1 U17179 ( .A(n20461), .ZN(n13813) );
  NAND2_X1 U17180 ( .A1(n13840), .A2(n13813), .ZN(n13819) );
  NAND2_X1 U17181 ( .A1(n13814), .A2(n13819), .ZN(P2_U2963) );
  AOI22_X1 U17182 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n13827), .B1(n13830), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13816) );
  NAND2_X1 U17183 ( .A1(n13816), .A2(n13815), .ZN(P2_U2976) );
  AOI22_X1 U17184 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13818) );
  NAND2_X1 U17185 ( .A1(n13818), .A2(n13817), .ZN(P2_U2956) );
  AOI22_X1 U17186 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13820) );
  NAND2_X1 U17187 ( .A1(n13820), .A2(n13819), .ZN(P2_U2978) );
  AOI22_X1 U17188 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n13822) );
  AOI22_X1 U17189 ( .A1(n15214), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n15215), .ZN(n20459) );
  INV_X1 U17190 ( .A(n20459), .ZN(n13821) );
  NAND2_X1 U17191 ( .A1(n13840), .A2(n13821), .ZN(n13831) );
  NAND2_X1 U17192 ( .A1(n13822), .A2(n13831), .ZN(P2_U2979) );
  AOI22_X1 U17193 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13824) );
  NAND2_X1 U17194 ( .A1(n13824), .A2(n13823), .ZN(P2_U2980) );
  AOI22_X1 U17195 ( .A1(P2_LWORD_REG_14__SCAN_IN), .A2(n13827), .B1(n13830), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n13826) );
  NAND2_X1 U17196 ( .A1(n13826), .A2(n13825), .ZN(P2_U2981) );
  AOI22_X1 U17197 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13827), .B1(n13830), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13829) );
  NAND2_X1 U17198 ( .A1(n13829), .A2(n13828), .ZN(P2_U2974) );
  AOI22_X1 U17199 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n13845), .B1(n13830), 
        .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n13832) );
  NAND2_X1 U17200 ( .A1(n13832), .A2(n13831), .ZN(P2_U2964) );
  INV_X1 U17201 ( .A(n13840), .ZN(n13917) );
  INV_X1 U17202 ( .A(n20441), .ZN(n14387) );
  INV_X1 U17203 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13833) );
  OAI222_X1 U17204 ( .A1(n13917), .A2(n14387), .B1(n13920), .B2(n13834), .C1(
        n13833), .C2(n13918), .ZN(P2_U2952) );
  NAND2_X1 U17205 ( .A1(n15215), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13836) );
  INV_X1 U17206 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17829) );
  OR2_X1 U17207 ( .A1(n15215), .A2(n17829), .ZN(n13835) );
  NAND2_X1 U17208 ( .A1(n13836), .A2(n13835), .ZN(n20463) );
  NAND2_X1 U17209 ( .A1(n13840), .A2(n20463), .ZN(n13847) );
  NAND2_X1 U17210 ( .A1(n13845), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13837) );
  OAI211_X1 U17211 ( .C1(n16495), .C2(n13920), .A(n13847), .B(n13837), .ZN(
        P2_U2962) );
  INV_X1 U17212 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20523) );
  NAND2_X1 U17213 ( .A1(n15215), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13839) );
  INV_X1 U17214 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17833) );
  OR2_X1 U17215 ( .A1(n15215), .A2(n17833), .ZN(n13838) );
  NAND2_X1 U17216 ( .A1(n13839), .A2(n13838), .ZN(n20469) );
  NAND2_X1 U17217 ( .A1(n13840), .A2(n20469), .ZN(n13843) );
  NAND2_X1 U17218 ( .A1(n13845), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13841) );
  OAI211_X1 U17219 ( .C1(n20523), .C2(n13920), .A(n13843), .B(n13841), .ZN(
        P2_U2975) );
  NAND2_X1 U17220 ( .A1(n13845), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13842) );
  OAI211_X1 U17221 ( .C1(n13844), .C2(n13920), .A(n13843), .B(n13842), .ZN(
        P2_U2960) );
  INV_X1 U17222 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20519) );
  NAND2_X1 U17223 ( .A1(n13845), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13846) );
  OAI211_X1 U17224 ( .C1(n20519), .C2(n13920), .A(n13847), .B(n13846), .ZN(
        P2_U2977) );
  MUX2_X1 U17225 ( .A(n20397), .B(n20403), .S(n20437), .Z(n13848) );
  OAI21_X1 U17226 ( .B1(n20428), .B2(n21207), .A(n13848), .ZN(P2_U2887) );
  OR2_X1 U17227 ( .A1(n17186), .A2(n21541), .ZN(n13849) );
  AOI21_X1 U17228 ( .B1(n17128), .B2(n12633), .A(n13849), .ZN(n13850) );
  NAND2_X1 U17229 ( .A1(n17170), .A2(n13850), .ZN(n13855) );
  OR2_X1 U17230 ( .A1(n13851), .A2(n14058), .ZN(n13852) );
  AND2_X1 U17231 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  OAI211_X1 U17232 ( .C1(n17170), .C2(n13856), .A(n13855), .B(n13854), .ZN(
        n13857) );
  INV_X1 U17233 ( .A(n13857), .ZN(n13863) );
  OAI21_X1 U17234 ( .B1(n13859), .B2(n21541), .A(n13858), .ZN(n13862) );
  NOR3_X1 U17235 ( .A1(n14116), .A2(n13860), .A3(n21541), .ZN(n13861) );
  AOI21_X1 U17236 ( .B1(n17170), .B2(n13862), .A(n13861), .ZN(n13992) );
  AND2_X1 U17237 ( .A1(n13863), .A2(n13992), .ZN(n17136) );
  NOR2_X1 U17238 ( .A1(n21438), .A2(n21441), .ZN(n14032) );
  NAND2_X1 U17239 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14032), .ZN(n17399) );
  INV_X1 U17240 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21255) );
  OAI22_X1 U17241 ( .A1(n17136), .A2(n21248), .B1(n17399), .B2(n21255), .ZN(
        n17391) );
  AND2_X1 U17242 ( .A1(n21439), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13864) );
  INV_X1 U17243 ( .A(n21526), .ZN(n13913) );
  NAND4_X1 U17244 ( .A1(n12633), .A2(n14116), .A3(n13989), .A4(n13866), .ZN(
        n13867) );
  NOR2_X1 U17245 ( .A1(n13867), .A2(n13883), .ZN(n14086) );
  OR2_X1 U17246 ( .A1(n13865), .A2(n14086), .ZN(n13874) );
  INV_X1 U17247 ( .A(n14112), .ZN(n13869) );
  INV_X1 U17248 ( .A(n13885), .ZN(n13884) );
  NAND3_X1 U17249 ( .A1(n13870), .A2(n13869), .A3(n13884), .ZN(n13871) );
  OAI21_X1 U17250 ( .B1(n17128), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13871), .ZN(n13872) );
  INV_X1 U17251 ( .A(n13872), .ZN(n13873) );
  NAND2_X1 U17252 ( .A1(n13874), .A2(n13873), .ZN(n17131) );
  NOR2_X1 U17253 ( .A1(n21438), .A2(n14158), .ZN(n13892) );
  INV_X1 U17254 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U17255 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13876), .B2(n13875), .ZN(
        n13893) );
  INV_X1 U17256 ( .A(n13893), .ZN(n13877) );
  AND2_X1 U17257 ( .A1(n13892), .A2(n13877), .ZN(n13879) );
  NOR3_X1 U17258 ( .A1(n14112), .A2(n13885), .A3(n14033), .ZN(n13878) );
  AOI211_X1 U17259 ( .C1(n17131), .C2(n21523), .A(n13879), .B(n13878), .ZN(
        n13881) );
  NAND2_X1 U17260 ( .A1(n13913), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13880) );
  OAI21_X1 U17261 ( .B1(n13913), .B2(n13881), .A(n13880), .ZN(P1_U3473) );
  OR2_X1 U17262 ( .A1(n16326), .A2(n14086), .ZN(n13890) );
  NAND2_X1 U17263 ( .A1(n13989), .A2(n13955), .ZN(n13882) );
  NOR2_X1 U17264 ( .A1(n13883), .A2(n13882), .ZN(n14097) );
  NAND2_X1 U17265 ( .A1(n13884), .A2(n10358), .ZN(n14092) );
  NAND2_X1 U17266 ( .A1(n13885), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14088) );
  AND2_X1 U17267 ( .A1(n14092), .A2(n14088), .ZN(n13891) );
  XNOR2_X1 U17268 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13887) );
  NAND2_X1 U17269 ( .A1(n13954), .A2(n13886), .ZN(n14093) );
  OAI22_X1 U17270 ( .A1(n17128), .A2(n13887), .B1(n13891), .B2(n14093), .ZN(
        n13888) );
  AOI21_X1 U17271 ( .B1(n14097), .B2(n13891), .A(n13888), .ZN(n13889) );
  AND2_X1 U17272 ( .A1(n13890), .A2(n13889), .ZN(n14104) );
  INV_X1 U17273 ( .A(n14104), .ZN(n13894) );
  INV_X1 U17274 ( .A(n14033), .ZN(n21521) );
  AOI222_X1 U17275 ( .A1(n13894), .A2(n21523), .B1(n13893), .B2(n13892), .C1(
        n21521), .C2(n13891), .ZN(n13896) );
  NAND2_X1 U17276 ( .A1(n13913), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13895) );
  OAI21_X1 U17277 ( .B1(n13913), .B2(n13896), .A(n13895), .ZN(P1_U3472) );
  MUX2_X1 U17278 ( .A(n9970), .B(n14878), .S(n17479), .Z(n13899) );
  OAI21_X1 U17279 ( .B1(n21190), .B2(n20428), .A(n13899), .ZN(P2_U2885) );
  INV_X1 U17280 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14952) );
  MUX2_X1 U17281 ( .A(n14952), .B(n16918), .S(n20437), .Z(n13902) );
  OAI21_X1 U17282 ( .B1(n16968), .B2(n20428), .A(n13902), .ZN(P2_U2886) );
  INV_X1 U17283 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14781) );
  NOR2_X1 U17284 ( .A1(n20437), .A2(n14781), .ZN(n13908) );
  AOI21_X1 U17285 ( .B1(n12900), .B2(n13216), .A(n13908), .ZN(n13909) );
  OAI21_X1 U17286 ( .B1(n20800), .B2(n20428), .A(n13909), .ZN(P2_U2884) );
  INV_X1 U17287 ( .A(n17128), .ZN(n13922) );
  AOI21_X1 U17288 ( .B1(n13922), .B2(n21523), .A(n13913), .ZN(n13914) );
  OAI22_X1 U17289 ( .A1(n10634), .A2(n14086), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13910), .ZN(n17130) );
  OAI22_X1 U17290 ( .A1(n21438), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14033), .ZN(n13911) );
  AOI21_X1 U17291 ( .B1(n17130), .B2(n21523), .A(n13911), .ZN(n13912) );
  OAI22_X1 U17292 ( .A1(n13914), .A2(n17127), .B1(n13913), .B2(n13912), .ZN(
        P1_U3474) );
  INV_X1 U17293 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13916) );
  INV_X1 U17294 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13915) );
  OAI222_X1 U17295 ( .A1(n13916), .A2(n13920), .B1(n13915), .B2(n13918), .C1(
        n13917), .C2(n14387), .ZN(P2_U2967) );
  INV_X1 U17296 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13919) );
  AOI22_X1 U17297 ( .A1(n15214), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15215), .ZN(n20450) );
  OAI222_X1 U17298 ( .A1(n13921), .A2(n13920), .B1(n13919), .B2(n13918), .C1(
        n13917), .C2(n20450), .ZN(P2_U2982) );
  INV_X1 U17299 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14486) );
  NAND3_X1 U17300 ( .A1(n17170), .A2(n13993), .A3(n13922), .ZN(n13923) );
  OAI21_X1 U17301 ( .B1(n13985), .B2(n17165), .A(n13923), .ZN(n13925) );
  NAND2_X1 U17302 ( .A1(n21392), .A2(n15100), .ZN(n14402) );
  INV_X1 U17303 ( .A(n14032), .ZN(n17396) );
  OR2_X1 U17304 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17396), .ZN(n21540) );
  INV_X2 U17305 ( .A(n21540), .ZN(n21410) );
  NOR2_X4 U17306 ( .A1(n21392), .A2(n21410), .ZN(n21407) );
  AOI22_X1 U17307 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n21407), .B1(n21410), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13926) );
  OAI21_X1 U17308 ( .B1(n14486), .B2(n14402), .A(n13926), .ZN(P1_U2910) );
  INV_X1 U17309 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14423) );
  AOI22_X1 U17310 ( .A1(n21410), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13927) );
  OAI21_X1 U17311 ( .B1(n14423), .B2(n14402), .A(n13927), .ZN(P1_U2908) );
  INV_X1 U17312 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14470) );
  AOI22_X1 U17313 ( .A1(n21410), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13928) );
  OAI21_X1 U17314 ( .B1(n14470), .B2(n14402), .A(n13928), .ZN(P1_U2911) );
  INV_X1 U17315 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U17316 ( .A1(n21410), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13929) );
  OAI21_X1 U17317 ( .B1(n14448), .B2(n14402), .A(n13929), .ZN(P1_U2913) );
  XNOR2_X1 U17318 ( .A(n13930), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13934) );
  OR2_X1 U17319 ( .A1(n9930), .A2(n13931), .ZN(n13932) );
  NAND2_X1 U17320 ( .A1(n13932), .A2(n13963), .ZN(n20342) );
  MUX2_X1 U17321 ( .A(n11874), .B(n20342), .S(n20437), .Z(n13933) );
  OAI21_X1 U17322 ( .B1(n13934), .B2(n20428), .A(n13933), .ZN(P2_U2880) );
  XNOR2_X1 U17323 ( .A(n21190), .B(n14882), .ZN(n13941) );
  XNOR2_X1 U17324 ( .A(n13935), .B(n13936), .ZN(n21201) );
  INV_X1 U17325 ( .A(n21201), .ZN(n13937) );
  NAND2_X1 U17326 ( .A1(n16968), .A2(n13937), .ZN(n13938) );
  OAI21_X1 U17327 ( .B1(n16968), .B2(n13937), .A(n13938), .ZN(n20494) );
  NOR2_X1 U17328 ( .A1(n20494), .A2(n20495), .ZN(n20493) );
  INV_X1 U17329 ( .A(n13938), .ZN(n13939) );
  NOR2_X1 U17330 ( .A1(n20493), .A2(n13939), .ZN(n13940) );
  NOR2_X1 U17331 ( .A1(n13940), .A2(n13941), .ZN(n14356) );
  AOI21_X1 U17332 ( .B1(n13941), .B2(n13940), .A(n14356), .ZN(n13944) );
  AOI22_X1 U17333 ( .A1(n20468), .A2(n20553), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n20491), .ZN(n13943) );
  INV_X1 U17334 ( .A(n14882), .ZN(n21192) );
  NAND2_X1 U17335 ( .A1(n21192), .A2(n20492), .ZN(n13942) );
  OAI211_X1 U17336 ( .C1(n13944), .C2(n20496), .A(n13943), .B(n13942), .ZN(
        P2_U2917) );
  NOR2_X1 U17337 ( .A1(n13945), .A2(n13946), .ZN(n13948) );
  INV_X1 U17338 ( .A(n13930), .ZN(n13947) );
  OAI211_X1 U17339 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13948), .A(
        n13947), .B(n20435), .ZN(n13950) );
  NAND2_X1 U17340 ( .A1(n13216), .A2(n20355), .ZN(n13949) );
  OAI211_X1 U17341 ( .C1(n13216), .C2(n20348), .A(n13950), .B(n13949), .ZN(
        P2_U2881) );
  INV_X1 U17342 ( .A(n13951), .ZN(n13952) );
  OAI21_X1 U17343 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13953), .A(
        n13952), .ZN(n21425) );
  INV_X1 U17344 ( .A(n13954), .ZN(n13957) );
  INV_X1 U17345 ( .A(n15373), .ZN(n15425) );
  AND3_X1 U17346 ( .A1(n15425), .A2(n10532), .A3(n10488), .ZN(n13990) );
  NAND3_X1 U17347 ( .A1(n13990), .A2(n15374), .A3(n13955), .ZN(n13956) );
  OAI21_X1 U17348 ( .B1(n17170), .B2(n13957), .A(n13956), .ZN(n13959) );
  INV_X1 U17349 ( .A(n13960), .ZN(n13961) );
  XNOR2_X1 U17350 ( .A(n13962), .B(n13961), .ZN(n15133) );
  INV_X1 U17351 ( .A(n15133), .ZN(n14165) );
  OAI222_X1 U17352 ( .A1(n21425), .A2(n15641), .B1(n12671), .B2(n21381), .C1(
        n17250), .C2(n14165), .ZN(P1_U2872) );
  NAND2_X1 U17353 ( .A1(n13964), .A2(n13963), .ZN(n13965) );
  INV_X1 U17354 ( .A(n17641), .ZN(n20331) );
  INV_X1 U17355 ( .A(n13967), .ZN(n13972) );
  INV_X1 U17356 ( .A(n13968), .ZN(n13971) );
  OAI211_X1 U17357 ( .C1(n13972), .C2(n13971), .A(n20435), .B(n10299), .ZN(
        n13974) );
  NAND2_X1 U17358 ( .A1(n17479), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13973) );
  OAI211_X1 U17359 ( .C1(n20331), .C2(n17479), .A(n13974), .B(n13973), .ZN(
        P2_U2879) );
  INV_X1 U17360 ( .A(n13975), .ZN(n13976) );
  AOI21_X1 U17361 ( .B1(n13977), .B2(n13995), .A(n13976), .ZN(n21358) );
  INV_X1 U17362 ( .A(n21358), .ZN(n14004) );
  OR2_X1 U17363 ( .A1(n13979), .A2(n13978), .ZN(n13980) );
  AND2_X1 U17364 ( .A1(n13980), .A2(n14151), .ZN(n21344) );
  INV_X1 U17365 ( .A(n21381), .ZN(n15643) );
  AOI22_X1 U17366 ( .A1(n21376), .A2(n21344), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n15643), .ZN(n13981) );
  OAI21_X1 U17367 ( .B1(n14004), .B2(n17250), .A(n13981), .ZN(P1_U2870) );
  INV_X1 U17368 ( .A(n13985), .ZN(n13983) );
  NAND2_X1 U17369 ( .A1(n21543), .A2(n21541), .ZN(n13982) );
  INV_X1 U17370 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n21394) );
  NOR3_X2 U17371 ( .A1(n13985), .A2(n13984), .A3(n21541), .ZN(n21422) );
  INV_X1 U17372 ( .A(DATAI_10_), .ZN(n13987) );
  NAND2_X1 U17373 ( .A1(n15371), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13986) );
  OAI21_X1 U17374 ( .B1(n15371), .B2(n13987), .A(n13986), .ZN(n15665) );
  NAND2_X1 U17375 ( .A1(n21422), .A2(n15665), .ZN(n14484) );
  NOR2_X1 U17376 ( .A1(n14483), .A2(n17165), .ZN(n21420) );
  NAND2_X1 U17377 ( .A1(n21420), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n13988) );
  OAI211_X1 U17378 ( .C1(n14553), .C2(n21394), .A(n14484), .B(n13988), .ZN(
        P1_U2962) );
  NAND2_X1 U17379 ( .A1(n9960), .A2(n13990), .ZN(n13991) );
  NAND2_X1 U17380 ( .A1(n13992), .A2(n13991), .ZN(n13994) );
  NAND2_X1 U17381 ( .A1(n10514), .A2(n15373), .ZN(n13998) );
  OAI21_X1 U17382 ( .B1(n13997), .B2(n13996), .A(n13995), .ZN(n15120) );
  INV_X1 U17383 ( .A(DATAI_1_), .ZN(n14000) );
  NAND2_X1 U17384 ( .A1(n15371), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13999) );
  OAI21_X1 U17385 ( .B1(n15371), .B2(n14000), .A(n13999), .ZN(n15376) );
  AOI22_X1 U17386 ( .A1(n15737), .A2(n15376), .B1(P1_EAX_REG_1__SCAN_IN), .B2(
        n15736), .ZN(n14001) );
  OAI21_X1 U17387 ( .B1(n15739), .B2(n15120), .A(n14001), .ZN(P1_U2903) );
  INV_X1 U17388 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n21409) );
  NAND2_X1 U17389 ( .A1(n14552), .A2(DATAI_2_), .ZN(n14003) );
  NAND2_X1 U17390 ( .A1(n15371), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14002) );
  AND2_X1 U17391 ( .A1(n14003), .A2(n14002), .ZN(n14457) );
  OAI222_X1 U17392 ( .A1(n15739), .A2(n14004), .B1(n15733), .B2(n21409), .C1(
        n15732), .C2(n14457), .ZN(P1_U2902) );
  XNOR2_X1 U17393 ( .A(n13970), .B(n20427), .ZN(n14010) );
  OR2_X1 U17394 ( .A1(n14006), .A2(n14005), .ZN(n14007) );
  AND2_X1 U17395 ( .A1(n14007), .A2(n16687), .ZN(n20316) );
  NOR2_X1 U17396 ( .A1(n13216), .A2(n10232), .ZN(n14008) );
  AOI21_X1 U17397 ( .B1(n20316), .B2(n13216), .A(n14008), .ZN(n14009) );
  OAI21_X1 U17398 ( .B1(n14010), .B2(n20428), .A(n14009), .ZN(P2_U2878) );
  NAND2_X1 U17399 ( .A1(n20800), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20700) );
  NOR2_X1 U17400 ( .A1(n20700), .A2(n20970), .ZN(n21176) );
  NOR2_X1 U17401 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20972), .ZN(
        n14019) );
  NOR2_X1 U17402 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12040), .ZN(n21237) );
  NOR2_X1 U17403 ( .A1(n14011), .A2(n21237), .ZN(n17729) );
  INV_X1 U17404 ( .A(n17729), .ZN(n21234) );
  AND2_X1 U17405 ( .A1(n21234), .A2(n21205), .ZN(n14012) );
  OAI21_X1 U17406 ( .B1(n21176), .B2(n14019), .A(n21023), .ZN(n14017) );
  INV_X1 U17407 ( .A(n14649), .ZN(n20868) );
  NAND2_X1 U17408 ( .A1(n12896), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20699) );
  INV_X1 U17409 ( .A(n20699), .ZN(n14379) );
  NAND2_X1 U17410 ( .A1(n20868), .A2(n14379), .ZN(n20771) );
  AND2_X1 U17411 ( .A1(n20771), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14013) );
  NAND2_X1 U17412 ( .A1(n14014), .A2(n14013), .ZN(n14021) );
  NAND2_X1 U17413 ( .A1(n20771), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14015) );
  NAND2_X1 U17414 ( .A1(n14021), .A2(n14015), .ZN(n14016) );
  OR2_X1 U17415 ( .A1(n14017), .A2(n14016), .ZN(n20765) );
  INV_X1 U17416 ( .A(n21207), .ZN(n20407) );
  INV_X1 U17417 ( .A(n20796), .ZN(n20759) );
  AOI22_X1 U17418 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20572), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20571), .ZN(n21006) );
  NOR2_X2 U17419 ( .A1(n20970), .A2(n20672), .ZN(n20764) );
  AOI22_X1 U17420 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20571), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n20572), .ZN(n21069) );
  AOI22_X1 U17421 ( .A1(n20759), .A2(n21066), .B1(n20764), .B2(n21003), .ZN(
        n14026) );
  INV_X1 U17422 ( .A(n14019), .ZN(n14023) );
  INV_X1 U17423 ( .A(n14020), .ZN(n20588) );
  INV_X1 U17424 ( .A(n14021), .ZN(n14022) );
  AOI211_X2 U17425 ( .C1(n14023), .C2(n21225), .A(n20588), .B(n14022), .ZN(
        n20763) );
  INV_X1 U17426 ( .A(n17484), .ZN(n20473) );
  NOR2_X2 U17427 ( .A1(n20473), .A2(n20977), .ZN(n21065) );
  INV_X1 U17428 ( .A(n20771), .ZN(n20774) );
  NOR2_X1 U17429 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20975), .ZN(n17735) );
  NOR2_X2 U17430 ( .A1(n20574), .A2(n11494), .ZN(n21064) );
  AOI22_X1 U17431 ( .A1(n20763), .A2(n21065), .B1(n20774), .B2(n21064), .ZN(
        n14025) );
  OAI211_X1 U17432 ( .C1(n20762), .C2(n14027), .A(n14026), .B(n14025), .ZN(
        P2_U3110) );
  NAND3_X1 U17433 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17143), .A3(
        n17132), .ZN(n14791) );
  INV_X1 U17434 ( .A(n14791), .ZN(n14035) );
  NOR2_X1 U17435 ( .A1(n16322), .A2(n14173), .ZN(n14560) );
  NAND2_X1 U17436 ( .A1(n14560), .A2(n14561), .ZN(n14038) );
  OR2_X1 U17437 ( .A1(n16326), .A2(n14113), .ZN(n14832) );
  INV_X1 U17438 ( .A(n14832), .ZN(n14031) );
  INV_X1 U17439 ( .A(n14030), .ZN(n14319) );
  NOR2_X1 U17440 ( .A1(n14318), .A2(n14791), .ZN(n14080) );
  AOI21_X1 U17441 ( .B1(n14031), .B2(n14319), .A(n14080), .ZN(n14037) );
  OAI211_X1 U17442 ( .C1(n14038), .C2(n21254), .A(n16320), .B(n14037), .ZN(
        n14034) );
  OAI21_X1 U17443 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_2__SCAN_IN), .A(n21439), .ZN(n21545) );
  OAI211_X1 U17444 ( .C1(n16320), .C2(n14035), .A(n14034), .B(n14702), .ZN(
        n14036) );
  INV_X1 U17445 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14041) );
  INV_X1 U17446 ( .A(n14865), .ZN(n14076) );
  NOR2_X2 U17447 ( .A1(n17306), .A2(n14552), .ZN(n14078) );
  NOR2_X2 U17448 ( .A1(n15371), .A2(n17306), .ZN(n14077) );
  AOI22_X1 U17449 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n14078), .B1(DATAI_17_), 
        .B2(n14077), .ZN(n15002) );
  INV_X1 U17450 ( .A(n15002), .ZN(n16339) );
  AND2_X1 U17451 ( .A1(n15376), .A2(n14637), .ZN(n16341) );
  OAI22_X1 U17452 ( .A1(n14037), .A2(n16334), .B1(n14791), .B2(n21441), .ZN(
        n14075) );
  AOI22_X1 U17453 ( .A1(n14076), .A2(n16339), .B1(n16341), .B2(n14075), .ZN(
        n14040) );
  NOR2_X2 U17454 ( .A1(n14038), .A2(n14562), .ZN(n14824) );
  AOI22_X1 U17455 ( .A1(DATAI_25_), .A2(n14077), .B1(BUF1_REG_25__SCAN_IN), 
        .B2(n14078), .ZN(n15012) );
  INV_X1 U17456 ( .A(n15012), .ZN(n16338) );
  NAND2_X1 U17457 ( .A1(n14079), .A2(n17165), .ZN(n15285) );
  AOI22_X1 U17458 ( .A1(n14824), .A2(n16338), .B1(n14080), .B2(n16340), .ZN(
        n14039) );
  OAI211_X1 U17459 ( .C1(n14084), .C2(n14041), .A(n14040), .B(n14039), .ZN(
        P1_U3074) );
  INV_X1 U17460 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14046) );
  AOI22_X1 U17461 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n14078), .B1(DATAI_22_), 
        .B2(n14077), .ZN(n15052) );
  INV_X1 U17462 ( .A(n15052), .ZN(n16356) );
  INV_X1 U17463 ( .A(DATAI_6_), .ZN(n14043) );
  NAND2_X1 U17464 ( .A1(n15371), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14042) );
  OAI21_X1 U17465 ( .B1(n15371), .B2(n14043), .A(n14042), .ZN(n15686) );
  AND2_X1 U17466 ( .A1(n15686), .A2(n14637), .ZN(n16362) );
  AOI22_X1 U17467 ( .A1(n14076), .A2(n16356), .B1(n16362), .B2(n14075), .ZN(
        n14045) );
  AOI22_X1 U17468 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n14078), .B1(DATAI_30_), 
        .B2(n14077), .ZN(n15054) );
  INV_X1 U17469 ( .A(n15054), .ZN(n16354) );
  NAND2_X1 U17470 ( .A1(n14079), .A2(n10488), .ZN(n15275) );
  AOI22_X1 U17471 ( .A1(n14824), .A2(n16354), .B1(n14080), .B2(n16360), .ZN(
        n14044) );
  OAI211_X1 U17472 ( .C1(n14084), .C2(n14046), .A(n14045), .B(n14044), .ZN(
        P1_U3079) );
  INV_X1 U17473 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U17474 ( .A1(DATAI_20_), .A2(n14077), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n14078), .ZN(n15046) );
  INV_X1 U17475 ( .A(n15046), .ZN(n16347) );
  INV_X1 U17476 ( .A(DATAI_4_), .ZN(n14048) );
  NAND2_X1 U17477 ( .A1(n15371), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14047) );
  OAI21_X1 U17478 ( .B1(n15371), .B2(n14048), .A(n14047), .ZN(n15698) );
  AND2_X1 U17479 ( .A1(n15698), .A2(n14637), .ZN(n16349) );
  AOI22_X1 U17480 ( .A1(n14076), .A2(n16347), .B1(n16349), .B2(n14075), .ZN(
        n14051) );
  AOI22_X1 U17481 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n14078), .B1(DATAI_28_), 
        .B2(n14077), .ZN(n15048) );
  INV_X1 U17482 ( .A(n15048), .ZN(n16346) );
  NAND2_X1 U17483 ( .A1(n14079), .A2(n14049), .ZN(n15280) );
  AOI22_X1 U17484 ( .A1(n14824), .A2(n16346), .B1(n14080), .B2(n16348), .ZN(
        n14050) );
  OAI211_X1 U17485 ( .C1(n14084), .C2(n14052), .A(n14051), .B(n14050), .ZN(
        P1_U3077) );
  INV_X1 U17486 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U17487 ( .A1(DATAI_23_), .A2(n14077), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n14078), .ZN(n15058) );
  INV_X1 U17488 ( .A(n15058), .ZN(n15289) );
  NAND2_X1 U17489 ( .A1(n14552), .A2(DATAI_7_), .ZN(n14054) );
  NAND2_X1 U17490 ( .A1(n15371), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14053) );
  AND2_X1 U17491 ( .A1(n14054), .A2(n14053), .ZN(n15681) );
  AOI22_X1 U17492 ( .A1(n14076), .A2(n15289), .B1(n14823), .B2(n14075), .ZN(
        n14056) );
  AOI22_X1 U17493 ( .A1(DATAI_31_), .A2(n14077), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n14078), .ZN(n15060) );
  INV_X1 U17494 ( .A(n15060), .ZN(n15293) );
  NAND2_X1 U17495 ( .A1(n14079), .A2(n15373), .ZN(n15291) );
  AOI22_X1 U17496 ( .A1(n14824), .A2(n15293), .B1(n14080), .B2(n15063), .ZN(
        n14055) );
  OAI211_X1 U17497 ( .C1(n14084), .C2(n14057), .A(n14056), .B(n14055), .ZN(
        P1_U3080) );
  INV_X1 U17498 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14061) );
  AOI22_X1 U17499 ( .A1(DATAI_18_), .A2(n14077), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n14078), .ZN(n15016) );
  INV_X1 U17500 ( .A(n15016), .ZN(n15311) );
  AOI22_X1 U17501 ( .A1(n14076), .A2(n15311), .B1(n14818), .B2(n14075), .ZN(
        n14060) );
  AOI22_X1 U17502 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n14078), .B1(DATAI_26_), 
        .B2(n14077), .ZN(n15018) );
  INV_X1 U17503 ( .A(n15018), .ZN(n15317) );
  NAND2_X1 U17504 ( .A1(n14079), .A2(n14058), .ZN(n15315) );
  AOI22_X1 U17505 ( .A1(n14824), .A2(n15317), .B1(n14080), .B2(n15021), .ZN(
        n14059) );
  OAI211_X1 U17506 ( .C1(n14084), .C2(n14061), .A(n14060), .B(n14059), .ZN(
        P1_U3075) );
  INV_X1 U17507 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14066) );
  AOI22_X1 U17508 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n14078), .B1(DATAI_21_), 
        .B2(n14077), .ZN(n15065) );
  INV_X1 U17509 ( .A(n15065), .ZN(n15296) );
  NAND2_X1 U17510 ( .A1(n14552), .A2(DATAI_5_), .ZN(n14063) );
  NAND2_X1 U17511 ( .A1(n15371), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14062) );
  AND2_X1 U17512 ( .A1(n14063), .A2(n14062), .ZN(n15694) );
  AOI22_X1 U17513 ( .A1(n14076), .A2(n15296), .B1(n14814), .B2(n14075), .ZN(
        n14065) );
  AOI22_X1 U17514 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n14078), .B1(DATAI_29_), 
        .B2(n14077), .ZN(n15067) );
  INV_X1 U17515 ( .A(n15067), .ZN(n15300) );
  NAND2_X1 U17516 ( .A1(n14079), .A2(n10487), .ZN(n15298) );
  AOI22_X1 U17517 ( .A1(n14824), .A2(n15300), .B1(n14080), .B2(n15070), .ZN(
        n14064) );
  OAI211_X1 U17518 ( .C1(n14084), .C2(n14066), .A(n14065), .B(n14064), .ZN(
        P1_U3078) );
  INV_X1 U17519 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14072) );
  AOI22_X1 U17520 ( .A1(DATAI_19_), .A2(n14077), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n14078), .ZN(n15072) );
  INV_X1 U17521 ( .A(n15072), .ZN(n15303) );
  NAND2_X1 U17522 ( .A1(n14552), .A2(DATAI_3_), .ZN(n14068) );
  NAND2_X1 U17523 ( .A1(n15371), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14067) );
  AND2_X1 U17524 ( .A1(n14068), .A2(n14067), .ZN(n15706) );
  AOI22_X1 U17525 ( .A1(n14076), .A2(n15303), .B1(n14810), .B2(n14075), .ZN(
        n14071) );
  AOI22_X1 U17526 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n14078), .B1(DATAI_27_), 
        .B2(n14077), .ZN(n15075) );
  INV_X1 U17527 ( .A(n15075), .ZN(n15307) );
  NAND2_X1 U17528 ( .A1(n14079), .A2(n14069), .ZN(n15305) );
  AOI22_X1 U17529 ( .A1(n14824), .A2(n15307), .B1(n14080), .B2(n15078), .ZN(
        n14070) );
  OAI211_X1 U17530 ( .C1(n14084), .C2(n14072), .A(n14071), .B(n14070), .ZN(
        P1_U3076) );
  INV_X1 U17531 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17532 ( .A1(DATAI_16_), .A2(n14077), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n14078), .ZN(n15023) );
  INV_X1 U17533 ( .A(n15023), .ZN(n15265) );
  NAND2_X1 U17534 ( .A1(n14552), .A2(DATAI_0_), .ZN(n14074) );
  NAND2_X1 U17535 ( .A1(n15371), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14073) );
  AND2_X1 U17536 ( .A1(n14074), .A2(n14073), .ZN(n14460) );
  AOI22_X1 U17537 ( .A1(n14076), .A2(n15265), .B1(n15271), .B2(n14075), .ZN(
        n14082) );
  AOI22_X1 U17538 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n14078), .B1(DATAI_24_), 
        .B2(n14077), .ZN(n15025) );
  INV_X1 U17539 ( .A(n15025), .ZN(n15266) );
  NAND2_X1 U17540 ( .A1(n14079), .A2(n15100), .ZN(n15269) );
  AOI22_X1 U17541 ( .A1(n14824), .A2(n15266), .B1(n14080), .B2(n15028), .ZN(
        n14081) );
  OAI211_X1 U17542 ( .C1(n14084), .C2(n14083), .A(n14082), .B(n14081), .ZN(
        P1_U3073) );
  INV_X1 U17543 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21415) );
  OAI222_X1 U17544 ( .A1(n15732), .A2(n14460), .B1(n15739), .B2(n14165), .C1(
        n21415), .C2(n15733), .ZN(P1_U2904) );
  NAND2_X1 U17545 ( .A1(n17136), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14101) );
  INV_X1 U17546 ( .A(n17136), .ZN(n14105) );
  INV_X1 U17547 ( .A(n14086), .ZN(n14087) );
  NAND2_X1 U17548 ( .A1(n15176), .A2(n14087), .ZN(n14099) );
  NAND2_X1 U17549 ( .A1(n14088), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14089) );
  NAND2_X1 U17550 ( .A1(n14090), .A2(n14089), .ZN(n21522) );
  XNOR2_X1 U17551 ( .A(n14091), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14095) );
  XNOR2_X1 U17552 ( .A(n14092), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14094) );
  OAI22_X1 U17553 ( .A1(n17128), .A2(n14095), .B1(n14094), .B2(n14093), .ZN(
        n14096) );
  AOI21_X1 U17554 ( .B1(n14097), .B2(n21522), .A(n14096), .ZN(n14098) );
  NAND2_X1 U17555 ( .A1(n14099), .A2(n14098), .ZN(n21524) );
  NAND2_X1 U17556 ( .A1(n14105), .A2(n21524), .ZN(n14100) );
  INV_X1 U17557 ( .A(n17142), .ZN(n17146) );
  NAND2_X1 U17558 ( .A1(n17146), .A2(n21438), .ZN(n14103) );
  NOR2_X1 U17559 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21438), .ZN(n14108) );
  NAND2_X1 U17560 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14108), .ZN(
        n14102) );
  NAND2_X1 U17561 ( .A1(n14103), .A2(n14102), .ZN(n14111) );
  NAND2_X1 U17562 ( .A1(n17136), .A2(n10358), .ZN(n14107) );
  NAND2_X1 U17563 ( .A1(n14105), .A2(n14104), .ZN(n14106) );
  AOI22_X1 U17564 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n14108), .B1(
        n21438), .B2(n17139), .ZN(n14109) );
  INV_X1 U17565 ( .A(n14109), .ZN(n14110) );
  NAND2_X1 U17566 ( .A1(n14111), .A2(n14110), .ZN(n17157) );
  NOR2_X1 U17567 ( .A1(n17157), .A2(n14112), .ZN(n14123) );
  NOR2_X1 U17568 ( .A1(n17136), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14117) );
  INV_X1 U17569 ( .A(n14113), .ZN(n14177) );
  INV_X1 U17570 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14114) );
  XNOR2_X1 U17571 ( .A(n14115), .B(n14114), .ZN(n21332) );
  OR2_X1 U17572 ( .A1(n21332), .A2(n14116), .ZN(n17389) );
  NAND2_X1 U17573 ( .A1(n14117), .A2(n17389), .ZN(n14120) );
  INV_X1 U17574 ( .A(n14117), .ZN(n14118) );
  NAND2_X1 U17575 ( .A1(n14118), .A2(n14114), .ZN(n14119) );
  OAI211_X1 U17576 ( .C1(n21438), .C2(n21255), .A(n14120), .B(n14119), .ZN(
        n17156) );
  INV_X1 U17577 ( .A(n17156), .ZN(n14122) );
  NOR3_X1 U17578 ( .A1(n14123), .A2(n14122), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n14121) );
  OAI21_X1 U17579 ( .B1(n14121), .B2(n17399), .A(n14564), .ZN(n21436) );
  NOR3_X1 U17580 ( .A1(n14123), .A2(n14122), .A3(n17396), .ZN(n17160) );
  AND2_X1 U17581 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n17400), .ZN(n16332) );
  OAI22_X1 U17582 ( .A1(n9807), .A2(n16334), .B1(n10634), .B2(n16332), .ZN(
        n14124) );
  OAI21_X1 U17583 ( .B1(n17160), .B2(n14124), .A(n21436), .ZN(n14125) );
  OAI21_X1 U17584 ( .B1(n21436), .B2(n14318), .A(n14125), .ZN(P1_U3478) );
  XNOR2_X1 U17585 ( .A(n9804), .B(n14126), .ZN(n14522) );
  OAI21_X1 U17586 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14617), .A(
        n15351), .ZN(n14132) );
  NAND3_X1 U17587 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17343), .A3(
        n11201), .ZN(n14130) );
  INV_X1 U17588 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21461) );
  NOR2_X1 U17589 ( .A1(n17352), .A2(n21461), .ZN(n14518) );
  AOI21_X1 U17590 ( .B1(n21427), .B2(n21344), .A(n14518), .ZN(n14129) );
  NAND3_X1 U17591 ( .A1(n14615), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n14145), .ZN(n14128) );
  NAND2_X1 U17592 ( .A1(n14615), .A2(n14149), .ZN(n14146) );
  NAND4_X1 U17593 ( .A1(n14130), .A2(n14129), .A3(n14128), .A4(n14146), .ZN(
        n14131) );
  AOI21_X1 U17594 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14132), .A(
        n14131), .ZN(n14133) );
  OAI21_X1 U17595 ( .B1(n17365), .B2(n14522), .A(n14133), .ZN(P1_U3029) );
  XOR2_X1 U17596 ( .A(n9805), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n14556) );
  XNOR2_X1 U17597 ( .A(n14136), .B(n14135), .ZN(n21374) );
  INV_X1 U17598 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21534) );
  OAI22_X1 U17599 ( .A1(n17364), .A2(n21374), .B1(n21534), .B2(n17352), .ZN(
        n14141) );
  NOR2_X1 U17600 ( .A1(n14138), .A2(n14137), .ZN(n14139) );
  OAI21_X1 U17601 ( .B1(n16220), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n15351), .ZN(n21431) );
  MUX2_X1 U17602 ( .A(n14139), .B(n21431), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n14140) );
  AOI211_X1 U17603 ( .C1(n21429), .C2(n14556), .A(n14141), .B(n14140), .ZN(
        n14142) );
  INV_X1 U17604 ( .A(n14142), .ZN(P1_U3030) );
  XNOR2_X1 U17605 ( .A(n14144), .B(n14143), .ZN(n14527) );
  OAI21_X1 U17606 ( .B1(n14617), .B2(n14145), .A(n15351), .ZN(n15383) );
  INV_X1 U17607 ( .A(n15383), .ZN(n14147) );
  NAND2_X1 U17608 ( .A1(n14147), .A2(n14146), .ZN(n14371) );
  NOR2_X1 U17609 ( .A1(n14149), .A2(n14148), .ZN(n14620) );
  AOI22_X1 U17610 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14371), .B1(
        n14620), .B2(n14368), .ZN(n14154) );
  NAND2_X1 U17611 ( .A1(n14151), .A2(n14150), .ZN(n14152) );
  AND2_X1 U17612 ( .A1(n14373), .A2(n14152), .ZN(n15173) );
  INV_X1 U17613 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21463) );
  NOR2_X1 U17614 ( .A1(n17352), .A2(n21463), .ZN(n14523) );
  AOI21_X1 U17615 ( .B1(n21427), .B2(n15173), .A(n14523), .ZN(n14153) );
  OAI211_X1 U17616 ( .C1(n17365), .C2(n14527), .A(n14154), .B(n14153), .ZN(
        P1_U3028) );
  INV_X1 U17617 ( .A(n14155), .ZN(n14159) );
  INV_X1 U17618 ( .A(n14156), .ZN(n14157) );
  AOI21_X1 U17619 ( .B1(n14159), .B2(n14158), .A(n14157), .ZN(n21428) );
  NAND2_X1 U17620 ( .A1(n17369), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n21434) );
  INV_X1 U17621 ( .A(n21434), .ZN(n14160) );
  AOI21_X1 U17622 ( .B1(n21428), .B2(n17267), .A(n14160), .ZN(n14164) );
  OAI21_X1 U17623 ( .B1(n14161), .B2(n14162), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14163) );
  OAI211_X1 U17624 ( .C1(n14165), .C2(n17306), .A(n14164), .B(n14163), .ZN(
        P1_U2999) );
  INV_X1 U17625 ( .A(n14166), .ZN(n14167) );
  NOR2_X1 U17626 ( .A1(n14168), .A2(n14167), .ZN(n14171) );
  INV_X1 U17627 ( .A(n14169), .ZN(n14170) );
  AOI21_X1 U17628 ( .B1(n14171), .B2(n13975), .A(n14170), .ZN(n15185) );
  INV_X1 U17629 ( .A(n15185), .ZN(n14252) );
  AOI22_X1 U17630 ( .A1(n21376), .A2(n15173), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n15643), .ZN(n14172) );
  OAI21_X1 U17631 ( .B1(n14252), .B2(n17250), .A(n14172), .ZN(P1_U2869) );
  INV_X1 U17632 ( .A(n16359), .ZN(n14201) );
  INV_X1 U17633 ( .A(n14173), .ZN(n14174) );
  NAND2_X1 U17634 ( .A1(n9830), .A2(n9807), .ZN(n14498) );
  NOR2_X2 U17635 ( .A1(n14325), .A2(n14498), .ZN(n16355) );
  INV_X1 U17636 ( .A(n14325), .ZN(n14176) );
  NAND2_X1 U17637 ( .A1(n9830), .A2(n14562), .ZN(n14487) );
  INV_X1 U17638 ( .A(n14487), .ZN(n14175) );
  NOR2_X1 U17639 ( .A1(n16326), .A2(n14177), .ZN(n15255) );
  OR2_X1 U17640 ( .A1(n10634), .A2(n14178), .ZN(n14705) );
  INV_X1 U17641 ( .A(n14705), .ZN(n14491) );
  AOI21_X1 U17642 ( .B1(n15255), .B2(n14491), .A(n16359), .ZN(n14183) );
  INV_X1 U17643 ( .A(n14183), .ZN(n14179) );
  NAND2_X1 U17644 ( .A1(n14179), .A2(n16320), .ZN(n14181) );
  INV_X1 U17645 ( .A(n14635), .ZN(n14185) );
  NAND2_X1 U17646 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14185), .ZN(n14180) );
  NAND2_X1 U17647 ( .A1(n14181), .A2(n14180), .ZN(n16361) );
  INV_X1 U17648 ( .A(n16361), .ZN(n14197) );
  OAI22_X1 U17649 ( .A1(n16337), .A2(n15023), .B1(n14197), .B2(n15030), .ZN(
        n14182) );
  AOI21_X1 U17650 ( .B1(n16355), .B2(n15266), .A(n14182), .ZN(n14187) );
  NAND2_X1 U17651 ( .A1(n9830), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16319) );
  OAI211_X1 U17652 ( .C1(n14325), .C2(n16319), .A(n16320), .B(n14183), .ZN(
        n14184) );
  OAI211_X1 U17653 ( .C1(n16320), .C2(n14185), .A(n14184), .B(n14702), .ZN(
        n16358) );
  NAND2_X1 U17654 ( .A1(n16358), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n14186) );
  OAI211_X1 U17655 ( .C1(n15269), .C2(n14201), .A(n14187), .B(n14186), .ZN(
        P1_U3153) );
  OAI22_X1 U17656 ( .A1(n16337), .A2(n15016), .B1(n14197), .B2(n15320), .ZN(
        n14188) );
  AOI21_X1 U17657 ( .B1(n16355), .B2(n15317), .A(n14188), .ZN(n14190) );
  NAND2_X1 U17658 ( .A1(n16358), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14189) );
  OAI211_X1 U17659 ( .C1(n14201), .C2(n15315), .A(n14190), .B(n14189), .ZN(
        P1_U3155) );
  OAI22_X1 U17660 ( .A1(n16337), .A2(n15072), .B1(n14197), .B2(n15309), .ZN(
        n14191) );
  AOI21_X1 U17661 ( .B1(n16355), .B2(n15307), .A(n14191), .ZN(n14193) );
  NAND2_X1 U17662 ( .A1(n16358), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14192) );
  OAI211_X1 U17663 ( .C1(n14201), .C2(n15305), .A(n14193), .B(n14192), .ZN(
        P1_U3156) );
  OAI22_X1 U17664 ( .A1(n16337), .A2(n15058), .B1(n14197), .B2(n15295), .ZN(
        n14194) );
  AOI21_X1 U17665 ( .B1(n16355), .B2(n15293), .A(n14194), .ZN(n14196) );
  NAND2_X1 U17666 ( .A1(n16358), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n14195) );
  OAI211_X1 U17667 ( .C1(n14201), .C2(n15291), .A(n14196), .B(n14195), .ZN(
        P1_U3160) );
  OAI22_X1 U17668 ( .A1(n16337), .A2(n15065), .B1(n14197), .B2(n15302), .ZN(
        n14198) );
  AOI21_X1 U17669 ( .B1(n16355), .B2(n15300), .A(n14198), .ZN(n14200) );
  NAND2_X1 U17670 ( .A1(n16358), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14199) );
  OAI211_X1 U17671 ( .C1(n14201), .C2(n15298), .A(n14200), .B(n14199), .ZN(
        P1_U3158) );
  NAND3_X1 U17672 ( .A1(n17143), .A2(n17138), .A3(n17132), .ZN(n15001) );
  INV_X1 U17673 ( .A(n15001), .ZN(n14207) );
  NAND2_X1 U17674 ( .A1(n14202), .A2(n16322), .ZN(n14499) );
  INV_X1 U17675 ( .A(n16326), .ZN(n21353) );
  OR2_X1 U17676 ( .A1(n15176), .A2(n21353), .ZN(n14998) );
  INV_X1 U17677 ( .A(n14998), .ZN(n14492) );
  NOR2_X1 U17678 ( .A1(n14318), .A2(n15001), .ZN(n14204) );
  AOI21_X1 U17679 ( .B1(n14492), .B2(n14319), .A(n14204), .ZN(n14205) );
  OAI211_X1 U17680 ( .C1(n14499), .C2(n21254), .A(n16320), .B(n14205), .ZN(
        n14203) );
  OAI211_X1 U17681 ( .C1(n16320), .C2(n14207), .A(n14203), .B(n14702), .ZN(
        n14250) );
  INV_X1 U17682 ( .A(n14204), .ZN(n14247) );
  INV_X1 U17683 ( .A(n14205), .ZN(n14206) );
  NAND2_X1 U17684 ( .A1(n14206), .A2(n16320), .ZN(n14209) );
  NAND2_X1 U17685 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14207), .ZN(n14208) );
  AND2_X1 U17686 ( .A1(n14209), .A2(n14208), .ZN(n14246) );
  OAI22_X1 U17687 ( .A1(n15315), .A2(n14247), .B1(n14246), .B2(n15320), .ZN(
        n14211) );
  OAI22_X1 U17688 ( .A1(n15016), .A2(n14772), .B1(n15073), .B2(n15018), .ZN(
        n14210) );
  AOI211_X1 U17689 ( .C1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .C2(n14250), .A(
        n14211), .B(n14210), .ZN(n14212) );
  INV_X1 U17690 ( .A(n14212), .ZN(P1_U3043) );
  OAI22_X1 U17691 ( .A1(n15269), .A2(n14247), .B1(n14246), .B2(n15030), .ZN(
        n14214) );
  OAI22_X1 U17692 ( .A1(n15023), .A2(n14772), .B1(n15073), .B2(n15025), .ZN(
        n14213) );
  AOI211_X1 U17693 ( .C1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .C2(n14250), .A(
        n14214), .B(n14213), .ZN(n14215) );
  INV_X1 U17694 ( .A(n14215), .ZN(P1_U3041) );
  INV_X1 U17695 ( .A(n16341), .ZN(n15288) );
  OAI22_X1 U17696 ( .A1(n15285), .A2(n14247), .B1(n15288), .B2(n14246), .ZN(
        n14217) );
  OAI22_X1 U17697 ( .A1(n15002), .A2(n14772), .B1(n15073), .B2(n15012), .ZN(
        n14216) );
  AOI211_X1 U17698 ( .C1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .C2(n14250), .A(
        n14217), .B(n14216), .ZN(n14218) );
  INV_X1 U17699 ( .A(n14218), .ZN(P1_U3042) );
  NAND3_X1 U17700 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n17138), .ZN(n14897) );
  INV_X1 U17701 ( .A(n14897), .ZN(n14224) );
  INV_X1 U17702 ( .A(n16322), .ZN(n14219) );
  AND2_X1 U17703 ( .A1(n15176), .A2(n16326), .ZN(n14895) );
  NOR2_X1 U17704 ( .A1(n14488), .A2(n17143), .ZN(n14221) );
  AOI21_X1 U17705 ( .B1(n14895), .B2(n14491), .A(n14221), .ZN(n14222) );
  OAI211_X1 U17706 ( .C1(n14282), .C2(n16319), .A(n16320), .B(n14222), .ZN(
        n14220) );
  OAI211_X1 U17707 ( .C1(n16320), .C2(n14224), .A(n14220), .B(n14702), .ZN(
        n14273) );
  INV_X1 U17708 ( .A(n14221), .ZN(n14269) );
  INV_X1 U17709 ( .A(n14222), .ZN(n14223) );
  NAND2_X1 U17710 ( .A1(n14223), .A2(n16320), .ZN(n14226) );
  NAND2_X1 U17711 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14224), .ZN(n14225) );
  AND2_X1 U17712 ( .A1(n14226), .A2(n14225), .ZN(n14268) );
  OAI22_X1 U17713 ( .A1(n15269), .A2(n14269), .B1(n14268), .B2(n15030), .ZN(
        n14229) );
  INV_X1 U17714 ( .A(n15318), .ZN(n14270) );
  INV_X1 U17715 ( .A(n14498), .ZN(n14227) );
  OAI22_X1 U17716 ( .A1(n14270), .A2(n15023), .B1(n15025), .B2(n14925), .ZN(
        n14228) );
  AOI211_X1 U17717 ( .C1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .C2(n14273), .A(
        n14229), .B(n14228), .ZN(n14230) );
  INV_X1 U17718 ( .A(n14230), .ZN(P1_U3121) );
  OAI22_X1 U17719 ( .A1(n15305), .A2(n14247), .B1(n14246), .B2(n15309), .ZN(
        n14232) );
  OAI22_X1 U17720 ( .A1(n15072), .A2(n14772), .B1(n15073), .B2(n15075), .ZN(
        n14231) );
  AOI211_X1 U17721 ( .C1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .C2(n14250), .A(
        n14232), .B(n14231), .ZN(n14233) );
  INV_X1 U17722 ( .A(n14233), .ZN(P1_U3044) );
  INV_X1 U17723 ( .A(n16349), .ZN(n15283) );
  OAI22_X1 U17724 ( .A1(n15280), .A2(n14247), .B1(n15283), .B2(n14246), .ZN(
        n14235) );
  OAI22_X1 U17725 ( .A1(n15046), .A2(n14772), .B1(n15073), .B2(n15048), .ZN(
        n14234) );
  AOI211_X1 U17726 ( .C1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .C2(n14250), .A(
        n14235), .B(n14234), .ZN(n14236) );
  INV_X1 U17727 ( .A(n14236), .ZN(P1_U3045) );
  OAI22_X1 U17728 ( .A1(n15298), .A2(n14247), .B1(n14246), .B2(n15302), .ZN(
        n14238) );
  OAI22_X1 U17729 ( .A1(n15065), .A2(n14772), .B1(n15073), .B2(n15067), .ZN(
        n14237) );
  AOI211_X1 U17730 ( .C1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .C2(n14250), .A(
        n14238), .B(n14237), .ZN(n14239) );
  INV_X1 U17731 ( .A(n14239), .ZN(P1_U3046) );
  OAI22_X1 U17732 ( .A1(n15291), .A2(n14247), .B1(n14246), .B2(n15295), .ZN(
        n14241) );
  OAI22_X1 U17733 ( .A1(n15058), .A2(n14772), .B1(n15073), .B2(n15060), .ZN(
        n14240) );
  AOI211_X1 U17734 ( .C1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .C2(n14250), .A(
        n14241), .B(n14240), .ZN(n14242) );
  INV_X1 U17735 ( .A(n14242), .ZN(P1_U3048) );
  OAI22_X1 U17736 ( .A1(n15315), .A2(n14269), .B1(n14268), .B2(n15320), .ZN(
        n14244) );
  OAI22_X1 U17737 ( .A1(n14270), .A2(n15016), .B1(n15018), .B2(n14925), .ZN(
        n14243) );
  AOI211_X1 U17738 ( .C1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .C2(n14273), .A(
        n14244), .B(n14243), .ZN(n14245) );
  INV_X1 U17739 ( .A(n14245), .ZN(P1_U3123) );
  INV_X1 U17740 ( .A(n16362), .ZN(n15278) );
  OAI22_X1 U17741 ( .A1(n15275), .A2(n14247), .B1(n15278), .B2(n14246), .ZN(
        n14249) );
  OAI22_X1 U17742 ( .A1(n15052), .A2(n14772), .B1(n15073), .B2(n15054), .ZN(
        n14248) );
  AOI211_X1 U17743 ( .C1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .C2(n14250), .A(
        n14249), .B(n14248), .ZN(n14251) );
  INV_X1 U17744 ( .A(n14251), .ZN(P1_U3047) );
  INV_X1 U17745 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n21406) );
  OAI222_X1 U17746 ( .A1(n15739), .A2(n14252), .B1(n15733), .B2(n21406), .C1(
        n15732), .C2(n15706), .ZN(P1_U2901) );
  OAI22_X1 U17747 ( .A1(n15291), .A2(n14269), .B1(n14268), .B2(n15295), .ZN(
        n14254) );
  OAI22_X1 U17748 ( .A1(n14270), .A2(n15058), .B1(n15060), .B2(n14925), .ZN(
        n14253) );
  AOI211_X1 U17749 ( .C1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .C2(n14273), .A(
        n14254), .B(n14253), .ZN(n14255) );
  INV_X1 U17750 ( .A(n14255), .ZN(P1_U3128) );
  OAI22_X1 U17751 ( .A1(n15305), .A2(n14269), .B1(n14268), .B2(n15309), .ZN(
        n14257) );
  OAI22_X1 U17752 ( .A1(n14270), .A2(n15072), .B1(n15075), .B2(n14925), .ZN(
        n14256) );
  AOI211_X1 U17753 ( .C1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .C2(n14273), .A(
        n14257), .B(n14256), .ZN(n14258) );
  INV_X1 U17754 ( .A(n14258), .ZN(P1_U3124) );
  OAI22_X1 U17755 ( .A1(n15298), .A2(n14269), .B1(n14268), .B2(n15302), .ZN(
        n14260) );
  OAI22_X1 U17756 ( .A1(n14270), .A2(n15065), .B1(n15067), .B2(n14925), .ZN(
        n14259) );
  AOI211_X1 U17757 ( .C1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .C2(n14273), .A(
        n14260), .B(n14259), .ZN(n14261) );
  INV_X1 U17758 ( .A(n14261), .ZN(P1_U3126) );
  OAI22_X1 U17759 ( .A1(n15280), .A2(n14269), .B1(n15283), .B2(n14268), .ZN(
        n14263) );
  OAI22_X1 U17760 ( .A1(n14270), .A2(n15046), .B1(n15048), .B2(n14925), .ZN(
        n14262) );
  AOI211_X1 U17761 ( .C1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .C2(n14273), .A(
        n14263), .B(n14262), .ZN(n14264) );
  INV_X1 U17762 ( .A(n14264), .ZN(P1_U3125) );
  OAI22_X1 U17763 ( .A1(n15275), .A2(n14269), .B1(n15278), .B2(n14268), .ZN(
        n14266) );
  OAI22_X1 U17764 ( .A1(n14270), .A2(n15052), .B1(n15054), .B2(n14925), .ZN(
        n14265) );
  AOI211_X1 U17765 ( .C1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .C2(n14273), .A(
        n14266), .B(n14265), .ZN(n14267) );
  INV_X1 U17766 ( .A(n14267), .ZN(P1_U3127) );
  OAI22_X1 U17767 ( .A1(n15285), .A2(n14269), .B1(n15288), .B2(n14268), .ZN(
        n14272) );
  OAI22_X1 U17768 ( .A1(n14270), .A2(n15002), .B1(n15012), .B2(n14925), .ZN(
        n14271) );
  AOI211_X1 U17769 ( .C1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .C2(n14273), .A(
        n14272), .B(n14271), .ZN(n14274) );
  INV_X1 U17770 ( .A(n14274), .ZN(P1_U3122) );
  NAND3_X1 U17771 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17138), .A3(
        n17132), .ZN(n14563) );
  INV_X1 U17772 ( .A(n14563), .ZN(n14279) );
  NOR2_X1 U17773 ( .A1(n14318), .A2(n14563), .ZN(n14276) );
  AOI21_X1 U17774 ( .B1(n14895), .B2(n14319), .A(n14276), .ZN(n14277) );
  OAI211_X1 U17775 ( .C1(n14282), .C2(n21254), .A(n16320), .B(n14277), .ZN(
        n14275) );
  OAI211_X1 U17776 ( .C1(n16320), .C2(n14279), .A(n14275), .B(n14702), .ZN(
        n14316) );
  INV_X1 U17777 ( .A(n14276), .ZN(n14312) );
  INV_X1 U17778 ( .A(n14277), .ZN(n14278) );
  NAND2_X1 U17779 ( .A1(n14278), .A2(n16320), .ZN(n14281) );
  NAND2_X1 U17780 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14279), .ZN(n14280) );
  OAI22_X1 U17781 ( .A1(n15315), .A2(n14312), .B1(n14311), .B2(n15320), .ZN(
        n14285) );
  INV_X1 U17782 ( .A(n14597), .ZN(n14313) );
  INV_X1 U17783 ( .A(n14324), .ZN(n14283) );
  OAI22_X1 U17784 ( .A1(n14313), .A2(n15018), .B1(n15016), .B2(n14926), .ZN(
        n14284) );
  AOI211_X1 U17785 ( .C1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .C2(n14316), .A(
        n14285), .B(n14284), .ZN(n14286) );
  INV_X1 U17786 ( .A(n14286), .ZN(P1_U3107) );
  OAI22_X1 U17787 ( .A1(n15269), .A2(n14312), .B1(n14311), .B2(n15030), .ZN(
        n14288) );
  OAI22_X1 U17788 ( .A1(n14313), .A2(n15025), .B1(n15023), .B2(n14926), .ZN(
        n14287) );
  AOI211_X1 U17789 ( .C1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .C2(n14316), .A(
        n14288), .B(n14287), .ZN(n14289) );
  INV_X1 U17790 ( .A(n14289), .ZN(P1_U3105) );
  XNOR2_X1 U17791 ( .A(n9925), .B(n20421), .ZN(n14295) );
  OR2_X1 U17792 ( .A1(n14291), .A2(n14290), .ZN(n14292) );
  AND2_X1 U17793 ( .A1(n14292), .A2(n17532), .ZN(n20294) );
  NOR2_X1 U17794 ( .A1(n13216), .A2(n20286), .ZN(n14293) );
  AOI21_X1 U17795 ( .B1(n20294), .B2(n13216), .A(n14293), .ZN(n14294) );
  OAI21_X1 U17796 ( .B1(n14295), .B2(n20428), .A(n14294), .ZN(P2_U2876) );
  OAI22_X1 U17797 ( .A1(n15280), .A2(n14312), .B1(n15283), .B2(n14311), .ZN(
        n14297) );
  OAI22_X1 U17798 ( .A1(n14313), .A2(n15048), .B1(n15046), .B2(n14926), .ZN(
        n14296) );
  AOI211_X1 U17799 ( .C1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .C2(n14316), .A(
        n14297), .B(n14296), .ZN(n14298) );
  INV_X1 U17800 ( .A(n14298), .ZN(P1_U3109) );
  OAI22_X1 U17801 ( .A1(n15285), .A2(n14312), .B1(n15288), .B2(n14311), .ZN(
        n14300) );
  OAI22_X1 U17802 ( .A1(n14313), .A2(n15012), .B1(n15002), .B2(n14926), .ZN(
        n14299) );
  AOI211_X1 U17803 ( .C1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .C2(n14316), .A(
        n14300), .B(n14299), .ZN(n14301) );
  INV_X1 U17804 ( .A(n14301), .ZN(P1_U3106) );
  OAI22_X1 U17805 ( .A1(n15275), .A2(n14312), .B1(n15278), .B2(n14311), .ZN(
        n14303) );
  OAI22_X1 U17806 ( .A1(n14313), .A2(n15054), .B1(n15052), .B2(n14926), .ZN(
        n14302) );
  AOI211_X1 U17807 ( .C1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .C2(n14316), .A(
        n14303), .B(n14302), .ZN(n14304) );
  INV_X1 U17808 ( .A(n14304), .ZN(P1_U3111) );
  OAI22_X1 U17809 ( .A1(n15291), .A2(n14312), .B1(n14311), .B2(n15295), .ZN(
        n14306) );
  OAI22_X1 U17810 ( .A1(n14313), .A2(n15060), .B1(n15058), .B2(n14926), .ZN(
        n14305) );
  AOI211_X1 U17811 ( .C1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .C2(n14316), .A(
        n14306), .B(n14305), .ZN(n14307) );
  INV_X1 U17812 ( .A(n14307), .ZN(P1_U3112) );
  OAI22_X1 U17813 ( .A1(n15298), .A2(n14312), .B1(n14311), .B2(n15302), .ZN(
        n14309) );
  OAI22_X1 U17814 ( .A1(n14313), .A2(n15067), .B1(n15065), .B2(n14926), .ZN(
        n14308) );
  AOI211_X1 U17815 ( .C1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .C2(n14316), .A(
        n14309), .B(n14308), .ZN(n14310) );
  INV_X1 U17816 ( .A(n14310), .ZN(P1_U3110) );
  OAI22_X1 U17817 ( .A1(n15305), .A2(n14312), .B1(n14311), .B2(n15309), .ZN(
        n14315) );
  OAI22_X1 U17818 ( .A1(n14313), .A2(n15075), .B1(n15072), .B2(n14926), .ZN(
        n14314) );
  AOI211_X1 U17819 ( .C1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .C2(n14316), .A(
        n14315), .B(n14314), .ZN(n14317) );
  INV_X1 U17820 ( .A(n14317), .ZN(P1_U3108) );
  NAND3_X1 U17821 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n17132), .ZN(n15257) );
  INV_X1 U17822 ( .A(n15257), .ZN(n14328) );
  NOR3_X1 U17823 ( .A1(n14325), .A2(n21254), .A3(n9830), .ZN(n16330) );
  INV_X1 U17824 ( .A(n16330), .ZN(n14320) );
  NOR2_X1 U17825 ( .A1(n14318), .A2(n15257), .ZN(n14410) );
  AOI21_X1 U17826 ( .B1(n15255), .B2(n14319), .A(n14410), .ZN(n14326) );
  NAND3_X1 U17827 ( .A1(n14320), .A2(n16320), .A3(n14326), .ZN(n14321) );
  OAI211_X1 U17828 ( .C1(n16320), .C2(n14328), .A(n14321), .B(n14702), .ZN(
        n14322) );
  INV_X1 U17829 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14334) );
  NOR2_X2 U17830 ( .A1(n14325), .A2(n14323), .ZN(n15312) );
  INV_X1 U17831 ( .A(n15312), .ZN(n14348) );
  NOR2_X2 U17832 ( .A1(n14325), .A2(n14324), .ZN(n14693) );
  INV_X1 U17833 ( .A(n14326), .ZN(n14327) );
  NAND2_X1 U17834 ( .A1(n14327), .A2(n16320), .ZN(n14330) );
  NAND2_X1 U17835 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14328), .ZN(n14329) );
  NAND2_X1 U17836 ( .A1(n14330), .A2(n14329), .ZN(n14409) );
  AOI22_X1 U17837 ( .A1(n14693), .A2(n15289), .B1(n14823), .B2(n14409), .ZN(
        n14331) );
  OAI21_X1 U17838 ( .B1(n15060), .B2(n14348), .A(n14331), .ZN(n14332) );
  AOI21_X1 U17839 ( .B1(n15063), .B2(n14410), .A(n14332), .ZN(n14333) );
  OAI21_X1 U17840 ( .B1(n14414), .B2(n14334), .A(n14333), .ZN(P1_U3144) );
  INV_X1 U17841 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U17842 ( .A1(n14693), .A2(n15311), .B1(n14818), .B2(n14409), .ZN(
        n14335) );
  OAI21_X1 U17843 ( .B1(n15018), .B2(n14348), .A(n14335), .ZN(n14336) );
  AOI21_X1 U17844 ( .B1(n15021), .B2(n14410), .A(n14336), .ZN(n14337) );
  OAI21_X1 U17845 ( .B1(n14414), .B2(n14338), .A(n14337), .ZN(P1_U3139) );
  INV_X1 U17846 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14342) );
  AOI22_X1 U17847 ( .A1(n14693), .A2(n15265), .B1(n15271), .B2(n14409), .ZN(
        n14339) );
  OAI21_X1 U17848 ( .B1(n15025), .B2(n14348), .A(n14339), .ZN(n14340) );
  AOI21_X1 U17849 ( .B1(n15028), .B2(n14410), .A(n14340), .ZN(n14341) );
  OAI21_X1 U17850 ( .B1(n14414), .B2(n14342), .A(n14341), .ZN(P1_U3137) );
  INV_X1 U17851 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14346) );
  AOI22_X1 U17852 ( .A1(n14693), .A2(n15303), .B1(n14810), .B2(n14409), .ZN(
        n14343) );
  OAI21_X1 U17853 ( .B1(n15075), .B2(n14348), .A(n14343), .ZN(n14344) );
  AOI21_X1 U17854 ( .B1(n15078), .B2(n14410), .A(n14344), .ZN(n14345) );
  OAI21_X1 U17855 ( .B1(n14414), .B2(n14346), .A(n14345), .ZN(P1_U3140) );
  AOI22_X1 U17856 ( .A1(n14693), .A2(n15296), .B1(n14814), .B2(n14409), .ZN(
        n14347) );
  OAI21_X1 U17857 ( .B1(n15067), .B2(n14348), .A(n14347), .ZN(n14349) );
  AOI21_X1 U17858 ( .B1(n15070), .B2(n14410), .A(n14349), .ZN(n14350) );
  OAI21_X1 U17859 ( .B1(n14414), .B2(n15940), .A(n14350), .ZN(P1_U3142) );
  INV_X1 U17860 ( .A(n14351), .ZN(n14352) );
  NAND2_X1 U17861 ( .A1(n14353), .A2(n14352), .ZN(n14354) );
  OAI21_X1 U17862 ( .B1(n14355), .B2(n14354), .A(n13945), .ZN(n20383) );
  AOI21_X1 U17863 ( .B1(n14882), .B2(n21190), .A(n14356), .ZN(n20487) );
  OR2_X1 U17864 ( .A1(n14358), .A2(n14357), .ZN(n14359) );
  NAND2_X1 U17865 ( .A1(n14359), .A2(n14360), .ZN(n21185) );
  XNOR2_X1 U17866 ( .A(n20800), .B(n21185), .ZN(n20486) );
  NOR2_X1 U17867 ( .A1(n20487), .A2(n20486), .ZN(n20485) );
  INV_X1 U17868 ( .A(n21185), .ZN(n20484) );
  NOR2_X1 U17869 ( .A1(n21181), .A2(n20484), .ZN(n14362) );
  XNOR2_X1 U17870 ( .A(n14361), .B(n14360), .ZN(n14943) );
  OAI21_X1 U17871 ( .B1(n20485), .B2(n14362), .A(n14943), .ZN(n20479) );
  XOR2_X1 U17872 ( .A(n20383), .B(n20479), .Z(n14365) );
  INV_X1 U17873 ( .A(n14943), .ZN(n20377) );
  AOI22_X1 U17874 ( .A1(n20492), .A2(n20377), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n20491), .ZN(n14364) );
  NAND2_X1 U17875 ( .A1(n20468), .A2(n17491), .ZN(n14363) );
  OAI211_X1 U17876 ( .C1(n14365), .C2(n20496), .A(n14364), .B(n14363), .ZN(
        P2_U2915) );
  XNOR2_X1 U17877 ( .A(n14366), .B(n14367), .ZN(n14634) );
  AOI21_X1 U17878 ( .B1(n14369), .B2(n14368), .A(n14618), .ZN(n14370) );
  AOI22_X1 U17879 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14371), .B1(
        n14620), .B2(n14370), .ZN(n14377) );
  AND2_X1 U17880 ( .A1(n14373), .A2(n14372), .ZN(n14374) );
  NOR2_X1 U17881 ( .A1(n14977), .A2(n14374), .ZN(n21370) );
  INV_X1 U17882 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n14375) );
  NOR2_X1 U17883 ( .A1(n17352), .A2(n14375), .ZN(n14631) );
  AOI21_X1 U17884 ( .B1(n21427), .B2(n21370), .A(n14631), .ZN(n14376) );
  OAI211_X1 U17885 ( .C1(n17365), .C2(n14634), .A(n14377), .B(n14376), .ZN(
        P1_U3027) );
  INV_X1 U17886 ( .A(n20594), .ZN(n14378) );
  OAI21_X1 U17887 ( .B1(n20715), .B2(n20764), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14383) );
  NAND2_X1 U17888 ( .A1(n20667), .A2(n14379), .ZN(n14386) );
  NOR2_X1 U17889 ( .A1(n20833), .A2(n20699), .ZN(n20742) );
  INV_X1 U17890 ( .A(n20742), .ZN(n14380) );
  AND2_X1 U17891 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n14380), .ZN(n14381) );
  NAND2_X1 U17892 ( .A1(n11704), .A2(n14381), .ZN(n14384) );
  OAI211_X1 U17893 ( .C1(n20975), .C2(n20742), .A(n14384), .B(n21023), .ZN(
        n14382) );
  AOI21_X1 U17894 ( .B1(n14383), .B2(n14386), .A(n14382), .ZN(n20729) );
  INV_X1 U17895 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14390) );
  INV_X1 U17896 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17819) );
  INV_X1 U17897 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19548) );
  OAI22_X2 U17898 ( .A1(n17819), .A2(n20579), .B1(n19548), .B2(n20577), .ZN(
        n21030) );
  AOI22_X1 U17899 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20572), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20571), .ZN(n21033) );
  INV_X1 U17900 ( .A(n21033), .ZN(n20944) );
  AOI22_X1 U17901 ( .A1(n20764), .A2(n21030), .B1(n20715), .B2(n20944), .ZN(
        n14389) );
  INV_X1 U17902 ( .A(n14384), .ZN(n14385) );
  AOI211_X2 U17903 ( .C1(n21225), .C2(n14386), .A(n20588), .B(n14385), .ZN(
        n20743) );
  NOR2_X2 U17904 ( .A1(n14387), .A2(n20977), .ZN(n21021) );
  NOR2_X2 U17905 ( .A1(n20574), .A2(n11463), .ZN(n21020) );
  AOI22_X1 U17906 ( .A1(n20743), .A2(n21021), .B1(n21020), .B2(n20742), .ZN(
        n14388) );
  OAI211_X1 U17907 ( .C1(n20729), .C2(n14390), .A(n14389), .B(n14388), .ZN(
        P2_U3096) );
  INV_X1 U17908 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U17909 ( .A1(n21410), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14391) );
  OAI21_X1 U17910 ( .B1(n14451), .B2(n14402), .A(n14391), .ZN(P1_U2912) );
  INV_X1 U17911 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U17912 ( .A1(n21410), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14392) );
  OAI21_X1 U17913 ( .B1(n14427), .B2(n14402), .A(n14392), .ZN(P1_U2906) );
  INV_X1 U17914 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14482) );
  AOI22_X1 U17915 ( .A1(n21410), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14393) );
  OAI21_X1 U17916 ( .B1(n14482), .B2(n14402), .A(n14393), .ZN(P1_U2916) );
  INV_X1 U17917 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U17918 ( .A1(n21410), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14394) );
  OAI21_X1 U17919 ( .B1(n14438), .B2(n14402), .A(n14394), .ZN(P1_U2907) );
  AOI22_X1 U17920 ( .A1(n21410), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14395) );
  OAI21_X1 U17921 ( .B1(n15693), .B2(n14402), .A(n14395), .ZN(P1_U2915) );
  INV_X1 U17922 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14474) );
  AOI22_X1 U17923 ( .A1(n21410), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14396) );
  OAI21_X1 U17924 ( .B1(n14474), .B2(n14402), .A(n14396), .ZN(P1_U2918) );
  INV_X1 U17925 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U17926 ( .A1(n21410), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14397) );
  OAI21_X1 U17927 ( .B1(n14431), .B2(n14402), .A(n14397), .ZN(P1_U2909) );
  INV_X1 U17928 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U17929 ( .A1(n21410), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14398) );
  OAI21_X1 U17930 ( .B1(n14479), .B2(n14402), .A(n14398), .ZN(P1_U2920) );
  AOI22_X1 U17931 ( .A1(n21410), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14399) );
  OAI21_X1 U17932 ( .B1(n15705), .B2(n14402), .A(n14399), .ZN(P1_U2917) );
  INV_X1 U17933 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14464) );
  AOI22_X1 U17934 ( .A1(n21410), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14400) );
  OAI21_X1 U17935 ( .B1(n14464), .B2(n14402), .A(n14400), .ZN(P1_U2914) );
  AOI22_X1 U17936 ( .A1(n21410), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14401) );
  OAI21_X1 U17937 ( .B1(n10895), .B2(n14402), .A(n14401), .ZN(P1_U2919) );
  INV_X1 U17938 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14405) );
  AOI22_X1 U17939 ( .A1(n15312), .A2(n16346), .B1(n14693), .B2(n16347), .ZN(
        n14404) );
  AOI22_X1 U17940 ( .A1(n16348), .A2(n14410), .B1(n16349), .B2(n14409), .ZN(
        n14403) );
  OAI211_X1 U17941 ( .C1(n14414), .C2(n14405), .A(n14404), .B(n14403), .ZN(
        P1_U3141) );
  INV_X1 U17942 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U17943 ( .A1(n15312), .A2(n16338), .B1(n14693), .B2(n16339), .ZN(
        n14407) );
  AOI22_X1 U17944 ( .A1(n16340), .A2(n14410), .B1(n16341), .B2(n14409), .ZN(
        n14406) );
  OAI211_X1 U17945 ( .C1(n14414), .C2(n14408), .A(n14407), .B(n14406), .ZN(
        P1_U3138) );
  INV_X1 U17946 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U17947 ( .A1(n15312), .A2(n16354), .B1(n14693), .B2(n16356), .ZN(
        n14412) );
  AOI22_X1 U17948 ( .A1(n16360), .A2(n14410), .B1(n16362), .B2(n14409), .ZN(
        n14411) );
  OAI211_X1 U17949 ( .C1(n14414), .C2(n14413), .A(n14412), .B(n14411), .ZN(
        P1_U3143) );
  AND2_X1 U17950 ( .A1(n14415), .A2(n14416), .ZN(n14418) );
  OR2_X1 U17951 ( .A1(n14418), .A2(n14417), .ZN(n14623) );
  XOR2_X1 U17952 ( .A(n14976), .B(n14977), .Z(n21318) );
  AOI22_X1 U17953 ( .A1(n21376), .A2(n21318), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n15643), .ZN(n14419) );
  OAI21_X1 U17954 ( .B1(n14623), .B2(n17250), .A(n14419), .ZN(P1_U2867) );
  INV_X1 U17955 ( .A(DATAI_12_), .ZN(n14421) );
  NAND2_X1 U17956 ( .A1(n15371), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14420) );
  OAI21_X1 U17957 ( .B1(n15371), .B2(n14421), .A(n14420), .ZN(n21416) );
  AOI22_X1 U17958 ( .A1(n21422), .A2(n21416), .B1(P1_UWORD_REG_12__SCAN_IN), 
        .B2(n14483), .ZN(n14422) );
  OAI21_X1 U17959 ( .B1(n14555), .B2(n14423), .A(n14422), .ZN(P1_U2949) );
  INV_X1 U17960 ( .A(DATAI_14_), .ZN(n14425) );
  NAND2_X1 U17961 ( .A1(n15371), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14424) );
  OAI21_X1 U17962 ( .B1(n15371), .B2(n14425), .A(n14424), .ZN(n21421) );
  AOI22_X1 U17963 ( .A1(n21422), .A2(n21421), .B1(P1_UWORD_REG_14__SCAN_IN), 
        .B2(n14483), .ZN(n14426) );
  OAI21_X1 U17964 ( .B1(n14555), .B2(n14427), .A(n14426), .ZN(P1_U2951) );
  INV_X1 U17965 ( .A(n21422), .ZN(n14554) );
  INV_X1 U17966 ( .A(DATAI_11_), .ZN(n14429) );
  NAND2_X1 U17967 ( .A1(n15371), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14428) );
  OAI21_X1 U17968 ( .B1(n15371), .B2(n14429), .A(n14428), .ZN(n15660) );
  INV_X1 U17969 ( .A(n15660), .ZN(n15333) );
  NOR2_X1 U17970 ( .A1(n14554), .A2(n15333), .ZN(n14452) );
  AOI21_X1 U17971 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n21419), .A(n14452), 
        .ZN(n14430) );
  OAI21_X1 U17972 ( .B1(n14431), .B2(n14555), .A(n14430), .ZN(P1_U2948) );
  INV_X1 U17973 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n21398) );
  INV_X1 U17974 ( .A(DATAI_8_), .ZN(n14433) );
  NAND2_X1 U17975 ( .A1(n15371), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14432) );
  OAI21_X1 U17976 ( .B1(n15371), .B2(n14433), .A(n14432), .ZN(n15676) );
  INV_X1 U17977 ( .A(n15676), .ZN(n15092) );
  NOR2_X1 U17978 ( .A1(n14554), .A2(n15092), .ZN(n14449) );
  AOI21_X1 U17979 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n21419), .A(n14449), 
        .ZN(n14434) );
  OAI21_X1 U17980 ( .B1(n21398), .B2(n14555), .A(n14434), .ZN(P1_U2960) );
  INV_X1 U17981 ( .A(DATAI_13_), .ZN(n14436) );
  NAND2_X1 U17982 ( .A1(n15371), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14435) );
  OAI21_X1 U17983 ( .B1(n15371), .B2(n14436), .A(n14435), .ZN(n15650) );
  INV_X1 U17984 ( .A(n15650), .ZN(n15731) );
  NOR2_X1 U17985 ( .A1(n14554), .A2(n15731), .ZN(n14442) );
  AOI21_X1 U17986 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n21419), .A(n14442), 
        .ZN(n14437) );
  OAI21_X1 U17987 ( .B1(n14438), .B2(n14555), .A(n14437), .ZN(P1_U2950) );
  NOR2_X1 U17988 ( .A1(n14554), .A2(n15694), .ZN(n14454) );
  AOI21_X1 U17989 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n21419), .A(n14454), 
        .ZN(n14439) );
  OAI21_X1 U17990 ( .B1(n10705), .B2(n14555), .A(n14439), .ZN(P1_U2957) );
  NOR2_X1 U17991 ( .A1(n14554), .A2(n15681), .ZN(n14446) );
  AOI21_X1 U17992 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n21419), .A(n14446), 
        .ZN(n14440) );
  OAI21_X1 U17993 ( .B1(n10733), .B2(n14555), .A(n14440), .ZN(P1_U2959) );
  NOR2_X1 U17994 ( .A1(n14554), .A2(n15706), .ZN(n14444) );
  AOI21_X1 U17995 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n21419), .A(n14444), 
        .ZN(n14441) );
  OAI21_X1 U17996 ( .B1(n21406), .B2(n14555), .A(n14441), .ZN(P1_U2955) );
  INV_X1 U17997 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n21387) );
  AOI21_X1 U17998 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n21419), .A(n14442), 
        .ZN(n14443) );
  OAI21_X1 U17999 ( .B1(n21387), .B2(n14555), .A(n14443), .ZN(P1_U2965) );
  AOI21_X1 U18000 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n14483), .A(n14444), 
        .ZN(n14445) );
  OAI21_X1 U18001 ( .B1(n15705), .B2(n14555), .A(n14445), .ZN(P1_U2940) );
  AOI21_X1 U18002 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n14483), .A(n14446), 
        .ZN(n14447) );
  OAI21_X1 U18003 ( .B1(n14448), .B2(n14555), .A(n14447), .ZN(P1_U2944) );
  AOI21_X1 U18004 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n14483), .A(n14449), 
        .ZN(n14450) );
  OAI21_X1 U18005 ( .B1(n14451), .B2(n14555), .A(n14450), .ZN(P1_U2945) );
  INV_X1 U18006 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n21391) );
  AOI21_X1 U18007 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n21419), .A(n14452), 
        .ZN(n14453) );
  OAI21_X1 U18008 ( .B1(n21391), .B2(n14555), .A(n14453), .ZN(P1_U2963) );
  AOI21_X1 U18009 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n14483), .A(n14454), 
        .ZN(n14455) );
  OAI21_X1 U18010 ( .B1(n15693), .B2(n14555), .A(n14455), .ZN(P1_U2942) );
  INV_X1 U18011 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n21401) );
  NAND2_X1 U18012 ( .A1(n21422), .A2(n15686), .ZN(n14462) );
  NAND2_X1 U18013 ( .A1(n14483), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n14456) );
  OAI211_X1 U18014 ( .C1(n14555), .C2(n21401), .A(n14462), .B(n14456), .ZN(
        P1_U2958) );
  NAND2_X1 U18015 ( .A1(n14483), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n14458) );
  INV_X1 U18016 ( .A(n14457), .ZN(n15712) );
  NAND2_X1 U18017 ( .A1(n21422), .A2(n15712), .ZN(n14472) );
  OAI211_X1 U18018 ( .C1(n14555), .C2(n21409), .A(n14458), .B(n14472), .ZN(
        P1_U2954) );
  INV_X1 U18019 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21404) );
  NAND2_X1 U18020 ( .A1(n21422), .A2(n15698), .ZN(n14480) );
  NAND2_X1 U18021 ( .A1(n14483), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n14459) );
  OAI211_X1 U18022 ( .C1(n14555), .C2(n21404), .A(n14480), .B(n14459), .ZN(
        P1_U2956) );
  NAND2_X1 U18023 ( .A1(n14483), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n14461) );
  INV_X1 U18024 ( .A(n14460), .ZN(n15718) );
  NAND2_X1 U18025 ( .A1(n21422), .A2(n15718), .ZN(n14477) );
  OAI211_X1 U18026 ( .C1(n14555), .C2(n21415), .A(n14461), .B(n14477), .ZN(
        P1_U2952) );
  NAND2_X1 U18027 ( .A1(n14483), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14463) );
  OAI211_X1 U18028 ( .C1(n14555), .C2(n14464), .A(n14463), .B(n14462), .ZN(
        P1_U2943) );
  INV_X1 U18029 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n21396) );
  INV_X1 U18030 ( .A(DATAI_9_), .ZN(n14466) );
  NAND2_X1 U18031 ( .A1(n15371), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14465) );
  OAI21_X1 U18032 ( .B1(n15371), .B2(n14466), .A(n14465), .ZN(n15671) );
  NAND2_X1 U18033 ( .A1(n21422), .A2(n15671), .ZN(n14468) );
  NAND2_X1 U18034 ( .A1(n21419), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n14467) );
  OAI211_X1 U18035 ( .C1(n14555), .C2(n21396), .A(n14468), .B(n14467), .ZN(
        P1_U2961) );
  NAND2_X1 U18036 ( .A1(n14483), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14469) );
  OAI211_X1 U18037 ( .C1(n14555), .C2(n14470), .A(n14469), .B(n14468), .ZN(
        P1_U2946) );
  INV_X1 U18038 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21412) );
  NAND2_X1 U18039 ( .A1(n21422), .A2(n15376), .ZN(n14475) );
  NAND2_X1 U18040 ( .A1(n14483), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n14471) );
  OAI211_X1 U18041 ( .C1(n14555), .C2(n21412), .A(n14475), .B(n14471), .ZN(
        P1_U2953) );
  NAND2_X1 U18042 ( .A1(n21419), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14473) );
  OAI211_X1 U18043 ( .C1(n14555), .C2(n14474), .A(n14473), .B(n14472), .ZN(
        P1_U2939) );
  NAND2_X1 U18044 ( .A1(n21419), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14476) );
  OAI211_X1 U18045 ( .C1(n14555), .C2(n10895), .A(n14476), .B(n14475), .ZN(
        P1_U2938) );
  NAND2_X1 U18046 ( .A1(n21419), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14478) );
  OAI211_X1 U18047 ( .C1(n14555), .C2(n14479), .A(n14478), .B(n14477), .ZN(
        P1_U2937) );
  NAND2_X1 U18048 ( .A1(n21419), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14481) );
  OAI211_X1 U18049 ( .C1(n14555), .C2(n14482), .A(n14481), .B(n14480), .ZN(
        P1_U2941) );
  NAND2_X1 U18050 ( .A1(n14483), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14485) );
  OAI211_X1 U18051 ( .C1(n14555), .C2(n14486), .A(n14485), .B(n14484), .ZN(
        P1_U2947) );
  OAI222_X1 U18052 ( .A1(n15739), .A2(n14623), .B1(n15733), .B2(n10705), .C1(
        n15732), .C2(n15694), .ZN(P1_U2899) );
  INV_X1 U18053 ( .A(n14488), .ZN(n14489) );
  NAND2_X1 U18054 ( .A1(n14489), .A2(n17143), .ZN(n14542) );
  INV_X1 U18055 ( .A(n14542), .ZN(n14490) );
  AOI21_X1 U18056 ( .B1(n14492), .B2(n14491), .A(n14490), .ZN(n14497) );
  NAND2_X1 U18057 ( .A1(n16319), .A2(n16320), .ZN(n16324) );
  NAND2_X1 U18058 ( .A1(n14499), .A2(n16320), .ZN(n14493) );
  NAND2_X1 U18059 ( .A1(n16324), .A2(n14493), .ZN(n14495) );
  NAND3_X1 U18060 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17143), .A3(
        n17138), .ZN(n14743) );
  AOI22_X1 U18061 ( .A1(n14497), .A2(n14495), .B1(n16334), .B2(n14743), .ZN(
        n14494) );
  NAND2_X1 U18062 ( .A1(n14702), .A2(n14494), .ZN(n14541) );
  INV_X1 U18063 ( .A(n14495), .ZN(n14496) );
  OAI22_X1 U18064 ( .A1(n14497), .A2(n14496), .B1(n21441), .B2(n14743), .ZN(
        n14540) );
  AOI22_X1 U18065 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14541), .B1(
        n16349), .B2(n14540), .ZN(n14502) );
  OAI22_X1 U18066 ( .A1(n14748), .A2(n15048), .B1(n15280), .B2(n14542), .ZN(
        n14500) );
  INV_X1 U18067 ( .A(n14500), .ZN(n14501) );
  OAI211_X1 U18068 ( .C1(n15046), .C2(n14789), .A(n14502), .B(n14501), .ZN(
        P1_U3061) );
  AOI22_X1 U18069 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14541), .B1(
        n16362), .B2(n14540), .ZN(n14505) );
  OAI22_X1 U18070 ( .A1(n14748), .A2(n15054), .B1(n15275), .B2(n14542), .ZN(
        n14503) );
  INV_X1 U18071 ( .A(n14503), .ZN(n14504) );
  OAI211_X1 U18072 ( .C1(n15052), .C2(n14789), .A(n14505), .B(n14504), .ZN(
        P1_U3063) );
  AOI22_X1 U18073 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14541), .B1(
        n16341), .B2(n14540), .ZN(n14508) );
  OAI22_X1 U18074 ( .A1(n14748), .A2(n15012), .B1(n15285), .B2(n14542), .ZN(
        n14506) );
  INV_X1 U18075 ( .A(n14506), .ZN(n14507) );
  OAI211_X1 U18076 ( .C1(n15002), .C2(n14789), .A(n14508), .B(n14507), .ZN(
        P1_U3058) );
  XNOR2_X1 U18077 ( .A(n14509), .B(n14602), .ZN(n14513) );
  INV_X1 U18078 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n15856) );
  OAI21_X1 U18079 ( .B1(n14510), .B2(n14511), .A(n14607), .ZN(n16870) );
  MUX2_X1 U18080 ( .A(n15856), .B(n16870), .S(n20437), .Z(n14512) );
  OAI21_X1 U18081 ( .B1(n14513), .B2(n20428), .A(n14512), .ZN(P2_U2874) );
  OAI21_X1 U18082 ( .B1(n14417), .B2(n14516), .A(n14515), .ZN(n21310) );
  AOI22_X1 U18083 ( .A1(n15737), .A2(n15686), .B1(P1_EAX_REG_6__SCAN_IN), .B2(
        n15736), .ZN(n14517) );
  OAI21_X1 U18084 ( .B1(n21310), .B2(n15739), .A(n14517), .ZN(P1_U2898) );
  INV_X1 U18085 ( .A(n17306), .ZN(n17298) );
  AOI21_X1 U18086 ( .B1(n14161), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14518), .ZN(n14519) );
  OAI21_X1 U18087 ( .B1(n17305), .B2(n21347), .A(n14519), .ZN(n14520) );
  AOI21_X1 U18088 ( .B1(n21358), .B2(n17298), .A(n14520), .ZN(n14521) );
  OAI21_X1 U18089 ( .B1(n17312), .B2(n14522), .A(n14521), .ZN(P1_U2997) );
  AOI21_X1 U18090 ( .B1(n14161), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n14523), .ZN(n14524) );
  OAI21_X1 U18091 ( .B1(n17305), .B2(n15174), .A(n14524), .ZN(n14525) );
  AOI21_X1 U18092 ( .B1(n15185), .B2(n17298), .A(n14525), .ZN(n14526) );
  OAI21_X1 U18093 ( .B1(n17312), .B2(n14527), .A(n14526), .ZN(P1_U2996) );
  AOI22_X1 U18094 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14541), .B1(
        n14814), .B2(n14540), .ZN(n14530) );
  OAI22_X1 U18095 ( .A1(n14748), .A2(n15067), .B1(n15298), .B2(n14542), .ZN(
        n14528) );
  INV_X1 U18096 ( .A(n14528), .ZN(n14529) );
  OAI211_X1 U18097 ( .C1(n15065), .C2(n14789), .A(n14530), .B(n14529), .ZN(
        P1_U3062) );
  AOI22_X1 U18098 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14541), .B1(
        n14810), .B2(n14540), .ZN(n14533) );
  OAI22_X1 U18099 ( .A1(n14748), .A2(n15075), .B1(n15305), .B2(n14542), .ZN(
        n14531) );
  INV_X1 U18100 ( .A(n14531), .ZN(n14532) );
  OAI211_X1 U18101 ( .C1(n15072), .C2(n14789), .A(n14533), .B(n14532), .ZN(
        P1_U3060) );
  AOI22_X1 U18102 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14541), .B1(
        n14818), .B2(n14540), .ZN(n14536) );
  OAI22_X1 U18103 ( .A1(n14748), .A2(n15018), .B1(n15315), .B2(n14542), .ZN(
        n14534) );
  INV_X1 U18104 ( .A(n14534), .ZN(n14535) );
  OAI211_X1 U18105 ( .C1(n15016), .C2(n14789), .A(n14536), .B(n14535), .ZN(
        P1_U3059) );
  AOI22_X1 U18106 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14541), .B1(
        n14823), .B2(n14540), .ZN(n14539) );
  OAI22_X1 U18107 ( .A1(n14748), .A2(n15060), .B1(n15291), .B2(n14542), .ZN(
        n14537) );
  INV_X1 U18108 ( .A(n14537), .ZN(n14538) );
  OAI211_X1 U18109 ( .C1(n15058), .C2(n14789), .A(n14539), .B(n14538), .ZN(
        P1_U3064) );
  AOI22_X1 U18110 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n14541), .B1(
        n15271), .B2(n14540), .ZN(n14545) );
  OAI22_X1 U18111 ( .A1(n14748), .A2(n15025), .B1(n15269), .B2(n14542), .ZN(
        n14543) );
  INV_X1 U18112 ( .A(n14543), .ZN(n14544) );
  OAI211_X1 U18113 ( .C1(n15023), .C2(n14789), .A(n14545), .B(n14544), .ZN(
        P1_U3057) );
  INV_X1 U18114 ( .A(n14415), .ZN(n14546) );
  AOI21_X1 U18115 ( .B1(n14547), .B2(n14169), .A(n14546), .ZN(n21371) );
  INV_X1 U18116 ( .A(n21371), .ZN(n14549) );
  AOI22_X1 U18117 ( .A1(n15737), .A2(n15698), .B1(P1_EAX_REG_4__SCAN_IN), .B2(
        n15736), .ZN(n14548) );
  OAI21_X1 U18118 ( .B1(n14549), .B2(n15739), .A(n14548), .ZN(P1_U2900) );
  INV_X1 U18119 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n15727) );
  INV_X1 U18120 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14550) );
  NOR2_X1 U18121 ( .A1(n14552), .A2(n14550), .ZN(n14551) );
  AOI21_X1 U18122 ( .B1(DATAI_15_), .B2(n14552), .A(n14551), .ZN(n15726) );
  INV_X1 U18123 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n21383) );
  OAI222_X1 U18124 ( .A1(n14555), .A2(n15727), .B1(n14554), .B2(n15726), .C1(
        n14553), .C2(n21383), .ZN(P1_U2967) );
  NAND2_X1 U18125 ( .A1(n14556), .A2(n17267), .ZN(n14559) );
  INV_X1 U18126 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15110) );
  OAI22_X1 U18127 ( .A1(n15759), .A2(n15110), .B1(n17352), .B2(n21534), .ZN(
        n14557) );
  AOI21_X1 U18128 ( .B1(n17296), .B2(n15110), .A(n14557), .ZN(n14558) );
  OAI211_X1 U18129 ( .C1(n15120), .C2(n17306), .A(n14559), .B(n14558), .ZN(
        P1_U2998) );
  INV_X1 U18130 ( .A(n14560), .ZN(n14703) );
  OAI21_X1 U18131 ( .B1(n14735), .B2(n14597), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14566) );
  NOR2_X1 U18132 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14563), .ZN(
        n14596) );
  AOI21_X1 U18133 ( .B1(n14895), .B2(n13865), .A(n14596), .ZN(n14567) );
  AND2_X1 U18134 ( .A1(n14569), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14833) );
  OAI21_X1 U18135 ( .B1(n17400), .B2(n14596), .A(n15008), .ZN(n14565) );
  INV_X1 U18136 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14576) );
  INV_X1 U18137 ( .A(n14567), .ZN(n14568) );
  NAND2_X1 U18138 ( .A1(n14568), .A2(n16320), .ZN(n14573) );
  INV_X1 U18139 ( .A(n14569), .ZN(n14570) );
  NAND2_X1 U18140 ( .A1(n14570), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14741) );
  INV_X1 U18141 ( .A(n14796), .ZN(n14571) );
  NAND2_X1 U18142 ( .A1(n14571), .A2(n14795), .ZN(n15261) );
  OR2_X1 U18143 ( .A1(n14741), .A2(n15261), .ZN(n14572) );
  NAND2_X1 U18144 ( .A1(n14573), .A2(n14572), .ZN(n14595) );
  AOI22_X1 U18145 ( .A1(n14735), .A2(n16338), .B1(n16341), .B2(n14595), .ZN(
        n14575) );
  AOI22_X1 U18146 ( .A1(n14597), .A2(n16339), .B1(n14596), .B2(n16340), .ZN(
        n14574) );
  OAI211_X1 U18147 ( .C1(n14601), .C2(n14576), .A(n14575), .B(n14574), .ZN(
        P1_U3098) );
  INV_X1 U18148 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14579) );
  AOI22_X1 U18149 ( .A1(n14735), .A2(n15300), .B1(n14814), .B2(n14595), .ZN(
        n14578) );
  AOI22_X1 U18150 ( .A1(n14597), .A2(n15296), .B1(n14596), .B2(n15070), .ZN(
        n14577) );
  OAI211_X1 U18151 ( .C1(n14601), .C2(n14579), .A(n14578), .B(n14577), .ZN(
        P1_U3102) );
  INV_X1 U18152 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14582) );
  AOI22_X1 U18153 ( .A1(n14735), .A2(n15293), .B1(n14823), .B2(n14595), .ZN(
        n14581) );
  AOI22_X1 U18154 ( .A1(n14597), .A2(n15289), .B1(n14596), .B2(n15063), .ZN(
        n14580) );
  OAI211_X1 U18155 ( .C1(n14601), .C2(n14582), .A(n14581), .B(n14580), .ZN(
        P1_U3104) );
  INV_X1 U18156 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U18157 ( .A1(n14735), .A2(n15317), .B1(n14818), .B2(n14595), .ZN(
        n14584) );
  AOI22_X1 U18158 ( .A1(n14597), .A2(n15311), .B1(n14596), .B2(n15021), .ZN(
        n14583) );
  OAI211_X1 U18159 ( .C1(n14601), .C2(n14585), .A(n14584), .B(n14583), .ZN(
        P1_U3099) );
  INV_X1 U18160 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14588) );
  AOI22_X1 U18161 ( .A1(n14735), .A2(n15266), .B1(n15271), .B2(n14595), .ZN(
        n14587) );
  AOI22_X1 U18162 ( .A1(n14597), .A2(n15265), .B1(n14596), .B2(n15028), .ZN(
        n14586) );
  OAI211_X1 U18163 ( .C1(n14601), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        P1_U3097) );
  INV_X1 U18164 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14591) );
  AOI22_X1 U18165 ( .A1(n14735), .A2(n16346), .B1(n16349), .B2(n14595), .ZN(
        n14590) );
  AOI22_X1 U18166 ( .A1(n14597), .A2(n16347), .B1(n14596), .B2(n16348), .ZN(
        n14589) );
  OAI211_X1 U18167 ( .C1(n14601), .C2(n14591), .A(n14590), .B(n14589), .ZN(
        P1_U3101) );
  INV_X1 U18168 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14594) );
  AOI22_X1 U18169 ( .A1(n14735), .A2(n15307), .B1(n14810), .B2(n14595), .ZN(
        n14593) );
  AOI22_X1 U18170 ( .A1(n14597), .A2(n15303), .B1(n14596), .B2(n15078), .ZN(
        n14592) );
  OAI211_X1 U18171 ( .C1(n14601), .C2(n14594), .A(n14593), .B(n14592), .ZN(
        P1_U3100) );
  INV_X1 U18172 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14600) );
  AOI22_X1 U18173 ( .A1(n14735), .A2(n16354), .B1(n16362), .B2(n14595), .ZN(
        n14599) );
  AOI22_X1 U18174 ( .A1(n14597), .A2(n16356), .B1(n14596), .B2(n16360), .ZN(
        n14598) );
  OAI211_X1 U18175 ( .C1(n14601), .C2(n14600), .A(n14599), .B(n14598), .ZN(
        P1_U3103) );
  AND2_X1 U18176 ( .A1(n14509), .A2(n14602), .ZN(n14605) );
  OAI211_X1 U18177 ( .C1(n14605), .C2(n14604), .A(n20435), .B(n14603), .ZN(
        n14611) );
  NAND2_X1 U18178 ( .A1(n14607), .A2(n14606), .ZN(n14608) );
  AND2_X1 U18179 ( .A1(n14609), .A2(n14608), .ZN(n20269) );
  NAND2_X1 U18180 ( .A1(n13216), .A2(n20269), .ZN(n14610) );
  OAI211_X1 U18181 ( .C1(n13216), .C2(n20266), .A(n14611), .B(n14610), .ZN(
        P2_U2873) );
  XNOR2_X1 U18182 ( .A(n14612), .B(n14613), .ZN(n14628) );
  INV_X1 U18183 ( .A(n14614), .ZN(n15384) );
  AOI21_X1 U18184 ( .B1(n14615), .B2(n15384), .A(n15383), .ZN(n14616) );
  OAI21_X1 U18185 ( .B1(n14617), .B2(n14618), .A(n14616), .ZN(n14962) );
  INV_X1 U18186 ( .A(n14618), .ZN(n14619) );
  NOR2_X1 U18187 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14619), .ZN(
        n14963) );
  AOI22_X1 U18188 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14962), .B1(
        n14963), .B2(n14620), .ZN(n14622) );
  INV_X1 U18189 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21467) );
  NOR2_X1 U18190 ( .A1(n17352), .A2(n21467), .ZN(n14624) );
  AOI21_X1 U18191 ( .B1(n21427), .B2(n21318), .A(n14624), .ZN(n14621) );
  OAI211_X1 U18192 ( .C1(n17365), .C2(n14628), .A(n14622), .B(n14621), .ZN(
        P1_U3026) );
  INV_X1 U18193 ( .A(n14623), .ZN(n21322) );
  AOI21_X1 U18194 ( .B1(n14161), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n14624), .ZN(n14625) );
  OAI21_X1 U18195 ( .B1(n17305), .B2(n21325), .A(n14625), .ZN(n14626) );
  AOI21_X1 U18196 ( .B1(n21322), .B2(n17298), .A(n14626), .ZN(n14627) );
  OAI21_X1 U18197 ( .B1(n17312), .B2(n14628), .A(n14627), .ZN(P1_U2994) );
  NAND2_X1 U18198 ( .A1(n21371), .A2(n17298), .ZN(n14633) );
  NOR2_X1 U18199 ( .A1(n15759), .A2(n14629), .ZN(n14630) );
  AOI211_X1 U18200 ( .C1(n17296), .C2(n21340), .A(n14631), .B(n14630), .ZN(
        n14632) );
  OAI211_X1 U18201 ( .C1(n14634), .C2(n17312), .A(n14633), .B(n14632), .ZN(
        P1_U2995) );
  NOR2_X1 U18202 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14635), .ZN(
        n14697) );
  INV_X1 U18203 ( .A(n14697), .ZN(n14678) );
  OAI21_X1 U18204 ( .B1(n14693), .B2(n16355), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14636) );
  INV_X1 U18205 ( .A(n13865), .ZN(n14997) );
  NAND2_X1 U18206 ( .A1(n15255), .A2(n14997), .ZN(n14639) );
  AOI21_X1 U18207 ( .B1(n14636), .B2(n14639), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n14638) );
  AND2_X1 U18208 ( .A1(n14637), .A2(n14741), .ZN(n15263) );
  NAND2_X1 U18209 ( .A1(n14796), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14641) );
  NAND2_X1 U18210 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14641), .ZN(n14901) );
  OAI211_X1 U18211 ( .C1(n14638), .C2(n14697), .A(n15263), .B(n14901), .ZN(
        n14684) );
  NAND2_X1 U18212 ( .A1(n14684), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14647) );
  INV_X1 U18213 ( .A(n14693), .ZN(n14644) );
  INV_X1 U18214 ( .A(n14639), .ZN(n14640) );
  NAND2_X1 U18215 ( .A1(n14640), .A2(n16320), .ZN(n14643) );
  INV_X1 U18216 ( .A(n14641), .ZN(n14896) );
  NAND2_X1 U18217 ( .A1(n14896), .A2(n14833), .ZN(n14642) );
  OAI22_X1 U18218 ( .A1(n14644), .A2(n15025), .B1(n14695), .B2(n15030), .ZN(
        n14645) );
  AOI21_X1 U18219 ( .B1(n16355), .B2(n15265), .A(n14645), .ZN(n14646) );
  OAI211_X1 U18220 ( .C1(n15269), .C2(n14678), .A(n14647), .B(n14646), .ZN(
        P1_U3145) );
  OAI21_X1 U18221 ( .B1(n20838), .B2(n20700), .A(n21177), .ZN(n14651) );
  NOR2_X1 U18222 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16970) );
  NAND2_X1 U18223 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16970), .ZN(
        n14654) );
  INV_X1 U18224 ( .A(n14648), .ZN(n14652) );
  INV_X1 U18225 ( .A(n16970), .ZN(n20619) );
  NOR2_X1 U18226 ( .A1(n20619), .A2(n14649), .ZN(n20660) );
  OAI21_X1 U18227 ( .B1(n14652), .B2(n20660), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14650) );
  OAI21_X1 U18228 ( .B1(n14651), .B2(n14654), .A(n14650), .ZN(n20662) );
  INV_X1 U18229 ( .A(n20662), .ZN(n14662) );
  INV_X1 U18230 ( .A(n21021), .ZN(n14661) );
  INV_X1 U18231 ( .A(n14651), .ZN(n14655) );
  AOI211_X1 U18232 ( .C1(n14652), .C2(n20975), .A(n21177), .B(n20660), .ZN(
        n14653) );
  INV_X1 U18233 ( .A(n20666), .ZN(n14659) );
  INV_X1 U18234 ( .A(n21030), .ZN(n14657) );
  NOR2_X2 U18235 ( .A1(n20838), .A2(n20672), .ZN(n20661) );
  AOI22_X1 U18236 ( .A1(n20944), .A2(n20661), .B1(n21020), .B2(n20660), .ZN(
        n14656) );
  OAI21_X1 U18237 ( .B1(n14657), .B2(n20698), .A(n14656), .ZN(n14658) );
  AOI21_X1 U18238 ( .B1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B2(n14659), .A(
        n14658), .ZN(n14660) );
  OAI21_X1 U18239 ( .B1(n14662), .B2(n14661), .A(n14660), .ZN(P2_U3072) );
  NOR2_X1 U18240 ( .A1(n15298), .A2(n14678), .ZN(n14666) );
  NAND2_X1 U18241 ( .A1(n16355), .A2(n15296), .ZN(n14664) );
  NAND2_X1 U18242 ( .A1(n14693), .A2(n15300), .ZN(n14663) );
  OAI211_X1 U18243 ( .C1(n14695), .C2(n15302), .A(n14664), .B(n14663), .ZN(
        n14665) );
  AOI211_X1 U18244 ( .C1(n14684), .C2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n14666), .B(n14665), .ZN(n14667) );
  INV_X1 U18245 ( .A(n14667), .ZN(P1_U3150) );
  NOR2_X1 U18246 ( .A1(n15291), .A2(n14678), .ZN(n14671) );
  NAND2_X1 U18247 ( .A1(n16355), .A2(n15289), .ZN(n14669) );
  NAND2_X1 U18248 ( .A1(n14693), .A2(n15293), .ZN(n14668) );
  OAI211_X1 U18249 ( .C1(n14695), .C2(n15295), .A(n14669), .B(n14668), .ZN(
        n14670) );
  AOI211_X1 U18250 ( .C1(n14684), .C2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n14671), .B(n14670), .ZN(n14672) );
  INV_X1 U18251 ( .A(n14672), .ZN(P1_U3152) );
  NOR2_X1 U18252 ( .A1(n15305), .A2(n14678), .ZN(n14676) );
  NAND2_X1 U18253 ( .A1(n16355), .A2(n15303), .ZN(n14674) );
  NAND2_X1 U18254 ( .A1(n14693), .A2(n15307), .ZN(n14673) );
  OAI211_X1 U18255 ( .C1(n14695), .C2(n15309), .A(n14674), .B(n14673), .ZN(
        n14675) );
  AOI211_X1 U18256 ( .C1(n14684), .C2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n14676), .B(n14675), .ZN(n14677) );
  INV_X1 U18257 ( .A(n14677), .ZN(P1_U3148) );
  NOR2_X1 U18258 ( .A1(n15315), .A2(n14678), .ZN(n14682) );
  NAND2_X1 U18259 ( .A1(n16355), .A2(n15311), .ZN(n14680) );
  NAND2_X1 U18260 ( .A1(n14693), .A2(n15317), .ZN(n14679) );
  OAI211_X1 U18261 ( .C1(n14695), .C2(n15320), .A(n14680), .B(n14679), .ZN(
        n14681) );
  AOI211_X1 U18262 ( .C1(n14684), .C2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n14682), .B(n14681), .ZN(n14683) );
  INV_X1 U18263 ( .A(n14683), .ZN(P1_U3147) );
  INV_X1 U18264 ( .A(n14684), .ZN(n14700) );
  INV_X1 U18265 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14688) );
  AOI22_X1 U18266 ( .A1(n14693), .A2(n16338), .B1(n16355), .B2(n16339), .ZN(
        n14685) );
  OAI21_X1 U18267 ( .B1(n14695), .B2(n15288), .A(n14685), .ZN(n14686) );
  AOI21_X1 U18268 ( .B1(n16340), .B2(n14697), .A(n14686), .ZN(n14687) );
  OAI21_X1 U18269 ( .B1(n14700), .B2(n14688), .A(n14687), .ZN(P1_U3146) );
  INV_X1 U18270 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14692) );
  AOI22_X1 U18271 ( .A1(n14693), .A2(n16346), .B1(n16355), .B2(n16347), .ZN(
        n14689) );
  OAI21_X1 U18272 ( .B1(n14695), .B2(n15283), .A(n14689), .ZN(n14690) );
  AOI21_X1 U18273 ( .B1(n16348), .B2(n14697), .A(n14690), .ZN(n14691) );
  OAI21_X1 U18274 ( .B1(n14700), .B2(n14692), .A(n14691), .ZN(P1_U3149) );
  INV_X1 U18275 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14699) );
  AOI22_X1 U18276 ( .A1(n14693), .A2(n16354), .B1(n16355), .B2(n16356), .ZN(
        n14694) );
  OAI21_X1 U18277 ( .B1(n14695), .B2(n15278), .A(n14694), .ZN(n14696) );
  AOI21_X1 U18278 ( .B1(n16360), .B2(n14697), .A(n14696), .ZN(n14698) );
  OAI21_X1 U18279 ( .B1(n14700), .B2(n14699), .A(n14698), .ZN(P1_U3151) );
  INV_X1 U18280 ( .A(n14701), .ZN(n14836) );
  INV_X1 U18281 ( .A(n14702), .ZN(n14707) );
  NOR2_X1 U18282 ( .A1(n14703), .A2(n16319), .ZN(n16331) );
  INV_X1 U18283 ( .A(n14704), .ZN(n14734) );
  OAI21_X1 U18284 ( .B1(n14832), .B2(n14705), .A(n14704), .ZN(n14709) );
  NOR3_X1 U18285 ( .A1(n16331), .A2(n16334), .A3(n14709), .ZN(n14706) );
  AOI211_X2 U18286 ( .C1(n16334), .C2(n14836), .A(n14707), .B(n14706), .ZN(
        n14739) );
  INV_X1 U18287 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14713) );
  INV_X1 U18288 ( .A(n14709), .ZN(n14710) );
  OAI22_X1 U18289 ( .A1(n14710), .A2(n16334), .B1(n14836), .B2(n21441), .ZN(
        n14732) );
  AOI22_X1 U18290 ( .A1(n14733), .A2(n15293), .B1(n14823), .B2(n14732), .ZN(
        n14712) );
  AOI22_X1 U18291 ( .A1(n14735), .A2(n15289), .B1(n14734), .B2(n15063), .ZN(
        n14711) );
  OAI211_X1 U18292 ( .C1(n14739), .C2(n14713), .A(n14712), .B(n14711), .ZN(
        P1_U3096) );
  INV_X1 U18293 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U18294 ( .A1(n14733), .A2(n16338), .B1(n16341), .B2(n14732), .ZN(
        n14715) );
  AOI22_X1 U18295 ( .A1(n14735), .A2(n16339), .B1(n14734), .B2(n16340), .ZN(
        n14714) );
  OAI211_X1 U18296 ( .C1(n14739), .C2(n14716), .A(n14715), .B(n14714), .ZN(
        P1_U3090) );
  INV_X1 U18297 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14719) );
  AOI22_X1 U18298 ( .A1(n14733), .A2(n15307), .B1(n14810), .B2(n14732), .ZN(
        n14718) );
  AOI22_X1 U18299 ( .A1(n14735), .A2(n15303), .B1(n14734), .B2(n15078), .ZN(
        n14717) );
  OAI211_X1 U18300 ( .C1(n14739), .C2(n14719), .A(n14718), .B(n14717), .ZN(
        P1_U3092) );
  INV_X1 U18301 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14722) );
  AOI22_X1 U18302 ( .A1(n14733), .A2(n16354), .B1(n16362), .B2(n14732), .ZN(
        n14721) );
  AOI22_X1 U18303 ( .A1(n14735), .A2(n16356), .B1(n14734), .B2(n16360), .ZN(
        n14720) );
  OAI211_X1 U18304 ( .C1(n14739), .C2(n14722), .A(n14721), .B(n14720), .ZN(
        P1_U3095) );
  INV_X1 U18305 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14725) );
  AOI22_X1 U18306 ( .A1(n14733), .A2(n15266), .B1(n15271), .B2(n14732), .ZN(
        n14724) );
  AOI22_X1 U18307 ( .A1(n14735), .A2(n15265), .B1(n14734), .B2(n15028), .ZN(
        n14723) );
  OAI211_X1 U18308 ( .C1(n14739), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        P1_U3089) );
  INV_X1 U18309 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14728) );
  AOI22_X1 U18310 ( .A1(n14733), .A2(n15300), .B1(n14814), .B2(n14732), .ZN(
        n14727) );
  AOI22_X1 U18311 ( .A1(n14735), .A2(n15296), .B1(n14734), .B2(n15070), .ZN(
        n14726) );
  OAI211_X1 U18312 ( .C1(n14739), .C2(n14728), .A(n14727), .B(n14726), .ZN(
        P1_U3094) );
  INV_X1 U18313 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14731) );
  AOI22_X1 U18314 ( .A1(n14733), .A2(n16346), .B1(n16349), .B2(n14732), .ZN(
        n14730) );
  AOI22_X1 U18315 ( .A1(n14735), .A2(n16347), .B1(n14734), .B2(n16348), .ZN(
        n14729) );
  OAI211_X1 U18316 ( .C1(n14739), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        P1_U3093) );
  INV_X1 U18317 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14738) );
  AOI22_X1 U18318 ( .A1(n14733), .A2(n15317), .B1(n14818), .B2(n14732), .ZN(
        n14737) );
  AOI22_X1 U18319 ( .A1(n14735), .A2(n15311), .B1(n14734), .B2(n15021), .ZN(
        n14736) );
  OAI211_X1 U18320 ( .C1(n14739), .C2(n14738), .A(n14737), .B(n14736), .ZN(
        P1_U3091) );
  NAND2_X1 U18321 ( .A1(n14772), .A2(n14748), .ZN(n14740) );
  AOI21_X1 U18322 ( .B1(n14740), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n16334), 
        .ZN(n14745) );
  NOR2_X1 U18323 ( .A1(n14998), .A2(n13865), .ZN(n14742) );
  INV_X1 U18324 ( .A(n14741), .ZN(n15000) );
  NAND2_X1 U18325 ( .A1(n14796), .A2(n17143), .ZN(n14746) );
  INV_X1 U18326 ( .A(n14746), .ZN(n14834) );
  AOI22_X1 U18327 ( .A1(n14745), .A2(n14742), .B1(n15000), .B2(n14834), .ZN(
        n14777) );
  INV_X1 U18328 ( .A(n14742), .ZN(n14744) );
  OR2_X1 U18329 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14743), .ZN(
        n14771) );
  AOI22_X1 U18330 ( .A1(n14745), .A2(n14744), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n14771), .ZN(n14747) );
  NAND2_X1 U18331 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14746), .ZN(n14840) );
  NAND3_X1 U18332 ( .A1(n15008), .A2(n14747), .A3(n14840), .ZN(n14770) );
  NAND2_X1 U18333 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14751) );
  OAI22_X1 U18334 ( .A1(n14772), .A2(n15060), .B1(n15291), .B2(n14771), .ZN(
        n14749) );
  AOI21_X1 U18335 ( .B1(n14774), .B2(n15289), .A(n14749), .ZN(n14750) );
  OAI211_X1 U18336 ( .C1(n14777), .C2(n15295), .A(n14751), .B(n14750), .ZN(
        P1_U3056) );
  NAND2_X1 U18337 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14754) );
  OAI22_X1 U18338 ( .A1(n14772), .A2(n15054), .B1(n15275), .B2(n14771), .ZN(
        n14752) );
  AOI21_X1 U18339 ( .B1(n14774), .B2(n16356), .A(n14752), .ZN(n14753) );
  OAI211_X1 U18340 ( .C1(n14777), .C2(n15278), .A(n14754), .B(n14753), .ZN(
        P1_U3055) );
  NAND2_X1 U18341 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14757) );
  OAI22_X1 U18342 ( .A1(n14772), .A2(n15018), .B1(n15315), .B2(n14771), .ZN(
        n14755) );
  AOI21_X1 U18343 ( .B1(n14774), .B2(n15311), .A(n14755), .ZN(n14756) );
  OAI211_X1 U18344 ( .C1(n14777), .C2(n15320), .A(n14757), .B(n14756), .ZN(
        P1_U3051) );
  NAND2_X1 U18345 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14760) );
  OAI22_X1 U18346 ( .A1(n14772), .A2(n15075), .B1(n15305), .B2(n14771), .ZN(
        n14758) );
  AOI21_X1 U18347 ( .B1(n14774), .B2(n15303), .A(n14758), .ZN(n14759) );
  OAI211_X1 U18348 ( .C1(n14777), .C2(n15309), .A(n14760), .B(n14759), .ZN(
        P1_U3052) );
  NAND2_X1 U18349 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n14763) );
  OAI22_X1 U18350 ( .A1(n14772), .A2(n15025), .B1(n15269), .B2(n14771), .ZN(
        n14761) );
  AOI21_X1 U18351 ( .B1(n14774), .B2(n15265), .A(n14761), .ZN(n14762) );
  OAI211_X1 U18352 ( .C1(n14777), .C2(n15030), .A(n14763), .B(n14762), .ZN(
        P1_U3049) );
  NAND2_X1 U18353 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14766) );
  OAI22_X1 U18354 ( .A1(n14772), .A2(n15012), .B1(n15285), .B2(n14771), .ZN(
        n14764) );
  AOI21_X1 U18355 ( .B1(n14774), .B2(n16339), .A(n14764), .ZN(n14765) );
  OAI211_X1 U18356 ( .C1(n14777), .C2(n15288), .A(n14766), .B(n14765), .ZN(
        P1_U3050) );
  NAND2_X1 U18357 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14769) );
  OAI22_X1 U18358 ( .A1(n14772), .A2(n15067), .B1(n15298), .B2(n14771), .ZN(
        n14767) );
  AOI21_X1 U18359 ( .B1(n14774), .B2(n15296), .A(n14767), .ZN(n14768) );
  OAI211_X1 U18360 ( .C1(n14777), .C2(n15302), .A(n14769), .B(n14768), .ZN(
        P1_U3054) );
  NAND2_X1 U18361 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14776) );
  OAI22_X1 U18362 ( .A1(n14772), .A2(n15048), .B1(n15280), .B2(n14771), .ZN(
        n14773) );
  AOI21_X1 U18363 ( .B1(n14774), .B2(n16347), .A(n14773), .ZN(n14775) );
  OAI211_X1 U18364 ( .C1(n14777), .C2(n15283), .A(n14776), .B(n14775), .ZN(
        P1_U3053) );
  NAND2_X1 U18365 ( .A1(n15196), .A2(n14778), .ZN(n14779) );
  XNOR2_X1 U18366 ( .A(n17581), .B(n14779), .ZN(n14780) );
  NAND2_X1 U18367 ( .A1(n14780), .A2(n20370), .ZN(n14788) );
  INV_X1 U18368 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n21118) );
  NAND2_X1 U18369 ( .A1(n20406), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n14783) );
  AOI22_X1 U18370 ( .A1(n20359), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20412), .ZN(n14782) );
  OAI211_X1 U18371 ( .C1(n14784), .C2(n20399), .A(n14783), .B(n14782), .ZN(
        n14786) );
  NOR2_X1 U18372 ( .A1(n21185), .A2(n20401), .ZN(n14785) );
  AOI211_X1 U18373 ( .C1(n20385), .C2(n12900), .A(n14786), .B(n14785), .ZN(
        n14787) );
  OAI211_X1 U18374 ( .C1(n20800), .C2(n20384), .A(n14788), .B(n14787), .ZN(
        P2_U2852) );
  OAI21_X1 U18375 ( .B1(n14824), .B2(n14826), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14790) );
  OAI21_X1 U18376 ( .B1(n14997), .B2(n14832), .A(n14790), .ZN(n14792) );
  NOR2_X1 U18377 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14791), .ZN(
        n14825) );
  AOI21_X1 U18378 ( .B1(n14792), .B2(n17400), .A(n14825), .ZN(n14794) );
  INV_X1 U18379 ( .A(n15263), .ZN(n14793) );
  INV_X1 U18380 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14800) );
  NAND2_X1 U18381 ( .A1(n13865), .A2(n16320), .ZN(n14797) );
  INV_X1 U18382 ( .A(n14833), .ZN(n15256) );
  OR2_X1 U18383 ( .A1(n14796), .A2(n14795), .ZN(n14999) );
  OAI22_X1 U18384 ( .A1(n14832), .A2(n14797), .B1(n15256), .B2(n14999), .ZN(
        n14822) );
  AOI22_X1 U18385 ( .A1(n14824), .A2(n16356), .B1(n16362), .B2(n14822), .ZN(
        n14799) );
  AOI22_X1 U18386 ( .A1(n14826), .A2(n16354), .B1(n16360), .B2(n14825), .ZN(
        n14798) );
  OAI211_X1 U18387 ( .C1(n14830), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        P1_U3071) );
  INV_X1 U18388 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14803) );
  AOI22_X1 U18389 ( .A1(n14824), .A2(n16347), .B1(n16349), .B2(n14822), .ZN(
        n14802) );
  AOI22_X1 U18390 ( .A1(n14826), .A2(n16346), .B1(n16348), .B2(n14825), .ZN(
        n14801) );
  OAI211_X1 U18391 ( .C1(n14830), .C2(n14803), .A(n14802), .B(n14801), .ZN(
        P1_U3069) );
  INV_X1 U18392 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14806) );
  AOI22_X1 U18393 ( .A1(n14824), .A2(n16339), .B1(n16341), .B2(n14822), .ZN(
        n14805) );
  AOI22_X1 U18394 ( .A1(n14826), .A2(n16338), .B1(n16340), .B2(n14825), .ZN(
        n14804) );
  OAI211_X1 U18395 ( .C1(n14830), .C2(n14806), .A(n14805), .B(n14804), .ZN(
        P1_U3066) );
  INV_X1 U18396 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U18397 ( .A1(n14824), .A2(n15265), .B1(n15271), .B2(n14822), .ZN(
        n14808) );
  AOI22_X1 U18398 ( .A1(n14826), .A2(n15266), .B1(n15028), .B2(n14825), .ZN(
        n14807) );
  OAI211_X1 U18399 ( .C1(n14830), .C2(n14809), .A(n14808), .B(n14807), .ZN(
        P1_U3065) );
  INV_X1 U18400 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14813) );
  AOI22_X1 U18401 ( .A1(n14824), .A2(n15303), .B1(n14810), .B2(n14822), .ZN(
        n14812) );
  AOI22_X1 U18402 ( .A1(n14826), .A2(n15307), .B1(n15078), .B2(n14825), .ZN(
        n14811) );
  OAI211_X1 U18403 ( .C1(n14830), .C2(n14813), .A(n14812), .B(n14811), .ZN(
        P1_U3068) );
  INV_X1 U18404 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14817) );
  AOI22_X1 U18405 ( .A1(n14824), .A2(n15296), .B1(n14814), .B2(n14822), .ZN(
        n14816) );
  AOI22_X1 U18406 ( .A1(n14826), .A2(n15300), .B1(n15070), .B2(n14825), .ZN(
        n14815) );
  OAI211_X1 U18407 ( .C1(n14830), .C2(n14817), .A(n14816), .B(n14815), .ZN(
        P1_U3070) );
  INV_X1 U18408 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14821) );
  AOI22_X1 U18409 ( .A1(n14824), .A2(n15311), .B1(n14818), .B2(n14822), .ZN(
        n14820) );
  AOI22_X1 U18410 ( .A1(n14826), .A2(n15317), .B1(n15021), .B2(n14825), .ZN(
        n14819) );
  OAI211_X1 U18411 ( .C1(n14830), .C2(n14821), .A(n14820), .B(n14819), .ZN(
        P1_U3067) );
  INV_X1 U18412 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14829) );
  AOI22_X1 U18413 ( .A1(n14824), .A2(n15289), .B1(n14823), .B2(n14822), .ZN(
        n14828) );
  AOI22_X1 U18414 ( .A1(n14826), .A2(n15293), .B1(n15063), .B2(n14825), .ZN(
        n14827) );
  OAI211_X1 U18415 ( .C1(n14830), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        P1_U3072) );
  NAND3_X1 U18416 ( .A1(n14865), .A2(n14864), .A3(n16320), .ZN(n14831) );
  NAND2_X1 U18417 ( .A1(n16320), .A2(n21254), .ZN(n15252) );
  NAND2_X1 U18418 ( .A1(n14831), .A2(n15252), .ZN(n14839) );
  NOR2_X1 U18419 ( .A1(n14832), .A2(n13865), .ZN(n14835) );
  AOI22_X1 U18420 ( .A1(n14839), .A2(n14835), .B1(n14834), .B2(n14833), .ZN(
        n14870) );
  INV_X1 U18421 ( .A(n14835), .ZN(n14838) );
  NOR2_X1 U18422 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14836), .ZN(
        n14867) );
  INV_X1 U18423 ( .A(n14867), .ZN(n14837) );
  AOI22_X1 U18424 ( .A1(n14839), .A2(n14838), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n14837), .ZN(n14841) );
  NAND3_X1 U18425 ( .A1(n15263), .A2(n14841), .A3(n14840), .ZN(n14863) );
  NAND2_X1 U18426 ( .A1(n14863), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n14844) );
  OAI22_X1 U18427 ( .A1(n15018), .A2(n14865), .B1(n14864), .B2(n15016), .ZN(
        n14842) );
  AOI21_X1 U18428 ( .B1(n15021), .B2(n14867), .A(n14842), .ZN(n14843) );
  OAI211_X1 U18429 ( .C1(n14870), .C2(n15320), .A(n14844), .B(n14843), .ZN(
        P1_U3083) );
  NAND2_X1 U18430 ( .A1(n14863), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14847) );
  OAI22_X1 U18431 ( .A1(n15054), .A2(n14865), .B1(n14864), .B2(n15052), .ZN(
        n14845) );
  AOI21_X1 U18432 ( .B1(n16360), .B2(n14867), .A(n14845), .ZN(n14846) );
  OAI211_X1 U18433 ( .C1(n14870), .C2(n15278), .A(n14847), .B(n14846), .ZN(
        P1_U3087) );
  NAND2_X1 U18434 ( .A1(n14863), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14850) );
  OAI22_X1 U18435 ( .A1(n15075), .A2(n14865), .B1(n14864), .B2(n15072), .ZN(
        n14848) );
  AOI21_X1 U18436 ( .B1(n15078), .B2(n14867), .A(n14848), .ZN(n14849) );
  OAI211_X1 U18437 ( .C1(n14870), .C2(n15309), .A(n14850), .B(n14849), .ZN(
        P1_U3084) );
  NAND2_X1 U18438 ( .A1(n14863), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14853) );
  OAI22_X1 U18439 ( .A1(n15025), .A2(n14865), .B1(n14864), .B2(n15023), .ZN(
        n14851) );
  AOI21_X1 U18440 ( .B1(n15028), .B2(n14867), .A(n14851), .ZN(n14852) );
  OAI211_X1 U18441 ( .C1(n14870), .C2(n15030), .A(n14853), .B(n14852), .ZN(
        P1_U3081) );
  NAND2_X1 U18442 ( .A1(n14863), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14856) );
  OAI22_X1 U18443 ( .A1(n15012), .A2(n14865), .B1(n14864), .B2(n15002), .ZN(
        n14854) );
  AOI21_X1 U18444 ( .B1(n16340), .B2(n14867), .A(n14854), .ZN(n14855) );
  OAI211_X1 U18445 ( .C1(n14870), .C2(n15288), .A(n14856), .B(n14855), .ZN(
        P1_U3082) );
  NAND2_X1 U18446 ( .A1(n14863), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14859) );
  OAI22_X1 U18447 ( .A1(n15048), .A2(n14865), .B1(n14864), .B2(n15046), .ZN(
        n14857) );
  AOI21_X1 U18448 ( .B1(n16348), .B2(n14867), .A(n14857), .ZN(n14858) );
  OAI211_X1 U18449 ( .C1(n14870), .C2(n15283), .A(n14859), .B(n14858), .ZN(
        P1_U3085) );
  NAND2_X1 U18450 ( .A1(n14863), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14862) );
  OAI22_X1 U18451 ( .A1(n15060), .A2(n14865), .B1(n14864), .B2(n15058), .ZN(
        n14860) );
  AOI21_X1 U18452 ( .B1(n15063), .B2(n14867), .A(n14860), .ZN(n14861) );
  OAI211_X1 U18453 ( .C1(n14870), .C2(n15295), .A(n14862), .B(n14861), .ZN(
        P1_U3088) );
  NAND2_X1 U18454 ( .A1(n14863), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14869) );
  OAI22_X1 U18455 ( .A1(n15067), .A2(n14865), .B1(n14864), .B2(n15065), .ZN(
        n14866) );
  AOI21_X1 U18456 ( .B1(n15070), .B2(n14867), .A(n14866), .ZN(n14868) );
  OAI211_X1 U18457 ( .C1(n14870), .C2(n15302), .A(n14869), .B(n14868), .ZN(
        P1_U3086) );
  XNOR2_X1 U18458 ( .A(n14603), .B(n14871), .ZN(n14873) );
  MUX2_X1 U18459 ( .A(n11912), .B(n17507), .S(n20437), .Z(n14872) );
  OAI21_X1 U18460 ( .B1(n14873), .B2(n20428), .A(n14872), .ZN(P2_U2872) );
  NOR2_X1 U18461 ( .A1(n12815), .A2(n14949), .ZN(n14875) );
  XNOR2_X1 U18462 ( .A(n14875), .B(n14874), .ZN(n14876) );
  NAND2_X1 U18463 ( .A1(n14876), .A2(n20370), .ZN(n14886) );
  OAI22_X1 U18464 ( .A1(n20396), .A2(n14878), .B1(n14877), .B2(n20380), .ZN(
        n14879) );
  AOI21_X1 U18465 ( .B1(n20328), .B2(n14880), .A(n14879), .ZN(n14881) );
  OAI21_X1 U18466 ( .B1(n20374), .B2(n21116), .A(n14881), .ZN(n14884) );
  NOR2_X1 U18467 ( .A1(n14882), .A2(n20401), .ZN(n14883) );
  AOI211_X1 U18468 ( .C1(n20385), .C2(n16946), .A(n14884), .B(n14883), .ZN(
        n14885) );
  OAI211_X1 U18469 ( .C1(n21190), .C2(n20384), .A(n14886), .B(n14885), .ZN(
        P2_U2853) );
  AOI21_X1 U18470 ( .B1(n14888), .B2(n14515), .A(n14887), .ZN(n21299) );
  INV_X1 U18471 ( .A(n21299), .ZN(n14892) );
  INV_X1 U18472 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14891) );
  OR2_X1 U18473 ( .A1(n14979), .A2(n14889), .ZN(n14890) );
  NAND2_X1 U18474 ( .A1(n15142), .A2(n14890), .ZN(n21295) );
  OAI222_X1 U18475 ( .A1(n14892), .A2(n17250), .B1(n21381), .B2(n14891), .C1(
        n21295), .C2(n15641), .ZN(P1_U2865) );
  OAI222_X1 U18476 ( .A1(n15739), .A2(n14892), .B1(n15733), .B2(n10733), .C1(
        n15732), .C2(n15681), .ZN(P1_U2897) );
  NAND2_X1 U18477 ( .A1(n14925), .A2(n16320), .ZN(n14894) );
  INV_X1 U18478 ( .A(n14926), .ZN(n14893) );
  OAI21_X1 U18479 ( .B1(n14894), .B2(n14893), .A(n15252), .ZN(n14900) );
  AND2_X1 U18480 ( .A1(n14895), .A2(n14997), .ZN(n14898) );
  OR2_X1 U18481 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14897), .ZN(
        n14924) );
  INV_X1 U18482 ( .A(n14898), .ZN(n14899) );
  AOI22_X1 U18483 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n14924), .B1(n14900), 
        .B2(n14899), .ZN(n14902) );
  NAND3_X1 U18484 ( .A1(n15008), .A2(n14902), .A3(n14901), .ZN(n14929) );
  NOR2_X1 U18485 ( .A1(n15291), .A2(n14924), .ZN(n14904) );
  OAI22_X1 U18486 ( .A1(n15060), .A2(n14926), .B1(n14925), .B2(n15058), .ZN(
        n14903) );
  AOI211_X1 U18487 ( .C1(n14929), .C2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n14904), .B(n14903), .ZN(n14905) );
  OAI21_X1 U18488 ( .B1(n14931), .B2(n15295), .A(n14905), .ZN(P1_U3120) );
  NOR2_X1 U18489 ( .A1(n15298), .A2(n14924), .ZN(n14907) );
  OAI22_X1 U18490 ( .A1(n15067), .A2(n14926), .B1(n14925), .B2(n15065), .ZN(
        n14906) );
  AOI211_X1 U18491 ( .C1(n14929), .C2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n14907), .B(n14906), .ZN(n14908) );
  OAI21_X1 U18492 ( .B1(n14931), .B2(n15302), .A(n14908), .ZN(P1_U3118) );
  NOR2_X1 U18493 ( .A1(n15305), .A2(n14924), .ZN(n14910) );
  OAI22_X1 U18494 ( .A1(n15075), .A2(n14926), .B1(n14925), .B2(n15072), .ZN(
        n14909) );
  AOI211_X1 U18495 ( .C1(n14929), .C2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n14910), .B(n14909), .ZN(n14911) );
  OAI21_X1 U18496 ( .B1(n14931), .B2(n15309), .A(n14911), .ZN(P1_U3116) );
  NOR2_X1 U18497 ( .A1(n15315), .A2(n14924), .ZN(n14913) );
  OAI22_X1 U18498 ( .A1(n15018), .A2(n14926), .B1(n14925), .B2(n15016), .ZN(
        n14912) );
  AOI211_X1 U18499 ( .C1(n14929), .C2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n14913), .B(n14912), .ZN(n14914) );
  OAI21_X1 U18500 ( .B1(n14931), .B2(n15320), .A(n14914), .ZN(P1_U3115) );
  NOR2_X1 U18501 ( .A1(n15275), .A2(n14924), .ZN(n14916) );
  OAI22_X1 U18502 ( .A1(n15054), .A2(n14926), .B1(n14925), .B2(n15052), .ZN(
        n14915) );
  AOI211_X1 U18503 ( .C1(n14929), .C2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n14916), .B(n14915), .ZN(n14917) );
  OAI21_X1 U18504 ( .B1(n14931), .B2(n15278), .A(n14917), .ZN(P1_U3119) );
  NOR2_X1 U18505 ( .A1(n15285), .A2(n14924), .ZN(n14919) );
  OAI22_X1 U18506 ( .A1(n15012), .A2(n14926), .B1(n14925), .B2(n15002), .ZN(
        n14918) );
  AOI211_X1 U18507 ( .C1(n14929), .C2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n14919), .B(n14918), .ZN(n14920) );
  OAI21_X1 U18508 ( .B1(n14931), .B2(n15288), .A(n14920), .ZN(P1_U3114) );
  NOR2_X1 U18509 ( .A1(n15280), .A2(n14924), .ZN(n14922) );
  OAI22_X1 U18510 ( .A1(n15048), .A2(n14926), .B1(n14925), .B2(n15046), .ZN(
        n14921) );
  AOI211_X1 U18511 ( .C1(n14929), .C2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n14922), .B(n14921), .ZN(n14923) );
  OAI21_X1 U18512 ( .B1(n14931), .B2(n15283), .A(n14923), .ZN(P1_U3117) );
  NOR2_X1 U18513 ( .A1(n15269), .A2(n14924), .ZN(n14928) );
  OAI22_X1 U18514 ( .A1(n15025), .A2(n14926), .B1(n14925), .B2(n15023), .ZN(
        n14927) );
  AOI211_X1 U18515 ( .C1(n14929), .C2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n14928), .B(n14927), .ZN(n14930) );
  OAI21_X1 U18516 ( .B1(n14931), .B2(n15030), .A(n14930), .ZN(P1_U3113) );
  XNOR2_X1 U18517 ( .A(n14932), .B(n14933), .ZN(n15088) );
  NOR2_X1 U18518 ( .A1(n14934), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15082) );
  INV_X1 U18519 ( .A(n15082), .ZN(n14936) );
  NAND3_X1 U18520 ( .A1(n14936), .A2(n12521), .A3(n14935), .ZN(n14948) );
  INV_X1 U18521 ( .A(n14937), .ZN(n14941) );
  INV_X1 U18522 ( .A(n14938), .ZN(n14940) );
  INV_X1 U18523 ( .A(n15231), .ZN(n14939) );
  OAI21_X1 U18524 ( .B1(n14941), .B2(n14940), .A(n14939), .ZN(n15083) );
  INV_X1 U18525 ( .A(n15083), .ZN(n20434) );
  AOI22_X1 U18526 ( .A1(n20376), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n17633), 
        .B2(n15942), .ZN(n14942) );
  OAI21_X1 U18527 ( .B1(n17671), .B2(n14943), .A(n14942), .ZN(n14946) );
  OAI21_X1 U18528 ( .B1(n17662), .B2(n17664), .A(n14944), .ZN(n15241) );
  NOR2_X1 U18529 ( .A1(n15241), .A2(n15942), .ZN(n14945) );
  AOI211_X1 U18530 ( .C1(n20434), .C2(n12878), .A(n14946), .B(n14945), .ZN(
        n14947) );
  OAI211_X1 U18531 ( .C1(n15088), .C2(n17681), .A(n14948), .B(n14947), .ZN(
        P2_U3042) );
  AOI211_X1 U18532 ( .C1(n20409), .C2(n14950), .A(n15194), .B(n14949), .ZN(
        n15193) );
  INV_X1 U18533 ( .A(n14951), .ZN(n20411) );
  INV_X1 U18534 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16707) );
  AOI22_X1 U18535 ( .A1(n15193), .A2(n20370), .B1(n20411), .B2(n16707), .ZN(
        n14959) );
  INV_X1 U18536 ( .A(n16709), .ZN(n14954) );
  OAI22_X1 U18537 ( .A1(n20396), .A2(n14952), .B1(n16707), .B2(n20380), .ZN(
        n14953) );
  AOI21_X1 U18538 ( .B1(n20328), .B2(n14954), .A(n14953), .ZN(n14956) );
  INV_X1 U18539 ( .A(n20401), .ZN(n20378) );
  NAND2_X1 U18540 ( .A1(n20378), .A2(n21201), .ZN(n14955) );
  OAI211_X1 U18541 ( .C1(n20374), .C2(n21114), .A(n14956), .B(n14955), .ZN(
        n14957) );
  AOI21_X1 U18542 ( .B1(n9818), .B2(n20385), .A(n14957), .ZN(n14958) );
  OAI211_X1 U18543 ( .C1(n20384), .C2(n16968), .A(n14959), .B(n14958), .ZN(
        P2_U2854) );
  XNOR2_X1 U18544 ( .A(n14960), .B(n14961), .ZN(n14972) );
  AOI211_X1 U18545 ( .C1(n14964), .C2(n14963), .A(n14982), .B(n14962), .ZN(
        n14980) );
  NOR2_X1 U18546 ( .A1(n16263), .A2(n14980), .ZN(n15140) );
  NOR2_X1 U18547 ( .A1(n17364), .A2(n21295), .ZN(n14966) );
  INV_X1 U18548 ( .A(n14981), .ZN(n17375) );
  NAND2_X1 U18549 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17375), .ZN(
        n15136) );
  INV_X1 U18550 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21470) );
  OR2_X1 U18551 ( .A1(n17352), .A2(n21470), .ZN(n14969) );
  OAI21_X1 U18552 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15136), .A(
        n14969), .ZN(n14965) );
  AOI211_X1 U18553 ( .C1(n15140), .C2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n14966), .B(n14965), .ZN(n14967) );
  OAI21_X1 U18554 ( .B1(n17365), .B2(n14972), .A(n14967), .ZN(P1_U3024) );
  NAND2_X1 U18555 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14968) );
  OAI211_X1 U18556 ( .C1(n17305), .C2(n21302), .A(n14969), .B(n14968), .ZN(
        n14970) );
  AOI21_X1 U18557 ( .B1(n21299), .B2(n17298), .A(n14970), .ZN(n14971) );
  OAI21_X1 U18558 ( .B1(n17312), .B2(n14972), .A(n14971), .ZN(P1_U2992) );
  XOR2_X1 U18559 ( .A(n14973), .B(n14974), .Z(n14986) );
  AOI21_X1 U18560 ( .B1(n14977), .B2(n14976), .A(n14975), .ZN(n14978) );
  OR2_X1 U18561 ( .A1(n14979), .A2(n14978), .ZN(n21305) );
  INV_X1 U18562 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21468) );
  OAI22_X1 U18563 ( .A1(n17364), .A2(n21305), .B1(n21468), .B2(n17352), .ZN(
        n14984) );
  AOI21_X1 U18564 ( .B1(n14982), .B2(n14981), .A(n14980), .ZN(n14983) );
  AOI211_X1 U18565 ( .C1(n14986), .C2(n21429), .A(n14984), .B(n14983), .ZN(
        n14985) );
  INV_X1 U18566 ( .A(n14985), .ZN(P1_U3025) );
  NAND2_X1 U18567 ( .A1(n14986), .A2(n17267), .ZN(n14990) );
  OAI22_X1 U18568 ( .A1(n15759), .A2(n14987), .B1(n17352), .B2(n21468), .ZN(
        n14988) );
  AOI21_X1 U18569 ( .B1(n17296), .B2(n21311), .A(n14988), .ZN(n14989) );
  OAI211_X1 U18570 ( .C1(n17306), .C2(n21310), .A(n14990), .B(n14989), .ZN(
        P1_U2993) );
  AOI21_X1 U18571 ( .B1(n14993), .B2(n14991), .A(n14992), .ZN(n14994) );
  INV_X1 U18572 ( .A(n14994), .ZN(n21278) );
  AOI22_X1 U18573 ( .A1(n15737), .A2(n15671), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15736), .ZN(n14995) );
  OAI21_X1 U18574 ( .B1(n21278), .B2(n15739), .A(n14995), .ZN(P1_U2895) );
  NAND3_X1 U18575 ( .A1(n16337), .A2(n15073), .A3(n16320), .ZN(n14996) );
  NAND2_X1 U18576 ( .A1(n14996), .A2(n15252), .ZN(n15005) );
  NOR2_X1 U18577 ( .A1(n14998), .A2(n14997), .ZN(n15003) );
  INV_X1 U18578 ( .A(n14999), .ZN(n15009) );
  NOR2_X1 U18579 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15001), .ZN(
        n15079) );
  NOR2_X1 U18580 ( .A1(n15073), .A2(n15002), .ZN(n15014) );
  INV_X1 U18581 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15011) );
  INV_X1 U18582 ( .A(n15079), .ZN(n15006) );
  INV_X1 U18583 ( .A(n15003), .ZN(n15004) );
  AOI22_X1 U18584 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15006), .B1(n15005), 
        .B2(n15004), .ZN(n15007) );
  OAI211_X1 U18585 ( .C1(n15009), .C2(n21441), .A(n15008), .B(n15007), .ZN(
        n15010) );
  OAI22_X1 U18586 ( .A1(n16337), .A2(n15012), .B1(n15011), .B2(n15074), .ZN(
        n15013) );
  AOI211_X1 U18587 ( .C1(n15079), .C2(n16340), .A(n15014), .B(n15013), .ZN(
        n15015) );
  OAI21_X1 U18588 ( .B1(n15081), .B2(n15288), .A(n15015), .ZN(P1_U3034) );
  NOR2_X1 U18589 ( .A1(n15073), .A2(n15016), .ZN(n15020) );
  INV_X1 U18590 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15017) );
  OAI22_X1 U18591 ( .A1(n16337), .A2(n15018), .B1(n15017), .B2(n15074), .ZN(
        n15019) );
  AOI211_X1 U18592 ( .C1(n15079), .C2(n15021), .A(n15020), .B(n15019), .ZN(
        n15022) );
  OAI21_X1 U18593 ( .B1(n15081), .B2(n15320), .A(n15022), .ZN(P1_U3035) );
  NOR2_X1 U18594 ( .A1(n15073), .A2(n15023), .ZN(n15027) );
  OAI22_X1 U18595 ( .A1(n16337), .A2(n15025), .B1(n15024), .B2(n15074), .ZN(
        n15026) );
  AOI211_X1 U18596 ( .C1(n15028), .C2(n15079), .A(n15027), .B(n15026), .ZN(
        n15029) );
  OAI21_X1 U18597 ( .B1(n15081), .B2(n15030), .A(n15029), .ZN(P1_U3033) );
  XOR2_X1 U18598 ( .A(n15031), .B(n15032), .Z(n20455) );
  INV_X1 U18599 ( .A(n15033), .ZN(n15040) );
  NAND2_X1 U18600 ( .A1(n20411), .A2(n17524), .ZN(n15039) );
  INV_X1 U18601 ( .A(n16870), .ZN(n17525) );
  AOI21_X1 U18602 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n20412), .A(
        n20376), .ZN(n15035) );
  NAND2_X1 U18603 ( .A1(n20359), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n15034) );
  OAI211_X1 U18604 ( .C1(n20374), .C2(n15036), .A(n15035), .B(n15034), .ZN(
        n15037) );
  AOI21_X1 U18605 ( .B1(n20385), .B2(n17525), .A(n15037), .ZN(n15038) );
  OAI211_X1 U18606 ( .C1(n15040), .C2(n20399), .A(n15039), .B(n15038), .ZN(
        n15044) );
  OR2_X1 U18607 ( .A1(n15194), .A2(n15041), .ZN(n20264) );
  AOI211_X1 U18608 ( .C1(n17524), .C2(n15042), .A(n21086), .B(n20264), .ZN(
        n15043) );
  AOI211_X1 U18609 ( .C1(n20455), .C2(n20378), .A(n15044), .B(n15043), .ZN(
        n15045) );
  INV_X1 U18610 ( .A(n15045), .ZN(P2_U2842) );
  NOR2_X1 U18611 ( .A1(n15073), .A2(n15046), .ZN(n15050) );
  INV_X1 U18612 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15047) );
  OAI22_X1 U18613 ( .A1(n16337), .A2(n15048), .B1(n15047), .B2(n15074), .ZN(
        n15049) );
  AOI211_X1 U18614 ( .C1(n15079), .C2(n16348), .A(n15050), .B(n15049), .ZN(
        n15051) );
  OAI21_X1 U18615 ( .B1(n15081), .B2(n15283), .A(n15051), .ZN(P1_U3037) );
  NOR2_X1 U18616 ( .A1(n15073), .A2(n15052), .ZN(n15056) );
  INV_X1 U18617 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15053) );
  OAI22_X1 U18618 ( .A1(n16337), .A2(n15054), .B1(n15053), .B2(n15074), .ZN(
        n15055) );
  AOI211_X1 U18619 ( .C1(n15079), .C2(n16360), .A(n15056), .B(n15055), .ZN(
        n15057) );
  OAI21_X1 U18620 ( .B1(n15081), .B2(n15278), .A(n15057), .ZN(P1_U3039) );
  NOR2_X1 U18621 ( .A1(n15073), .A2(n15058), .ZN(n15062) );
  OAI22_X1 U18622 ( .A1(n16337), .A2(n15060), .B1(n15059), .B2(n15074), .ZN(
        n15061) );
  AOI211_X1 U18623 ( .C1(n15079), .C2(n15063), .A(n15062), .B(n15061), .ZN(
        n15064) );
  OAI21_X1 U18624 ( .B1(n15081), .B2(n15295), .A(n15064), .ZN(P1_U3040) );
  NOR2_X1 U18625 ( .A1(n15073), .A2(n15065), .ZN(n15069) );
  INV_X1 U18626 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15066) );
  OAI22_X1 U18627 ( .A1(n16337), .A2(n15067), .B1(n15066), .B2(n15074), .ZN(
        n15068) );
  AOI211_X1 U18628 ( .C1(n15079), .C2(n15070), .A(n15069), .B(n15068), .ZN(
        n15071) );
  OAI21_X1 U18629 ( .B1(n15081), .B2(n15302), .A(n15071), .ZN(P1_U3038) );
  NOR2_X1 U18630 ( .A1(n15073), .A2(n15072), .ZN(n15077) );
  OAI22_X1 U18631 ( .A1(n16337), .A2(n15075), .B1(n10642), .B2(n15074), .ZN(
        n15076) );
  AOI211_X1 U18632 ( .C1(n15079), .C2(n15078), .A(n15077), .B(n15076), .ZN(
        n15080) );
  OAI21_X1 U18633 ( .B1(n15081), .B2(n15309), .A(n15080), .ZN(P1_U3036) );
  NOR2_X1 U18634 ( .A1(n15082), .A2(n17566), .ZN(n15086) );
  OAI22_X1 U18635 ( .A1(n12303), .A2(n20324), .B1(n17571), .B2(n20386), .ZN(
        n15085) );
  OAI22_X1 U18636 ( .A1(n15083), .A2(n17577), .B1(n17596), .B2(n20379), .ZN(
        n15084) );
  AOI211_X1 U18637 ( .C1(n15086), .C2(n14935), .A(n15085), .B(n15084), .ZN(
        n15087) );
  OAI21_X1 U18638 ( .B1(n15088), .B2(n17572), .A(n15087), .ZN(P2_U3010) );
  INV_X1 U18639 ( .A(n14991), .ZN(n15089) );
  AOI21_X1 U18640 ( .B1(n15091), .B2(n15090), .A(n15089), .ZN(n21363) );
  INV_X1 U18641 ( .A(n21363), .ZN(n15093) );
  OAI222_X1 U18642 ( .A1(n15739), .A2(n15093), .B1(n15733), .B2(n21398), .C1(
        n15732), .C2(n15092), .ZN(P1_U2896) );
  INV_X1 U18643 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15095) );
  INV_X1 U18644 ( .A(n15094), .ZN(n15160) );
  XNOR2_X1 U18645 ( .A(n15161), .B(n15160), .ZN(n17381) );
  OAI222_X1 U18646 ( .A1(n17250), .A2(n21278), .B1(n15095), .B2(n21381), .C1(
        n15641), .C2(n17381), .ZN(P1_U2863) );
  AND2_X1 U18647 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21439), .ZN(n15097) );
  NAND3_X1 U18648 ( .A1(n21438), .A2(n21441), .A3(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n17172) );
  INV_X1 U18649 ( .A(n17172), .ZN(n15096) );
  AOI22_X1 U18650 ( .A1(n10631), .A2(n15097), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15096), .ZN(n15098) );
  AND2_X1 U18651 ( .A1(n21452), .A2(n21254), .ZN(n17163) );
  NAND2_X1 U18652 ( .A1(n17165), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n15102) );
  NAND2_X1 U18653 ( .A1(n15101), .A2(n17163), .ZN(n15152) );
  INV_X1 U18654 ( .A(n15102), .ZN(n15103) );
  NAND2_X1 U18655 ( .A1(n15117), .A2(n15104), .ZN(n21346) );
  NOR2_X2 U18656 ( .A1(n15164), .A2(n17400), .ZN(n21331) );
  NAND2_X1 U18657 ( .A1(n21331), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15112) );
  INV_X1 U18658 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15107) );
  NAND2_X1 U18659 ( .A1(n15430), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15109) );
  NAND2_X1 U18660 ( .A1(n21339), .A2(n15110), .ZN(n15111) );
  OAI211_X1 U18661 ( .C1(n21346), .C2(n13865), .A(n15112), .B(n15111), .ZN(
        n15115) );
  OR2_X1 U18662 ( .A1(n15153), .A2(n15152), .ZN(n15129) );
  INV_X1 U18663 ( .A(n15155), .ZN(n15113) );
  AOI21_X1 U18664 ( .B1(n15129), .B2(n21534), .A(n15113), .ZN(n15114) );
  AOI211_X1 U18665 ( .C1(n21343), .C2(P1_EBX_REG_1__SCAN_IN), .A(n15115), .B(
        n15114), .ZN(n15122) );
  NAND2_X1 U18666 ( .A1(n15117), .A2(n15116), .ZN(n15119) );
  NOR2_X1 U18667 ( .A1(n15430), .A2(n21438), .ZN(n15118) );
  NAND2_X1 U18668 ( .A1(n15119), .A2(n21277), .ZN(n21357) );
  INV_X1 U18669 ( .A(n15120), .ZN(n21378) );
  NAND2_X1 U18670 ( .A1(n21357), .A2(n21378), .ZN(n15121) );
  OAI211_X1 U18671 ( .C1(n21374), .C2(n21296), .A(n15122), .B(n15121), .ZN(
        P1_U2839) );
  XNOR2_X1 U18672 ( .A(n15124), .B(n15123), .ZN(n15147) );
  NAND2_X1 U18673 ( .A1(n21363), .A2(n17298), .ZN(n15128) );
  INV_X1 U18674 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15125) );
  NOR2_X1 U18675 ( .A1(n17352), .A2(n15125), .ZN(n15144) );
  INV_X1 U18676 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21283) );
  NOR2_X1 U18677 ( .A1(n15759), .A2(n21283), .ZN(n15126) );
  AOI211_X1 U18678 ( .C1(n17296), .C2(n21285), .A(n15144), .B(n15126), .ZN(
        n15127) );
  OAI211_X1 U18679 ( .C1(n15147), .C2(n17312), .A(n15128), .B(n15127), .ZN(
        P1_U2991) );
  INV_X1 U18680 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n15135) );
  OAI21_X1 U18681 ( .B1(n21331), .B2(n21339), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15130) );
  OAI21_X1 U18682 ( .B1(n21346), .B2(n10634), .A(n15130), .ZN(n15132) );
  OAI22_X1 U18683 ( .A1(n21425), .A2(n21296), .B1(n21308), .B2(n12671), .ZN(
        n15131) );
  AOI211_X1 U18684 ( .C1(n21357), .C2(n15133), .A(n15132), .B(n15131), .ZN(
        n15134) );
  OAI21_X1 U18685 ( .B1(n21292), .B2(n15135), .A(n15134), .ZN(P1_U2840) );
  AOI221_X1 U18686 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15138), .C2(n15137), .A(
        n15136), .ZN(n15139) );
  AOI21_X1 U18687 ( .B1(n15140), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n15139), .ZN(n15146) );
  INV_X1 U18688 ( .A(n15161), .ZN(n15141) );
  AOI21_X1 U18689 ( .B1(n15143), .B2(n15142), .A(n15141), .ZN(n21362) );
  AOI21_X1 U18690 ( .B1(n21427), .B2(n21362), .A(n15144), .ZN(n15145) );
  OAI211_X1 U18691 ( .C1(n17365), .C2(n15147), .A(n15146), .B(n15145), .ZN(
        P1_U3023) );
  OR2_X1 U18692 ( .A1(n14992), .A2(n15148), .ZN(n15149) );
  NAND2_X1 U18693 ( .A1(n15150), .A2(n15149), .ZN(n17307) );
  AOI22_X1 U18694 ( .A1(n15737), .A2(n15665), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15736), .ZN(n15151) );
  OAI21_X1 U18695 ( .B1(n17307), .B2(n15739), .A(n15151), .ZN(P1_U2894) );
  NAND2_X1 U18696 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .ZN(n15154) );
  NAND2_X1 U18697 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21321), .ZN(n21315) );
  INV_X1 U18698 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21474) );
  NOR2_X1 U18699 ( .A1(n21276), .A2(n21474), .ZN(n15157) );
  NAND2_X1 U18700 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15326) );
  NAND3_X1 U18701 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(n15181), .ZN(n21316) );
  NOR3_X2 U18702 ( .A1(n21468), .A2(n21467), .A3(n21316), .ZN(n21303) );
  NAND3_X1 U18703 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_8__SCAN_IN), 
        .A3(n21303), .ZN(n21271) );
  OAI21_X1 U18704 ( .B1(n15326), .B2(n21271), .A(n21317), .ZN(n15156) );
  INV_X1 U18705 ( .A(n15156), .ZN(n15327) );
  MUX2_X1 U18706 ( .A(n15157), .B(n15327), .S(P1_REIP_REG_10__SCAN_IN), .Z(
        n15158) );
  INV_X1 U18707 ( .A(n15158), .ZN(n15170) );
  OAI21_X1 U18708 ( .B1(n15161), .B2(n15160), .A(n15159), .ZN(n15162) );
  INV_X1 U18709 ( .A(n15162), .ZN(n15163) );
  OR2_X1 U18710 ( .A1(n15163), .A2(n15360), .ZN(n15171) );
  INV_X1 U18711 ( .A(n15171), .ZN(n15389) );
  AOI22_X1 U18712 ( .A1(n21345), .A2(n15389), .B1(n21343), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n15166) );
  NOR2_X1 U18713 ( .A1(n15165), .A2(n15164), .ZN(n21330) );
  OAI211_X1 U18714 ( .C1(n21349), .C2(n15167), .A(n15166), .B(n21273), .ZN(
        n15168) );
  AOI21_X1 U18715 ( .B1(n21339), .B2(n17303), .A(n15168), .ZN(n15169) );
  OAI211_X1 U18716 ( .C1(n21277), .C2(n17307), .A(n15170), .B(n15169), .ZN(
        P1_U2830) );
  INV_X1 U18717 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15172) );
  OAI222_X1 U18718 ( .A1(n17307), .A2(n17250), .B1(n15172), .B2(n21381), .C1(
        n15171), .C2(n15641), .ZN(P1_U2862) );
  NAND2_X1 U18719 ( .A1(n21345), .A2(n15173), .ZN(n15180) );
  NAND2_X1 U18720 ( .A1(n21343), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n15179) );
  INV_X1 U18721 ( .A(n15174), .ZN(n15175) );
  AOI22_X1 U18722 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n21331), .B1(
        n21339), .B2(n15175), .ZN(n15178) );
  INV_X1 U18723 ( .A(n15176), .ZN(n16333) );
  OR2_X1 U18724 ( .A1(n21346), .A2(n16333), .ZN(n15177) );
  NAND4_X1 U18725 ( .A1(n15180), .A2(n15179), .A3(n15178), .A4(n15177), .ZN(
        n15184) );
  INV_X1 U18726 ( .A(n15181), .ZN(n15182) );
  NAND2_X1 U18727 ( .A1(n21317), .A2(n15182), .ZN(n21361) );
  NOR2_X1 U18728 ( .A1(n21361), .A2(n21463), .ZN(n15183) );
  AOI211_X1 U18729 ( .C1(n15185), .C2(n21357), .A(n15184), .B(n15183), .ZN(
        n15186) );
  OAI21_X1 U18730 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n21326), .A(n15186), .ZN(
        P1_U2837) );
  INV_X1 U18731 ( .A(n12236), .ZN(n16929) );
  NAND2_X1 U18732 ( .A1(n9818), .A2(n16964), .ZN(n15192) );
  INV_X1 U18733 ( .A(n15187), .ZN(n15188) );
  OR2_X1 U18734 ( .A1(n15189), .A2(n15188), .ZN(n16926) );
  OAI21_X1 U18735 ( .B1(n15190), .B2(n11600), .A(n16926), .ZN(n15191) );
  OAI211_X1 U18736 ( .C1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n16929), .A(
        n15192), .B(n15191), .ZN(n17695) );
  AOI21_X1 U18737 ( .B1(n15194), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15193), .ZN(n16948) );
  AOI221_X1 U18738 ( .B1(n15196), .B2(n15195), .C1(n15194), .C2(n13684), .A(
        n12040), .ZN(n16947) );
  AOI222_X1 U18739 ( .A1(n17695), .A2(n21082), .B1(n16948), .B2(n16947), .C1(
        n17730), .C2(n21197), .ZN(n15210) );
  NOR2_X1 U18740 ( .A1(n17682), .A2(n21205), .ZN(n17736) );
  INV_X1 U18741 ( .A(n15197), .ZN(n15198) );
  NOR2_X1 U18742 ( .A1(n15199), .A2(n15198), .ZN(n15200) );
  NAND2_X1 U18743 ( .A1(n15201), .A2(n15200), .ZN(n15206) );
  INV_X1 U18744 ( .A(n15202), .ZN(n15204) );
  AND4_X1 U18745 ( .A1(n15206), .A2(n15205), .A3(n15204), .A4(n15203), .ZN(
        n17720) );
  NOR2_X1 U18746 ( .A1(n17720), .A2(n15207), .ZN(n15208) );
  AOI211_X1 U18747 ( .C1(P2_FLUSH_REG_SCAN_IN), .C2(n17736), .A(n17735), .B(
        n15208), .ZN(n16966) );
  NAND2_X1 U18748 ( .A1(n16966), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15209) );
  OAI21_X1 U18749 ( .B1(n15210), .B2(n16966), .A(n15209), .ZN(P2_U3600) );
  NOR2_X1 U18750 ( .A1(n15211), .A2(n15212), .ZN(n15213) );
  OR2_X1 U18751 ( .A1(n9905), .A2(n15213), .ZN(n16470) );
  INV_X1 U18752 ( .A(n16470), .ZN(n15222) );
  NAND2_X1 U18753 ( .A1(n20443), .A2(BUF1_REG_17__SCAN_IN), .ZN(n15220) );
  NAND2_X1 U18754 ( .A1(n20444), .A2(BUF2_REG_17__SCAN_IN), .ZN(n15219) );
  AOI22_X1 U18755 ( .A1(n20442), .A2(n15217), .B1(n20491), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15218) );
  NAND3_X1 U18756 ( .A1(n15220), .A2(n15219), .A3(n15218), .ZN(n15221) );
  AOI21_X1 U18757 ( .B1(n15222), .B2(n20477), .A(n15221), .ZN(n15223) );
  OAI21_X1 U18758 ( .B1(n16832), .B2(n16543), .A(n15223), .ZN(P2_U2902) );
  NAND2_X1 U18759 ( .A1(n15225), .A2(n15224), .ZN(n15226) );
  XNOR2_X1 U18760 ( .A(n15227), .B(n15226), .ZN(n17574) );
  OAI211_X1 U18761 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n17633), .B(n15228), .ZN(n15239) );
  OAI21_X1 U18762 ( .B1(n9931), .B2(n15230), .A(n15229), .ZN(n20482) );
  INV_X1 U18763 ( .A(n20482), .ZN(n15237) );
  NOR2_X1 U18764 ( .A1(n15232), .A2(n15231), .ZN(n15233) );
  OR2_X1 U18765 ( .A1(n15234), .A2(n15233), .ZN(n20367) );
  OAI22_X1 U18766 ( .A1(n17672), .A2(n20367), .B1(n20324), .B2(n15235), .ZN(
        n15236) );
  AOI21_X1 U18767 ( .B1(n15237), .B2(n17637), .A(n15236), .ZN(n15238) );
  OAI211_X1 U18768 ( .C1(n15241), .C2(n15240), .A(n15239), .B(n15238), .ZN(
        n15245) );
  XNOR2_X1 U18769 ( .A(n15243), .B(n15242), .ZN(n17573) );
  NOR2_X1 U18770 ( .A1(n17573), .A2(n17681), .ZN(n15244) );
  AOI211_X1 U18771 ( .C1(n12521), .C2(n17574), .A(n15245), .B(n15244), .ZN(
        n15246) );
  INV_X1 U18772 ( .A(n15246), .ZN(P2_U3041) );
  NAND2_X1 U18773 ( .A1(n17369), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n17382) );
  OAI21_X1 U18774 ( .B1(n15759), .B2(n21275), .A(n17382), .ZN(n15247) );
  AOI21_X1 U18775 ( .B1(n17296), .B2(n21281), .A(n15247), .ZN(n15251) );
  XNOR2_X1 U18776 ( .A(n16288), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15249) );
  XNOR2_X1 U18777 ( .A(n15248), .B(n15249), .ZN(n17385) );
  NAND2_X1 U18778 ( .A1(n17385), .A2(n17267), .ZN(n15250) );
  OAI211_X1 U18779 ( .C1(n21278), .C2(n17306), .A(n15251), .B(n15250), .ZN(
        P1_U2990) );
  NOR3_X1 U18780 ( .A1(n15318), .A2(n15312), .A3(n16334), .ZN(n15254) );
  INV_X1 U18781 ( .A(n15252), .ZN(n15253) );
  NOR2_X1 U18782 ( .A1(n15254), .A2(n15253), .ZN(n15258) );
  NAND2_X1 U18783 ( .A1(n15255), .A2(n13865), .ZN(n15259) );
  OAI22_X1 U18784 ( .A1(n15258), .A2(n15259), .B1(n15256), .B2(n15261), .ZN(
        n15273) );
  NOR2_X1 U18785 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15257), .ZN(
        n15264) );
  INV_X1 U18786 ( .A(n15264), .ZN(n15314) );
  INV_X1 U18787 ( .A(n15258), .ZN(n15260) );
  AOI22_X1 U18788 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15261), .B1(n15260), 
        .B2(n15259), .ZN(n15262) );
  OAI211_X1 U18789 ( .C1(n15264), .C2(n17400), .A(n15263), .B(n15262), .ZN(
        n15310) );
  AOI22_X1 U18790 ( .A1(n15312), .A2(n15265), .B1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n15310), .ZN(n15268) );
  NAND2_X1 U18791 ( .A1(n15318), .A2(n15266), .ZN(n15267) );
  OAI211_X1 U18792 ( .C1(n15269), .C2(n15314), .A(n15268), .B(n15267), .ZN(
        n15270) );
  AOI21_X1 U18793 ( .B1(n15273), .B2(n15271), .A(n15270), .ZN(n15272) );
  INV_X1 U18794 ( .A(n15272), .ZN(P1_U3129) );
  AOI22_X1 U18795 ( .A1(n15312), .A2(n16356), .B1(
        P1_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n15310), .ZN(n15274) );
  OAI21_X1 U18796 ( .B1(n15275), .B2(n15314), .A(n15274), .ZN(n15276) );
  AOI21_X1 U18797 ( .B1(n15318), .B2(n16354), .A(n15276), .ZN(n15277) );
  OAI21_X1 U18798 ( .B1(n15321), .B2(n15278), .A(n15277), .ZN(P1_U3135) );
  AOI22_X1 U18799 ( .A1(n15312), .A2(n16347), .B1(
        P1_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n15310), .ZN(n15279) );
  OAI21_X1 U18800 ( .B1(n15280), .B2(n15314), .A(n15279), .ZN(n15281) );
  AOI21_X1 U18801 ( .B1(n15318), .B2(n16346), .A(n15281), .ZN(n15282) );
  OAI21_X1 U18802 ( .B1(n15321), .B2(n15283), .A(n15282), .ZN(P1_U3133) );
  AOI22_X1 U18803 ( .A1(n15312), .A2(n16339), .B1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n15310), .ZN(n15284) );
  OAI21_X1 U18804 ( .B1(n15285), .B2(n15314), .A(n15284), .ZN(n15286) );
  AOI21_X1 U18805 ( .B1(n15318), .B2(n16338), .A(n15286), .ZN(n15287) );
  OAI21_X1 U18806 ( .B1(n15321), .B2(n15288), .A(n15287), .ZN(P1_U3130) );
  AOI22_X1 U18807 ( .A1(n15312), .A2(n15289), .B1(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n15310), .ZN(n15290) );
  OAI21_X1 U18808 ( .B1(n15291), .B2(n15314), .A(n15290), .ZN(n15292) );
  AOI21_X1 U18809 ( .B1(n15318), .B2(n15293), .A(n15292), .ZN(n15294) );
  OAI21_X1 U18810 ( .B1(n15321), .B2(n15295), .A(n15294), .ZN(P1_U3136) );
  AOI22_X1 U18811 ( .A1(n15312), .A2(n15296), .B1(
        P1_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n15310), .ZN(n15297) );
  OAI21_X1 U18812 ( .B1(n15298), .B2(n15314), .A(n15297), .ZN(n15299) );
  AOI21_X1 U18813 ( .B1(n15318), .B2(n15300), .A(n15299), .ZN(n15301) );
  OAI21_X1 U18814 ( .B1(n15321), .B2(n15302), .A(n15301), .ZN(P1_U3134) );
  AOI22_X1 U18815 ( .A1(n15312), .A2(n15303), .B1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n15310), .ZN(n15304) );
  OAI21_X1 U18816 ( .B1(n15305), .B2(n15314), .A(n15304), .ZN(n15306) );
  AOI21_X1 U18817 ( .B1(n15318), .B2(n15307), .A(n15306), .ZN(n15308) );
  OAI21_X1 U18818 ( .B1(n15321), .B2(n15309), .A(n15308), .ZN(P1_U3132) );
  AOI22_X1 U18819 ( .A1(n15312), .A2(n15311), .B1(
        P1_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n15310), .ZN(n15313) );
  OAI21_X1 U18820 ( .B1(n15315), .B2(n15314), .A(n15313), .ZN(n15316) );
  AOI21_X1 U18821 ( .B1(n15318), .B2(n15317), .A(n15316), .ZN(n15319) );
  OAI21_X1 U18822 ( .B1(n15321), .B2(n15320), .A(n15319), .ZN(P1_U3131) );
  OAI21_X1 U18823 ( .B1(n15322), .B2(n15324), .A(n15323), .ZN(n16176) );
  INV_X1 U18824 ( .A(n16172), .ZN(n15331) );
  XNOR2_X1 U18825 ( .A(n15360), .B(n15359), .ZN(n15334) );
  INV_X1 U18826 ( .A(n15334), .ZN(n17374) );
  AOI22_X1 U18827 ( .A1(n21345), .A2(n17374), .B1(n21343), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15325) );
  OAI211_X1 U18828 ( .C1(n21349), .C2(n10782), .A(n15325), .B(n21273), .ZN(
        n15330) );
  NOR2_X1 U18829 ( .A1(n21276), .A2(n15326), .ZN(n15328) );
  MUX2_X1 U18830 ( .A(n15328), .B(n15327), .S(P1_REIP_REG_11__SCAN_IN), .Z(
        n15329) );
  AOI211_X1 U18831 ( .C1(n21339), .C2(n15331), .A(n15330), .B(n15329), .ZN(
        n15332) );
  OAI21_X1 U18832 ( .B1(n21277), .B2(n16176), .A(n15332), .ZN(P1_U2829) );
  OAI222_X1 U18833 ( .A1(n15739), .A2(n16176), .B1(n15733), .B2(n21391), .C1(
        n15732), .C2(n15333), .ZN(P1_U2893) );
  INV_X1 U18834 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15890) );
  OAI222_X1 U18835 ( .A1(n17250), .A2(n16176), .B1(n21381), .B2(n15890), .C1(
        n15641), .C2(n15334), .ZN(P1_U2861) );
  NAND2_X1 U18836 ( .A1(n15335), .A2(n15336), .ZN(n15583) );
  INV_X1 U18837 ( .A(n15583), .ZN(n15559) );
  AOI21_X1 U18838 ( .B1(n15335), .B2(n15735), .A(n15337), .ZN(n15338) );
  NOR2_X1 U18839 ( .A1(n15559), .A2(n15338), .ZN(n17293) );
  INV_X1 U18840 ( .A(n17293), .ZN(n15734) );
  OR2_X1 U18841 ( .A1(n15362), .A2(n15339), .ZN(n15340) );
  NAND2_X1 U18842 ( .A1(n15589), .A2(n15340), .ZN(n17363) );
  INV_X1 U18843 ( .A(n17363), .ZN(n15341) );
  AOI22_X1 U18844 ( .A1(n21376), .A2(n15341), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n15643), .ZN(n15342) );
  OAI21_X1 U18845 ( .B1(n15734), .B2(n17250), .A(n15342), .ZN(P1_U2859) );
  OAI21_X1 U18846 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n16288), .ZN(n15344) );
  OAI21_X1 U18847 ( .B1(n15343), .B2(n15345), .A(n15344), .ZN(n15348) );
  INV_X1 U18848 ( .A(n17289), .ZN(n15346) );
  OAI21_X1 U18849 ( .B1(n15356), .B2(n10274), .A(n15346), .ZN(n15347) );
  NOR2_X1 U18850 ( .A1(n15348), .A2(n15347), .ZN(n17288) );
  AOI21_X1 U18851 ( .B1(n15348), .B2(n15347), .A(n17288), .ZN(n17302) );
  NAND3_X1 U18852 ( .A1(n15353), .A2(n15356), .A3(n17354), .ZN(n15366) );
  OAI21_X1 U18853 ( .B1(n15350), .B2(n15355), .A(n15349), .ZN(n15352) );
  OAI211_X1 U18854 ( .C1(n16220), .C2(n15353), .A(n15352), .B(n15351), .ZN(
        n15354) );
  INV_X1 U18855 ( .A(n15354), .ZN(n17380) );
  NOR2_X1 U18856 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15355), .ZN(
        n17376) );
  NAND2_X1 U18857 ( .A1(n17376), .A2(n17343), .ZN(n15357) );
  AOI21_X1 U18858 ( .B1(n17380), .B2(n15357), .A(n15356), .ZN(n15364) );
  AOI21_X1 U18859 ( .B1(n15360), .B2(n15359), .A(n15358), .ZN(n15361) );
  OR2_X1 U18860 ( .A1(n15362), .A2(n15361), .ZN(n17244) );
  INV_X1 U18861 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21479) );
  OAI22_X1 U18862 ( .A1(n17364), .A2(n17244), .B1(n21479), .B2(n17352), .ZN(
        n15363) );
  NOR2_X1 U18863 ( .A1(n15364), .A2(n15363), .ZN(n15365) );
  OAI211_X1 U18864 ( .C1(n17302), .C2(n17365), .A(n15366), .B(n15365), .ZN(
        P1_U3019) );
  OAI21_X1 U18865 ( .B1(n15369), .B2(n15368), .A(n15634), .ZN(n17230) );
  NOR2_X2 U18866 ( .A1(n15370), .A2(n15371), .ZN(n15723) );
  INV_X1 U18867 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20550) );
  INV_X1 U18868 ( .A(n15370), .ZN(n15372) );
  AND2_X1 U18869 ( .A1(n15374), .A2(n15373), .ZN(n15375) );
  AOI22_X1 U18870 ( .A1(n15719), .A2(n15376), .B1(n15736), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n15377) );
  OAI21_X1 U18871 ( .B1(n20550), .B2(n15721), .A(n15377), .ZN(n15378) );
  AOI21_X1 U18872 ( .B1(n15723), .B2(DATAI_17_), .A(n15378), .ZN(n15379) );
  OAI21_X1 U18873 ( .B1(n17230), .B2(n15739), .A(n15379), .ZN(P1_U2887) );
  XNOR2_X1 U18874 ( .A(n16167), .B(n11272), .ZN(n15381) );
  INV_X1 U18875 ( .A(n15343), .ZN(n16156) );
  NOR2_X1 U18876 ( .A1(n16156), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15380) );
  MUX2_X1 U18877 ( .A(n15381), .B(n15380), .S(n10274), .Z(n15382) );
  NOR3_X1 U18878 ( .A1(n15343), .A2(n16288), .A3(n11272), .ZN(n16169) );
  OR2_X1 U18879 ( .A1(n15382), .A2(n16169), .ZN(n17311) );
  NOR2_X1 U18880 ( .A1(n15384), .A2(n15383), .ZN(n15385) );
  AOI21_X1 U18881 ( .B1(n15385), .B2(n15386), .A(n16263), .ZN(n17384) );
  INV_X1 U18882 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15387) );
  NAND2_X1 U18883 ( .A1(n15386), .A2(n17375), .ZN(n17388) );
  AOI221_X1 U18884 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n15387), .C2(n11272), .A(
        n17388), .ZN(n15388) );
  AOI21_X1 U18885 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17384), .A(
        n15388), .ZN(n15391) );
  AOI22_X1 U18886 ( .A1(n21427), .A2(n15389), .B1(n17369), .B2(
        P1_REIP_REG_10__SCAN_IN), .ZN(n15390) );
  OAI211_X1 U18887 ( .C1(n17311), .C2(n17365), .A(n15391), .B(n15390), .ZN(
        P1_U3021) );
  NAND2_X1 U18888 ( .A1(n15404), .A2(n19987), .ZN(n15392) );
  NAND2_X1 U18889 ( .A1(n15393), .A2(n15392), .ZN(n19986) );
  NOR2_X1 U18890 ( .A1(n20154), .A2(n19986), .ZN(n15403) );
  NAND2_X1 U18891 ( .A1(n19981), .A2(n20206), .ZN(n15400) );
  NOR2_X1 U18892 ( .A1(n19555), .A2(n18794), .ZN(n18795) );
  INV_X1 U18893 ( .A(n17086), .ZN(n19978) );
  OAI211_X1 U18894 ( .C1(n15398), .C2(n15397), .A(n15396), .B(n15395), .ZN(
        n17088) );
  AOI21_X1 U18895 ( .B1(n19978), .B2(n16987), .A(n17088), .ZN(n15399) );
  OAI211_X1 U18896 ( .C1(n15400), .C2(n18730), .A(n15399), .B(n17191), .ZN(
        n20013) );
  INV_X1 U18897 ( .A(n20013), .ZN(n20024) );
  NAND2_X1 U18898 ( .A1(n15401), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19551) );
  INV_X1 U18899 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19540) );
  NAND3_X1 U18900 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n20151)
         );
  OR2_X1 U18901 ( .A1(n19540), .A2(n20151), .ZN(n15402) );
  OAI211_X1 U18902 ( .C1(n20202), .C2(n20024), .A(n19551), .B(n15402), .ZN(
        n20182) );
  MUX2_X1 U18903 ( .A(n15403), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n20185), .Z(P3_U3284) );
  NAND3_X1 U18904 ( .A1(n9850), .A2(n15404), .A3(n19987), .ZN(n19539) );
  NOR2_X1 U18905 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n19539), .ZN(n15405) );
  OAI21_X1 U18906 ( .B1(n15405), .B2(n20151), .A(n19651), .ZN(n19546) );
  INV_X1 U18907 ( .A(n19546), .ZN(n15406) );
  NAND2_X1 U18908 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n19121) );
  AOI22_X1 U18909 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n20201), .B2(n19121), .ZN(n17078) );
  NOR2_X1 U18910 ( .A1(n15406), .A2(n17078), .ZN(n15408) );
  NOR2_X1 U18911 ( .A1(n20153), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19588) );
  OR2_X1 U18912 ( .A1(n19588), .A2(n15406), .ZN(n17076) );
  OR2_X1 U18913 ( .A1(n19608), .A2(n17076), .ZN(n15407) );
  MUX2_X1 U18914 ( .A(n15408), .B(n15407), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  XOR2_X1 U18915 ( .A(n13945), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n15411)
         );
  INV_X1 U18916 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n15409) );
  MUX2_X1 U18917 ( .A(n15409), .B(n20367), .S(n20437), .Z(n15410) );
  OAI21_X1 U18918 ( .B1(n15411), .B2(n20428), .A(n15410), .ZN(P2_U2882) );
  AOI22_X1 U18919 ( .A1(n20444), .A2(BUF2_REG_30__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n15414) );
  AOI22_X1 U18920 ( .A1(n20442), .A2(n15412), .B1(n20491), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n15413) );
  OAI211_X1 U18921 ( .C1(n15415), .C2(n16543), .A(n15414), .B(n15413), .ZN(
        n15416) );
  AOI21_X1 U18922 ( .B1(n15417), .B2(n20477), .A(n15416), .ZN(n15418) );
  INV_X1 U18923 ( .A(n15418), .ZN(P2_U2889) );
  INV_X1 U18924 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17802) );
  AOI22_X1 U18925 ( .A1(n10753), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n15421), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15422) );
  INV_X1 U18926 ( .A(n15422), .ZN(n15423) );
  NAND3_X1 U18927 ( .A1(n15434), .A2(n15425), .A3(n15733), .ZN(n15427) );
  AOI22_X1 U18928 ( .A1(n15723), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15736), .ZN(n15426) );
  OAI211_X1 U18929 ( .C1(n15721), .C2(n17802), .A(n15427), .B(n15426), .ZN(
        P1_U2873) );
  AOI21_X1 U18930 ( .B1(n14161), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15428), .ZN(n15429) );
  OAI21_X1 U18931 ( .B1(n17305), .B2(n15430), .A(n15429), .ZN(n15431) );
  AOI21_X1 U18932 ( .B1(n15434), .B2(n17298), .A(n15431), .ZN(n15432) );
  OAI21_X1 U18933 ( .B1(n15433), .B2(n17312), .A(n15432), .ZN(P1_U2968) );
  INV_X1 U18934 ( .A(n15434), .ZN(n15447) );
  INV_X1 U18935 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21486) );
  NAND2_X1 U18936 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15443) );
  NAND3_X1 U18937 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .ZN(n15442) );
  NOR3_X1 U18938 ( .A1(n21479), .A2(n15442), .A3(n21271), .ZN(n17240) );
  NAND3_X1 U18939 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n17240), .ZN(n15561) );
  NOR3_X1 U18940 ( .A1(n21486), .A2(n15443), .A3(n15561), .ZN(n17210) );
  NAND4_X1 U18941 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .A4(n17210), .ZN(n15554) );
  NAND2_X1 U18942 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n17195) );
  INV_X1 U18943 ( .A(n17195), .ZN(n15435) );
  NAND2_X1 U18944 ( .A1(n15435), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15436) );
  NOR2_X1 U18945 ( .A1(n15554), .A2(n15436), .ZN(n15517) );
  AND3_X1 U18946 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_24__SCAN_IN), .ZN(n15437) );
  NAND2_X1 U18947 ( .A1(n15517), .A2(n15437), .ZN(n15484) );
  NAND2_X1 U18948 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n15438) );
  NAND2_X1 U18949 ( .A1(n15439), .A2(n21317), .ZN(n15463) );
  INV_X1 U18950 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n15445) );
  INV_X1 U18951 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21509) );
  OAI21_X1 U18952 ( .B1(n15445), .B2(n21509), .A(n21317), .ZN(n15440) );
  NAND2_X1 U18953 ( .A1(n15463), .A2(n15440), .ZN(n15457) );
  AOI22_X1 U18954 ( .A1(n21343), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n21331), .ZN(n15441) );
  INV_X1 U18955 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21481) );
  NAND2_X1 U18956 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n17216) );
  NAND2_X1 U18957 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n15444) );
  NOR3_X1 U18958 ( .A1(n15456), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n15445), 
        .ZN(n15446) );
  INV_X1 U18959 ( .A(n15474), .ZN(n15448) );
  OAI22_X1 U18960 ( .A1(n15450), .A2(n12759), .B1(n15449), .B2(n15448), .ZN(
        n15451) );
  XOR2_X1 U18961 ( .A(n15452), .B(n15451), .Z(n15599) );
  INV_X1 U18962 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15600) );
  AOI22_X1 U18963 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21331), .B1(
        n21339), .B2(n15453), .ZN(n15454) );
  OAI21_X1 U18964 ( .B1(n21308), .B2(n15600), .A(n15454), .ZN(n15455) );
  AOI21_X1 U18965 ( .B1(n15599), .B2(n21345), .A(n15455), .ZN(n15460) );
  INV_X1 U18966 ( .A(n15456), .ZN(n15458) );
  OAI21_X1 U18967 ( .B1(n15458), .B2(P1_REIP_REG_30__SCAN_IN), .A(n15457), 
        .ZN(n15459) );
  OAI211_X1 U18968 ( .C1(n15649), .C2(n21277), .A(n15460), .B(n15459), .ZN(
        P1_U2810) );
  AOI21_X1 U18969 ( .B1(n15461), .B2(n15462), .A(n15420), .ZN(n15748) );
  INV_X1 U18970 ( .A(n15748), .ZN(n15655) );
  INV_X1 U18971 ( .A(n15463), .ZN(n15479) );
  OAI21_X1 U18972 ( .B1(n15474), .B2(n15465), .A(n15464), .ZN(n17314) );
  OAI22_X1 U18973 ( .A1(n11131), .A2(n21349), .B1(n21348), .B2(n15746), .ZN(
        n15466) );
  AOI21_X1 U18974 ( .B1(n21343), .B2(P1_EBX_REG_29__SCAN_IN), .A(n15466), .ZN(
        n15467) );
  OAI21_X1 U18975 ( .B1(n17314), .B2(n21296), .A(n15467), .ZN(n15468) );
  AOI21_X1 U18976 ( .B1(n15479), .B2(P1_REIP_REG_29__SCAN_IN), .A(n15468), 
        .ZN(n15470) );
  NAND3_X1 U18977 ( .A1(n9858), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n21509), 
        .ZN(n15469) );
  OAI211_X1 U18978 ( .C1(n15655), .C2(n21277), .A(n15470), .B(n15469), .ZN(
        P1_U2811) );
  OAI21_X1 U18979 ( .B1(n15471), .B2(n15472), .A(n15461), .ZN(n15763) );
  AND2_X1 U18980 ( .A1(n15487), .A2(n15473), .ZN(n15475) );
  OR2_X1 U18981 ( .A1(n15475), .A2(n15474), .ZN(n17323) );
  AOI22_X1 U18982 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n21331), .B1(
        n21339), .B2(n15761), .ZN(n15477) );
  NAND2_X1 U18983 ( .A1(n21343), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n15476) );
  OAI211_X1 U18984 ( .C1(n17323), .C2(n21296), .A(n15477), .B(n15476), .ZN(
        n15478) );
  AOI21_X1 U18985 ( .B1(n15479), .B2(P1_REIP_REG_28__SCAN_IN), .A(n15478), 
        .ZN(n15481) );
  INV_X1 U18986 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21505) );
  NAND2_X1 U18987 ( .A1(n9858), .A2(n21505), .ZN(n15480) );
  OAI211_X1 U18988 ( .C1(n15763), .C2(n21277), .A(n15481), .B(n15480), .ZN(
        P1_U2812) );
  INV_X1 U18989 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21503) );
  NAND2_X1 U18990 ( .A1(n21503), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15494) );
  INV_X1 U18991 ( .A(n15482), .ZN(n15496) );
  AOI21_X1 U18992 ( .B1(n15483), .B2(n15496), .A(n15471), .ZN(n15770) );
  NAND2_X1 U18993 ( .A1(n15770), .A2(n21312), .ZN(n15493) );
  AND2_X1 U18994 ( .A1(n15484), .A2(n21317), .ZN(n15503) );
  NAND2_X1 U18995 ( .A1(n9851), .A2(n15485), .ZN(n15486) );
  NAND2_X1 U18996 ( .A1(n15487), .A2(n15486), .ZN(n16188) );
  INV_X1 U18997 ( .A(n15768), .ZN(n15488) );
  AOI22_X1 U18998 ( .A1(n15488), .A2(n21339), .B1(n21331), .B2(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15490) );
  NAND2_X1 U18999 ( .A1(n21343), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n15489) );
  OAI211_X1 U19000 ( .C1(n16188), .C2(n21296), .A(n15490), .B(n15489), .ZN(
        n15491) );
  AOI21_X1 U19001 ( .B1(n15503), .B2(P1_REIP_REG_27__SCAN_IN), .A(n15491), 
        .ZN(n15492) );
  OAI211_X1 U19002 ( .C1(n15506), .C2(n15494), .A(n15493), .B(n15492), .ZN(
        P1_U2813) );
  AOI21_X1 U19003 ( .B1(n15497), .B2(n15507), .A(n15482), .ZN(n16106) );
  NAND2_X1 U19004 ( .A1(n16106), .A2(n21312), .ZN(n15505) );
  NAND2_X1 U19005 ( .A1(n9910), .A2(n15498), .ZN(n15499) );
  NAND2_X1 U19006 ( .A1(n9851), .A2(n15499), .ZN(n17332) );
  AOI22_X1 U19007 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n21331), .B1(
        n21339), .B2(n16102), .ZN(n15501) );
  NAND2_X1 U19008 ( .A1(n21343), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n15500) );
  OAI211_X1 U19009 ( .C1(n17332), .C2(n21296), .A(n15501), .B(n15500), .ZN(
        n15502) );
  AOI21_X1 U19010 ( .B1(n15503), .B2(P1_REIP_REG_26__SCAN_IN), .A(n15502), 
        .ZN(n15504) );
  OAI211_X1 U19011 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(n15506), .A(n15505), 
        .B(n15504), .ZN(P1_U2814) );
  OAI21_X1 U19012 ( .B1(n15509), .B2(n15508), .A(n15507), .ZN(n16115) );
  OR2_X1 U19013 ( .A1(n15522), .A2(n15510), .ZN(n15511) );
  NAND2_X1 U19014 ( .A1(n9910), .A2(n15511), .ZN(n15604) );
  INV_X1 U19015 ( .A(n15604), .ZN(n16199) );
  INV_X1 U19016 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15605) );
  INV_X1 U19017 ( .A(n16117), .ZN(n15512) );
  AOI22_X1 U19018 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n21331), .B1(
        n21339), .B2(n15512), .ZN(n15513) );
  OAI21_X1 U19019 ( .B1(n21308), .B2(n15605), .A(n15513), .ZN(n15515) );
  INV_X1 U19020 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21497) );
  NOR3_X1 U19021 ( .A1(n15516), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n21497), 
        .ZN(n15514) );
  AOI211_X1 U19022 ( .C1(n16199), .C2(n21345), .A(n15515), .B(n15514), .ZN(
        n15519) );
  NOR2_X1 U19023 ( .A1(n15516), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15529) );
  OAI21_X1 U19024 ( .B1(n15529), .B2(n10338), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15518) );
  OAI211_X1 U19025 ( .C1(n16115), .C2(n21277), .A(n15519), .B(n15518), .ZN(
        P1_U2815) );
  XNOR2_X1 U19026 ( .A(n10278), .B(n15521), .ZN(n16125) );
  INV_X1 U19027 ( .A(n15522), .ZN(n15523) );
  OAI21_X1 U19028 ( .B1(n15524), .B2(n15537), .A(n15523), .ZN(n17346) );
  INV_X1 U19029 ( .A(n15525), .ZN(n16127) );
  OAI22_X1 U19030 ( .A1(n15526), .A2(n21349), .B1(n21348), .B2(n16127), .ZN(
        n15527) );
  AOI21_X1 U19031 ( .B1(n21343), .B2(P1_EBX_REG_24__SCAN_IN), .A(n15527), .ZN(
        n15528) );
  OAI21_X1 U19032 ( .B1(n17346), .B2(n21296), .A(n15528), .ZN(n15530) );
  AOI211_X1 U19033 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n10338), .A(n15530), 
        .B(n15529), .ZN(n15531) );
  OAI21_X1 U19034 ( .B1(n16125), .B2(n21277), .A(n15531), .ZN(P1_U2816) );
  AOI21_X1 U19035 ( .B1(n15533), .B2(n15532), .A(n15520), .ZN(n16135) );
  INV_X1 U19036 ( .A(n16135), .ZN(n15685) );
  INV_X1 U19037 ( .A(n15534), .ZN(n16133) );
  OAI22_X1 U19038 ( .A1(n15535), .A2(n21349), .B1(n21348), .B2(n16133), .ZN(
        n15540) );
  AND2_X1 U19039 ( .A1(n15612), .A2(n15536), .ZN(n15538) );
  OR2_X1 U19040 ( .A1(n15538), .A2(n15537), .ZN(n15607) );
  NOR2_X1 U19041 ( .A1(n15607), .A2(n21296), .ZN(n15539) );
  AOI211_X1 U19042 ( .C1(n21343), .C2(P1_EBX_REG_23__SCAN_IN), .A(n15540), .B(
        n15539), .ZN(n15543) );
  OAI21_X1 U19043 ( .B1(n15541), .B2(P1_REIP_REG_23__SCAN_IN), .A(n10338), 
        .ZN(n15542) );
  OAI211_X1 U19044 ( .C1(n15685), .C2(n21277), .A(n15543), .B(n15542), .ZN(
        P1_U2817) );
  INV_X1 U19045 ( .A(n15544), .ZN(n15548) );
  INV_X1 U19046 ( .A(n15545), .ZN(n15547) );
  AOI21_X1 U19047 ( .B1(n15548), .B2(n15547), .A(n15546), .ZN(n16146) );
  INV_X1 U19048 ( .A(n16146), .ZN(n15701) );
  NOR2_X1 U19049 ( .A1(n15630), .A2(n15549), .ZN(n15550) );
  OR2_X1 U19050 ( .A1(n15618), .A2(n15550), .ZN(n16245) );
  INV_X1 U19051 ( .A(n16245), .ZN(n15553) );
  AOI22_X1 U19052 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n21331), .B1(
        n21339), .B2(n16141), .ZN(n15551) );
  OAI21_X1 U19053 ( .B1(n21308), .B2(n15623), .A(n15551), .ZN(n15552) );
  AOI21_X1 U19054 ( .B1(n21345), .B2(n15553), .A(n15552), .ZN(n15557) );
  AND2_X1 U19055 ( .A1(n21317), .A2(n15554), .ZN(n17202) );
  OAI21_X1 U19056 ( .B1(n15555), .B2(P1_REIP_REG_20__SCAN_IN), .A(n17202), 
        .ZN(n15556) );
  OAI211_X1 U19057 ( .C1(n15701), .C2(n21277), .A(n15557), .B(n15556), .ZN(
        P1_U2820) );
  NAND2_X1 U19058 ( .A1(n15559), .A2(n15558), .ZN(n15571) );
  XOR2_X1 U19059 ( .A(n15560), .B(n15571), .Z(n17279) );
  AND2_X1 U19060 ( .A1(n21317), .A2(n15561), .ZN(n15585) );
  NOR2_X1 U19061 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15566), .ZN(n15579) );
  OAI21_X1 U19062 ( .B1(n15585), .B2(n15579), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15570) );
  OAI21_X1 U19063 ( .B1(n9902), .B2(n15562), .A(n16278), .ZN(n16295) );
  INV_X1 U19064 ( .A(n16295), .ZN(n15563) );
  AOI22_X1 U19065 ( .A1(n21345), .A2(n15563), .B1(n21343), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n15564) );
  OAI211_X1 U19066 ( .C1(n21349), .C2(n15565), .A(n15564), .B(n21273), .ZN(
        n15568) );
  INV_X1 U19067 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21484) );
  NOR3_X1 U19068 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n15566), .A3(n21484), 
        .ZN(n15567) );
  AOI211_X1 U19069 ( .C1(n21339), .C2(n17278), .A(n15568), .B(n15567), .ZN(
        n15569) );
  OAI211_X1 U19070 ( .C1(n15725), .C2(n21277), .A(n15570), .B(n15569), .ZN(
        P1_U2824) );
  OR2_X1 U19071 ( .A1(n15583), .A2(n15584), .ZN(n15581) );
  INV_X1 U19072 ( .A(n15571), .ZN(n15572) );
  AOI21_X1 U19073 ( .B1(n15573), .B2(n15581), .A(n15572), .ZN(n17284) );
  INV_X1 U19074 ( .A(n17284), .ZN(n15728) );
  AND2_X1 U19075 ( .A1(n15587), .A2(n15574), .ZN(n15575) );
  OR2_X1 U19076 ( .A1(n15575), .A2(n9902), .ZN(n16303) );
  AOI21_X1 U19077 ( .B1(n21331), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n21330), .ZN(n15577) );
  AOI22_X1 U19078 ( .A1(n21343), .A2(P1_EBX_REG_15__SCAN_IN), .B1(n21339), 
        .B2(n17283), .ZN(n15576) );
  OAI211_X1 U19079 ( .C1(n21296), .C2(n16303), .A(n15577), .B(n15576), .ZN(
        n15578) );
  AOI211_X1 U19080 ( .C1(n15585), .C2(P1_REIP_REG_15__SCAN_IN), .A(n15579), 
        .B(n15578), .ZN(n15580) );
  OAI21_X1 U19081 ( .B1(n15728), .B2(n21277), .A(n15580), .ZN(P1_U2825) );
  INV_X1 U19082 ( .A(n15581), .ZN(n15582) );
  AOI21_X1 U19083 ( .B1(n15584), .B2(n15583), .A(n15582), .ZN(n16165) );
  INV_X1 U19084 ( .A(n16165), .ZN(n15730) );
  OAI21_X1 U19085 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n15586), .A(n15585), 
        .ZN(n15596) );
  INV_X1 U19086 ( .A(n16163), .ZN(n15594) );
  INV_X1 U19087 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15592) );
  INV_X1 U19088 ( .A(n15587), .ZN(n15588) );
  AOI21_X1 U19089 ( .B1(n15590), .B2(n15589), .A(n15588), .ZN(n17357) );
  AOI22_X1 U19090 ( .A1(n21345), .A2(n17357), .B1(n21343), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n15591) );
  OAI211_X1 U19091 ( .C1(n21349), .C2(n15592), .A(n15591), .B(n21273), .ZN(
        n15593) );
  AOI21_X1 U19092 ( .B1(n21339), .B2(n15594), .A(n15593), .ZN(n15595) );
  OAI211_X1 U19093 ( .C1(n15730), .C2(n21277), .A(n15596), .B(n15595), .ZN(
        P1_U2826) );
  INV_X1 U19094 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15597) );
  OAI22_X1 U19095 ( .A1(n15598), .A2(n15641), .B1(n21381), .B2(n15597), .ZN(
        P1_U2841) );
  INV_X1 U19096 ( .A(n15599), .ZN(n16181) );
  OAI222_X1 U19097 ( .A1(n15641), .A2(n16181), .B1(n15600), .B2(n21381), .C1(
        n15649), .C2(n17250), .ZN(P1_U2842) );
  OAI222_X1 U19098 ( .A1(n15655), .A2(n17250), .B1(n15601), .B2(n21381), .C1(
        n17314), .C2(n15641), .ZN(P1_U2843) );
  INV_X1 U19099 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15602) );
  OAI222_X1 U19100 ( .A1(n17323), .A2(n15641), .B1(n15602), .B2(n21381), .C1(
        n15763), .C2(n17250), .ZN(P1_U2844) );
  INV_X1 U19101 ( .A(n15770), .ZN(n15664) );
  INV_X1 U19102 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15603) );
  OAI222_X1 U19103 ( .A1(n15664), .A2(n17250), .B1(n15603), .B2(n21381), .C1(
        n16188), .C2(n15641), .ZN(P1_U2845) );
  INV_X1 U19104 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15953) );
  INV_X1 U19105 ( .A(n16106), .ZN(n15670) );
  OAI222_X1 U19106 ( .A1(n17332), .A2(n15641), .B1(n15953), .B2(n21381), .C1(
        n15670), .C2(n17250), .ZN(P1_U2846) );
  OAI222_X1 U19107 ( .A1(n16115), .A2(n17250), .B1(n15605), .B2(n21381), .C1(
        n15604), .C2(n15641), .ZN(P1_U2847) );
  INV_X1 U19108 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15606) );
  OAI222_X1 U19109 ( .A1(n16125), .A2(n17250), .B1(n15606), .B2(n21381), .C1(
        n17346), .C2(n15641), .ZN(P1_U2848) );
  INV_X1 U19110 ( .A(n15607), .ZN(n16203) );
  AOI22_X1 U19111 ( .A1(n16203), .A2(n21376), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n15643), .ZN(n15608) );
  OAI21_X1 U19112 ( .B1(n15685), .B2(n17250), .A(n15608), .ZN(P1_U2849) );
  XOR2_X1 U19113 ( .A(n15611), .B(n15610), .Z(n17258) );
  INV_X1 U19114 ( .A(n17258), .ZN(n15689) );
  INV_X1 U19115 ( .A(n15612), .ZN(n15613) );
  AOI21_X1 U19116 ( .B1(n15614), .B2(n15620), .A(n15613), .ZN(n17194) );
  AOI22_X1 U19117 ( .A1(n17194), .A2(n21376), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n15643), .ZN(n15615) );
  OAI21_X1 U19118 ( .B1(n15689), .B2(n17250), .A(n15615), .ZN(P1_U2850) );
  OAI21_X1 U19119 ( .B1(n15546), .B2(n15616), .A(n15610), .ZN(n17203) );
  OR2_X1 U19120 ( .A1(n15618), .A2(n15617), .ZN(n15619) );
  NAND2_X1 U19121 ( .A1(n15620), .A2(n15619), .ZN(n17204) );
  INV_X1 U19122 ( .A(n17204), .ZN(n15621) );
  AOI22_X1 U19123 ( .A1(n15621), .A2(n21376), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n15643), .ZN(n15622) );
  OAI21_X1 U19124 ( .B1(n17203), .B2(n17250), .A(n15622), .ZN(P1_U2851) );
  OAI22_X1 U19125 ( .A1(n16245), .A2(n15641), .B1(n15623), .B2(n21381), .ZN(
        n15624) );
  INV_X1 U19126 ( .A(n15624), .ZN(n15625) );
  OAI21_X1 U19127 ( .B1(n15701), .B2(n17250), .A(n15625), .ZN(P1_U2852) );
  AND2_X1 U19128 ( .A1(n15627), .A2(n15626), .ZN(n15628) );
  OR2_X1 U19129 ( .A1(n15628), .A2(n15544), .ZN(n17215) );
  AND2_X1 U19130 ( .A1(n15637), .A2(n15629), .ZN(n15631) );
  OR2_X1 U19131 ( .A1(n15631), .A2(n15630), .ZN(n17220) );
  OAI22_X1 U19132 ( .A1(n17220), .A2(n15641), .B1(n17212), .B2(n21381), .ZN(
        n15632) );
  INV_X1 U19133 ( .A(n15632), .ZN(n15633) );
  OAI21_X1 U19134 ( .B1(n17215), .B2(n17250), .A(n15633), .ZN(P1_U2853) );
  XOR2_X1 U19135 ( .A(n15635), .B(n15634), .Z(n17225) );
  INV_X1 U19136 ( .A(n17225), .ZN(n15717) );
  OAI21_X1 U19137 ( .B1(n16278), .B2(n16279), .A(n15636), .ZN(n15638) );
  AND2_X1 U19138 ( .A1(n15638), .A2(n15637), .ZN(n17224) );
  AOI22_X1 U19139 ( .A1(n17224), .A2(n21376), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n15643), .ZN(n15639) );
  OAI21_X1 U19140 ( .B1(n15717), .B2(n17250), .A(n15639), .ZN(P1_U2854) );
  OAI222_X1 U19141 ( .A1(n15725), .A2(n17250), .B1(n15640), .B2(n21381), .C1(
        n16295), .C2(n15641), .ZN(P1_U2856) );
  INV_X1 U19142 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15642) );
  OAI222_X1 U19143 ( .A1(n15728), .A2(n17250), .B1(n21381), .B2(n15642), .C1(
        n16303), .C2(n15641), .ZN(P1_U2857) );
  AOI22_X1 U19144 ( .A1(n21376), .A2(n17357), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n15643), .ZN(n15644) );
  OAI21_X1 U19145 ( .B1(n15730), .B2(n17250), .A(n15644), .ZN(P1_U2858) );
  INV_X1 U19146 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n15646) );
  AOI22_X1 U19147 ( .A1(n15719), .A2(n21421), .B1(n15736), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n15645) );
  OAI21_X1 U19148 ( .B1(n15646), .B2(n15721), .A(n15645), .ZN(n15647) );
  AOI21_X1 U19149 ( .B1(n15723), .B2(DATAI_30_), .A(n15647), .ZN(n15648) );
  OAI21_X1 U19150 ( .B1(n15649), .B2(n15739), .A(n15648), .ZN(P1_U2874) );
  INV_X1 U19151 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n15652) );
  AOI22_X1 U19152 ( .A1(n15719), .A2(n15650), .B1(n15736), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n15651) );
  OAI21_X1 U19153 ( .B1(n15652), .B2(n15721), .A(n15651), .ZN(n15653) );
  AOI21_X1 U19154 ( .B1(n15723), .B2(DATAI_29_), .A(n15653), .ZN(n15654) );
  OAI21_X1 U19155 ( .B1(n15655), .B2(n15739), .A(n15654), .ZN(P1_U2875) );
  INV_X1 U19156 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U19157 ( .A1(n15719), .A2(n21416), .B1(n15736), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n15656) );
  OAI21_X1 U19158 ( .B1(n15657), .B2(n15721), .A(n15656), .ZN(n15658) );
  AOI21_X1 U19159 ( .B1(n15723), .B2(DATAI_28_), .A(n15658), .ZN(n15659) );
  OAI21_X1 U19160 ( .B1(n15763), .B2(n15739), .A(n15659), .ZN(P1_U2876) );
  AOI22_X1 U19161 ( .A1(n15719), .A2(n15660), .B1(n15736), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n15661) );
  OAI21_X1 U19162 ( .B1(n17807), .B2(n15721), .A(n15661), .ZN(n15662) );
  AOI21_X1 U19163 ( .B1(n15723), .B2(DATAI_27_), .A(n15662), .ZN(n15663) );
  OAI21_X1 U19164 ( .B1(n15664), .B2(n15739), .A(n15663), .ZN(P1_U2877) );
  INV_X1 U19165 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n15667) );
  AOI22_X1 U19166 ( .A1(n15719), .A2(n15665), .B1(n15736), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n15666) );
  OAI21_X1 U19167 ( .B1(n15721), .B2(n15667), .A(n15666), .ZN(n15668) );
  AOI21_X1 U19168 ( .B1(n15723), .B2(DATAI_26_), .A(n15668), .ZN(n15669) );
  OAI21_X1 U19169 ( .B1(n15670), .B2(n15739), .A(n15669), .ZN(P1_U2878) );
  INV_X1 U19170 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n15673) );
  AOI22_X1 U19171 ( .A1(n15719), .A2(n15671), .B1(n15736), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n15672) );
  OAI21_X1 U19172 ( .B1(n15721), .B2(n15673), .A(n15672), .ZN(n15674) );
  AOI21_X1 U19173 ( .B1(n15723), .B2(DATAI_25_), .A(n15674), .ZN(n15675) );
  OAI21_X1 U19174 ( .B1(n16115), .B2(n15739), .A(n15675), .ZN(P1_U2879) );
  INV_X1 U19175 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n15678) );
  AOI22_X1 U19176 ( .A1(n15719), .A2(n15676), .B1(n15736), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n15677) );
  OAI21_X1 U19177 ( .B1(n15721), .B2(n15678), .A(n15677), .ZN(n15679) );
  AOI21_X1 U19178 ( .B1(n15723), .B2(DATAI_24_), .A(n15679), .ZN(n15680) );
  OAI21_X1 U19179 ( .B1(n16125), .B2(n15739), .A(n15680), .ZN(P1_U2880) );
  INV_X1 U19180 ( .A(n15721), .ZN(n15709) );
  INV_X1 U19181 ( .A(n15719), .ZN(n15707) );
  OAI22_X1 U19182 ( .A1(n15707), .A2(n15681), .B1(n15733), .B2(n14448), .ZN(
        n15682) );
  AOI21_X1 U19183 ( .B1(n15709), .B2(BUF1_REG_23__SCAN_IN), .A(n15682), .ZN(
        n15684) );
  NAND2_X1 U19184 ( .A1(n15723), .A2(DATAI_23_), .ZN(n15683) );
  OAI211_X1 U19185 ( .C1(n15685), .C2(n15739), .A(n15684), .B(n15683), .ZN(
        P1_U2881) );
  INV_X1 U19186 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n15688) );
  AOI22_X1 U19187 ( .A1(n15719), .A2(n15686), .B1(n15736), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n15687) );
  OAI21_X1 U19188 ( .B1(n15721), .B2(n15688), .A(n15687), .ZN(n15691) );
  NOR2_X1 U19189 ( .A1(n15689), .A2(n15739), .ZN(n15690) );
  AOI211_X1 U19190 ( .C1(n15723), .C2(DATAI_22_), .A(n15691), .B(n15690), .ZN(
        n15692) );
  INV_X1 U19191 ( .A(n15692), .ZN(P1_U2882) );
  OAI22_X1 U19192 ( .A1(n15707), .A2(n15694), .B1(n15733), .B2(n15693), .ZN(
        n15695) );
  AOI21_X1 U19193 ( .B1(n15709), .B2(BUF1_REG_21__SCAN_IN), .A(n15695), .ZN(
        n15697) );
  NAND2_X1 U19194 ( .A1(n15723), .A2(DATAI_21_), .ZN(n15696) );
  OAI211_X1 U19195 ( .C1(n17203), .C2(n15739), .A(n15697), .B(n15696), .ZN(
        P1_U2883) );
  INV_X1 U19196 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n15700) );
  AOI22_X1 U19197 ( .A1(n15719), .A2(n15698), .B1(n15736), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n15699) );
  OAI21_X1 U19198 ( .B1(n15721), .B2(n15700), .A(n15699), .ZN(n15703) );
  NOR2_X1 U19199 ( .A1(n15701), .A2(n15739), .ZN(n15702) );
  AOI211_X1 U19200 ( .C1(n15723), .C2(DATAI_20_), .A(n15703), .B(n15702), .ZN(
        n15704) );
  INV_X1 U19201 ( .A(n15704), .ZN(P1_U2884) );
  OAI22_X1 U19202 ( .A1(n15707), .A2(n15706), .B1(n15733), .B2(n15705), .ZN(
        n15708) );
  AOI21_X1 U19203 ( .B1(n15709), .B2(BUF1_REG_19__SCAN_IN), .A(n15708), .ZN(
        n15711) );
  NAND2_X1 U19204 ( .A1(n15723), .A2(DATAI_19_), .ZN(n15710) );
  OAI211_X1 U19205 ( .C1(n17215), .C2(n15739), .A(n15711), .B(n15710), .ZN(
        P1_U2885) );
  INV_X1 U19206 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n15714) );
  AOI22_X1 U19207 ( .A1(n15719), .A2(n15712), .B1(n15736), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n15713) );
  OAI21_X1 U19208 ( .B1(n15721), .B2(n15714), .A(n15713), .ZN(n15715) );
  AOI21_X1 U19209 ( .B1(n15723), .B2(DATAI_18_), .A(n15715), .ZN(n15716) );
  OAI21_X1 U19210 ( .B1(n15717), .B2(n15739), .A(n15716), .ZN(P1_U2886) );
  AOI22_X1 U19211 ( .A1(n15719), .A2(n15718), .B1(n15736), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n15720) );
  OAI21_X1 U19212 ( .B1(n15721), .B2(n17819), .A(n15720), .ZN(n15722) );
  AOI21_X1 U19213 ( .B1(n15723), .B2(DATAI_16_), .A(n15722), .ZN(n15724) );
  OAI21_X1 U19214 ( .B1(n15725), .B2(n15739), .A(n15724), .ZN(P1_U2888) );
  OAI222_X1 U19215 ( .A1(n15739), .A2(n15728), .B1(n15733), .B2(n15727), .C1(
        n15732), .C2(n15726), .ZN(P1_U2889) );
  AOI22_X1 U19216 ( .A1(n15737), .A2(n21421), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15736), .ZN(n15729) );
  OAI21_X1 U19217 ( .B1(n15730), .B2(n15739), .A(n15729), .ZN(P1_U2890) );
  OAI222_X1 U19218 ( .A1(n15739), .A2(n15734), .B1(n15733), .B2(n21387), .C1(
        n15732), .C2(n15731), .ZN(P1_U2891) );
  XOR2_X1 U19219 ( .A(n15735), .B(n15335), .Z(n17299) );
  INV_X1 U19220 ( .A(n17299), .ZN(n15740) );
  AOI22_X1 U19221 ( .A1(n15737), .A2(n21416), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15736), .ZN(n15738) );
  OAI21_X1 U19222 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(P1_U2892) );
  NAND2_X1 U19223 ( .A1(n15742), .A2(n15741), .ZN(n15743) );
  AOI22_X1 U19224 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_29__SCAN_IN), .ZN(n15745) );
  OAI21_X1 U19225 ( .B1(n17305), .B2(n15746), .A(n15745), .ZN(n15747) );
  AOI21_X1 U19226 ( .B1(n15748), .B2(n17298), .A(n15747), .ZN(n15749) );
  OAI21_X1 U19227 ( .B1(n15750), .B2(n17312), .A(n15749), .ZN(P1_U2970) );
  MUX2_X1 U19228 ( .A(n15754), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .S(
        n16288), .Z(n15755) );
  OAI22_X1 U19229 ( .A1(n15759), .A2(n15758), .B1(n17352), .B2(n21505), .ZN(
        n15760) );
  AOI21_X1 U19230 ( .B1(n17296), .B2(n15761), .A(n15760), .ZN(n15762) );
  MUX2_X1 U19231 ( .A(n15765), .B(n15764), .S(n16288), .Z(n15766) );
  XNOR2_X1 U19232 ( .A(n15766), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16194) );
  NOR2_X1 U19233 ( .A1(n17352), .A2(n21503), .ZN(n16189) );
  AOI21_X1 U19234 ( .B1(n14161), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16189), .ZN(n15767) );
  OAI21_X1 U19235 ( .B1(n17305), .B2(n15768), .A(n15767), .ZN(n15769) );
  AOI21_X1 U19236 ( .B1(n15770), .B2(n17298), .A(n15769), .ZN(n15771) );
  OAI21_X1 U19237 ( .B1(n16194), .B2(n17312), .A(n15771), .ZN(P1_U2972) );
  AOI22_X1 U19238 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(keyinput178), .B1(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput221), .ZN(n15772) );
  OAI221_X1 U19239 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(keyinput178), .C1(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(keyinput221), .A(n15772), .ZN(
        n15779) );
  AOI22_X1 U19240 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(keyinput172), 
        .B1(P2_EBX_REG_20__SCAN_IN), .B2(keyinput185), .ZN(n15773) );
  OAI221_X1 U19241 ( .B1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B2(keyinput172), 
        .C1(P2_EBX_REG_20__SCAN_IN), .C2(keyinput185), .A(n15773), .ZN(n15778)
         );
  AOI22_X1 U19242 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(keyinput142), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(keyinput167), .ZN(n15774) );
  OAI221_X1 U19243 ( .B1(P3_EAX_REG_17__SCAN_IN), .B2(keyinput142), .C1(
        P2_REIP_REG_1__SCAN_IN), .C2(keyinput167), .A(n15774), .ZN(n15777) );
  AOI22_X1 U19244 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput243), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(keyinput206), .ZN(n15775) );
  OAI221_X1 U19245 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput243), .C1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .C2(keyinput206), .A(n15775), .ZN(
        n15776) );
  NOR4_X1 U19246 ( .A1(n15779), .A2(n15778), .A3(n15777), .A4(n15776), .ZN(
        n15807) );
  AOI22_X1 U19247 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(keyinput189), .B1(
        P2_INSTQUEUE_REG_7__4__SCAN_IN), .B2(keyinput169), .ZN(n15780) );
  OAI221_X1 U19248 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(keyinput189), .C1(
        P2_INSTQUEUE_REG_7__4__SCAN_IN), .C2(keyinput169), .A(n15780), .ZN(
        n15787) );
  AOI22_X1 U19249 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(keyinput171), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput132), .ZN(n15781) );
  OAI221_X1 U19250 ( .B1(P1_DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput171), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput132), .A(n15781), .ZN(n15786)
         );
  AOI22_X1 U19251 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(keyinput208), .B1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(keyinput177), .ZN(n15782) );
  OAI221_X1 U19252 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(keyinput208), .C1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .C2(keyinput177), .A(n15782), .ZN(
        n15785) );
  AOI22_X1 U19253 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(keyinput146), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(keyinput160), .ZN(n15783) );
  OAI221_X1 U19254 ( .B1(P2_BE_N_REG_2__SCAN_IN), .B2(keyinput146), .C1(
        P1_ADDRESS_REG_22__SCAN_IN), .C2(keyinput160), .A(n15783), .ZN(n15784)
         );
  NOR4_X1 U19255 ( .A1(n15787), .A2(n15786), .A3(n15785), .A4(n15784), .ZN(
        n15806) );
  AOI22_X1 U19256 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(keyinput222), .B1(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput203), .ZN(n15788) );
  OAI221_X1 U19257 ( .B1(P2_LWORD_REG_9__SCAN_IN), .B2(keyinput222), .C1(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(keyinput203), .A(n15788), .ZN(
        n15795) );
  AOI22_X1 U19258 ( .A1(P2_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput197), .B1(
        READY21_REG_SCAN_IN), .B2(keyinput136), .ZN(n15789) );
  OAI221_X1 U19259 ( .B1(P2_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput197), .C1(
        READY21_REG_SCAN_IN), .C2(keyinput136), .A(n15789), .ZN(n15794) );
  AOI22_X1 U19260 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(keyinput207), 
        .B1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B2(keyinput158), .ZN(n15790) );
  OAI221_X1 U19261 ( .B1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B2(keyinput207), 
        .C1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .C2(keyinput158), .A(n15790), 
        .ZN(n15793) );
  AOI22_X1 U19262 ( .A1(P3_UWORD_REG_5__SCAN_IN), .A2(keyinput151), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(keyinput242), .ZN(n15791) );
  OAI221_X1 U19263 ( .B1(P3_UWORD_REG_5__SCAN_IN), .B2(keyinput151), .C1(
        P2_EBX_REG_5__SCAN_IN), .C2(keyinput242), .A(n15791), .ZN(n15792) );
  NOR4_X1 U19264 ( .A1(n15795), .A2(n15794), .A3(n15793), .A4(n15792), .ZN(
        n15805) );
  AOI22_X1 U19265 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(keyinput251), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(keyinput205), .ZN(n15796) );
  OAI221_X1 U19266 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(keyinput251), .C1(
        P1_DATAO_REG_26__SCAN_IN), .C2(keyinput205), .A(n15796), .ZN(n15803)
         );
  AOI22_X1 U19267 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput138), .B1(
        DATAI_13_), .B2(keyinput250), .ZN(n15797) );
  OAI221_X1 U19268 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput138), .C1(
        DATAI_13_), .C2(keyinput250), .A(n15797), .ZN(n15802) );
  AOI22_X1 U19269 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput214), 
        .B1(P1_DATAO_REG_13__SCAN_IN), .B2(keyinput141), .ZN(n15798) );
  OAI221_X1 U19270 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput214), 
        .C1(P1_DATAO_REG_13__SCAN_IN), .C2(keyinput141), .A(n15798), .ZN(
        n15801) );
  AOI22_X1 U19271 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(keyinput238), 
        .B1(P3_LWORD_REG_15__SCAN_IN), .B2(keyinput179), .ZN(n15799) );
  OAI221_X1 U19272 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput238), 
        .C1(P3_LWORD_REG_15__SCAN_IN), .C2(keyinput179), .A(n15799), .ZN(
        n15800) );
  NOR4_X1 U19273 ( .A1(n15803), .A2(n15802), .A3(n15801), .A4(n15800), .ZN(
        n15804) );
  NAND4_X1 U19274 ( .A1(n15807), .A2(n15806), .A3(n15805), .A4(n15804), .ZN(
        n15930) );
  AOI22_X1 U19275 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(keyinput218), .B1(
        P1_EAX_REG_8__SCAN_IN), .B2(keyinput161), .ZN(n15808) );
  OAI221_X1 U19276 ( .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput218), .C1(
        P1_EAX_REG_8__SCAN_IN), .C2(keyinput161), .A(n15808), .ZN(n15815) );
  AOI22_X1 U19277 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(keyinput235), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(keyinput188), .ZN(n15809) );
  OAI221_X1 U19278 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(keyinput235), .C1(
        P3_EAX_REG_21__SCAN_IN), .C2(keyinput188), .A(n15809), .ZN(n15814) );
  AOI22_X1 U19279 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(keyinput204), 
        .B1(P3_LWORD_REG_13__SCAN_IN), .B2(keyinput201), .ZN(n15810) );
  OAI221_X1 U19280 ( .B1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput204), 
        .C1(P3_LWORD_REG_13__SCAN_IN), .C2(keyinput201), .A(n15810), .ZN(
        n15813) );
  AOI22_X1 U19281 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(keyinput210), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(keyinput156), .ZN(n15811) );
  OAI221_X1 U19282 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(keyinput210), .C1(
        P2_EBX_REG_11__SCAN_IN), .C2(keyinput156), .A(n15811), .ZN(n15812) );
  NOR4_X1 U19283 ( .A1(n15815), .A2(n15814), .A3(n15813), .A4(n15812), .ZN(
        n15843) );
  AOI22_X1 U19284 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(keyinput176), 
        .B1(P2_EAX_REG_29__SCAN_IN), .B2(keyinput202), .ZN(n15816) );
  OAI221_X1 U19285 ( .B1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(keyinput176), 
        .C1(P2_EAX_REG_29__SCAN_IN), .C2(keyinput202), .A(n15816), .ZN(n15823)
         );
  AOI22_X1 U19286 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(keyinput149), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(keyinput226), .ZN(n15817) );
  OAI221_X1 U19287 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(keyinput149), .C1(
        P1_ADDRESS_REG_8__SCAN_IN), .C2(keyinput226), .A(n15817), .ZN(n15822)
         );
  AOI22_X1 U19288 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(keyinput215), 
        .B1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput131), .ZN(n15818) );
  OAI221_X1 U19289 ( .B1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B2(keyinput215), 
        .C1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .C2(keyinput131), .A(n15818), 
        .ZN(n15821) );
  AOI22_X1 U19290 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(keyinput192), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(keyinput223), .ZN(n15819) );
  OAI221_X1 U19291 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(keyinput192), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(keyinput223), .A(n15819), .ZN(n15820) );
  NOR4_X1 U19292 ( .A1(n15823), .A2(n15822), .A3(n15821), .A4(n15820), .ZN(
        n15842) );
  AOI22_X1 U19293 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput230), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput245), .ZN(n15824) );
  OAI221_X1 U19294 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput230), .C1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput245), .A(n15824), .ZN(
        n15831) );
  AOI22_X1 U19295 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(keyinput184), 
        .B1(P3_EAX_REG_22__SCAN_IN), .B2(keyinput157), .ZN(n15825) );
  OAI221_X1 U19296 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(keyinput184), 
        .C1(P3_EAX_REG_22__SCAN_IN), .C2(keyinput157), .A(n15825), .ZN(n15830)
         );
  AOI22_X1 U19297 ( .A1(P1_DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput211), .B1(
        P1_EAX_REG_13__SCAN_IN), .B2(keyinput135), .ZN(n15826) );
  OAI221_X1 U19298 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput211), .C1(
        P1_EAX_REG_13__SCAN_IN), .C2(keyinput135), .A(n15826), .ZN(n15829) );
  AOI22_X1 U19299 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput162), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(keyinput239), .ZN(n15827) );
  OAI221_X1 U19300 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput162), .C1(
        P1_ADDRESS_REG_11__SCAN_IN), .C2(keyinput239), .A(n15827), .ZN(n15828)
         );
  NOR4_X1 U19301 ( .A1(n15831), .A2(n15830), .A3(n15829), .A4(n15828), .ZN(
        n15841) );
  AOI22_X1 U19302 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(keyinput254), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(keyinput148), .ZN(n15832) );
  OAI221_X1 U19303 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput254), .C1(
        P1_REIP_REG_10__SCAN_IN), .C2(keyinput148), .A(n15832), .ZN(n15839) );
  AOI22_X1 U19304 ( .A1(P2_EBX_REG_3__SCAN_IN), .A2(keyinput247), .B1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(keyinput209), .ZN(n15833) );
  OAI221_X1 U19305 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(keyinput247), .C1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .C2(keyinput209), .A(n15833), .ZN(
        n15838) );
  AOI22_X1 U19306 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput253), .B1(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput168), .ZN(n15834) );
  OAI221_X1 U19307 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput253), .C1(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput168), .A(n15834), 
        .ZN(n15837) );
  AOI22_X1 U19308 ( .A1(BUF1_REG_21__SCAN_IN), .A2(keyinput155), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput154), .ZN(n15835) );
  OAI221_X1 U19309 ( .B1(BUF1_REG_21__SCAN_IN), .B2(keyinput155), .C1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(keyinput154), .A(n15835), 
        .ZN(n15836) );
  NOR4_X1 U19310 ( .A1(n15839), .A2(n15838), .A3(n15837), .A4(n15836), .ZN(
        n15840) );
  NAND4_X1 U19311 ( .A1(n15843), .A2(n15842), .A3(n15841), .A4(n15840), .ZN(
        n15929) );
  AOI22_X1 U19312 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(keyinput186), 
        .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput219), .ZN(n15844) );
  OAI221_X1 U19313 ( .B1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B2(keyinput186), 
        .C1(P1_EBX_REG_5__SCAN_IN), .C2(keyinput219), .A(n15844), .ZN(n15852)
         );
  AOI22_X1 U19314 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(keyinput255), .B1(
        BUF2_REG_14__SCAN_IN), .B2(keyinput163), .ZN(n15845) );
  OAI221_X1 U19315 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(keyinput255), .C1(
        BUF2_REG_14__SCAN_IN), .C2(keyinput163), .A(n15845), .ZN(n15851) );
  INV_X1 U19316 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n15847) );
  AOI22_X1 U19317 ( .A1(keyinput150), .A2(P3_ADDRESS_REG_10__SCAN_IN), .B1(
        n15847), .B2(keyinput134), .ZN(n15846) );
  OAI221_X1 U19318 ( .B1(keyinput150), .B2(P3_ADDRESS_REG_10__SCAN_IN), .C1(
        n15847), .C2(keyinput134), .A(n15846), .ZN(n15850) );
  INV_X1 U19319 ( .A(P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21093) );
  AOI22_X1 U19320 ( .A1(n21093), .A2(keyinput236), .B1(keyinput145), .B2(
        n19456), .ZN(n15848) );
  OAI221_X1 U19321 ( .B1(n21093), .B2(keyinput236), .C1(n19456), .C2(
        keyinput145), .A(n15848), .ZN(n15849) );
  NOR4_X1 U19322 ( .A1(n15852), .A2(n15851), .A3(n15850), .A4(n15849), .ZN(
        n15884) );
  AOI22_X1 U19323 ( .A1(n15942), .A2(keyinput128), .B1(keyinput183), .B2(
        n20160), .ZN(n15853) );
  OAI221_X1 U19324 ( .B1(n15942), .B2(keyinput128), .C1(n20160), .C2(
        keyinput183), .A(n15853), .ZN(n15861) );
  AOI22_X1 U19325 ( .A1(n17879), .A2(keyinput139), .B1(n21463), .B2(
        keyinput194), .ZN(n15854) );
  OAI221_X1 U19326 ( .B1(n17879), .B2(keyinput139), .C1(n21463), .C2(
        keyinput194), .A(n15854), .ZN(n15860) );
  INV_X1 U19327 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n20531) );
  AOI22_X1 U19328 ( .A1(n20531), .A2(keyinput144), .B1(n15856), .B2(
        keyinput225), .ZN(n15855) );
  OAI221_X1 U19329 ( .B1(n20531), .B2(keyinput144), .C1(n15856), .C2(
        keyinput225), .A(n15855), .ZN(n15859) );
  INV_X1 U19330 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n18739) );
  AOI22_X1 U19331 ( .A1(n18739), .A2(keyinput175), .B1(n21415), .B2(
        keyinput224), .ZN(n15857) );
  OAI221_X1 U19332 ( .B1(n18739), .B2(keyinput175), .C1(n21415), .C2(
        keyinput224), .A(n15857), .ZN(n15858) );
  NOR4_X1 U19333 ( .A1(n15861), .A2(n15860), .A3(n15859), .A4(n15858), .ZN(
        n15883) );
  AOI22_X1 U19334 ( .A1(n15667), .A2(keyinput166), .B1(n11729), .B2(
        keyinput231), .ZN(n15862) );
  OAI221_X1 U19335 ( .B1(n15667), .B2(keyinput166), .C1(n11729), .C2(
        keyinput231), .A(n15862), .ZN(n15869) );
  INV_X1 U19336 ( .A(P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n21091) );
  AOI22_X1 U19337 ( .A1(n21091), .A2(keyinput165), .B1(n16191), .B2(
        keyinput216), .ZN(n15863) );
  OAI221_X1 U19338 ( .B1(n21091), .B2(keyinput165), .C1(n16191), .C2(
        keyinput216), .A(n15863), .ZN(n15868) );
  INV_X1 U19339 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21471) );
  AOI22_X1 U19340 ( .A1(n21394), .A2(keyinput241), .B1(n21471), .B2(
        keyinput133), .ZN(n15864) );
  OAI221_X1 U19341 ( .B1(n21394), .B2(keyinput241), .C1(n21471), .C2(
        keyinput133), .A(n15864), .ZN(n15867) );
  INV_X1 U19342 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18288) );
  INV_X1 U19343 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18487) );
  AOI22_X1 U19344 ( .A1(n18288), .A2(keyinput187), .B1(keyinput248), .B2(
        n18487), .ZN(n15865) );
  OAI221_X1 U19345 ( .B1(n18288), .B2(keyinput187), .C1(n18487), .C2(
        keyinput248), .A(n15865), .ZN(n15866) );
  NOR4_X1 U19346 ( .A1(n15869), .A2(n15868), .A3(n15867), .A4(n15866), .ZN(
        n15882) );
  INV_X1 U19347 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15871) );
  AOI22_X1 U19348 ( .A1(n15872), .A2(keyinput234), .B1(keyinput195), .B2(
        n15871), .ZN(n15870) );
  OAI221_X1 U19349 ( .B1(n15872), .B2(keyinput234), .C1(n15871), .C2(
        keyinput195), .A(n15870), .ZN(n15880) );
  INV_X1 U19350 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15874) );
  INV_X1 U19351 ( .A(P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21089) );
  AOI22_X1 U19352 ( .A1(n15874), .A2(keyinput143), .B1(keyinput252), .B2(
        n21089), .ZN(n15873) );
  OAI221_X1 U19353 ( .B1(n15874), .B2(keyinput143), .C1(n21089), .C2(
        keyinput252), .A(n15873), .ZN(n15879) );
  AOI22_X1 U19354 ( .A1(n17030), .A2(keyinput193), .B1(n16707), .B2(
        keyinput174), .ZN(n15875) );
  OAI221_X1 U19355 ( .B1(n17030), .B2(keyinput193), .C1(n16707), .C2(
        keyinput174), .A(n15875), .ZN(n15878) );
  INV_X1 U19356 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n18760) );
  AOI22_X1 U19357 ( .A1(n18760), .A2(keyinput220), .B1(n11708), .B2(
        keyinput237), .ZN(n15876) );
  OAI221_X1 U19358 ( .B1(n18760), .B2(keyinput220), .C1(n11708), .C2(
        keyinput237), .A(n15876), .ZN(n15877) );
  NOR4_X1 U19359 ( .A1(n15880), .A2(n15879), .A3(n15878), .A4(n15877), .ZN(
        n15881) );
  NAND4_X1 U19360 ( .A1(n15884), .A2(n15883), .A3(n15882), .A4(n15881), .ZN(
        n15928) );
  INV_X1 U19361 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15987) );
  AOI22_X1 U19362 ( .A1(n13804), .A2(keyinput153), .B1(keyinput227), .B2(
        n15987), .ZN(n15885) );
  OAI221_X1 U19363 ( .B1(n13804), .B2(keyinput153), .C1(n15987), .C2(
        keyinput227), .A(n15885), .ZN(n15894) );
  INV_X1 U19364 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20140) );
  AOI22_X1 U19365 ( .A1(n14738), .A2(keyinput229), .B1(keyinput129), .B2(
        n20140), .ZN(n15886) );
  OAI221_X1 U19366 ( .B1(n14738), .B2(keyinput229), .C1(n20140), .C2(
        keyinput129), .A(n15886), .ZN(n15893) );
  INV_X1 U19367 ( .A(READY11_REG_SCAN_IN), .ZN(n15888) );
  AOI22_X1 U19368 ( .A1(n15888), .A2(keyinput198), .B1(keyinput244), .B2(
        n20026), .ZN(n15887) );
  OAI221_X1 U19369 ( .B1(n15888), .B2(keyinput198), .C1(n20026), .C2(
        keyinput244), .A(n15887), .ZN(n15892) );
  AOI22_X1 U19370 ( .A1(n15955), .A2(keyinput173), .B1(n15890), .B2(
        keyinput232), .ZN(n15889) );
  OAI221_X1 U19371 ( .B1(n15955), .B2(keyinput173), .C1(n15890), .C2(
        keyinput232), .A(n15889), .ZN(n15891) );
  NOR4_X1 U19372 ( .A1(n15894), .A2(n15893), .A3(n15892), .A4(n15891), .ZN(
        n15926) );
  INV_X1 U19373 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n17483) );
  INV_X1 U19374 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n20508) );
  AOI22_X1 U19375 ( .A1(n17483), .A2(keyinput180), .B1(keyinput213), .B2(
        n20508), .ZN(n15895) );
  OAI221_X1 U19376 ( .B1(n17483), .B2(keyinput180), .C1(n20508), .C2(
        keyinput213), .A(n15895), .ZN(n15904) );
  AOI22_X1 U19377 ( .A1(n12320), .A2(keyinput152), .B1(keyinput147), .B2(
        n18073), .ZN(n15896) );
  OAI221_X1 U19378 ( .B1(n12320), .B2(keyinput152), .C1(n18073), .C2(
        keyinput147), .A(n15896), .ZN(n15903) );
  INV_X1 U19379 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15899) );
  AOI22_X1 U19380 ( .A1(n15899), .A2(keyinput240), .B1(keyinput164), .B2(
        n15898), .ZN(n15897) );
  OAI221_X1 U19381 ( .B1(n15899), .B2(keyinput240), .C1(n15898), .C2(
        keyinput164), .A(n15897), .ZN(n15902) );
  AOI22_X1 U19382 ( .A1(n10705), .A2(keyinput200), .B1(n15997), .B2(
        keyinput190), .ZN(n15900) );
  OAI221_X1 U19383 ( .B1(n10705), .B2(keyinput200), .C1(n15997), .C2(
        keyinput190), .A(n15900), .ZN(n15901) );
  NOR4_X1 U19384 ( .A1(n15904), .A2(n15903), .A3(n15902), .A4(n15901), .ZN(
        n15925) );
  INV_X1 U19385 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21466) );
  INV_X1 U19386 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20521) );
  AOI22_X1 U19387 ( .A1(n21466), .A2(keyinput170), .B1(n20521), .B2(
        keyinput191), .ZN(n15905) );
  OAI221_X1 U19388 ( .B1(n21466), .B2(keyinput170), .C1(n20521), .C2(
        keyinput191), .A(n15905), .ZN(n15914) );
  INV_X1 U19389 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17883) );
  INV_X1 U19390 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15907) );
  AOI22_X1 U19391 ( .A1(n17883), .A2(keyinput181), .B1(keyinput249), .B2(
        n15907), .ZN(n15906) );
  OAI221_X1 U19392 ( .B1(n17883), .B2(keyinput181), .C1(n15907), .C2(
        keyinput249), .A(n15906), .ZN(n15913) );
  INV_X1 U19393 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n21152) );
  AOI22_X1 U19394 ( .A1(n17138), .A2(keyinput233), .B1(n21152), .B2(
        keyinput140), .ZN(n15908) );
  OAI221_X1 U19395 ( .B1(n17138), .B2(keyinput233), .C1(n21152), .C2(
        keyinput140), .A(n15908), .ZN(n15912) );
  INV_X1 U19396 ( .A(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15910) );
  INV_X1 U19397 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n16467) );
  AOI22_X1 U19398 ( .A1(n15910), .A2(keyinput196), .B1(n16467), .B2(
        keyinput182), .ZN(n15909) );
  OAI221_X1 U19399 ( .B1(n15910), .B2(keyinput196), .C1(n16467), .C2(
        keyinput182), .A(n15909), .ZN(n15911) );
  NOR4_X1 U19400 ( .A1(n15914), .A2(n15913), .A3(n15912), .A4(n15911), .ZN(
        n15924) );
  INV_X1 U19401 ( .A(P3_DATAO_REG_19__SCAN_IN), .ZN(n18752) );
  AOI22_X1 U19402 ( .A1(n18752), .A2(keyinput130), .B1(n15953), .B2(
        keyinput228), .ZN(n15915) );
  OAI221_X1 U19403 ( .B1(n18752), .B2(keyinput130), .C1(n15953), .C2(
        keyinput228), .A(n15915), .ZN(n15922) );
  INV_X1 U19404 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n18737) );
  AOI22_X1 U19405 ( .A1(n15940), .A2(keyinput137), .B1(keyinput212), .B2(
        n18737), .ZN(n15916) );
  OAI221_X1 U19406 ( .B1(n15940), .B2(keyinput137), .C1(n18737), .C2(
        keyinput212), .A(n15916), .ZN(n15921) );
  INV_X1 U19407 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21487) );
  INV_X1 U19408 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15950) );
  AOI22_X1 U19409 ( .A1(n21487), .A2(keyinput199), .B1(keyinput159), .B2(
        n15950), .ZN(n15917) );
  OAI221_X1 U19410 ( .B1(n21487), .B2(keyinput199), .C1(n15950), .C2(
        keyinput159), .A(n15917), .ZN(n15920) );
  AOI22_X1 U19411 ( .A1(n16713), .A2(keyinput246), .B1(keyinput217), .B2(
        n18454), .ZN(n15918) );
  OAI221_X1 U19412 ( .B1(n16713), .B2(keyinput246), .C1(n18454), .C2(
        keyinput217), .A(n15918), .ZN(n15919) );
  NOR4_X1 U19413 ( .A1(n15922), .A2(n15921), .A3(n15920), .A4(n15919), .ZN(
        n15923) );
  NAND4_X1 U19414 ( .A1(n15926), .A2(n15925), .A3(n15924), .A4(n15923), .ZN(
        n15927) );
  NOR4_X1 U19415 ( .A1(n15930), .A2(n15929), .A3(n15928), .A4(n15927), .ZN(
        n16095) );
  AOI22_X1 U19416 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(keyinput120), 
        .B1(DATAI_13_), .B2(keyinput122), .ZN(n15931) );
  OAI221_X1 U19417 ( .B1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput120), 
        .C1(DATAI_13_), .C2(keyinput122), .A(n15931), .ZN(n15938) );
  AOI22_X1 U19418 ( .A1(P3_DATAO_REG_16__SCAN_IN), .A2(keyinput92), .B1(
        P2_LWORD_REG_9__SCAN_IN), .B2(keyinput94), .ZN(n15932) );
  OAI221_X1 U19419 ( .B1(P3_DATAO_REG_16__SCAN_IN), .B2(keyinput92), .C1(
        P2_LWORD_REG_9__SCAN_IN), .C2(keyinput94), .A(n15932), .ZN(n15937) );
  INV_X1 U19420 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U19421 ( .A1(n16713), .A2(keyinput118), .B1(keyinput57), .B2(n17476), .ZN(n15933) );
  OAI221_X1 U19422 ( .B1(n16713), .B2(keyinput118), .C1(n17476), .C2(
        keyinput57), .A(n15933), .ZN(n15936) );
  INV_X1 U19423 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n18510) );
  AOI22_X1 U19424 ( .A1(n18288), .A2(keyinput59), .B1(n18510), .B2(keyinput107), .ZN(n15934) );
  OAI221_X1 U19425 ( .B1(n18288), .B2(keyinput59), .C1(n18510), .C2(
        keyinput107), .A(n15934), .ZN(n15935) );
  NOR4_X1 U19426 ( .A1(n15938), .A2(n15937), .A3(n15936), .A4(n15935), .ZN(
        n15972) );
  AOI22_X1 U19427 ( .A1(n21394), .A2(keyinput113), .B1(n15940), .B2(keyinput9), 
        .ZN(n15939) );
  OAI221_X1 U19428 ( .B1(n21394), .B2(keyinput113), .C1(n15940), .C2(keyinput9), .A(n15939), .ZN(n15948) );
  AOI22_X1 U19429 ( .A1(n15942), .A2(keyinput0), .B1(keyinput5), .B2(n21471), 
        .ZN(n15941) );
  OAI221_X1 U19430 ( .B1(n15942), .B2(keyinput0), .C1(n21471), .C2(keyinput5), 
        .A(n15941), .ZN(n15947) );
  INV_X1 U19431 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20568) );
  INV_X1 U19432 ( .A(P3_LWORD_REG_13__SCAN_IN), .ZN(n18766) );
  AOI22_X1 U19433 ( .A1(n20568), .A2(keyinput27), .B1(n18766), .B2(keyinput73), 
        .ZN(n15943) );
  OAI221_X1 U19434 ( .B1(n20568), .B2(keyinput27), .C1(n18766), .C2(keyinput73), .A(n15943), .ZN(n15946) );
  INV_X1 U19435 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21473) );
  INV_X1 U19436 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n20813) );
  AOI22_X1 U19437 ( .A1(n21473), .A2(keyinput98), .B1(n20813), .B2(keyinput3), 
        .ZN(n15944) );
  OAI221_X1 U19438 ( .B1(n21473), .B2(keyinput98), .C1(n20813), .C2(keyinput3), 
        .A(n15944), .ZN(n15945) );
  NOR4_X1 U19439 ( .A1(n15948), .A2(n15947), .A3(n15946), .A4(n15945), .ZN(
        n15971) );
  AOI22_X1 U19440 ( .A1(n12996), .A2(keyinput41), .B1(keyinput31), .B2(n15950), 
        .ZN(n15949) );
  OAI221_X1 U19441 ( .B1(n12996), .B2(keyinput41), .C1(n15950), .C2(keyinput31), .A(n15949), .ZN(n15959) );
  INV_X1 U19442 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21478) );
  AOI22_X1 U19443 ( .A1(n18108), .A2(keyinput123), .B1(n21478), .B2(
        keyinput111), .ZN(n15951) );
  OAI221_X1 U19444 ( .B1(n18108), .B2(keyinput123), .C1(n21478), .C2(
        keyinput111), .A(n15951), .ZN(n15958) );
  INV_X1 U19445 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18748) );
  AOI22_X1 U19446 ( .A1(n15953), .A2(keyinput100), .B1(keyinput60), .B2(n18748), .ZN(n15952) );
  OAI221_X1 U19447 ( .B1(n15953), .B2(keyinput100), .C1(n18748), .C2(
        keyinput60), .A(n15952), .ZN(n15957) );
  INV_X1 U19448 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18799) );
  AOI22_X1 U19449 ( .A1(n18799), .A2(keyinput14), .B1(keyinput45), .B2(n15955), 
        .ZN(n15954) );
  OAI221_X1 U19450 ( .B1(n18799), .B2(keyinput14), .C1(n15955), .C2(keyinput45), .A(n15954), .ZN(n15956) );
  NOR4_X1 U19451 ( .A1(n15959), .A2(n15958), .A3(n15957), .A4(n15956), .ZN(
        n15970) );
  AOI22_X1 U19452 ( .A1(n17228), .A2(keyinput117), .B1(keyinput2), .B2(n18752), 
        .ZN(n15960) );
  OAI221_X1 U19453 ( .B1(n17228), .B2(keyinput117), .C1(n18752), .C2(keyinput2), .A(n15960), .ZN(n15968) );
  AOI22_X1 U19454 ( .A1(n17030), .A2(keyinput65), .B1(n12320), .B2(keyinput24), 
        .ZN(n15961) );
  OAI221_X1 U19455 ( .B1(n17030), .B2(keyinput65), .C1(n12320), .C2(keyinput24), .A(n15961), .ZN(n15967) );
  AOI22_X1 U19456 ( .A1(n20508), .A2(keyinput85), .B1(n15963), .B2(keyinput78), 
        .ZN(n15962) );
  OAI221_X1 U19457 ( .B1(n20508), .B2(keyinput85), .C1(n15963), .C2(keyinput78), .A(n15962), .ZN(n15966) );
  AOI22_X1 U19458 ( .A1(n20140), .A2(keyinput1), .B1(n21474), .B2(keyinput127), 
        .ZN(n15964) );
  OAI221_X1 U19459 ( .B1(n20140), .B2(keyinput1), .C1(n21474), .C2(keyinput127), .A(n15964), .ZN(n15965) );
  NOR4_X1 U19460 ( .A1(n15968), .A2(n15967), .A3(n15966), .A4(n15965), .ZN(
        n15969) );
  NAND4_X1 U19461 ( .A1(n15972), .A2(n15971), .A3(n15970), .A4(n15969), .ZN(
        n16094) );
  INV_X1 U19462 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n15974) );
  AOI22_X1 U19463 ( .A1(n21398), .A2(keyinput33), .B1(keyinput13), .B2(n15974), 
        .ZN(n15973) );
  OAI221_X1 U19464 ( .B1(n21398), .B2(keyinput33), .C1(n15974), .C2(keyinput13), .A(n15973), .ZN(n15984) );
  AOI22_X1 U19465 ( .A1(n15667), .A2(keyinput38), .B1(n15976), .B2(keyinput48), 
        .ZN(n15975) );
  OAI221_X1 U19466 ( .B1(n15667), .B2(keyinput38), .C1(n15976), .C2(keyinput48), .A(n15975), .ZN(n15983) );
  INV_X1 U19467 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n15978) );
  AOI22_X1 U19468 ( .A1(n15978), .A2(keyinput83), .B1(n16707), .B2(keyinput46), 
        .ZN(n15977) );
  OAI221_X1 U19469 ( .B1(n15978), .B2(keyinput83), .C1(n16707), .C2(keyinput46), .A(n15977), .ZN(n15982) );
  INV_X1 U19470 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15980) );
  AOI22_X1 U19471 ( .A1(n17871), .A2(keyinput102), .B1(keyinput58), .B2(n15980), .ZN(n15979) );
  OAI221_X1 U19472 ( .B1(n17871), .B2(keyinput102), .C1(n15980), .C2(
        keyinput58), .A(n15979), .ZN(n15981) );
  NOR4_X1 U19473 ( .A1(n15984), .A2(n15983), .A3(n15982), .A4(n15981), .ZN(
        n16017) );
  INV_X1 U19474 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18746) );
  INV_X1 U19475 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n21496) );
  AOI22_X1 U19476 ( .A1(n18746), .A2(keyinput29), .B1(n21496), .B2(keyinput32), 
        .ZN(n15985) );
  OAI221_X1 U19477 ( .B1(n18746), .B2(keyinput29), .C1(n21496), .C2(keyinput32), .A(n15985), .ZN(n15994) );
  AOI22_X1 U19478 ( .A1(n15987), .A2(keyinput99), .B1(n13684), .B2(keyinput93), 
        .ZN(n15986) );
  OAI221_X1 U19479 ( .B1(n15987), .B2(keyinput99), .C1(n13684), .C2(keyinput93), .A(n15986), .ZN(n15993) );
  AOI22_X1 U19480 ( .A1(n18454), .A2(keyinput89), .B1(n17483), .B2(keyinput52), 
        .ZN(n15988) );
  OAI221_X1 U19481 ( .B1(n18454), .B2(keyinput89), .C1(n17483), .C2(keyinput52), .A(n15988), .ZN(n15992) );
  INV_X1 U19482 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n15990) );
  AOI22_X1 U19483 ( .A1(n20521), .A2(keyinput63), .B1(keyinput90), .B2(n15990), 
        .ZN(n15989) );
  OAI221_X1 U19484 ( .B1(n20521), .B2(keyinput63), .C1(n15990), .C2(keyinput90), .A(n15989), .ZN(n15991) );
  NOR4_X1 U19485 ( .A1(n15994), .A2(n15993), .A3(n15992), .A4(n15991), .ZN(
        n16016) );
  AOI22_X1 U19486 ( .A1(n16191), .A2(keyinput88), .B1(keyinput110), .B2(n13343), .ZN(n15995) );
  OAI221_X1 U19487 ( .B1(n16191), .B2(keyinput88), .C1(n13343), .C2(
        keyinput110), .A(n15995), .ZN(n16004) );
  AOI22_X1 U19488 ( .A1(n15997), .A2(keyinput62), .B1(n11729), .B2(keyinput103), .ZN(n15996) );
  OAI221_X1 U19489 ( .B1(n15997), .B2(keyinput62), .C1(n11729), .C2(
        keyinput103), .A(n15996), .ZN(n16003) );
  AOI22_X1 U19490 ( .A1(n20531), .A2(keyinput16), .B1(n16475), .B2(keyinput74), 
        .ZN(n15998) );
  OAI221_X1 U19491 ( .B1(n20531), .B2(keyinput16), .C1(n16475), .C2(keyinput74), .A(n15998), .ZN(n16002) );
  INV_X1 U19492 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16000) );
  AOI22_X1 U19493 ( .A1(n16000), .A2(keyinput30), .B1(n14738), .B2(keyinput101), .ZN(n15999) );
  OAI221_X1 U19494 ( .B1(n16000), .B2(keyinput30), .C1(n14738), .C2(
        keyinput101), .A(n15999), .ZN(n16001) );
  NOR4_X1 U19495 ( .A1(n16004), .A2(n16003), .A3(n16002), .A4(n16001), .ZN(
        n16015) );
  INV_X1 U19496 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20094) );
  AOI22_X1 U19497 ( .A1(n21487), .A2(keyinput71), .B1(keyinput22), .B2(n20094), 
        .ZN(n16005) );
  OAI221_X1 U19498 ( .B1(n21487), .B2(keyinput71), .C1(n20094), .C2(keyinput22), .A(n16005), .ZN(n16013) );
  AOI22_X1 U19499 ( .A1(n16007), .A2(keyinput40), .B1(keyinput19), .B2(n18073), 
        .ZN(n16006) );
  OAI221_X1 U19500 ( .B1(n16007), .B2(keyinput40), .C1(n18073), .C2(keyinput19), .A(n16006), .ZN(n16012) );
  INV_X1 U19501 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21516) );
  AOI22_X1 U19502 ( .A1(n21516), .A2(keyinput34), .B1(n17869), .B2(keyinput4), 
        .ZN(n16008) );
  OAI221_X1 U19503 ( .B1(n21516), .B2(keyinput34), .C1(n17869), .C2(keyinput4), 
        .A(n16008), .ZN(n16011) );
  INV_X1 U19504 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n20504) );
  INV_X1 U19505 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n18843) );
  AOI22_X1 U19506 ( .A1(n20504), .A2(keyinput115), .B1(n18843), .B2(keyinput35), .ZN(n16009) );
  OAI221_X1 U19507 ( .B1(n20504), .B2(keyinput115), .C1(n18843), .C2(
        keyinput35), .A(n16009), .ZN(n16010) );
  NOR4_X1 U19508 ( .A1(n16013), .A2(n16012), .A3(n16011), .A4(n16010), .ZN(
        n16014) );
  NAND4_X1 U19509 ( .A1(n16017), .A2(n16016), .A3(n16015), .A4(n16014), .ZN(
        n16093) );
  OAI22_X1 U19510 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(keyinput97), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput105), .ZN(n16018) );
  AOI221_X1 U19511 ( .B1(P2_EBX_REG_13__SCAN_IN), .B2(keyinput97), .C1(
        keyinput105), .C2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n16018), 
        .ZN(n16025) );
  OAI22_X1 U19512 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(keyinput109), 
        .B1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B2(keyinput44), .ZN(n16019) );
  AOI221_X1 U19513 ( .B1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput109), 
        .C1(keyinput44), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(n16019), .ZN(
        n16024) );
  OAI22_X1 U19514 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(keyinput82), .B1(
        keyinput87), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16020) );
  AOI221_X1 U19515 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(keyinput82), .C1(
        P1_INSTQUEUE_REG_9__2__SCAN_IN), .C2(keyinput87), .A(n16020), .ZN(
        n16023) );
  OAI22_X1 U19516 ( .A1(P2_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput69), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(keyinput53), .ZN(n16021) );
  AOI221_X1 U19517 ( .B1(P2_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput69), .C1(
        keyinput53), .C2(P1_DATAO_REG_31__SCAN_IN), .A(n16021), .ZN(n16022) );
  NAND4_X1 U19518 ( .A1(n16025), .A2(n16024), .A3(n16023), .A4(n16022), .ZN(
        n16053) );
  OAI22_X1 U19519 ( .A1(READY21_REG_SCAN_IN), .A2(keyinput8), .B1(
        P3_REIP_REG_15__SCAN_IN), .B2(keyinput50), .ZN(n16026) );
  AOI221_X1 U19520 ( .B1(READY21_REG_SCAN_IN), .B2(keyinput8), .C1(keyinput50), 
        .C2(P3_REIP_REG_15__SCAN_IN), .A(n16026), .ZN(n16033) );
  OAI22_X1 U19521 ( .A1(P1_EAX_REG_0__SCAN_IN), .A2(keyinput96), .B1(
        keyinput64), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16027) );
  AOI221_X1 U19522 ( .B1(P1_EAX_REG_0__SCAN_IN), .B2(keyinput96), .C1(
        P3_EBX_REG_18__SCAN_IN), .C2(keyinput64), .A(n16027), .ZN(n16032) );
  OAI22_X1 U19523 ( .A1(P3_LWORD_REG_15__SCAN_IN), .A2(keyinput51), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(keyinput55), .ZN(n16028) );
  AOI221_X1 U19524 ( .B1(P3_LWORD_REG_15__SCAN_IN), .B2(keyinput51), .C1(
        keyinput55), .C2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n16028), .ZN(
        n16031) );
  OAI22_X1 U19525 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(keyinput12), .B1(
        keyinput43), .B2(P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16029) );
  AOI221_X1 U19526 ( .B1(P2_ADDRESS_REG_24__SCAN_IN), .B2(keyinput12), .C1(
        P1_DATAWIDTH_REG_14__SCAN_IN), .C2(keyinput43), .A(n16029), .ZN(n16030) );
  NAND4_X1 U19527 ( .A1(n16033), .A2(n16032), .A3(n16031), .A4(n16030), .ZN(
        n16052) );
  OAI22_X1 U19528 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(keyinput81), .B1(
        P1_EBX_REG_1__SCAN_IN), .B2(keyinput126), .ZN(n16034) );
  AOI221_X1 U19529 ( .B1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(keyinput81), 
        .C1(keyinput126), .C2(P1_EBX_REG_1__SCAN_IN), .A(n16034), .ZN(n16041)
         );
  OAI22_X1 U19530 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(keyinput77), .B1(
        P3_INSTQUEUE_REG_15__4__SCAN_IN), .B2(keyinput112), .ZN(n16035) );
  AOI221_X1 U19531 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(keyinput77), .C1(
        keyinput112), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(n16035), .ZN(
        n16040) );
  OAI22_X1 U19532 ( .A1(P3_MORE_REG_SCAN_IN), .A2(keyinput6), .B1(keyinput121), 
        .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16036) );
  AOI221_X1 U19533 ( .B1(P3_MORE_REG_SCAN_IN), .B2(keyinput6), .C1(
        P3_INSTQUEUE_REG_2__5__SCAN_IN), .C2(keyinput121), .A(n16036), .ZN(
        n16039) );
  OAI22_X1 U19534 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(keyinput79), .B1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput17), .ZN(n16037) );
  AOI221_X1 U19535 ( .B1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B2(keyinput79), 
        .C1(keyinput17), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16037), 
        .ZN(n16038) );
  NAND4_X1 U19536 ( .A1(n16041), .A2(n16040), .A3(n16039), .A4(n16038), .ZN(
        n16051) );
  OAI22_X1 U19537 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(keyinput68), 
        .B1(keyinput26), .B2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16042)
         );
  AOI221_X1 U19538 ( .B1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput68), 
        .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(keyinput26), .A(n16042), 
        .ZN(n16049) );
  OAI22_X1 U19539 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(keyinput39), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(keyinput61), .ZN(n16043) );
  AOI221_X1 U19540 ( .B1(P2_REIP_REG_1__SCAN_IN), .B2(keyinput39), .C1(
        keyinput61), .C2(P1_LWORD_REG_9__SCAN_IN), .A(n16043), .ZN(n16048) );
  OAI22_X1 U19541 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(keyinput114), .B1(
        P1_EAX_REG_5__SCAN_IN), .B2(keyinput72), .ZN(n16044) );
  AOI221_X1 U19542 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(keyinput114), .C1(
        keyinput72), .C2(P1_EAX_REG_5__SCAN_IN), .A(n16044), .ZN(n16047) );
  OAI22_X1 U19543 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(keyinput75), 
        .B1(keyinput42), .B2(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n16045) );
  AOI221_X1 U19544 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput75), 
        .C1(P1_ADDRESS_REG_4__SCAN_IN), .C2(keyinput42), .A(n16045), .ZN(
        n16046) );
  NAND4_X1 U19545 ( .A1(n16049), .A2(n16048), .A3(n16047), .A4(n16046), .ZN(
        n16050) );
  NOR4_X1 U19546 ( .A1(n16053), .A2(n16052), .A3(n16051), .A4(n16050), .ZN(
        n16091) );
  OAI22_X1 U19547 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(keyinput91), .B1(
        keyinput11), .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n16054) );
  AOI221_X1 U19548 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput91), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput11), .A(n16054), .ZN(n16061) );
  OAI22_X1 U19549 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(keyinput54), .B1(
        keyinput23), .B2(P3_UWORD_REG_5__SCAN_IN), .ZN(n16055) );
  AOI221_X1 U19550 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(keyinput54), .C1(
        P3_UWORD_REG_5__SCAN_IN), .C2(keyinput23), .A(n16055), .ZN(n16060) );
  OAI22_X1 U19551 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(keyinput66), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(keyinput36), .ZN(n16056) );
  AOI221_X1 U19552 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(keyinput66), .C1(
        keyinput36), .C2(P2_UWORD_REG_14__SCAN_IN), .A(n16056), .ZN(n16059) );
  OAI22_X1 U19553 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(keyinput21), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput125), .ZN(n16057) );
  AOI221_X1 U19554 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(keyinput21), .C1(
        keyinput125), .C2(P1_READREQUEST_REG_SCAN_IN), .A(n16057), .ZN(n16058)
         );
  NAND4_X1 U19555 ( .A1(n16061), .A2(n16060), .A3(n16059), .A4(n16058), .ZN(
        n16089) );
  OAI22_X1 U19556 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(keyinput95), .B1(
        P2_DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput124), .ZN(n16062) );
  AOI221_X1 U19557 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput95), .C1(
        keyinput124), .C2(P2_DATAWIDTH_REG_13__SCAN_IN), .A(n16062), .ZN(
        n16069) );
  OAI22_X1 U19558 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(keyinput49), 
        .B1(BUF2_REG_9__SCAN_IN), .B2(keyinput25), .ZN(n16063) );
  AOI221_X1 U19559 ( .B1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(keyinput49), 
        .C1(keyinput25), .C2(BUF2_REG_9__SCAN_IN), .A(n16063), .ZN(n16068) );
  OAI22_X1 U19560 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(keyinput80), .B1(
        keyinput18), .B2(P2_BE_N_REG_2__SCAN_IN), .ZN(n16064) );
  AOI221_X1 U19561 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(keyinput80), .C1(
        P2_BE_N_REG_2__SCAN_IN), .C2(keyinput18), .A(n16064), .ZN(n16067) );
  OAI22_X1 U19562 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(keyinput106), 
        .B1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B2(keyinput67), .ZN(n16065) );
  AOI221_X1 U19563 ( .B1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput106), 
        .C1(keyinput67), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(n16065), 
        .ZN(n16066) );
  NAND4_X1 U19564 ( .A1(n16069), .A2(n16068), .A3(n16067), .A4(n16066), .ZN(
        n16088) );
  OAI22_X1 U19565 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(keyinput28), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(keyinput116), .ZN(n16070) );
  AOI221_X1 U19566 ( .B1(P2_EBX_REG_11__SCAN_IN), .B2(keyinput28), .C1(
        keyinput116), .C2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n16070), 
        .ZN(n16077) );
  OAI22_X1 U19567 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput10), .B1(
        P3_DATAO_REG_27__SCAN_IN), .B2(keyinput47), .ZN(n16071) );
  AOI221_X1 U19568 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput10), .C1(
        keyinput47), .C2(P3_DATAO_REG_27__SCAN_IN), .A(n16071), .ZN(n16076) );
  OAI22_X1 U19569 ( .A1(P1_EAX_REG_13__SCAN_IN), .A2(keyinput7), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput86), .ZN(n16072) );
  AOI221_X1 U19570 ( .B1(P1_EAX_REG_13__SCAN_IN), .B2(keyinput7), .C1(
        keyinput86), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n16072), .ZN(
        n16075) );
  OAI22_X1 U19571 ( .A1(READY11_REG_SCAN_IN), .A2(keyinput70), .B1(keyinput108), .B2(P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16073) );
  AOI221_X1 U19572 ( .B1(READY11_REG_SCAN_IN), .B2(keyinput70), .C1(
        P2_DATAWIDTH_REG_2__SCAN_IN), .C2(keyinput108), .A(n16073), .ZN(n16074) );
  NAND4_X1 U19573 ( .A1(n16077), .A2(n16076), .A3(n16075), .A4(n16074), .ZN(
        n16087) );
  OAI22_X1 U19574 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput104), .B1(
        P3_DATAO_REG_28__SCAN_IN), .B2(keyinput84), .ZN(n16078) );
  AOI221_X1 U19575 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput104), .C1(
        keyinput84), .C2(P3_DATAO_REG_28__SCAN_IN), .A(n16078), .ZN(n16085) );
  OAI22_X1 U19576 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(keyinput15), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(keyinput76), .ZN(n16079) );
  AOI221_X1 U19577 ( .B1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B2(keyinput15), 
        .C1(keyinput76), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(n16079), .ZN(
        n16084) );
  OAI22_X1 U19578 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(keyinput20), .B1(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(keyinput56), .ZN(n16080) );
  AOI221_X1 U19579 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(keyinput20), .C1(
        keyinput56), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n16080), .ZN(
        n16083) );
  OAI22_X1 U19580 ( .A1(P2_EBX_REG_3__SCAN_IN), .A2(keyinput119), .B1(
        P2_DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput37), .ZN(n16081) );
  AOI221_X1 U19581 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(keyinput119), .C1(
        keyinput37), .C2(P2_DATAWIDTH_REG_4__SCAN_IN), .A(n16081), .ZN(n16082)
         );
  NAND4_X1 U19582 ( .A1(n16085), .A2(n16084), .A3(n16083), .A4(n16082), .ZN(
        n16086) );
  NOR4_X1 U19583 ( .A1(n16089), .A2(n16088), .A3(n16087), .A4(n16086), .ZN(
        n16090) );
  NAND2_X1 U19584 ( .A1(n16091), .A2(n16090), .ZN(n16092) );
  NOR4_X1 U19585 ( .A1(n16095), .A2(n16094), .A3(n16093), .A4(n16092), .ZN(
        n16109) );
  INV_X1 U19586 ( .A(n16096), .ZN(n16097) );
  NAND2_X1 U19587 ( .A1(n10274), .A2(n16097), .ZN(n16099) );
  AOI21_X1 U19588 ( .B1(n16100), .B2(n16099), .A(n16098), .ZN(n16101) );
  XNOR2_X1 U19589 ( .A(n16101), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17331) );
  INV_X1 U19590 ( .A(n16102), .ZN(n16104) );
  AOI22_X1 U19591 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n16103) );
  OAI21_X1 U19592 ( .B1(n17305), .B2(n16104), .A(n16103), .ZN(n16105) );
  AOI21_X1 U19593 ( .B1(n16106), .B2(n17298), .A(n16105), .ZN(n16107) );
  OAI21_X1 U19594 ( .B1(n17312), .B2(n17331), .A(n16107), .ZN(n16108) );
  XOR2_X1 U19595 ( .A(n16109), .B(n16108), .Z(P1_U2973) );
  AOI22_X1 U19596 ( .A1(n16112), .A2(n16111), .B1(n16110), .B2(n10274), .ZN(
        n16113) );
  NOR2_X1 U19597 ( .A1(n16113), .A2(n16098), .ZN(n16114) );
  XNOR2_X1 U19598 ( .A(n16114), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16201) );
  INV_X1 U19599 ( .A(n16115), .ZN(n16119) );
  AOI22_X1 U19600 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n16116) );
  OAI21_X1 U19601 ( .B1(n17305), .B2(n16117), .A(n16116), .ZN(n16118) );
  AOI21_X1 U19602 ( .B1(n16119), .B2(n17298), .A(n16118), .ZN(n16120) );
  OAI21_X1 U19603 ( .B1(n17312), .B2(n16201), .A(n16120), .ZN(P1_U2974) );
  AOI21_X1 U19604 ( .B1(n16288), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16121), .ZN(n16122) );
  AOI21_X1 U19605 ( .B1(n10274), .B2(n16207), .A(n16122), .ZN(n16124) );
  XNOR2_X1 U19606 ( .A(n10274), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16123) );
  XNOR2_X1 U19607 ( .A(n16124), .B(n16123), .ZN(n17344) );
  INV_X1 U19608 ( .A(n16125), .ZN(n16129) );
  AOI22_X1 U19609 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n16126) );
  OAI21_X1 U19610 ( .B1(n17305), .B2(n16127), .A(n16126), .ZN(n16128) );
  AOI21_X1 U19611 ( .B1(n16129), .B2(n17298), .A(n16128), .ZN(n16130) );
  OAI21_X1 U19612 ( .B1(n17344), .B2(n17312), .A(n16130), .ZN(P1_U2975) );
  XNOR2_X1 U19613 ( .A(n16288), .B(n16207), .ZN(n16131) );
  XNOR2_X1 U19614 ( .A(n16121), .B(n16131), .ZN(n16211) );
  INV_X1 U19615 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21495) );
  NOR2_X1 U19616 ( .A1(n17352), .A2(n21495), .ZN(n16202) );
  AOI21_X1 U19617 ( .B1(n14161), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16202), .ZN(n16132) );
  OAI21_X1 U19618 ( .B1(n17305), .B2(n16133), .A(n16132), .ZN(n16134) );
  AOI21_X1 U19619 ( .B1(n16135), .B2(n17298), .A(n16134), .ZN(n16136) );
  OAI21_X1 U19620 ( .B1(n16211), .B2(n17312), .A(n16136), .ZN(P1_U2976) );
  NAND2_X1 U19621 ( .A1(n16137), .A2(n10274), .ZN(n16234) );
  INV_X1 U19622 ( .A(n11281), .ZN(n16139) );
  INV_X1 U19623 ( .A(n16138), .ZN(n16252) );
  NAND3_X1 U19624 ( .A1(n16139), .A2(n16253), .A3(n16252), .ZN(n16233) );
  NAND2_X1 U19625 ( .A1(n16234), .A2(n16233), .ZN(n16140) );
  XNOR2_X1 U19626 ( .A(n16140), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16251) );
  INV_X1 U19627 ( .A(n16141), .ZN(n16144) );
  INV_X1 U19628 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n16142) );
  NOR2_X1 U19629 ( .A1(n17352), .A2(n16142), .ZN(n16247) );
  AOI21_X1 U19630 ( .B1(n14161), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16247), .ZN(n16143) );
  OAI21_X1 U19631 ( .B1(n17305), .B2(n16144), .A(n16143), .ZN(n16145) );
  AOI21_X1 U19632 ( .B1(n16146), .B2(n17298), .A(n16145), .ZN(n16147) );
  OAI21_X1 U19633 ( .B1(n17312), .B2(n16251), .A(n16147), .ZN(P1_U2979) );
  OAI21_X1 U19634 ( .B1(n11281), .B2(n16149), .A(n16148), .ZN(n16271) );
  NAND2_X1 U19635 ( .A1(n17225), .A2(n17298), .ZN(n16154) );
  INV_X1 U19636 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n16150) );
  NOR2_X1 U19637 ( .A1(n17352), .A2(n16150), .ZN(n16266) );
  INV_X1 U19638 ( .A(n17221), .ZN(n16151) );
  NOR2_X1 U19639 ( .A1(n17305), .A2(n16151), .ZN(n16152) );
  AOI211_X1 U19640 ( .C1(n14161), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16266), .B(n16152), .ZN(n16153) );
  OAI211_X1 U19641 ( .C1(n17312), .C2(n16271), .A(n16154), .B(n16153), .ZN(
        P1_U2981) );
  INV_X1 U19642 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U19643 ( .A1(n16288), .A2(n17353), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n10274), .ZN(n16161) );
  NOR2_X1 U19644 ( .A1(n16156), .A2(n16155), .ZN(n16273) );
  INV_X1 U19645 ( .A(n16157), .ZN(n16159) );
  OAI21_X1 U19646 ( .B1(n16273), .B2(n16159), .A(n16158), .ZN(n16160) );
  XOR2_X1 U19647 ( .A(n16161), .B(n16160), .Z(n17356) );
  AOI22_X1 U19648 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16162) );
  OAI21_X1 U19649 ( .B1(n17305), .B2(n16163), .A(n16162), .ZN(n16164) );
  AOI21_X1 U19650 ( .B1(n16165), .B2(n17298), .A(n16164), .ZN(n16166) );
  OAI21_X1 U19651 ( .B1(n17312), .B2(n17356), .A(n16166), .ZN(P1_U2985) );
  NOR3_X1 U19652 ( .A1(n16167), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n10274), .ZN(n16168) );
  NOR2_X1 U19653 ( .A1(n16169), .A2(n16168), .ZN(n16170) );
  XOR2_X1 U19654 ( .A(n11273), .B(n16170), .Z(n17377) );
  NAND2_X1 U19655 ( .A1(n17377), .A2(n17267), .ZN(n16175) );
  INV_X1 U19656 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n16171) );
  NOR2_X1 U19657 ( .A1(n17352), .A2(n16171), .ZN(n17373) );
  NOR2_X1 U19658 ( .A1(n17305), .A2(n16172), .ZN(n16173) );
  AOI211_X1 U19659 ( .C1(n14161), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17373), .B(n16173), .ZN(n16174) );
  OAI211_X1 U19660 ( .C1(n17306), .C2(n16176), .A(n16175), .B(n16174), .ZN(
        P1_U2988) );
  INV_X1 U19661 ( .A(n16177), .ZN(n16186) );
  NAND2_X1 U19662 ( .A1(n16179), .A2(n16178), .ZN(n16183) );
  OAI21_X1 U19663 ( .B1(n16181), .B2(n17364), .A(n16180), .ZN(n16182) );
  AOI21_X1 U19664 ( .B1(n16184), .B2(n16183), .A(n16182), .ZN(n16185) );
  OAI21_X1 U19665 ( .B1(n16186), .B2(n17365), .A(n16185), .ZN(P1_U3001) );
  INV_X1 U19666 ( .A(n16187), .ZN(n17326) );
  NOR2_X1 U19667 ( .A1(n16188), .A2(n17364), .ZN(n16190) );
  AOI211_X1 U19668 ( .C1(n17326), .C2(n16191), .A(n16190), .B(n16189), .ZN(
        n16193) );
  NAND2_X1 U19669 ( .A1(n17321), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16192) );
  OAI211_X1 U19670 ( .C1(n16194), .C2(n17365), .A(n16193), .B(n16192), .ZN(
        P1_U3004) );
  NAND2_X1 U19671 ( .A1(n17369), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16195) );
  OAI221_X1 U19672 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17335), 
        .C1(n16197), .C2(n16196), .A(n16195), .ZN(n16198) );
  AOI21_X1 U19673 ( .B1(n16199), .B2(n21427), .A(n16198), .ZN(n16200) );
  OAI21_X1 U19674 ( .B1(n16201), .B2(n17365), .A(n16200), .ZN(P1_U3006) );
  AOI21_X1 U19675 ( .B1(n16203), .B2(n21427), .A(n16202), .ZN(n16206) );
  NOR2_X1 U19676 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n16204), .ZN(
        n17342) );
  NAND2_X1 U19677 ( .A1(n17375), .A2(n17342), .ZN(n16205) );
  OAI211_X1 U19678 ( .C1(n16208), .C2(n16207), .A(n16206), .B(n16205), .ZN(
        n16209) );
  INV_X1 U19679 ( .A(n16209), .ZN(n16210) );
  OAI21_X1 U19680 ( .B1(n16211), .B2(n17365), .A(n16210), .ZN(P1_U3008) );
  INV_X1 U19681 ( .A(n16212), .ZN(n16213) );
  NOR2_X1 U19682 ( .A1(n16214), .A2(n16213), .ZN(n16215) );
  XNOR2_X1 U19683 ( .A(n16215), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17261) );
  INV_X1 U19684 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n16224) );
  NAND2_X1 U19685 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16216), .ZN(
        n16217) );
  OAI22_X1 U19686 ( .A1(n16220), .A2(n16219), .B1(n16218), .B2(n16217), .ZN(
        n16243) );
  AOI21_X1 U19687 ( .B1(n21432), .B2(n16221), .A(n16243), .ZN(n17372) );
  NOR3_X1 U19688 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17372), .A3(
        n16222), .ZN(n16237) );
  OAI21_X1 U19689 ( .B1(n16239), .B2(n16237), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16223) );
  OAI21_X1 U19690 ( .B1(n17352), .B2(n16224), .A(n16223), .ZN(n16225) );
  AOI21_X1 U19691 ( .B1(n17194), .B2(n21427), .A(n16225), .ZN(n16232) );
  INV_X1 U19692 ( .A(n17372), .ZN(n16226) );
  NAND2_X1 U19693 ( .A1(n16227), .A2(n16226), .ZN(n16257) );
  INV_X1 U19694 ( .A(n16257), .ZN(n16230) );
  NAND4_X1 U19695 ( .A1(n16230), .A2(n16229), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(n16228), .ZN(n16231) );
  OAI211_X1 U19696 ( .C1(n17261), .C2(n17365), .A(n16232), .B(n16231), .ZN(
        P1_U3009) );
  AOI22_X1 U19697 ( .A1(n16234), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n11282), .B2(n16233), .ZN(n16236) );
  XNOR2_X1 U19698 ( .A(n16236), .B(n16235), .ZN(n17262) );
  INV_X1 U19699 ( .A(n17262), .ZN(n16241) );
  OAI22_X1 U19700 ( .A1(n17204), .A2(n17364), .B1(n17352), .B2(n21492), .ZN(
        n16238) );
  AOI211_X1 U19701 ( .C1(n16239), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16238), .B(n16237), .ZN(n16240) );
  OAI21_X1 U19702 ( .B1(n16241), .B2(n17365), .A(n16240), .ZN(P1_U3010) );
  NAND2_X1 U19703 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16242) );
  OAI21_X1 U19704 ( .B1(n16243), .B2(n21432), .A(n16242), .ZN(n16244) );
  NAND2_X1 U19705 ( .A1(n16244), .A2(n16256), .ZN(n16249) );
  OAI21_X1 U19706 ( .B1(n16253), .B2(n16257), .A(n11282), .ZN(n16248) );
  NOR2_X1 U19707 ( .A1(n16245), .A2(n17364), .ZN(n16246) );
  AOI211_X1 U19708 ( .C1(n16249), .C2(n16248), .A(n16247), .B(n16246), .ZN(
        n16250) );
  OAI21_X1 U19709 ( .B1(n16251), .B2(n17365), .A(n16250), .ZN(P1_U3011) );
  MUX2_X1 U19710 ( .A(n10274), .B(n16252), .S(n16148), .Z(n16254) );
  XNOR2_X1 U19711 ( .A(n16254), .B(n16253), .ZN(n17268) );
  INV_X1 U19712 ( .A(n17268), .ZN(n16261) );
  INV_X1 U19713 ( .A(n17220), .ZN(n16259) );
  NAND2_X1 U19714 ( .A1(n17369), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n16255) );
  OAI221_X1 U19715 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16257), 
        .C1(n16253), .C2(n16256), .A(n16255), .ZN(n16258) );
  AOI21_X1 U19716 ( .B1(n16259), .B2(n21427), .A(n16258), .ZN(n16260) );
  OAI21_X1 U19717 ( .B1(n16261), .B2(n17365), .A(n16260), .ZN(P1_U3012) );
  OAI21_X1 U19718 ( .B1(n17353), .B2(n17368), .A(n16262), .ZN(n16307) );
  OAI21_X1 U19719 ( .B1(n16263), .B2(n16267), .A(n16307), .ZN(n16281) );
  INV_X1 U19720 ( .A(n17224), .ZN(n16264) );
  NOR2_X1 U19721 ( .A1(n17364), .A2(n16264), .ZN(n16265) );
  AOI211_X1 U19722 ( .C1(n16281), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16266), .B(n16265), .ZN(n16270) );
  NAND3_X1 U19723 ( .A1(n17355), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17354), .ZN(n16302) );
  NOR2_X1 U19724 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16302), .ZN(
        n16268) );
  NAND2_X1 U19725 ( .A1(n16268), .A2(n16267), .ZN(n16269) );
  OAI211_X1 U19726 ( .C1(n16271), .C2(n17365), .A(n16270), .B(n16269), .ZN(
        P1_U3013) );
  AOI21_X1 U19727 ( .B1(n16274), .B2(n16273), .A(n16272), .ZN(n16276) );
  NOR2_X1 U19728 ( .A1(n10274), .A2(n16276), .ZN(n16275) );
  AOI22_X1 U19729 ( .A1(n10274), .A2(n16276), .B1(n16296), .B2(n16275), .ZN(
        n16277) );
  XNOR2_X1 U19730 ( .A(n16280), .B(n16277), .ZN(n17277) );
  XOR2_X1 U19731 ( .A(n16279), .B(n16278), .Z(n17251) );
  AOI22_X1 U19732 ( .A1(n17251), .A2(n21427), .B1(n17369), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16284) );
  OAI21_X1 U19733 ( .B1(n16300), .B2(n16302), .A(n16280), .ZN(n16282) );
  NAND2_X1 U19734 ( .A1(n16282), .A2(n16281), .ZN(n16283) );
  OAI211_X1 U19735 ( .C1(n17277), .C2(n17365), .A(n16284), .B(n16283), .ZN(
        P1_U3014) );
  NOR2_X1 U19736 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16293) );
  OR2_X1 U19737 ( .A1(n16285), .A2(n15343), .ZN(n16287) );
  AND2_X1 U19738 ( .A1(n16287), .A2(n16286), .ZN(n16309) );
  INV_X1 U19739 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16315) );
  MUX2_X1 U19740 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n16315), .S(
        n16288), .Z(n16308) );
  NOR2_X1 U19741 ( .A1(n16293), .A2(n16311), .ZN(n16292) );
  INV_X1 U19742 ( .A(n16289), .ZN(n16290) );
  OAI22_X1 U19743 ( .A1(n16292), .A2(n16291), .B1(n16311), .B2(n16290), .ZN(
        n17282) );
  NOR2_X1 U19744 ( .A1(n16293), .A2(n16302), .ZN(n16299) );
  INV_X1 U19745 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n16294) );
  OAI22_X1 U19746 ( .A1(n17364), .A2(n16295), .B1(n17352), .B2(n16294), .ZN(
        n16298) );
  NOR2_X1 U19747 ( .A1(n16307), .A2(n16296), .ZN(n16297) );
  AOI211_X1 U19748 ( .C1(n16300), .C2(n16299), .A(n16298), .B(n16297), .ZN(
        n16301) );
  OAI21_X1 U19749 ( .B1(n17282), .B2(n17365), .A(n16301), .ZN(P1_U3015) );
  INV_X1 U19750 ( .A(n16302), .ZN(n16314) );
  INV_X1 U19751 ( .A(n16303), .ZN(n16305) );
  NOR2_X1 U19752 ( .A1(n17352), .A2(n21484), .ZN(n16304) );
  AOI21_X1 U19753 ( .B1(n21427), .B2(n16305), .A(n16304), .ZN(n16306) );
  OAI21_X1 U19754 ( .B1(n16307), .B2(n16315), .A(n16306), .ZN(n16313) );
  NOR2_X1 U19755 ( .A1(n16309), .A2(n16308), .ZN(n16310) );
  NOR2_X1 U19756 ( .A1(n16311), .A2(n16310), .ZN(n17287) );
  NOR2_X1 U19757 ( .A1(n17287), .A2(n17365), .ZN(n16312) );
  AOI211_X1 U19758 ( .C1(n16315), .C2(n16314), .A(n16313), .B(n16312), .ZN(
        n16316) );
  INV_X1 U19759 ( .A(n16316), .ZN(P1_U3016) );
  NOR2_X1 U19760 ( .A1(n9830), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16317) );
  OAI22_X1 U19761 ( .A1(n16324), .A2(n16317), .B1(n13865), .B2(n16332), .ZN(
        n16318) );
  MUX2_X1 U19762 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n16318), .S(
        n21436), .Z(P1_U3477) );
  INV_X1 U19763 ( .A(n16319), .ZN(n16321) );
  NAND2_X1 U19764 ( .A1(n16321), .A2(n16320), .ZN(n16323) );
  MUX2_X1 U19765 ( .A(n16324), .B(n16323), .S(n16322), .Z(n16325) );
  OAI21_X1 U19766 ( .B1(n16332), .B2(n16326), .A(n16325), .ZN(n16327) );
  MUX2_X1 U19767 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n16327), .S(
        n21436), .Z(P1_U3476) );
  NOR2_X1 U19768 ( .A1(n14202), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16329) );
  NOR4_X1 U19769 ( .A1(n16331), .A2(n16330), .A3(n16329), .A4(n16328), .ZN(
        n16335) );
  OAI22_X1 U19770 ( .A1(n16335), .A2(n16334), .B1(n16333), .B2(n16332), .ZN(
        n16336) );
  MUX2_X1 U19771 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n16336), .S(
        n21436), .Z(P1_U3475) );
  INV_X1 U19772 ( .A(n16337), .ZN(n16357) );
  AOI22_X1 U19773 ( .A1(n16357), .A2(n16339), .B1(n16355), .B2(n16338), .ZN(
        n16345) );
  NAND2_X1 U19774 ( .A1(n16358), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n16344) );
  NAND2_X1 U19775 ( .A1(n16340), .A2(n16359), .ZN(n16343) );
  NAND2_X1 U19776 ( .A1(n16341), .A2(n16361), .ZN(n16342) );
  NAND4_X1 U19777 ( .A1(n16345), .A2(n16344), .A3(n16343), .A4(n16342), .ZN(
        P1_U3154) );
  AOI22_X1 U19778 ( .A1(n16357), .A2(n16347), .B1(n16355), .B2(n16346), .ZN(
        n16353) );
  NAND2_X1 U19779 ( .A1(n16358), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n16352) );
  NAND2_X1 U19780 ( .A1(n16348), .A2(n16359), .ZN(n16351) );
  NAND2_X1 U19781 ( .A1(n16349), .A2(n16361), .ZN(n16350) );
  NAND4_X1 U19782 ( .A1(n16353), .A2(n16352), .A3(n16351), .A4(n16350), .ZN(
        P1_U3157) );
  AOI22_X1 U19783 ( .A1(n16357), .A2(n16356), .B1(n16355), .B2(n16354), .ZN(
        n16366) );
  NAND2_X1 U19784 ( .A1(n16358), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n16365) );
  NAND2_X1 U19785 ( .A1(n16360), .A2(n16359), .ZN(n16364) );
  NAND2_X1 U19786 ( .A1(n16362), .A2(n16361), .ZN(n16363) );
  NAND4_X1 U19787 ( .A1(n16366), .A2(n16365), .A3(n16364), .A4(n16363), .ZN(
        P1_U3159) );
  NAND4_X1 U19788 ( .A1(n17402), .A2(n20370), .A3(n15196), .A4(n16367), .ZN(
        n16374) );
  AOI22_X1 U19789 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n20412), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n20406), .ZN(n16368) );
  INV_X1 U19790 ( .A(n16368), .ZN(n16371) );
  INV_X1 U19791 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n17464) );
  OAI22_X1 U19792 ( .A1(n16369), .A2(n20401), .B1(n17464), .B2(n20396), .ZN(
        n16370) );
  AOI211_X1 U19793 ( .C1(n16372), .C2(n20328), .A(n16371), .B(n16370), .ZN(
        n16373) );
  OAI211_X1 U19794 ( .C1(n17465), .C2(n20402), .A(n16374), .B(n16373), .ZN(
        P2_U2824) );
  XOR2_X1 U19795 ( .A(n16376), .B(n16389), .Z(n16806) );
  INV_X1 U19796 ( .A(n16806), .ZN(n16544) );
  NAND2_X1 U19797 ( .A1(n16393), .A2(n16377), .ZN(n16378) );
  NAND2_X1 U19798 ( .A1(n16379), .A2(n16378), .ZN(n16803) );
  INV_X1 U19799 ( .A(n16803), .ZN(n16464) );
  NAND2_X1 U19800 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n20359), .ZN(n16380) );
  OAI211_X1 U19801 ( .C1(n16638), .C2(n20380), .A(n20347), .B(n16380), .ZN(
        n16381) );
  AOI21_X1 U19802 ( .B1(n20328), .B2(n16382), .A(n16381), .ZN(n16383) );
  OAI21_X1 U19803 ( .B1(n21141), .B2(n20374), .A(n16383), .ZN(n16387) );
  AOI211_X1 U19804 ( .C1(n16640), .C2(n16385), .A(n16384), .B(n21086), .ZN(
        n16386) );
  AOI211_X1 U19805 ( .C1(n16464), .C2(n20385), .A(n16387), .B(n16386), .ZN(
        n16388) );
  OAI21_X1 U19806 ( .B1(n16544), .B2(n20401), .A(n16388), .ZN(P2_U2836) );
  AOI21_X1 U19807 ( .B1(n16390), .B2(n13641), .A(n16375), .ZN(n17497) );
  INV_X1 U19808 ( .A(n17497), .ZN(n16403) );
  OR2_X1 U19809 ( .A1(n13643), .A2(n16391), .ZN(n16392) );
  NAND2_X1 U19810 ( .A1(n16393), .A2(n16392), .ZN(n17480) );
  AOI22_X1 U19811 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n20412), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n20406), .ZN(n16394) );
  NAND2_X1 U19812 ( .A1(n20347), .A2(n16394), .ZN(n16395) );
  AOI21_X1 U19813 ( .B1(n20359), .B2(P2_EBX_REG_18__SCAN_IN), .A(n16395), .ZN(
        n16396) );
  OAI21_X1 U19814 ( .B1(n17480), .B2(n20402), .A(n16396), .ZN(n16400) );
  AOI211_X1 U19815 ( .C1(n16652), .C2(n16398), .A(n16397), .B(n21086), .ZN(
        n16399) );
  AOI211_X1 U19816 ( .C1(n16401), .C2(n20328), .A(n16400), .B(n16399), .ZN(
        n16402) );
  OAI21_X1 U19817 ( .B1(n16403), .B2(n20401), .A(n16402), .ZN(P2_U2837) );
  NAND2_X1 U19818 ( .A1(n16405), .A2(n16404), .ZN(n16406) );
  NAND2_X1 U19819 ( .A1(n12523), .A2(n16406), .ZN(n17409) );
  OR2_X1 U19820 ( .A1(n16408), .A2(n16407), .ZN(n16471) );
  NAND3_X1 U19821 ( .A1(n16471), .A2(n16409), .A3(n20435), .ZN(n16411) );
  NAND2_X1 U19822 ( .A1(n17479), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16410) );
  OAI211_X1 U19823 ( .C1(n17479), .C2(n17409), .A(n16411), .B(n16410), .ZN(
        P2_U2858) );
  INV_X1 U19824 ( .A(n16412), .ZN(n16414) );
  XNOR2_X1 U19825 ( .A(n16416), .B(n16415), .ZN(n16486) );
  NOR2_X1 U19826 ( .A1(n17417), .A2(n17479), .ZN(n16417) );
  AOI21_X1 U19827 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n17479), .A(n16417), .ZN(
        n16418) );
  OAI21_X1 U19828 ( .B1(n16486), .B2(n20428), .A(n16418), .ZN(P2_U2859) );
  OAI21_X1 U19830 ( .B1(n9870), .B2(n16421), .A(n16420), .ZN(n16492) );
  NOR2_X1 U19831 ( .A1(n16554), .A2(n17479), .ZN(n16422) );
  AOI21_X1 U19832 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n17479), .A(n16422), .ZN(
        n16423) );
  OAI21_X1 U19833 ( .B1(n16492), .B2(n20428), .A(n16423), .ZN(P2_U2860) );
  CLKBUF_X1 U19834 ( .A(n16424), .Z(n16427) );
  OAI21_X1 U19835 ( .B1(n16427), .B2(n16426), .A(n16425), .ZN(n16500) );
  OR2_X1 U19836 ( .A1(n16437), .A2(n16428), .ZN(n16429) );
  NAND2_X1 U19837 ( .A1(n12876), .A2(n16429), .ZN(n17429) );
  NOR2_X1 U19838 ( .A1(n17429), .A2(n17479), .ZN(n16430) );
  AOI21_X1 U19839 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n17479), .A(n16430), .ZN(
        n16431) );
  OAI21_X1 U19840 ( .B1(n16500), .B2(n20428), .A(n16431), .ZN(P2_U2861) );
  OAI21_X1 U19841 ( .B1(n16432), .B2(n16434), .A(n16433), .ZN(n16509) );
  NOR2_X1 U19842 ( .A1(n16448), .A2(n16435), .ZN(n16436) );
  OR2_X1 U19843 ( .A1(n16437), .A2(n16436), .ZN(n16740) );
  NOR2_X1 U19844 ( .A1(n16740), .A2(n17479), .ZN(n16438) );
  AOI21_X1 U19845 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n17479), .A(n16438), .ZN(
        n16439) );
  OAI21_X1 U19846 ( .B1(n16509), .B2(n20428), .A(n16439), .ZN(P2_U2862) );
  AOI21_X1 U19847 ( .B1(n16440), .B2(n16443), .A(n16442), .ZN(n16444) );
  XOR2_X1 U19848 ( .A(n16445), .B(n16444), .Z(n16518) );
  AND2_X1 U19849 ( .A1(n16447), .A2(n16446), .ZN(n16449) );
  OR2_X1 U19850 ( .A1(n16449), .A2(n16448), .ZN(n17454) );
  NOR2_X1 U19851 ( .A1(n17454), .A2(n17479), .ZN(n16450) );
  AOI21_X1 U19852 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n17479), .A(n16450), .ZN(
        n16451) );
  OAI21_X1 U19853 ( .B1(n16518), .B2(n20428), .A(n16451), .ZN(P2_U2863) );
  OR2_X1 U19854 ( .A1(n16455), .A2(n16456), .ZN(n16457) );
  AND2_X1 U19855 ( .A1(n16453), .A2(n16457), .ZN(n16534) );
  NAND2_X1 U19856 ( .A1(n16534), .A2(n20435), .ZN(n16460) );
  INV_X1 U19857 ( .A(n16790), .ZN(n16458) );
  NAND2_X1 U19858 ( .A1(n16458), .A2(n13216), .ZN(n16459) );
  OAI211_X1 U19859 ( .C1(n13216), .C2(n11916), .A(n16460), .B(n16459), .ZN(
        P2_U2866) );
  NAND2_X1 U19860 ( .A1(n16461), .A2(n16462), .ZN(n16463) );
  AND2_X1 U19861 ( .A1(n9901), .A2(n16463), .ZN(n16541) );
  NAND2_X1 U19862 ( .A1(n16541), .A2(n20435), .ZN(n16466) );
  NAND2_X1 U19863 ( .A1(n16464), .A2(n13216), .ZN(n16465) );
  OAI211_X1 U19864 ( .C1(n20437), .C2(n16467), .A(n16466), .B(n16465), .ZN(
        P2_U2868) );
  MUX2_X1 U19865 ( .A(n16659), .B(n16468), .S(n17479), .Z(n16469) );
  OAI21_X1 U19866 ( .B1(n16470), .B2(n20428), .A(n16469), .ZN(P2_U2870) );
  NAND3_X1 U19867 ( .A1(n16471), .A2(n16409), .A3(n20477), .ZN(n16480) );
  NOR2_X1 U19868 ( .A1(n12578), .A2(n16472), .ZN(n16473) );
  INV_X1 U19869 ( .A(n17414), .ZN(n16477) );
  OAI22_X1 U19870 ( .A1(n16523), .A2(n20456), .B1(n20475), .B2(n16475), .ZN(
        n16476) );
  AOI21_X1 U19871 ( .B1(n20492), .B2(n16477), .A(n16476), .ZN(n16479) );
  AOI22_X1 U19872 ( .A1(n20444), .A2(BUF2_REG_29__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n16478) );
  NAND3_X1 U19873 ( .A1(n16480), .A2(n16479), .A3(n16478), .ZN(P2_U2890) );
  INV_X1 U19874 ( .A(n17416), .ZN(n16483) );
  OAI22_X1 U19875 ( .A1(n16523), .A2(n20459), .B1(n20475), .B2(n16481), .ZN(
        n16482) );
  AOI21_X1 U19876 ( .B1(n20492), .B2(n16483), .A(n16482), .ZN(n16485) );
  AOI22_X1 U19877 ( .A1(n20444), .A2(BUF2_REG_28__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16484) );
  OAI211_X1 U19878 ( .C1(n16486), .C2(n20496), .A(n16485), .B(n16484), .ZN(
        P2_U2891) );
  OAI22_X1 U19879 ( .A1(n16523), .A2(n20461), .B1(n20475), .B2(n16487), .ZN(
        n16488) );
  AOI21_X1 U19880 ( .B1(n20492), .B2(n16489), .A(n16488), .ZN(n16491) );
  AOI22_X1 U19881 ( .A1(n20444), .A2(BUF2_REG_27__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16490) );
  OAI211_X1 U19882 ( .C1(n16492), .C2(n20496), .A(n16491), .B(n16490), .ZN(
        P2_U2892) );
  NAND2_X1 U19883 ( .A1(n16503), .A2(n16493), .ZN(n16494) );
  AND2_X1 U19884 ( .A1(n9864), .A2(n16494), .ZN(n17430) );
  INV_X1 U19885 ( .A(n20463), .ZN(n16496) );
  OAI22_X1 U19886 ( .A1(n16523), .A2(n16496), .B1(n20475), .B2(n16495), .ZN(
        n16497) );
  AOI21_X1 U19887 ( .B1(n20492), .B2(n17430), .A(n16497), .ZN(n16499) );
  AOI22_X1 U19888 ( .A1(n20444), .A2(BUF2_REG_26__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16498) );
  OAI211_X1 U19889 ( .C1(n16500), .C2(n20496), .A(n16499), .B(n16498), .ZN(
        P2_U2893) );
  NAND2_X1 U19890 ( .A1(n16513), .A2(n16501), .ZN(n16502) );
  NAND2_X1 U19891 ( .A1(n16503), .A2(n16502), .ZN(n17451) );
  INV_X1 U19892 ( .A(n17451), .ZN(n16506) );
  OAI22_X1 U19893 ( .A1(n16523), .A2(n20466), .B1(n20475), .B2(n16504), .ZN(
        n16505) );
  AOI21_X1 U19894 ( .B1(n20492), .B2(n16506), .A(n16505), .ZN(n16508) );
  AOI22_X1 U19895 ( .A1(n20444), .A2(BUF2_REG_25__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n16507) );
  OAI211_X1 U19896 ( .C1(n16509), .C2(n20496), .A(n16508), .B(n16507), .ZN(
        P2_U2894) );
  OR2_X1 U19897 ( .A1(n16511), .A2(n16510), .ZN(n16512) );
  AND2_X1 U19898 ( .A1(n16513), .A2(n16512), .ZN(n17452) );
  INV_X1 U19899 ( .A(n20469), .ZN(n16514) );
  OAI22_X1 U19900 ( .A1(n16523), .A2(n16514), .B1(n20475), .B2(n13844), .ZN(
        n16515) );
  AOI21_X1 U19901 ( .B1(n20492), .B2(n17452), .A(n16515), .ZN(n16517) );
  AOI22_X1 U19902 ( .A1(n20444), .A2(BUF2_REG_24__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16516) );
  OAI211_X1 U19903 ( .C1(n16518), .C2(n20496), .A(n16517), .B(n16516), .ZN(
        P2_U2895) );
  AOI21_X1 U19904 ( .B1(n16519), .B2(n16521), .A(n16520), .ZN(n17466) );
  INV_X1 U19905 ( .A(n17466), .ZN(n16528) );
  INV_X1 U19906 ( .A(n16766), .ZN(n16525) );
  OAI22_X1 U19907 ( .A1(n16523), .A2(n20576), .B1(n20475), .B2(n16522), .ZN(
        n16524) );
  AOI21_X1 U19908 ( .B1(n20492), .B2(n16525), .A(n16524), .ZN(n16527) );
  AOI22_X1 U19909 ( .A1(n20444), .A2(BUF2_REG_23__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16526) );
  OAI211_X1 U19910 ( .C1(n16528), .C2(n20496), .A(n16527), .B(n16526), .ZN(
        P2_U2896) );
  NAND2_X1 U19911 ( .A1(n20443), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16532) );
  NAND2_X1 U19912 ( .A1(n20444), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16531) );
  AOI22_X1 U19913 ( .A1(n20442), .A2(n16529), .B1(n20491), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16530) );
  NAND3_X1 U19914 ( .A1(n16532), .A2(n16531), .A3(n16530), .ZN(n16533) );
  AOI21_X1 U19915 ( .B1(n16534), .B2(n20477), .A(n16533), .ZN(n16535) );
  OAI21_X1 U19916 ( .B1(n16794), .B2(n16543), .A(n16535), .ZN(P2_U2898) );
  NAND2_X1 U19917 ( .A1(n20443), .A2(BUF1_REG_19__SCAN_IN), .ZN(n16539) );
  NAND2_X1 U19918 ( .A1(n20444), .A2(BUF2_REG_19__SCAN_IN), .ZN(n16538) );
  AOI22_X1 U19919 ( .A1(n20442), .A2(n16536), .B1(n20491), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16537) );
  NAND3_X1 U19920 ( .A1(n16539), .A2(n16538), .A3(n16537), .ZN(n16540) );
  AOI21_X1 U19921 ( .B1(n16541), .B2(n20477), .A(n16540), .ZN(n16542) );
  OAI21_X1 U19922 ( .B1(n16544), .B2(n16543), .A(n16542), .ZN(P2_U2900) );
  NAND2_X1 U19923 ( .A1(n16546), .A2(n16545), .ZN(n16548) );
  XOR2_X1 U19924 ( .A(n16548), .B(n9798), .Z(n16728) );
  AOI21_X1 U19925 ( .B1(n16717), .B2(n12559), .A(n12519), .ZN(n16726) );
  NAND2_X1 U19926 ( .A1(n20376), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16720) );
  OAI21_X1 U19927 ( .B1(n17596), .B2(n16549), .A(n16720), .ZN(n16550) );
  AOI21_X1 U19928 ( .B1(n17582), .B2(n17403), .A(n16550), .ZN(n16551) );
  OAI21_X1 U19929 ( .B1(n17409), .B2(n17577), .A(n16551), .ZN(n16552) );
  AOI21_X1 U19930 ( .B1(n16726), .B2(n12599), .A(n16552), .ZN(n16553) );
  OAI21_X1 U19931 ( .B1(n16728), .B2(n17572), .A(n16553), .ZN(P2_U2985) );
  NAND2_X1 U19932 ( .A1(n17582), .A2(n16555), .ZN(n16557) );
  OAI211_X1 U19933 ( .C1(n17596), .C2(n16558), .A(n16557), .B(n16556), .ZN(
        n16561) );
  NOR3_X1 U19934 ( .A1(n16559), .A2(n12558), .A3(n17566), .ZN(n16560) );
  AOI211_X1 U19935 ( .C1(n17591), .C2(n12879), .A(n16561), .B(n16560), .ZN(
        n16562) );
  OAI21_X1 U19936 ( .B1(n16563), .B2(n17572), .A(n16562), .ZN(P2_U2987) );
  INV_X1 U19937 ( .A(n16577), .ZN(n16565) );
  AOI21_X1 U19938 ( .B1(n16564), .B2(n16576), .A(n16565), .ZN(n16567) );
  MUX2_X1 U19939 ( .A(n16567), .B(n16576), .S(n16566), .Z(n16569) );
  NAND2_X1 U19940 ( .A1(n16569), .A2(n16568), .ZN(n16739) );
  INV_X1 U19941 ( .A(n16580), .ZN(n16570) );
  AOI21_X1 U19942 ( .B1(n16729), .B2(n16570), .A(n9865), .ZN(n16737) );
  NOR2_X1 U19943 ( .A1(n17429), .A2(n17577), .ZN(n16574) );
  NAND2_X1 U19944 ( .A1(n20376), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16731) );
  NAND2_X1 U19945 ( .A1(n17564), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16571) );
  OAI211_X1 U19946 ( .C1(n17571), .C2(n16572), .A(n16731), .B(n16571), .ZN(
        n16573) );
  AOI211_X1 U19947 ( .C1(n16737), .C2(n12599), .A(n16574), .B(n16573), .ZN(
        n16575) );
  OAI21_X1 U19948 ( .B1(n17572), .B2(n16739), .A(n16575), .ZN(P2_U2988) );
  NAND2_X1 U19949 ( .A1(n16577), .A2(n16576), .ZN(n16578) );
  XNOR2_X1 U19950 ( .A(n16564), .B(n16578), .ZN(n16751) );
  AOI21_X1 U19951 ( .B1(n16747), .B2(n16579), .A(n16580), .ZN(n16749) );
  NAND2_X1 U19952 ( .A1(n20376), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16741) );
  OAI21_X1 U19953 ( .B1(n17596), .B2(n16581), .A(n16741), .ZN(n16582) );
  AOI21_X1 U19954 ( .B1(n17582), .B2(n17447), .A(n16582), .ZN(n16583) );
  OAI21_X1 U19955 ( .B1(n16740), .B2(n17577), .A(n16583), .ZN(n16584) );
  AOI21_X1 U19956 ( .B1(n16749), .B2(n12599), .A(n16584), .ZN(n16585) );
  OAI21_X1 U19957 ( .B1(n17572), .B2(n16751), .A(n16585), .ZN(P2_U2989) );
  INV_X1 U19958 ( .A(n16586), .ZN(n16587) );
  OAI21_X1 U19959 ( .B1(n16587), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16579), .ZN(n16761) );
  XNOR2_X1 U19960 ( .A(n16589), .B(n16754), .ZN(n16590) );
  XNOR2_X1 U19961 ( .A(n9809), .B(n16590), .ZN(n16759) );
  OAI22_X1 U19962 ( .A1(n12471), .A2(n20347), .B1(n17571), .B2(n16591), .ZN(
        n16592) );
  AOI21_X1 U19963 ( .B1(n17564), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16592), .ZN(n16593) );
  OAI21_X1 U19964 ( .B1(n17454), .B2(n17577), .A(n16593), .ZN(n16594) );
  AOI21_X1 U19965 ( .B1(n16759), .B2(n17592), .A(n16594), .ZN(n16595) );
  OAI21_X1 U19966 ( .B1(n16761), .B2(n17566), .A(n16595), .ZN(P2_U2990) );
  INV_X1 U19967 ( .A(n16596), .ZN(n16610) );
  NOR2_X1 U19968 ( .A1(n16610), .A2(n16776), .ZN(n16609) );
  OAI21_X1 U19969 ( .B1(n16609), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16586), .ZN(n16772) );
  XOR2_X1 U19970 ( .A(n16597), .B(n16598), .Z(n16769) );
  NAND2_X1 U19971 ( .A1(n20376), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16765) );
  OAI21_X1 U19972 ( .B1(n17596), .B2(n16599), .A(n16765), .ZN(n16600) );
  AOI21_X1 U19973 ( .B1(n17582), .B2(n16601), .A(n16600), .ZN(n16602) );
  OAI21_X1 U19974 ( .B1(n17468), .B2(n17577), .A(n16602), .ZN(n16603) );
  AOI21_X1 U19975 ( .B1(n16769), .B2(n17592), .A(n16603), .ZN(n16604) );
  OAI21_X1 U19976 ( .B1(n16772), .B2(n17566), .A(n16604), .ZN(P2_U2991) );
  NAND2_X1 U19977 ( .A1(n16606), .A2(n16605), .ZN(n16608) );
  XOR2_X1 U19978 ( .A(n16608), .B(n16607), .Z(n16784) );
  INV_X1 U19979 ( .A(n16609), .ZN(n16774) );
  NAND2_X1 U19980 ( .A1(n16610), .A2(n16776), .ZN(n16773) );
  NAND3_X1 U19981 ( .A1(n16774), .A2(n12599), .A3(n16773), .ZN(n16618) );
  OAI22_X1 U19982 ( .A1(n17121), .A2(n20324), .B1(n17571), .B2(n16611), .ZN(
        n16616) );
  OR2_X1 U19983 ( .A1(n16613), .A2(n16612), .ZN(n16614) );
  NAND2_X1 U19984 ( .A1(n13667), .A2(n16614), .ZN(n17471) );
  NOR2_X1 U19985 ( .A1(n17471), .A2(n17577), .ZN(n16615) );
  AOI211_X1 U19986 ( .C1(n17564), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16616), .B(n16615), .ZN(n16617) );
  OAI211_X1 U19987 ( .C1(n16784), .C2(n17572), .A(n16618), .B(n16617), .ZN(
        P2_U2992) );
  NAND2_X1 U19988 ( .A1(n16622), .A2(n16621), .ZN(n16623) );
  AOI21_X1 U19989 ( .B1(n16637), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16624) );
  NOR2_X1 U19990 ( .A1(n16624), .A2(n16596), .ZN(n16796) );
  NAND2_X1 U19991 ( .A1(n20376), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16789) );
  OAI21_X1 U19992 ( .B1(n17596), .B2(n16625), .A(n16789), .ZN(n16626) );
  AOI21_X1 U19993 ( .B1(n17582), .B2(n16627), .A(n16626), .ZN(n16628) );
  OAI21_X1 U19994 ( .B1(n16790), .B2(n17577), .A(n16628), .ZN(n16629) );
  AOI21_X1 U19995 ( .B1(n16796), .B2(n12599), .A(n16629), .ZN(n16630) );
  OAI21_X1 U19996 ( .B1(n16798), .B2(n17572), .A(n16630), .ZN(P2_U2993) );
  NAND2_X1 U19997 ( .A1(n16632), .A2(n16631), .ZN(n16636) );
  INV_X1 U19998 ( .A(n16646), .ZN(n16633) );
  NOR2_X1 U19999 ( .A1(n16634), .A2(n16633), .ZN(n16635) );
  XOR2_X1 U20000 ( .A(n16636), .B(n16635), .Z(n16810) );
  AOI21_X1 U20001 ( .B1(n16799), .B2(n16644), .A(n16637), .ZN(n16807) );
  NAND2_X1 U20002 ( .A1(n20376), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16802) );
  OAI21_X1 U20003 ( .B1(n17596), .B2(n16638), .A(n16802), .ZN(n16639) );
  AOI21_X1 U20004 ( .B1(n16640), .B2(n17582), .A(n16639), .ZN(n16641) );
  OAI21_X1 U20005 ( .B1(n17577), .B2(n16803), .A(n16641), .ZN(n16642) );
  AOI21_X1 U20006 ( .B1(n16807), .B2(n12599), .A(n16642), .ZN(n16643) );
  OAI21_X1 U20007 ( .B1(n16810), .B2(n17572), .A(n16643), .ZN(P2_U2995) );
  OAI21_X1 U20008 ( .B1(n16662), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16644), .ZN(n16821) );
  NAND2_X1 U20009 ( .A1(n16646), .A2(n16645), .ZN(n16647) );
  XNOR2_X1 U20010 ( .A(n16648), .B(n16647), .ZN(n16811) );
  NAND2_X1 U20011 ( .A1(n16811), .A2(n17592), .ZN(n16654) );
  NAND2_X1 U20012 ( .A1(n20376), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16816) );
  OAI21_X1 U20013 ( .B1(n17596), .B2(n16649), .A(n16816), .ZN(n16651) );
  NOR2_X1 U20014 ( .A1(n17480), .A2(n17577), .ZN(n16650) );
  AOI211_X1 U20015 ( .C1(n17582), .C2(n16652), .A(n16651), .B(n16650), .ZN(
        n16653) );
  OAI211_X1 U20016 ( .C1(n17566), .C2(n16821), .A(n16654), .B(n16653), .ZN(
        P2_U2996) );
  NAND2_X1 U20017 ( .A1(n16656), .A2(n16655), .ZN(n16657) );
  XNOR2_X1 U20018 ( .A(n16658), .B(n16657), .ZN(n16838) );
  INV_X1 U20019 ( .A(n16659), .ZN(n16830) );
  NOR2_X1 U20020 ( .A1(n20347), .A2(n21137), .ZN(n16829) );
  AOI21_X1 U20021 ( .B1(n17564), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16829), .ZN(n16660) );
  OAI21_X1 U20022 ( .B1(n17571), .B2(n16661), .A(n16660), .ZN(n16664) );
  INV_X1 U20023 ( .A(n16822), .ZN(n16828) );
  AOI211_X1 U20024 ( .C1(n16834), .C2(n16828), .A(n17566), .B(n16662), .ZN(
        n16663) );
  AOI211_X1 U20025 ( .C1(n16830), .C2(n17591), .A(n16664), .B(n16663), .ZN(
        n16665) );
  OAI21_X1 U20026 ( .B1(n16838), .B2(n17572), .A(n16665), .ZN(P2_U2997) );
  AND2_X1 U20027 ( .A1(n16667), .A2(n16666), .ZN(n16669) );
  OR2_X1 U20028 ( .A1(n16669), .A2(n16668), .ZN(n16843) );
  INV_X1 U20029 ( .A(n16843), .ZN(n20418) );
  NAND2_X1 U20030 ( .A1(n20376), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16841) );
  NAND2_X1 U20031 ( .A1(n17564), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16670) );
  OAI211_X1 U20032 ( .C1(n17571), .C2(n16671), .A(n16841), .B(n16670), .ZN(
        n16676) );
  AND2_X1 U20033 ( .A1(n16674), .A2(n16673), .ZN(n16844) );
  NOR3_X1 U20034 ( .A1(n16672), .A2(n16844), .A3(n17572), .ZN(n16675) );
  AOI211_X1 U20035 ( .C1(n20418), .C2(n17591), .A(n16676), .B(n16675), .ZN(
        n16678) );
  OAI211_X1 U20036 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n9857), .A(
        n16828), .B(n12599), .ZN(n16677) );
  NAND2_X1 U20037 ( .A1(n16678), .A2(n16677), .ZN(P2_U2998) );
  AOI21_X1 U20038 ( .B1(n16680), .B2(n16679), .A(n9832), .ZN(n17629) );
  NAND2_X1 U20039 ( .A1(n16681), .A2(n16897), .ZN(n16686) );
  INV_X1 U20040 ( .A(n16682), .ZN(n16683) );
  NOR2_X1 U20041 ( .A1(n16684), .A2(n16683), .ZN(n16685) );
  XNOR2_X1 U20042 ( .A(n16686), .B(n16685), .ZN(n17632) );
  AOI21_X1 U20043 ( .B1(n16688), .B2(n16687), .A(n14290), .ZN(n20431) );
  AOI22_X1 U20044 ( .A1(n17591), .A2(n20431), .B1(n17564), .B2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16691) );
  INV_X1 U20045 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n21128) );
  OAI22_X1 U20046 ( .A1(n21128), .A2(n20347), .B1(n17571), .B2(n20304), .ZN(
        n16689) );
  INV_X1 U20047 ( .A(n16689), .ZN(n16690) );
  OAI211_X1 U20048 ( .C1(n17632), .C2(n17572), .A(n16691), .B(n16690), .ZN(
        n16692) );
  AOI21_X1 U20049 ( .B1(n17629), .B2(n12599), .A(n16692), .ZN(n16693) );
  INV_X1 U20050 ( .A(n16693), .ZN(P2_U3004) );
  XNOR2_X1 U20051 ( .A(n16695), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16696) );
  XNOR2_X1 U20052 ( .A(n16694), .B(n16696), .ZN(n17652) );
  OAI22_X1 U20053 ( .A1(n16697), .A2(n17596), .B1(n21123), .B2(n20347), .ZN(
        n16699) );
  NOR2_X1 U20054 ( .A1(n17577), .A2(n20342), .ZN(n16698) );
  AOI211_X1 U20055 ( .C1(n17582), .C2(n20337), .A(n16699), .B(n16698), .ZN(
        n16706) );
  AND2_X1 U20056 ( .A1(n16700), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16701) );
  AOI21_X1 U20057 ( .B1(n16703), .B2(n16702), .A(n16701), .ZN(n17555) );
  NAND2_X1 U20058 ( .A1(n17553), .A2(n17552), .ZN(n16704) );
  XNOR2_X1 U20059 ( .A(n17555), .B(n16704), .ZN(n17651) );
  OR2_X1 U20060 ( .A1(n17651), .A2(n17572), .ZN(n16705) );
  OAI211_X1 U20061 ( .C1(n17652), .C2(n17566), .A(n16706), .B(n16705), .ZN(
        P2_U3007) );
  AOI22_X1 U20062 ( .A1(n9818), .A2(n17591), .B1(n17582), .B2(n16707), .ZN(
        n16716) );
  OAI21_X1 U20063 ( .B1(n16709), .B2(n10342), .A(n16708), .ZN(n16710) );
  XNOR2_X1 U20064 ( .A(n16710), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16920) );
  AOI22_X1 U20065 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17564), .B1(
        n17592), .B2(n16920), .ZN(n16715) );
  NAND2_X1 U20066 ( .A1(n20376), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n16916) );
  AOI21_X1 U20067 ( .B1(n16713), .B2(n16712), .A(n16711), .ZN(n16914) );
  NAND2_X1 U20068 ( .A1(n12599), .A2(n16914), .ZN(n16714) );
  NAND4_X1 U20069 ( .A1(n16716), .A2(n16715), .A3(n16916), .A4(n16714), .ZN(
        P2_U3013) );
  NAND4_X1 U20070 ( .A1(n16718), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A4(n16717), .ZN(n16719) );
  OAI211_X1 U20071 ( .C1(n17671), .C2(n17414), .A(n16720), .B(n16719), .ZN(
        n16721) );
  INV_X1 U20072 ( .A(n16721), .ZN(n16724) );
  NAND2_X1 U20073 ( .A1(n16722), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16723) );
  OAI211_X1 U20074 ( .C1(n17409), .C2(n17672), .A(n16724), .B(n16723), .ZN(
        n16725) );
  AOI21_X1 U20075 ( .B1(n16726), .B2(n12521), .A(n16725), .ZN(n16727) );
  OAI21_X1 U20076 ( .B1(n16728), .B2(n17681), .A(n16727), .ZN(P2_U3017) );
  NOR2_X1 U20077 ( .A1(n16746), .A2(n16729), .ZN(n16736) );
  OAI21_X1 U20078 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n16730), .ZN(n16732) );
  OAI21_X1 U20079 ( .B1(n16742), .B2(n16732), .A(n16731), .ZN(n16733) );
  AOI21_X1 U20080 ( .B1(n17637), .B2(n17430), .A(n16733), .ZN(n16734) );
  OAI21_X1 U20081 ( .B1(n17429), .B2(n17672), .A(n16734), .ZN(n16735) );
  AOI211_X1 U20082 ( .C1(n16737), .C2(n12521), .A(n16736), .B(n16735), .ZN(
        n16738) );
  OAI21_X1 U20083 ( .B1(n17681), .B2(n16739), .A(n16738), .ZN(P2_U3020) );
  INV_X1 U20084 ( .A(n16740), .ZN(n17443) );
  NOR2_X1 U20085 ( .A1(n17671), .A2(n17451), .ZN(n16744) );
  OAI21_X1 U20086 ( .B1(n16742), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16741), .ZN(n16743) );
  AOI211_X1 U20087 ( .C1(n17443), .C2(n12878), .A(n16744), .B(n16743), .ZN(
        n16745) );
  OAI21_X1 U20088 ( .B1(n16747), .B2(n16746), .A(n16745), .ZN(n16748) );
  AOI21_X1 U20089 ( .B1(n16749), .B2(n12521), .A(n16748), .ZN(n16750) );
  OAI21_X1 U20090 ( .B1(n17681), .B2(n16751), .A(n16750), .ZN(P2_U3021) );
  AOI21_X1 U20091 ( .B1(n16754), .B2(n16753), .A(n16752), .ZN(n16756) );
  NOR2_X1 U20092 ( .A1(n20324), .A2(n12471), .ZN(n16755) );
  AOI211_X1 U20093 ( .C1(n17637), .C2(n17452), .A(n16756), .B(n16755), .ZN(
        n16757) );
  OAI21_X1 U20094 ( .B1(n17454), .B2(n17672), .A(n16757), .ZN(n16758) );
  AOI21_X1 U20095 ( .B1(n16759), .B2(n17639), .A(n16758), .ZN(n16760) );
  OAI21_X1 U20096 ( .B1(n16761), .B2(n17669), .A(n16760), .ZN(P2_U3022) );
  NOR2_X1 U20097 ( .A1(n16839), .A2(n16762), .ZN(n16777) );
  OAI211_X1 U20098 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16777), .B(n16763), .ZN(
        n16764) );
  OAI211_X1 U20099 ( .C1(n17671), .C2(n16766), .A(n16765), .B(n16764), .ZN(
        n16768) );
  NOR2_X1 U20100 ( .A1(n17468), .A2(n17672), .ZN(n16767) );
  AOI211_X1 U20101 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n16792), .A(
        n16768), .B(n16767), .ZN(n16771) );
  NAND2_X1 U20102 ( .A1(n16769), .A2(n17639), .ZN(n16770) );
  OAI211_X1 U20103 ( .C1(n16772), .C2(n17669), .A(n16771), .B(n16770), .ZN(
        P2_U3023) );
  NAND3_X1 U20104 ( .A1(n16774), .A2(n12521), .A3(n16773), .ZN(n16783) );
  OAI21_X1 U20105 ( .B1(n16775), .B2(n13653), .A(n13670), .ZN(n17485) );
  NAND2_X1 U20106 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n20376), .ZN(n16779) );
  NAND2_X1 U20107 ( .A1(n16777), .A2(n16776), .ZN(n16778) );
  OAI211_X1 U20108 ( .C1(n17671), .C2(n17485), .A(n16779), .B(n16778), .ZN(
        n16781) );
  NOR2_X1 U20109 ( .A1(n17471), .A2(n17672), .ZN(n16780) );
  AOI211_X1 U20110 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n16792), .A(
        n16781), .B(n16780), .ZN(n16782) );
  OAI211_X1 U20111 ( .C1(n16784), .C2(n17681), .A(n16783), .B(n16782), .ZN(
        P2_U3024) );
  INV_X1 U20112 ( .A(n16785), .ZN(n16786) );
  NAND3_X1 U20113 ( .A1(n16800), .A2(n16787), .A3(n16786), .ZN(n16788) );
  OAI211_X1 U20114 ( .C1(n16790), .C2(n17672), .A(n16789), .B(n16788), .ZN(
        n16791) );
  AOI21_X1 U20115 ( .B1(n16792), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16791), .ZN(n16793) );
  OAI21_X1 U20116 ( .B1(n16794), .B2(n17671), .A(n16793), .ZN(n16795) );
  AOI21_X1 U20117 ( .B1(n16796), .B2(n12521), .A(n16795), .ZN(n16797) );
  OAI21_X1 U20118 ( .B1(n16798), .B2(n17681), .A(n16797), .ZN(P2_U3025) );
  NOR2_X1 U20119 ( .A1(n16812), .A2(n16799), .ZN(n16805) );
  NAND2_X1 U20120 ( .A1(n16800), .A2(n16799), .ZN(n16801) );
  OAI211_X1 U20121 ( .C1(n16803), .C2(n17672), .A(n16802), .B(n16801), .ZN(
        n16804) );
  AOI211_X1 U20122 ( .C1(n16806), .C2(n17637), .A(n16805), .B(n16804), .ZN(
        n16809) );
  NAND2_X1 U20123 ( .A1(n16807), .A2(n12521), .ZN(n16808) );
  OAI211_X1 U20124 ( .C1(n16810), .C2(n17681), .A(n16809), .B(n16808), .ZN(
        P2_U3027) );
  NAND2_X1 U20125 ( .A1(n16811), .A2(n17639), .ZN(n16820) );
  NOR2_X1 U20126 ( .A1(n16812), .A2(n16814), .ZN(n16818) );
  NAND3_X1 U20127 ( .A1(n16857), .A2(n16814), .A3(n16813), .ZN(n16815) );
  OAI211_X1 U20128 ( .C1(n17480), .C2(n17672), .A(n16816), .B(n16815), .ZN(
        n16817) );
  AOI211_X1 U20129 ( .C1(n17497), .C2(n17637), .A(n16818), .B(n16817), .ZN(
        n16819) );
  OAI211_X1 U20130 ( .C1(n16821), .C2(n17669), .A(n16820), .B(n16819), .ZN(
        P2_U3028) );
  AOI21_X1 U20131 ( .B1(n17669), .B2(n16823), .A(n16822), .ZN(n16824) );
  AOI211_X1 U20132 ( .C1(n16825), .C2(n16862), .A(n16861), .B(n16824), .ZN(
        n16849) );
  OAI21_X1 U20133 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17675), .A(
        n16849), .ZN(n16826) );
  NAND2_X1 U20134 ( .A1(n16826), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16837) );
  NAND3_X1 U20135 ( .A1(n16857), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16827) );
  OAI21_X1 U20136 ( .B1(n16828), .B2(n17669), .A(n16827), .ZN(n16835) );
  AOI21_X1 U20137 ( .B1(n16830), .B2(n12878), .A(n16829), .ZN(n16831) );
  OAI21_X1 U20138 ( .B1(n16832), .B2(n17671), .A(n16831), .ZN(n16833) );
  AOI21_X1 U20139 ( .B1(n16835), .B2(n16834), .A(n16833), .ZN(n16836) );
  OAI211_X1 U20140 ( .C1(n16838), .C2(n17681), .A(n16837), .B(n16836), .ZN(
        P2_U3029) );
  INV_X1 U20141 ( .A(n9857), .ZN(n17504) );
  OAI22_X1 U20142 ( .A1(n17504), .A2(n17669), .B1(n16862), .B2(n16839), .ZN(
        n16847) );
  AOI21_X1 U20143 ( .B1(n16840), .B2(n13624), .A(n13640), .ZN(n20446) );
  NAND2_X1 U20144 ( .A1(n20446), .A2(n17637), .ZN(n16842) );
  OAI211_X1 U20145 ( .C1(n17672), .C2(n16843), .A(n16842), .B(n16841), .ZN(
        n16846) );
  NOR3_X1 U20146 ( .A1(n16672), .A2(n16844), .A3(n17681), .ZN(n16845) );
  AOI211_X1 U20147 ( .C1(n10092), .C2(n16847), .A(n16846), .B(n16845), .ZN(
        n16848) );
  OAI21_X1 U20148 ( .B1(n16849), .B2(n10092), .A(n16848), .ZN(P2_U3030) );
  INV_X1 U20149 ( .A(n17515), .ZN(n16851) );
  OR2_X1 U20150 ( .A1(n16850), .A2(n16851), .ZN(n16855) );
  NAND2_X1 U20151 ( .A1(n16853), .A2(n16852), .ZN(n16854) );
  XNOR2_X1 U20152 ( .A(n16855), .B(n16854), .ZN(n17502) );
  INV_X1 U20153 ( .A(n17502), .ZN(n16865) );
  NOR2_X1 U20154 ( .A1(n12438), .A2(n20324), .ZN(n16856) );
  AOI21_X1 U20155 ( .B1(n16857), .B2(n16862), .A(n16856), .ZN(n16858) );
  OAI21_X1 U20156 ( .B1(n17672), .B2(n17507), .A(n16858), .ZN(n16860) );
  NOR2_X1 U20157 ( .A1(n20451), .A2(n17671), .ZN(n16859) );
  AOI211_X1 U20158 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16861), .A(
        n16860), .B(n16859), .ZN(n16864) );
  NAND2_X1 U20159 ( .A1(n12613), .A2(n16862), .ZN(n17503) );
  NAND3_X1 U20160 ( .A1(n17504), .A2(n12521), .A3(n17503), .ZN(n16863) );
  OAI211_X1 U20161 ( .C1(n16865), .C2(n17681), .A(n16864), .B(n16863), .ZN(
        P2_U3031) );
  NAND2_X1 U20162 ( .A1(n16867), .A2(n16866), .ZN(n16869) );
  XOR2_X1 U20163 ( .A(n16869), .B(n16868), .Z(n17526) );
  INV_X1 U20164 ( .A(n17526), .ZN(n16876) );
  OAI22_X1 U20165 ( .A1(n17672), .A2(n16870), .B1(n15036), .B2(n20347), .ZN(
        n16872) );
  AOI21_X1 U20166 ( .B1(n17619), .B2(n11910), .A(n17616), .ZN(n17603) );
  NAND2_X1 U20167 ( .A1(n17619), .A2(n11953), .ZN(n17602) );
  OAI22_X1 U20168 ( .A1(n17603), .A2(n11953), .B1(n11910), .B2(n17602), .ZN(
        n16871) );
  AOI211_X1 U20169 ( .C1(n20455), .C2(n17637), .A(n16872), .B(n16871), .ZN(
        n16875) );
  OAI21_X1 U20170 ( .B1(n9859), .B2(n11910), .A(n11953), .ZN(n16873) );
  OR2_X1 U20171 ( .A1(n9859), .A2(n17614), .ZN(n17512) );
  NAND2_X1 U20172 ( .A1(n17527), .A2(n12521), .ZN(n16874) );
  OAI211_X1 U20173 ( .C1(n16876), .C2(n17681), .A(n16875), .B(n16874), .ZN(
        P2_U3033) );
  OAI21_X1 U20174 ( .B1(n9832), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n9859), .ZN(n17541) );
  NOR2_X1 U20175 ( .A1(n9868), .A2(n16877), .ZN(n16881) );
  NOR2_X1 U20176 ( .A1(n16879), .A2(n16878), .ZN(n16880) );
  XNOR2_X1 U20177 ( .A(n16881), .B(n16880), .ZN(n17543) );
  OAI21_X1 U20178 ( .B1(n16884), .B2(n16883), .A(n16882), .ZN(n20462) );
  INV_X1 U20179 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n21130) );
  NOR2_X1 U20180 ( .A1(n21130), .A2(n20347), .ZN(n16889) );
  XNOR2_X1 U20181 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16887) );
  OAI21_X1 U20182 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17675), .A(
        n16909), .ZN(n17628) );
  INV_X1 U20183 ( .A(n17628), .ZN(n16885) );
  OAI22_X1 U20184 ( .A1(n16887), .A2(n17625), .B1(n16886), .B2(n16885), .ZN(
        n16888) );
  AOI211_X1 U20185 ( .C1(n12878), .C2(n20294), .A(n16889), .B(n16888), .ZN(
        n16890) );
  OAI21_X1 U20186 ( .B1(n20462), .B2(n17671), .A(n16890), .ZN(n16891) );
  AOI21_X1 U20187 ( .B1(n17543), .B2(n17639), .A(n16891), .ZN(n16892) );
  OAI21_X1 U20188 ( .B1(n17541), .B2(n17669), .A(n16892), .ZN(P2_U3035) );
  INV_X1 U20189 ( .A(n16893), .ZN(n16895) );
  INV_X1 U20190 ( .A(n16679), .ZN(n16894) );
  AOI21_X1 U20191 ( .B1(n16895), .B2(n16908), .A(n16894), .ZN(n17547) );
  INV_X1 U20192 ( .A(n17547), .ZN(n16913) );
  INV_X1 U20193 ( .A(n16897), .ZN(n16898) );
  NOR2_X1 U20194 ( .A1(n16899), .A2(n16898), .ZN(n16900) );
  XNOR2_X1 U20195 ( .A(n16896), .B(n16900), .ZN(n17546) );
  OAI21_X1 U20196 ( .B1(n16901), .B2(n16903), .A(n16902), .ZN(n20467) );
  NOR2_X1 U20197 ( .A1(n20467), .A2(n17671), .ZN(n16911) );
  INV_X1 U20198 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n21126) );
  NOR2_X1 U20199 ( .A1(n21126), .A2(n20347), .ZN(n16904) );
  AOI21_X1 U20200 ( .B1(n16905), .B2(n16908), .A(n16904), .ZN(n16907) );
  NAND2_X1 U20201 ( .A1(n12878), .A2(n20316), .ZN(n16906) );
  OAI211_X1 U20202 ( .C1(n16909), .C2(n16908), .A(n16907), .B(n16906), .ZN(
        n16910) );
  AOI211_X1 U20203 ( .C1(n17546), .C2(n17639), .A(n16911), .B(n16910), .ZN(
        n16912) );
  OAI21_X1 U20204 ( .B1(n16913), .B2(n17669), .A(n16912), .ZN(P2_U3037) );
  INV_X1 U20205 ( .A(n17670), .ZN(n16915) );
  AOI22_X1 U20206 ( .A1(n16915), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n12521), .B2(n16914), .ZN(n16917) );
  OAI211_X1 U20207 ( .C1(n17672), .C2(n16918), .A(n16917), .B(n16916), .ZN(
        n16919) );
  INV_X1 U20208 ( .A(n16919), .ZN(n16925) );
  AOI22_X1 U20209 ( .A1(n17639), .A2(n16920), .B1(n17637), .B2(n21201), .ZN(
        n16924) );
  OAI211_X1 U20210 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n16922), .B(n16921), .ZN(n16923) );
  NAND3_X1 U20211 ( .A1(n16925), .A2(n16924), .A3(n16923), .ZN(P2_U3045) );
  INV_X1 U20212 ( .A(n16964), .ZN(n16931) );
  INV_X1 U20213 ( .A(n16926), .ZN(n16928) );
  MUX2_X1 U20214 ( .A(n16929), .B(n16928), .S(n16927), .Z(n16930) );
  OAI21_X1 U20215 ( .B1(n20403), .B2(n16931), .A(n16930), .ZN(n17694) );
  AOI21_X1 U20216 ( .B1(n17694), .B2(n20975), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n16933) );
  OAI22_X1 U20217 ( .A1(n16947), .A2(n16933), .B1(n16932), .B2(n16965), .ZN(
        n16934) );
  INV_X1 U20218 ( .A(n16966), .ZN(n17084) );
  MUX2_X1 U20219 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n16934), .S(
        n17084), .Z(P2_U3601) );
  INV_X1 U20220 ( .A(n21082), .ZN(n21179) );
  INV_X1 U20221 ( .A(n16936), .ZN(n16937) );
  NAND2_X1 U20222 ( .A1(n12236), .A2(n16937), .ZN(n16953) );
  NAND2_X1 U20223 ( .A1(n16952), .A2(n12234), .ZN(n16940) );
  NOR2_X1 U20224 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16938) );
  OR2_X1 U20225 ( .A1(n16935), .A2(n16938), .ZN(n16951) );
  NOR2_X1 U20226 ( .A1(n16951), .A2(n16939), .ZN(n16941) );
  NAND2_X1 U20227 ( .A1(n16940), .A2(n16941), .ZN(n16944) );
  OR2_X1 U20228 ( .A1(n17708), .A2(n17704), .ZN(n16959) );
  INV_X1 U20229 ( .A(n16941), .ZN(n16942) );
  NAND2_X1 U20230 ( .A1(n16959), .A2(n16942), .ZN(n16943) );
  OAI211_X1 U20231 ( .C1(n16935), .C2(n16953), .A(n16944), .B(n16943), .ZN(
        n16945) );
  AOI21_X1 U20232 ( .B1(n16946), .B2(n16964), .A(n16945), .ZN(n17688) );
  INV_X1 U20233 ( .A(n16947), .ZN(n16949) );
  OAI222_X1 U20234 ( .A1(n21190), .A2(n16965), .B1(n21179), .B2(n17688), .C1(
        n16949), .C2(n16948), .ZN(n16950) );
  MUX2_X1 U20235 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16950), .S(
        n17084), .Z(P2_U3599) );
  INV_X1 U20236 ( .A(n16951), .ZN(n16958) );
  NAND3_X1 U20237 ( .A1(n16952), .A2(n16958), .A3(n12234), .ZN(n16955) );
  INV_X1 U20238 ( .A(n16953), .ZN(n16954) );
  AOI21_X1 U20239 ( .B1(n16955), .B2(n13041), .A(n16954), .ZN(n16961) );
  NAND2_X1 U20240 ( .A1(n12236), .A2(n16936), .ZN(n16956) );
  NAND2_X1 U20241 ( .A1(n16956), .A2(n13041), .ZN(n16957) );
  AOI21_X1 U20242 ( .B1(n16959), .B2(n16958), .A(n16957), .ZN(n16960) );
  MUX2_X1 U20243 ( .A(n16961), .B(n16960), .S(n17691), .Z(n16962) );
  INV_X1 U20244 ( .A(n16962), .ZN(n16963) );
  AOI21_X1 U20245 ( .B1(n13907), .B2(n16964), .A(n16963), .ZN(n17690) );
  OAI22_X1 U20246 ( .A1(n20800), .A2(n16965), .B1(n17690), .B2(n21179), .ZN(
        n16967) );
  MUX2_X1 U20247 ( .A(n16967), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16966), .Z(P2_U3596) );
  INV_X1 U20248 ( .A(n20810), .ZN(n20768) );
  NOR2_X2 U20249 ( .A1(n20768), .A2(n20672), .ZN(n20607) );
  OAI21_X1 U20250 ( .B1(n21075), .B2(n20607), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16969) );
  NAND2_X1 U20251 ( .A1(n16969), .A2(n21177), .ZN(n16974) );
  NAND2_X1 U20252 ( .A1(n16970), .A2(n21203), .ZN(n20591) );
  NOR2_X1 U20253 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20591), .ZN(
        n20575) );
  INV_X1 U20254 ( .A(n20575), .ZN(n16971) );
  AND2_X1 U20255 ( .A1(n21019), .A2(n16971), .ZN(n16977) );
  INV_X1 U20256 ( .A(n16972), .ZN(n16975) );
  OAI21_X1 U20257 ( .B1(n16975), .B2(n20575), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16973) );
  OAI21_X1 U20258 ( .B1(n16974), .B2(n16977), .A(n16973), .ZN(n20581) );
  INV_X1 U20259 ( .A(n16974), .ZN(n16978) );
  AOI211_X1 U20260 ( .C1(n16975), .C2(n20975), .A(n21177), .B(n20575), .ZN(
        n16976) );
  AOI22_X1 U20261 ( .A1(n21066), .A2(n20607), .B1(n21064), .B2(n20575), .ZN(
        n16980) );
  NAND2_X1 U20262 ( .A1(n21003), .A2(n21075), .ZN(n16979) );
  OAI211_X1 U20263 ( .C1(n20585), .C2(n16981), .A(n16980), .B(n16979), .ZN(
        n16982) );
  AOI21_X1 U20264 ( .B1(n21065), .B2(n20581), .A(n16982), .ZN(n16983) );
  INV_X1 U20265 ( .A(n16983), .ZN(P2_U3054) );
  INV_X1 U20266 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n18279) );
  INV_X1 U20267 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n18277) );
  INV_X1 U20268 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n18557) );
  INV_X1 U20269 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n18561) );
  NOR2_X1 U20270 ( .A1(n18624), .A2(n16984), .ZN(n16985) );
  NAND4_X1 U20271 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .A4(n18424), .ZN(n18384) );
  NAND2_X1 U20272 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n18341), .ZN(n18335) );
  NAND2_X1 U20273 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n18331), .ZN(n17061) );
  INV_X1 U20274 ( .A(n18577), .ZN(n18578) );
  NOR2_X2 U20275 ( .A1(n19584), .A2(n18578), .ZN(n18579) );
  NOR2_X1 U20276 ( .A1(n18579), .A2(n18319), .ZN(n18320) );
  AOI22_X1 U20277 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n9794), .B1(
        P3_INSTQUEUE_REG_10__4__SCAN_IN), .B2(n9793), .ZN(n16991) );
  AOI22_X1 U20278 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16990) );
  AOI22_X1 U20279 ( .A1(n18519), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20280 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16988) );
  NAND4_X1 U20281 ( .A1(n16991), .A2(n16990), .A3(n16989), .A4(n16988), .ZN(
        n16997) );
  AOI22_X1 U20282 ( .A1(n18520), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20283 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20284 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18533), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20285 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18503), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16992) );
  NAND4_X1 U20286 ( .A1(n16995), .A2(n16994), .A3(n16993), .A4(n16992), .ZN(
        n16996) );
  OR2_X1 U20287 ( .A1(n16997), .A2(n16996), .ZN(n18323) );
  AOI22_X1 U20288 ( .A1(n18520), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20289 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9794), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20290 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20291 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18534), .B1(
        n18472), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16998) );
  NAND4_X1 U20292 ( .A1(n17001), .A2(n17000), .A3(n16999), .A4(n16998), .ZN(
        n17007) );
  AOI22_X1 U20293 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18473), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17005) );
  AOI22_X1 U20294 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20295 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18519), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20296 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17002) );
  NAND4_X1 U20297 ( .A1(n17005), .A2(n17004), .A3(n17003), .A4(n17002), .ZN(
        n17006) );
  NOR2_X1 U20298 ( .A1(n17007), .A2(n17006), .ZN(n18332) );
  AOI22_X1 U20299 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20300 ( .A1(n18519), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20301 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20302 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17008) );
  NAND4_X1 U20303 ( .A1(n17011), .A2(n17010), .A3(n17009), .A4(n17008), .ZN(
        n17017) );
  AOI22_X1 U20304 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18503), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20305 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20306 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20307 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17012) );
  NAND4_X1 U20308 ( .A1(n17015), .A2(n17014), .A3(n17013), .A4(n17012), .ZN(
        n17016) );
  NOR2_X1 U20309 ( .A1(n17017), .A2(n17016), .ZN(n18343) );
  AOI22_X1 U20310 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17067), .ZN(n17021) );
  AOI22_X1 U20311 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n18518), .ZN(n17020) );
  AOI22_X1 U20312 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9794), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20313 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18534), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17018) );
  NAND4_X1 U20314 ( .A1(n17021), .A2(n17020), .A3(n17019), .A4(n17018), .ZN(
        n17027) );
  AOI22_X1 U20315 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n13311), .ZN(n17025) );
  AOI22_X1 U20316 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20317 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18455), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20318 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18473), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17066), .ZN(n17022) );
  NAND4_X1 U20319 ( .A1(n17025), .A2(n17024), .A3(n17023), .A4(n17022), .ZN(
        n17026) );
  NOR2_X1 U20320 ( .A1(n17027), .A2(n17026), .ZN(n18342) );
  NOR2_X1 U20321 ( .A1(n18343), .A2(n18342), .ZN(n18338) );
  AOI22_X1 U20322 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18473), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20323 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20324 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17028) );
  OAI21_X1 U20325 ( .B1(n17030), .B2(n17029), .A(n17028), .ZN(n17036) );
  AOI22_X1 U20326 ( .A1(n13259), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20327 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20328 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18472), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20329 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17031) );
  NAND4_X1 U20330 ( .A1(n17034), .A2(n17033), .A3(n17032), .A4(n17031), .ZN(
        n17035) );
  AOI211_X1 U20331 ( .C1(n13311), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n17036), .B(n17035), .ZN(n17037) );
  NAND3_X1 U20332 ( .A1(n17039), .A2(n17038), .A3(n17037), .ZN(n18337) );
  NAND2_X1 U20333 ( .A1(n18338), .A2(n18337), .ZN(n18336) );
  NOR2_X1 U20334 ( .A1(n18332), .A2(n18336), .ZN(n18329) );
  AOI22_X1 U20335 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20336 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20337 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17040) );
  OAI21_X1 U20338 ( .B1(n18487), .B2(n18453), .A(n17040), .ZN(n17046) );
  AOI22_X1 U20339 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20340 ( .A1(n18519), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20341 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18503), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20342 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17041) );
  NAND4_X1 U20343 ( .A1(n17044), .A2(n17043), .A3(n17042), .A4(n17041), .ZN(
        n17045) );
  AOI211_X1 U20344 ( .C1(n9793), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n17046), .B(n17045), .ZN(n17047) );
  NAND3_X1 U20345 ( .A1(n17049), .A2(n17048), .A3(n17047), .ZN(n18328) );
  NAND2_X1 U20346 ( .A1(n18329), .A2(n18328), .ZN(n18327) );
  INV_X1 U20347 ( .A(n18327), .ZN(n18324) );
  NAND2_X1 U20348 ( .A1(n18323), .A2(n18324), .ZN(n18322) );
  AOI22_X1 U20349 ( .A1(n18520), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20350 ( .A1(n13259), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20351 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n9794), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17051) );
  AOI22_X1 U20352 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18534), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17050) );
  NAND4_X1 U20353 ( .A1(n17053), .A2(n17052), .A3(n17051), .A4(n17050), .ZN(
        n17059) );
  AOI22_X1 U20354 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20355 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20356 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20357 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17054) );
  NAND4_X1 U20358 ( .A1(n17057), .A2(n17056), .A3(n17055), .A4(n17054), .ZN(
        n17058) );
  NOR2_X1 U20359 ( .A1(n17059), .A2(n17058), .ZN(n18315) );
  XOR2_X1 U20360 ( .A(n18322), .B(n18315), .Z(n18596) );
  AOI22_X1 U20361 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18320), .B1(n18579), 
        .B2(n18596), .ZN(n17060) );
  OAI21_X1 U20362 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17061), .A(n17060), .ZN(
        P3_U2675) );
  AOI22_X1 U20363 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20364 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18503), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20365 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17063) );
  AOI22_X1 U20366 ( .A1(n13259), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17062) );
  NAND4_X1 U20367 ( .A1(n17065), .A2(n17064), .A3(n17063), .A4(n17062), .ZN(
        n17073) );
  AOI22_X1 U20368 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20369 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20370 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20371 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18533), .B1(
        n18519), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17068) );
  NAND4_X1 U20372 ( .A1(n17071), .A2(n17070), .A3(n17069), .A4(n17068), .ZN(
        n17072) );
  NOR2_X1 U20373 ( .A1(n17073), .A2(n17072), .ZN(n18677) );
  NOR2_X1 U20374 ( .A1(n18624), .A2(n17074), .ZN(n18481) );
  NOR2_X1 U20375 ( .A1(n18579), .A2(n9927), .ZN(n18465) );
  OAI21_X1 U20376 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n18481), .A(n18465), .ZN(
        n17075) );
  OAI21_X1 U20377 ( .B1(n18677), .B2(n18570), .A(n17075), .ZN(P3_U2690) );
  NAND2_X1 U20378 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19697) );
  INV_X1 U20379 ( .A(n19121), .ZN(n19165) );
  NOR2_X1 U20380 ( .A1(n19542), .A2(n19165), .ZN(n17077) );
  AOI221_X1 U20381 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19697), .C1(n17077), 
        .C2(n19697), .A(n17076), .ZN(n19545) );
  NOR2_X1 U20382 ( .A1(n17078), .A2(n20021), .ZN(n17079) );
  OAI21_X1 U20383 ( .B1(n17079), .B2(n19608), .A(n19546), .ZN(n19543) );
  AOI22_X1 U20384 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19545), .B1(
        n19543), .B2(n20026), .ZN(P3_U2865) );
  INV_X1 U20385 ( .A(n17712), .ZN(n17080) );
  NOR4_X1 U20386 ( .A1(n15199), .A2(n17080), .A3(n11624), .A4(n21179), .ZN(
        n17081) );
  NAND2_X1 U20387 ( .A1(n17084), .A2(n17081), .ZN(n17082) );
  OAI21_X1 U20388 ( .B1(n17084), .B2(n17083), .A(n17082), .ZN(P2_U3595) );
  INV_X1 U20389 ( .A(n17085), .ZN(n19982) );
  AOI211_X1 U20390 ( .C1(n19568), .C2(n17087), .A(n19559), .B(n17086), .ZN(
        n17089) );
  AOI21_X1 U20391 ( .B1(n20205), .B2(n19559), .A(n17091), .ZN(n17093) );
  AOI21_X1 U20392 ( .B1(n17093), .B2(n17092), .A(n10001), .ZN(n17892) );
  INV_X1 U20393 ( .A(n17094), .ZN(n17095) );
  NAND3_X1 U20394 ( .A1(n19981), .A2(n17892), .A3(n17095), .ZN(n17096) );
  NOR2_X1 U20395 ( .A1(n18698), .A2(n19983), .ZN(n19381) );
  NAND2_X1 U20396 ( .A1(n19466), .A2(n19381), .ZN(n19439) );
  INV_X1 U20397 ( .A(n19439), .ZN(n19251) );
  NOR2_X1 U20398 ( .A1(n19511), .A2(n19533), .ZN(n19374) );
  INV_X1 U20399 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n19232) );
  NOR2_X1 U20400 ( .A1(n19219), .A2(n19232), .ZN(n17779) );
  NOR3_X1 U20401 ( .A1(n19488), .A2(n19496), .A3(n19480), .ZN(n19322) );
  OAI21_X1 U20402 ( .B1(n20181), .B2(n9952), .A(n19507), .ZN(n19504) );
  NAND2_X1 U20403 ( .A1(n19322), .A2(n19504), .ZN(n19444) );
  NOR2_X1 U20404 ( .A1(n19456), .A2(n19468), .ZN(n19450) );
  NAND2_X1 U20405 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19450), .ZN(
        n19324) );
  NOR2_X1 U20406 ( .A1(n19444), .A2(n19324), .ZN(n19337) );
  NAND3_X1 U20407 ( .A1(n18959), .A2(n17100), .A3(n19337), .ZN(n19319) );
  NOR2_X1 U20408 ( .A1(n17098), .A2(n19319), .ZN(n19259) );
  INV_X1 U20409 ( .A(n17099), .ZN(n17740) );
  NOR2_X1 U20410 ( .A1(n19507), .A2(n9952), .ZN(n19483) );
  AND2_X1 U20411 ( .A1(n19483), .A2(n19322), .ZN(n19446) );
  NAND2_X1 U20412 ( .A1(n19446), .A2(n19450), .ZN(n19428) );
  NOR2_X1 U20413 ( .A1(n19449), .A2(n19428), .ZN(n19378) );
  NAND2_X1 U20414 ( .A1(n17100), .A2(n19378), .ZN(n19317) );
  INV_X1 U20415 ( .A(n19317), .ZN(n19277) );
  NAND2_X1 U20416 ( .A1(n17740), .A2(n19277), .ZN(n19220) );
  INV_X1 U20417 ( .A(n19220), .ZN(n17101) );
  INV_X1 U20418 ( .A(n20016), .ZN(n19988) );
  INV_X1 U20419 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19289) );
  INV_X1 U20420 ( .A(n17100), .ZN(n19326) );
  NAND2_X1 U20421 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19378), .ZN(
        n19429) );
  NOR2_X1 U20422 ( .A1(n19326), .A2(n19429), .ZN(n19338) );
  NAND2_X1 U20423 ( .A1(n18926), .A2(n19338), .ZN(n19281) );
  NOR2_X1 U20424 ( .A1(n19289), .A2(n19281), .ZN(n17105) );
  AOI222_X1 U20425 ( .A1(n19259), .A2(n19977), .B1(n17101), .B2(n19988), .C1(
        n17105), .C2(n20014), .ZN(n17102) );
  INV_X1 U20426 ( .A(n17102), .ZN(n19243) );
  NAND4_X1 U20427 ( .A1(n19466), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17779), .A4(n19243), .ZN(n17767) );
  OAI21_X1 U20428 ( .B1(n19536), .B2(n17792), .A(n17767), .ZN(n17103) );
  AOI21_X1 U20429 ( .B1(n17794), .B2(n19251), .A(n17103), .ZN(n17185) );
  INV_X1 U20430 ( .A(n19419), .ZN(n17108) );
  INV_X1 U20431 ( .A(n17104), .ZN(n17107) );
  INV_X1 U20432 ( .A(n20014), .ZN(n19427) );
  AOI21_X1 U20433 ( .B1(n19244), .B2(n19259), .A(n20009), .ZN(n19242) );
  AOI21_X1 U20434 ( .B1(n19977), .B2(n19221), .A(n19242), .ZN(n19223) );
  OAI221_X1 U20435 ( .B1(n19427), .B2(n17105), .C1(n19427), .C2(n17779), .A(
        n19223), .ZN(n17106) );
  AOI221_X1 U20436 ( .B1(n17107), .B2(n19988), .C1(n19317), .C2(n19988), .A(
        n17106), .ZN(n17179) );
  OAI21_X1 U20437 ( .B1(n17108), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17179), .ZN(n17791) );
  NOR2_X1 U20438 ( .A1(n19364), .A2(n19533), .ZN(n17772) );
  INV_X1 U20439 ( .A(n17772), .ZN(n19520) );
  INV_X1 U20440 ( .A(n17109), .ZN(n17761) );
  AOI22_X1 U20441 ( .A1(n19374), .A2(n17756), .B1(n19251), .B2(n17761), .ZN(
        n17182) );
  OAI211_X1 U20442 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n19520), .A(
        n17182), .B(n19497), .ZN(n17110) );
  AOI21_X1 U20443 ( .B1(n19466), .B2(n17791), .A(n17110), .ZN(n17115) );
  NOR2_X1 U20444 ( .A1(n17112), .A2(n17111), .ZN(n17113) );
  XNOR2_X1 U20445 ( .A(n17113), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17760) );
  AOI22_X1 U20446 ( .A1(n9790), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n19443), 
        .B2(n17760), .ZN(n17114) );
  OAI221_X1 U20447 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17185), 
        .C1(n17758), .C2(n17115), .A(n17114), .ZN(P3_U2833) );
  OAI22_X1 U20448 ( .A1(n17471), .A2(n20402), .B1(n20401), .B2(n17485), .ZN(
        n17116) );
  INV_X1 U20449 ( .A(n17116), .ZN(n17126) );
  AOI211_X1 U20450 ( .C1(n17119), .C2(n17118), .A(n17117), .B(n21086), .ZN(
        n17124) );
  INV_X1 U20451 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n17120) );
  OAI222_X1 U20452 ( .A1(n17122), .A2(n20399), .B1(n20374), .B2(n17121), .C1(
        n20396), .C2(n17120), .ZN(n17123) );
  AOI211_X1 U20453 ( .C1(n20412), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17124), .B(n17123), .ZN(n17125) );
  NAND2_X1 U20454 ( .A1(n17126), .A2(n17125), .ZN(P2_U2833) );
  OAI21_X1 U20455 ( .B1(n17128), .B2(n17127), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17129) );
  OR2_X1 U20456 ( .A1(n17130), .A2(n17129), .ZN(n17133) );
  OAI21_X1 U20457 ( .B1(n17133), .B2(n17132), .A(n17131), .ZN(n17135) );
  INV_X1 U20458 ( .A(n17133), .ZN(n17134) );
  OAI22_X1 U20459 ( .A1(n17136), .A2(n17135), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17134), .ZN(n17137) );
  AOI21_X1 U20460 ( .B1(n17139), .B2(n17138), .A(n17137), .ZN(n17141) );
  NOR2_X1 U20461 ( .A1(n17139), .A2(n17138), .ZN(n17140) );
  OR2_X1 U20462 ( .A1(n17141), .A2(n17140), .ZN(n17145) );
  NAND2_X1 U20463 ( .A1(n17145), .A2(n17142), .ZN(n17144) );
  NAND2_X1 U20464 ( .A1(n17144), .A2(n17143), .ZN(n17149) );
  INV_X1 U20465 ( .A(n17145), .ZN(n17147) );
  NAND2_X1 U20466 ( .A1(n17147), .A2(n17146), .ZN(n17148) );
  NAND2_X1 U20467 ( .A1(n17149), .A2(n17148), .ZN(n17159) );
  INV_X1 U20468 ( .A(n17150), .ZN(n17151) );
  NOR2_X1 U20469 ( .A1(n17152), .A2(n17151), .ZN(n17155) );
  OAI21_X1 U20470 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n17153), .ZN(n17154) );
  NAND4_X1 U20471 ( .A1(n17157), .A2(n17156), .A3(n17155), .A4(n17154), .ZN(
        n17158) );
  AOI21_X1 U20472 ( .B1(n17159), .B2(n21437), .A(n17158), .ZN(n17169) );
  INV_X1 U20473 ( .A(n17169), .ZN(n17161) );
  AOI21_X1 U20474 ( .B1(n17162), .B2(n17161), .A(n17160), .ZN(n17175) );
  INV_X1 U20475 ( .A(n17163), .ZN(n17164) );
  NOR4_X1 U20476 ( .A1(n12774), .A2(n17165), .A3(n17186), .A4(n17164), .ZN(
        n17166) );
  AOI221_X1 U20477 ( .B1(n17168), .B2(n17167), .C1(n21452), .C2(n17167), .A(
        n17166), .ZN(n17395) );
  OAI221_X1 U20478 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n17169), 
        .A(n17395), .ZN(n17171) );
  AND2_X1 U20479 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17171), .ZN(n17401) );
  OAI211_X1 U20480 ( .C1(n21452), .C2(P1_STATE2_REG_2__SCAN_IN), .A(n17172), 
        .B(n17401), .ZN(n17398) );
  INV_X1 U20481 ( .A(n17398), .ZN(n17174) );
  OAI21_X1 U20482 ( .B1(n17172), .B2(n10053), .A(n17171), .ZN(n17173) );
  AOI22_X1 U20483 ( .A1(n17175), .A2(n17174), .B1(n21439), .B2(n17173), .ZN(
        P1_U3161) );
  NAND2_X1 U20484 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17751), .ZN(
        n17741) );
  NAND2_X1 U20485 ( .A1(n17177), .A2(n17176), .ZN(n17178) );
  XNOR2_X1 U20486 ( .A(n17178), .B(n17751), .ZN(n17748) );
  OAI21_X1 U20487 ( .B1(n17179), .B2(n19533), .A(n19497), .ZN(n17180) );
  AOI21_X1 U20488 ( .B1(n17772), .B2(n17181), .A(n17180), .ZN(n17769) );
  AOI21_X1 U20489 ( .B1(n17769), .B2(n17182), .A(n17751), .ZN(n17183) );
  AOI21_X1 U20490 ( .B1(n19443), .B2(n17748), .A(n17183), .ZN(n17184) );
  NAND2_X1 U20491 ( .A1(n9790), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17743) );
  OAI211_X1 U20492 ( .C1(n17185), .C2(n17741), .A(n17184), .B(n17743), .ZN(
        P3_U2832) );
  INV_X1 U20493 ( .A(HOLD), .ZN(n21444) );
  NOR2_X1 U20494 ( .A1(n10503), .A2(n21444), .ZN(n21446) );
  INV_X1 U20495 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21547) );
  NOR2_X1 U20496 ( .A1(n12634), .A2(n21547), .ZN(n21451) );
  AOI21_X1 U20497 ( .B1(HOLD), .B2(P1_STATE_REG_1__SCAN_IN), .A(n21451), .ZN(
        n17187) );
  NAND2_X1 U20498 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21541), .ZN(n21458) );
  OAI211_X1 U20499 ( .C1(n21446), .C2(n17187), .A(n17186), .B(n21458), .ZN(
        P1_U3195) );
  AND2_X1 U20500 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n21407), .ZN(P1_U2905)
         );
  NOR2_X1 U20501 ( .A1(n21226), .A2(n17682), .ZN(n21081) );
  AOI22_X1 U20502 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21081), .B1(
        P2_STATEBS16_REG_SCAN_IN), .B2(n21237), .ZN(n17188) );
  AOI21_X1 U20503 ( .B1(n17188), .B2(n21225), .A(n17736), .ZN(P2_U3178) );
  INV_X1 U20504 ( .A(n17725), .ZN(n21220) );
  AOI221_X1 U20505 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17736), .C1(n21220), .C2(
        n17736), .A(n21023), .ZN(n21210) );
  INV_X1 U20506 ( .A(n21210), .ZN(n21211) );
  NOR2_X1 U20507 ( .A1(n17701), .A2(n21211), .ZN(P2_U3047) );
  OR3_X1 U20508 ( .A1(n17189), .A2(n18732), .A3(n19555), .ZN(n17190) );
  NAND2_X1 U20509 ( .A1(n19584), .A2(n18724), .ZN(n18668) );
  INV_X1 U20510 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18793) );
  AOI22_X1 U20511 ( .A1(n18723), .A2(BUF2_REG_0__SCAN_IN), .B1(n18722), .B2(
        n17192), .ZN(n17193) );
  OAI221_X1 U20512 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n18668), .C1(n18793), 
        .C2(n18724), .A(n17193), .ZN(P3_U2735) );
  AOI22_X1 U20513 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n21331), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n17202), .ZN(n17199) );
  AOI22_X1 U20514 ( .A1(n21343), .A2(P1_EBX_REG_22__SCAN_IN), .B1(n21339), 
        .B2(n17257), .ZN(n17198) );
  AOI22_X1 U20515 ( .A1(n17258), .A2(n21312), .B1(n21345), .B2(n17194), .ZN(
        n17197) );
  OAI211_X1 U20516 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(P1_REIP_REG_21__SCAN_IN), .A(n10025), .B(n17195), .ZN(n17196) );
  NAND4_X1 U20517 ( .A1(n17199), .A2(n17198), .A3(n17197), .A4(n17196), .ZN(
        P1_U2818) );
  INV_X1 U20518 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17209) );
  OAI22_X1 U20519 ( .A1(n21308), .A2(n17200), .B1(n21348), .B2(n17266), .ZN(
        n17201) );
  AOI21_X1 U20520 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n17202), .A(n17201), 
        .ZN(n17208) );
  INV_X1 U20521 ( .A(n17203), .ZN(n17263) );
  OAI22_X1 U20522 ( .A1(n17205), .A2(P1_REIP_REG_21__SCAN_IN), .B1(n17204), 
        .B2(n21296), .ZN(n17206) );
  AOI21_X1 U20523 ( .B1(n17263), .B2(n21312), .A(n17206), .ZN(n17207) );
  OAI211_X1 U20524 ( .C1(n17209), .C2(n21349), .A(n17208), .B(n17207), .ZN(
        P1_U2819) );
  NOR2_X1 U20525 ( .A1(n21292), .A2(n17210), .ZN(n17231) );
  INV_X1 U20526 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17211) );
  OAI21_X1 U20527 ( .B1(n21349), .B2(n17211), .A(n21273), .ZN(n17214) );
  OAI22_X1 U20528 ( .A1(n21308), .A2(n17212), .B1(n21348), .B2(n17272), .ZN(
        n17213) );
  AOI211_X1 U20529 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(n17231), .A(n17214), 
        .B(n17213), .ZN(n17219) );
  INV_X1 U20530 ( .A(n17215), .ZN(n17269) );
  INV_X1 U20531 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21490) );
  AOI21_X1 U20532 ( .B1(n21490), .B2(n16150), .A(n9908), .ZN(n17217) );
  AOI22_X1 U20533 ( .A1(n17269), .A2(n21312), .B1(n17217), .B2(n17216), .ZN(
        n17218) );
  OAI211_X1 U20534 ( .C1(n21296), .C2(n17220), .A(n17219), .B(n17218), .ZN(
        P1_U2821) );
  AOI22_X1 U20535 ( .A1(n21343), .A2(P1_EBX_REG_18__SCAN_IN), .B1(n17221), 
        .B2(n21339), .ZN(n17222) );
  OAI211_X1 U20536 ( .C1(n21349), .C2(n10900), .A(n17222), .B(n21273), .ZN(
        n17223) );
  AOI21_X1 U20537 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n17231), .A(n17223), 
        .ZN(n17227) );
  AOI22_X1 U20538 ( .A1(n17225), .A2(n21312), .B1(n21345), .B2(n17224), .ZN(
        n17226) );
  OAI211_X1 U20539 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n9908), .A(n17227), .B(
        n17226), .ZN(P1_U2822) );
  OAI22_X1 U20540 ( .A1(n21308), .A2(n17253), .B1(n21349), .B2(n17228), .ZN(
        n17229) );
  AOI21_X1 U20541 ( .B1(n17273), .B2(n21339), .A(n17229), .ZN(n17235) );
  INV_X1 U20542 ( .A(n17230), .ZN(n17274) );
  AOI22_X1 U20543 ( .A1(n17274), .A2(n21312), .B1(n21345), .B2(n17251), .ZN(
        n17234) );
  OAI21_X1 U20544 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n17232), .A(n17231), 
        .ZN(n17233) );
  NAND4_X1 U20545 ( .A1(n17235), .A2(n17234), .A3(n21273), .A4(n17233), .ZN(
        P1_U2823) );
  OAI21_X1 U20546 ( .B1(n21349), .B2(n17236), .A(n21273), .ZN(n17239) );
  OAI22_X1 U20547 ( .A1(n17363), .A2(n21296), .B1(n21308), .B2(n17237), .ZN(
        n17238) );
  AOI211_X1 U20548 ( .C1(n17292), .C2(n21339), .A(n17239), .B(n17238), .ZN(
        n17242) );
  AOI22_X1 U20549 ( .A1(n17293), .A2(n21312), .B1(n10337), .B2(
        P1_REIP_REG_13__SCAN_IN), .ZN(n17241) );
  OAI211_X1 U20550 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n17243), .A(n17242), 
        .B(n17241), .ZN(P1_U2827) );
  AOI22_X1 U20551 ( .A1(n21343), .A2(P1_EBX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n21331), .ZN(n17249) );
  INV_X1 U20552 ( .A(n17244), .ZN(n17254) );
  AOI21_X1 U20553 ( .B1(n21345), .B2(n17254), .A(n21330), .ZN(n17248) );
  INV_X1 U20554 ( .A(n17245), .ZN(n17297) );
  AOI22_X1 U20555 ( .A1(n17299), .A2(n21312), .B1(n17297), .B2(n21339), .ZN(
        n17247) );
  OAI21_X1 U20556 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n9867), .A(n10337), .ZN(
        n17246) );
  NAND4_X1 U20557 ( .A1(n17249), .A2(n17248), .A3(n17247), .A4(n17246), .ZN(
        P1_U2828) );
  INV_X1 U20558 ( .A(n17250), .ZN(n21377) );
  AOI22_X1 U20559 ( .A1(n17274), .A2(n21377), .B1(n21376), .B2(n17251), .ZN(
        n17252) );
  OAI21_X1 U20560 ( .B1(n21381), .B2(n17253), .A(n17252), .ZN(P1_U2855) );
  AOI22_X1 U20561 ( .A1(n17299), .A2(n21377), .B1(n21376), .B2(n17254), .ZN(
        n17255) );
  OAI21_X1 U20562 ( .B1(n21381), .B2(n17256), .A(n17255), .ZN(P1_U2860) );
  AOI22_X1 U20563 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n17260) );
  AOI22_X1 U20564 ( .A1(n17298), .A2(n17258), .B1(n17296), .B2(n17257), .ZN(
        n17259) );
  OAI211_X1 U20565 ( .C1(n17312), .C2(n17261), .A(n17260), .B(n17259), .ZN(
        P1_U2977) );
  AOI22_X1 U20566 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n17265) );
  AOI22_X1 U20567 ( .A1(n17263), .A2(n17298), .B1(n17267), .B2(n17262), .ZN(
        n17264) );
  OAI211_X1 U20568 ( .C1(n17305), .C2(n17266), .A(n17265), .B(n17264), .ZN(
        P1_U2978) );
  AOI22_X1 U20569 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20570 ( .A1(n17269), .A2(n17298), .B1(n17268), .B2(n17267), .ZN(
        n17270) );
  OAI211_X1 U20571 ( .C1(n17305), .C2(n17272), .A(n17271), .B(n17270), .ZN(
        P1_U2980) );
  AOI22_X1 U20572 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20573 ( .A1(n17274), .A2(n17298), .B1(n17273), .B2(n17296), .ZN(
        n17275) );
  OAI211_X1 U20574 ( .C1(n17312), .C2(n17277), .A(n17276), .B(n17275), .ZN(
        P1_U2982) );
  AOI22_X1 U20575 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20576 ( .A1(n17279), .A2(n17298), .B1(n17296), .B2(n17278), .ZN(
        n17280) );
  OAI211_X1 U20577 ( .C1(n17312), .C2(n17282), .A(n17281), .B(n17280), .ZN(
        P1_U2983) );
  AOI22_X1 U20578 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20579 ( .A1(n17284), .A2(n17298), .B1(n17296), .B2(n17283), .ZN(
        n17285) );
  OAI211_X1 U20580 ( .C1(n17287), .C2(n17312), .A(n17286), .B(n17285), .ZN(
        P1_U2984) );
  NOR2_X1 U20581 ( .A1(n17289), .A2(n17288), .ZN(n17291) );
  XOR2_X1 U20582 ( .A(n17291), .B(n17290), .Z(n17366) );
  AOI22_X1 U20583 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U20584 ( .A1(n17293), .A2(n17298), .B1(n17292), .B2(n17296), .ZN(
        n17294) );
  OAI211_X1 U20585 ( .C1(n17312), .C2(n17366), .A(n17295), .B(n17294), .ZN(
        P1_U2986) );
  AOI22_X1 U20586 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20587 ( .A1(n17299), .A2(n17298), .B1(n17297), .B2(n17296), .ZN(
        n17300) );
  OAI211_X1 U20588 ( .C1(n17302), .C2(n17312), .A(n17301), .B(n17300), .ZN(
        P1_U2987) );
  AOI22_X1 U20589 ( .A1(n14161), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n17369), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n17310) );
  INV_X1 U20590 ( .A(n17303), .ZN(n17304) );
  OAI22_X1 U20591 ( .A1(n17307), .A2(n17306), .B1(n17305), .B2(n17304), .ZN(
        n17308) );
  INV_X1 U20592 ( .A(n17308), .ZN(n17309) );
  OAI211_X1 U20593 ( .C1(n17312), .C2(n17311), .A(n17310), .B(n17309), .ZN(
        P1_U2989) );
  AOI22_X1 U20594 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n17369), .B1(n17313), 
        .B2(n17319), .ZN(n17318) );
  INV_X1 U20595 ( .A(n17314), .ZN(n17315) );
  OAI211_X1 U20596 ( .C1(n17320), .C2(n17319), .A(n17318), .B(n17317), .ZN(
        P1_U3002) );
  AOI22_X1 U20597 ( .A1(n17322), .A2(n21429), .B1(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17321), .ZN(n17330) );
  NAND2_X1 U20598 ( .A1(n17369), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n17329) );
  INV_X1 U20599 ( .A(n17323), .ZN(n17324) );
  NAND2_X1 U20600 ( .A1(n17324), .A2(n21427), .ZN(n17328) );
  OAI211_X1 U20601 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n17326), .B(n17325), .ZN(
        n17327) );
  NAND4_X1 U20602 ( .A1(n17330), .A2(n17329), .A3(n17328), .A4(n17327), .ZN(
        P1_U3003) );
  INV_X1 U20603 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21501) );
  INV_X1 U20604 ( .A(n17331), .ZN(n17334) );
  INV_X1 U20605 ( .A(n17332), .ZN(n17333) );
  AOI22_X1 U20606 ( .A1(n17334), .A2(n21429), .B1(n21427), .B2(n17333), .ZN(
        n17340) );
  NOR2_X1 U20607 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17335), .ZN(
        n17337) );
  OAI22_X1 U20608 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17338), .B1(
        n17337), .B2(n17336), .ZN(n17339) );
  OAI211_X1 U20609 ( .C1(n21501), .C2(n17352), .A(n17340), .B(n17339), .ZN(
        P1_U3005) );
  INV_X1 U20610 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17348) );
  AOI21_X1 U20611 ( .B1(n17343), .B2(n17342), .A(n17341), .ZN(n17345) );
  OAI222_X1 U20612 ( .A1(n17346), .A2(n17364), .B1(n17348), .B2(n17345), .C1(
        n17365), .C2(n17344), .ZN(n17347) );
  INV_X1 U20613 ( .A(n17347), .ZN(n17351) );
  NAND3_X1 U20614 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17349), .A3(
        n17348), .ZN(n17350) );
  OAI211_X1 U20615 ( .C1(n21497), .C2(n17352), .A(n17351), .B(n17350), .ZN(
        P1_U3007) );
  NOR2_X1 U20616 ( .A1(n17353), .A2(n17368), .ZN(n17362) );
  AOI21_X1 U20617 ( .B1(n17355), .B2(n17354), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17361) );
  INV_X1 U20618 ( .A(n17356), .ZN(n17358) );
  AOI22_X1 U20619 ( .A1(n17358), .A2(n21429), .B1(n21427), .B2(n17357), .ZN(
        n17360) );
  NAND2_X1 U20620 ( .A1(n17369), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n17359) );
  OAI211_X1 U20621 ( .C1(n17362), .C2(n17361), .A(n17360), .B(n17359), .ZN(
        P1_U3017) );
  OAI22_X1 U20622 ( .A1(n17366), .A2(n17365), .B1(n17364), .B2(n17363), .ZN(
        n17367) );
  AOI21_X1 U20623 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17368), .A(
        n17367), .ZN(n17371) );
  NAND2_X1 U20624 ( .A1(n17369), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n17370) );
  OAI211_X1 U20625 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n17372), .A(
        n17371), .B(n17370), .ZN(P1_U3018) );
  AOI21_X1 U20626 ( .B1(n21427), .B2(n17374), .A(n17373), .ZN(n17379) );
  AOI22_X1 U20627 ( .A1(n17377), .A2(n21429), .B1(n17376), .B2(n17375), .ZN(
        n17378) );
  OAI211_X1 U20628 ( .C1(n17380), .C2(n11273), .A(n17379), .B(n17378), .ZN(
        P1_U3020) );
  INV_X1 U20629 ( .A(n17381), .ZN(n21272) );
  INV_X1 U20630 ( .A(n17382), .ZN(n17383) );
  AOI21_X1 U20631 ( .B1(n21427), .B2(n21272), .A(n17383), .ZN(n17387) );
  AOI22_X1 U20632 ( .A1(n17385), .A2(n21429), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17384), .ZN(n17386) );
  OAI211_X1 U20633 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17388), .A(
        n17387), .B(n17386), .ZN(P1_U3022) );
  INV_X1 U20634 ( .A(n17389), .ZN(n17390) );
  NAND3_X1 U20635 ( .A1(n17391), .A2(n17390), .A3(n21523), .ZN(n17392) );
  OAI21_X1 U20636 ( .B1(n21526), .B2(n14114), .A(n17392), .ZN(P1_U3468) );
  NAND4_X1 U20637 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n21441), .A4(n21452), .ZN(n17393) );
  AND2_X1 U20638 ( .A1(n17394), .A2(n17393), .ZN(n21440) );
  AOI21_X1 U20639 ( .B1(n21440), .B2(n17396), .A(n17395), .ZN(n17397) );
  AOI21_X1 U20640 ( .B1(n21438), .B2(n17398), .A(n17397), .ZN(P1_U3162) );
  OAI21_X1 U20641 ( .B1(n17401), .B2(n17400), .A(n17399), .ZN(P1_U3466) );
  INV_X1 U20642 ( .A(n17402), .ZN(n17412) );
  AOI21_X1 U20643 ( .B1(n17404), .B2(n17403), .A(n21086), .ZN(n17411) );
  AOI22_X1 U20644 ( .A1(n20359), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20412), .ZN(n17405) );
  OAI21_X1 U20645 ( .B1(n20374), .B2(n21159), .A(n17405), .ZN(n17406) );
  AOI21_X1 U20646 ( .B1(n17407), .B2(n20328), .A(n17406), .ZN(n17408) );
  OAI21_X1 U20647 ( .B1(n17409), .B2(n20402), .A(n17408), .ZN(n17410) );
  OAI21_X1 U20648 ( .B1(n17414), .B2(n20401), .A(n17413), .ZN(P2_U2826) );
  AOI22_X1 U20649 ( .A1(n17415), .A2(n20328), .B1(P2_REIP_REG_28__SCAN_IN), 
        .B2(n20406), .ZN(n17426) );
  AOI22_X1 U20650 ( .A1(n20359), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20412), .ZN(n17425) );
  OAI22_X1 U20651 ( .A1(n17417), .A2(n20402), .B1(n20401), .B2(n17416), .ZN(
        n17418) );
  INV_X1 U20652 ( .A(n17418), .ZN(n17424) );
  AOI21_X1 U20653 ( .B1(n17421), .B2(n17420), .A(n17419), .ZN(n17422) );
  NAND2_X1 U20654 ( .A1(n20370), .A2(n17422), .ZN(n17423) );
  NAND4_X1 U20655 ( .A1(n17426), .A2(n17425), .A3(n17424), .A4(n17423), .ZN(
        P2_U2827) );
  INV_X1 U20656 ( .A(n17427), .ZN(n17428) );
  AOI22_X1 U20657 ( .A1(n17428), .A2(n20328), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n20359), .ZN(n17439) );
  AOI22_X1 U20658 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20412), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n20406), .ZN(n17438) );
  INV_X1 U20659 ( .A(n17429), .ZN(n17431) );
  AOI22_X1 U20660 ( .A1(n17431), .A2(n20385), .B1(n20378), .B2(n17430), .ZN(
        n17437) );
  AOI21_X1 U20661 ( .B1(n17434), .B2(n17433), .A(n17432), .ZN(n17435) );
  NAND2_X1 U20662 ( .A1(n20370), .A2(n17435), .ZN(n17436) );
  NAND4_X1 U20663 ( .A1(n17439), .A2(n17438), .A3(n17437), .A4(n17436), .ZN(
        P2_U2829) );
  AOI22_X1 U20664 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20412), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n20406), .ZN(n17440) );
  OAI21_X1 U20665 ( .B1(n20396), .B2(n17441), .A(n17440), .ZN(n17442) );
  AOI21_X1 U20666 ( .B1(n17443), .B2(n20385), .A(n17442), .ZN(n17444) );
  OAI21_X1 U20667 ( .B1(n17445), .B2(n20399), .A(n17444), .ZN(n17449) );
  AOI211_X1 U20668 ( .C1(n17447), .C2(n17446), .A(n9896), .B(n21086), .ZN(
        n17448) );
  NOR2_X1 U20669 ( .A1(n17449), .A2(n17448), .ZN(n17450) );
  OAI21_X1 U20670 ( .B1(n17451), .B2(n20401), .A(n17450), .ZN(P2_U2830) );
  AOI22_X1 U20671 ( .A1(n9834), .A2(n20328), .B1(P2_REIP_REG_24__SCAN_IN), 
        .B2(n20406), .ZN(n17463) );
  AOI22_X1 U20672 ( .A1(n20359), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20412), .ZN(n17462) );
  INV_X1 U20673 ( .A(n17452), .ZN(n17453) );
  OAI22_X1 U20674 ( .A1(n17454), .A2(n20402), .B1(n20401), .B2(n17453), .ZN(
        n17455) );
  INV_X1 U20675 ( .A(n17455), .ZN(n17461) );
  AOI21_X1 U20676 ( .B1(n17458), .B2(n17457), .A(n17456), .ZN(n17459) );
  NAND2_X1 U20677 ( .A1(n20370), .A2(n17459), .ZN(n17460) );
  NAND4_X1 U20678 ( .A1(n17463), .A2(n17462), .A3(n17461), .A4(n17460), .ZN(
        P2_U2831) );
  AOI22_X1 U20679 ( .A1(n20437), .A2(n17465), .B1(n17464), .B2(n17479), .ZN(
        P2_U2856) );
  AOI22_X1 U20680 ( .A1(n17466), .A2(n20435), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n17479), .ZN(n17467) );
  OAI21_X1 U20681 ( .B1(n17479), .B2(n17468), .A(n17467), .ZN(P2_U2864) );
  AOI21_X1 U20682 ( .B1(n17470), .B2(n16453), .A(n17469), .ZN(n17487) );
  INV_X1 U20683 ( .A(n17471), .ZN(n17472) );
  AOI22_X1 U20684 ( .A1(n17487), .A2(n20435), .B1(n13216), .B2(n17472), .ZN(
        n17473) );
  OAI21_X1 U20685 ( .B1(n20437), .B2(n17120), .A(n17473), .ZN(P2_U2865) );
  AOI21_X1 U20686 ( .B1(n17474), .B2(n9901), .A(n16455), .ZN(n17492) );
  AOI22_X1 U20687 ( .A1(n17492), .A2(n20435), .B1(n13216), .B2(n20245), .ZN(
        n17475) );
  OAI21_X1 U20688 ( .B1(n20437), .B2(n17476), .A(n17475), .ZN(P2_U2867) );
  OR2_X1 U20689 ( .A1(n9905), .A2(n17477), .ZN(n17478) );
  AND2_X1 U20690 ( .A1(n16461), .A2(n17478), .ZN(n17496) );
  NOR2_X1 U20691 ( .A1(n17480), .A2(n17479), .ZN(n17481) );
  AOI21_X1 U20692 ( .B1(n17496), .B2(n20435), .A(n17481), .ZN(n17482) );
  OAI21_X1 U20693 ( .B1(n20437), .B2(n17483), .A(n17482), .ZN(P2_U2869) );
  AOI22_X1 U20694 ( .A1(n20442), .A2(n17484), .B1(n20491), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n17490) );
  AOI22_X1 U20695 ( .A1(n20444), .A2(BUF2_REG_22__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n17489) );
  INV_X1 U20696 ( .A(n17485), .ZN(n17486) );
  AOI22_X1 U20697 ( .A1(n17487), .A2(n20477), .B1(n20492), .B2(n17486), .ZN(
        n17488) );
  NAND3_X1 U20698 ( .A1(n17490), .A2(n17489), .A3(n17488), .ZN(P2_U2897) );
  AOI22_X1 U20699 ( .A1(n20442), .A2(n17491), .B1(n20491), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n17495) );
  AOI22_X1 U20700 ( .A1(n20444), .A2(BUF2_REG_20__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U20701 ( .A1(n10332), .A2(n20492), .B1(n20477), .B2(n17492), .ZN(
        n17493) );
  NAND3_X1 U20702 ( .A1(n17495), .A2(n17494), .A3(n17493), .ZN(P2_U2899) );
  AOI22_X1 U20703 ( .A1(n20442), .A2(n20553), .B1(n20491), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U20704 ( .A1(n20444), .A2(BUF2_REG_18__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n17499) );
  AOI22_X1 U20705 ( .A1(n17497), .A2(n20492), .B1(n20477), .B2(n17496), .ZN(
        n17498) );
  NAND3_X1 U20706 ( .A1(n17500), .A2(n17499), .A3(n17498), .ZN(P2_U2901) );
  AOI22_X1 U20707 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n20376), .B1(n17582), 
        .B2(n17501), .ZN(n17510) );
  NAND2_X1 U20708 ( .A1(n17502), .A2(n17592), .ZN(n17506) );
  NAND3_X1 U20709 ( .A1(n17504), .A2(n12599), .A3(n17503), .ZN(n17505) );
  OAI211_X1 U20710 ( .C1(n17577), .C2(n17507), .A(n17506), .B(n17505), .ZN(
        n17508) );
  INV_X1 U20711 ( .A(n17508), .ZN(n17509) );
  OAI211_X1 U20712 ( .C1(n17511), .C2(n17596), .A(n17510), .B(n17509), .ZN(
        P2_U2999) );
  AOI22_X1 U20713 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17564), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n20376), .ZN(n17523) );
  NAND2_X1 U20714 ( .A1(n17512), .A2(n17601), .ZN(n17513) );
  AND2_X1 U20715 ( .A1(n17513), .A2(n12613), .ZN(n17606) );
  INV_X1 U20716 ( .A(n17606), .ZN(n17520) );
  NAND2_X1 U20717 ( .A1(n16850), .A2(n17515), .ZN(n17519) );
  AND2_X1 U20718 ( .A1(n17515), .A2(n17514), .ZN(n17516) );
  OR2_X1 U20719 ( .A1(n17517), .A2(n17516), .ZN(n17518) );
  NAND2_X1 U20720 ( .A1(n17519), .A2(n17518), .ZN(n17609) );
  OAI22_X1 U20721 ( .A1(n17520), .A2(n17566), .B1(n17609), .B2(n17572), .ZN(
        n17521) );
  AOI21_X1 U20722 ( .B1(n17591), .B2(n20269), .A(n17521), .ZN(n17522) );
  OAI211_X1 U20723 ( .C1(n17571), .C2(n20263), .A(n17523), .B(n17522), .ZN(
        P2_U3000) );
  AOI22_X1 U20724 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n20376), .B1(n17582), 
        .B2(n17524), .ZN(n17529) );
  AOI222_X1 U20725 ( .A1(n12599), .A2(n17527), .B1(n17526), .B2(n17592), .C1(
        n17591), .C2(n17525), .ZN(n17528) );
  OAI211_X1 U20726 ( .C1(n17530), .C2(n17596), .A(n17529), .B(n17528), .ZN(
        P2_U3001) );
  AOI22_X1 U20727 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17564), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n20376), .ZN(n17540) );
  AND2_X1 U20728 ( .A1(n17532), .A2(n17531), .ZN(n17533) );
  XNOR2_X1 U20729 ( .A(n9859), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17617) );
  XOR2_X1 U20730 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17535), .Z(
        n17536) );
  XNOR2_X1 U20731 ( .A(n17534), .B(n17536), .ZN(n17618) );
  AOI22_X1 U20732 ( .A1(n17617), .A2(n12599), .B1(n17592), .B2(n17618), .ZN(
        n17537) );
  INV_X1 U20733 ( .A(n17537), .ZN(n17538) );
  AOI21_X1 U20734 ( .B1(n17591), .B2(n10334), .A(n17538), .ZN(n17539) );
  OAI211_X1 U20735 ( .C1(n17571), .C2(n20274), .A(n17540), .B(n17539), .ZN(
        P2_U3002) );
  AOI22_X1 U20736 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n20376), .B1(n17582), 
        .B2(n20293), .ZN(n17545) );
  INV_X1 U20737 ( .A(n17541), .ZN(n17542) );
  AOI222_X1 U20738 ( .A1(n17543), .A2(n17592), .B1(n17591), .B2(n20294), .C1(
        n12599), .C2(n17542), .ZN(n17544) );
  OAI211_X1 U20739 ( .C1(n20287), .C2(n17596), .A(n17545), .B(n17544), .ZN(
        P2_U3003) );
  AOI22_X1 U20740 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n20376), .B1(n17582), 
        .B2(n20315), .ZN(n17549) );
  AOI222_X1 U20741 ( .A1(n17547), .A2(n12599), .B1(n17592), .B2(n17546), .C1(
        n17591), .C2(n20316), .ZN(n17548) );
  OAI211_X1 U20742 ( .C1(n20309), .C2(n17596), .A(n17549), .B(n17548), .ZN(
        P2_U3005) );
  AOI22_X1 U20743 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17564), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n20376), .ZN(n17563) );
  XOR2_X1 U20744 ( .A(n17550), .B(n17551), .Z(n17642) );
  INV_X1 U20745 ( .A(n17552), .ZN(n17554) );
  OAI21_X1 U20746 ( .B1(n17555), .B2(n17554), .A(n17553), .ZN(n17559) );
  NAND2_X1 U20747 ( .A1(n17557), .A2(n17556), .ZN(n17558) );
  XNOR2_X1 U20748 ( .A(n17559), .B(n17558), .ZN(n17640) );
  AOI22_X1 U20749 ( .A1(n17642), .A2(n12599), .B1(n17592), .B2(n17640), .ZN(
        n17560) );
  INV_X1 U20750 ( .A(n17560), .ZN(n17561) );
  AOI21_X1 U20751 ( .B1(n17591), .B2(n17641), .A(n17561), .ZN(n17562) );
  OAI211_X1 U20752 ( .C1(n17571), .C2(n20321), .A(n17563), .B(n17562), .ZN(
        P2_U3006) );
  AOI22_X1 U20753 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17564), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n20376), .ZN(n17570) );
  OAI22_X1 U20754 ( .A1(n17567), .A2(n17566), .B1(n17572), .B2(n17565), .ZN(
        n17568) );
  AOI21_X1 U20755 ( .B1(n17591), .B2(n20355), .A(n17568), .ZN(n17569) );
  OAI211_X1 U20756 ( .C1(n17571), .C2(n20353), .A(n17570), .B(n17569), .ZN(
        P2_U3008) );
  AOI22_X1 U20757 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n20376), .B1(n17582), 
        .B2(n20366), .ZN(n17580) );
  OR2_X1 U20758 ( .A1(n17573), .A2(n17572), .ZN(n17576) );
  NAND2_X1 U20759 ( .A1(n17574), .A2(n12599), .ZN(n17575) );
  OAI211_X1 U20760 ( .C1(n17577), .C2(n20367), .A(n17576), .B(n17575), .ZN(
        n17578) );
  INV_X1 U20761 ( .A(n17578), .ZN(n17579) );
  OAI211_X1 U20762 ( .C1(n20373), .C2(n17596), .A(n17580), .B(n17579), .ZN(
        P2_U3009) );
  AOI22_X1 U20763 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n20376), .B1(n17582), 
        .B2(n17581), .ZN(n17595) );
  NAND2_X1 U20764 ( .A1(n17584), .A2(n17583), .ZN(n17586) );
  XNOR2_X1 U20765 ( .A(n17586), .B(n17585), .ZN(n17667) );
  INV_X1 U20766 ( .A(n17667), .ZN(n17593) );
  INV_X1 U20767 ( .A(n17587), .ZN(n17588) );
  AND2_X1 U20768 ( .A1(n17590), .A2(n17589), .ZN(n17661) );
  AOI222_X1 U20769 ( .A1(n17593), .A2(n17592), .B1(n12599), .B2(n17661), .C1(
        n12900), .C2(n17591), .ZN(n17594) );
  OAI211_X1 U20770 ( .C1(n17597), .C2(n17596), .A(n17595), .B(n17594), .ZN(
        P2_U3011) );
  NAND2_X1 U20771 ( .A1(n17619), .A2(n17601), .ZN(n17613) );
  AOI21_X1 U20772 ( .B1(n17600), .B2(n17599), .A(n17598), .ZN(n20452) );
  AOI21_X1 U20773 ( .B1(n17603), .B2(n17602), .A(n17601), .ZN(n17605) );
  NOR2_X1 U20774 ( .A1(n20347), .A2(n12083), .ZN(n17604) );
  AOI211_X1 U20775 ( .C1(n20452), .C2(n17637), .A(n17605), .B(n17604), .ZN(
        n17612) );
  NAND2_X1 U20776 ( .A1(n12878), .A2(n20269), .ZN(n17608) );
  NAND2_X1 U20777 ( .A1(n17606), .A2(n12521), .ZN(n17607) );
  OAI211_X1 U20778 ( .C1(n17609), .C2(n17681), .A(n17608), .B(n17607), .ZN(
        n17610) );
  INV_X1 U20779 ( .A(n17610), .ZN(n17611) );
  OAI211_X1 U20780 ( .C1(n17614), .C2(n17613), .A(n17612), .B(n17611), .ZN(
        P2_U3032) );
  AOI21_X1 U20781 ( .B1(n16882), .B2(n17615), .A(n15031), .ZN(n20458) );
  AOI22_X1 U20782 ( .A1(n20458), .A2(n17637), .B1(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17616), .ZN(n17623) );
  AOI222_X1 U20783 ( .A1(n17618), .A2(n17639), .B1(n12878), .B2(n10334), .C1(
        n12521), .C2(n17617), .ZN(n17622) );
  NAND2_X1 U20784 ( .A1(n17619), .A2(n11910), .ZN(n17621) );
  NAND2_X1 U20785 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n20376), .ZN(n17620) );
  NAND4_X1 U20786 ( .A1(n17623), .A2(n17622), .A3(n17621), .A4(n17620), .ZN(
        P2_U3034) );
  NOR2_X1 U20787 ( .A1(n21128), .A2(n20347), .ZN(n17627) );
  XNOR2_X1 U20788 ( .A(n16902), .B(n17624), .ZN(n20465) );
  OAI22_X1 U20789 ( .A1(n20465), .A2(n17671), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17625), .ZN(n17626) );
  AOI211_X1 U20790 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17628), .A(
        n17627), .B(n17626), .ZN(n17631) );
  AOI22_X1 U20791 ( .A1(n17629), .A2(n12521), .B1(n12878), .B2(n20431), .ZN(
        n17630) );
  OAI211_X1 U20792 ( .C1(n17632), .C2(n17681), .A(n17631), .B(n17630), .ZN(
        P2_U3036) );
  NAND2_X1 U20793 ( .A1(n17634), .A2(n17633), .ZN(n17658) );
  OAI21_X1 U20794 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17658), .A(
        n17656), .ZN(n17638) );
  AOI21_X1 U20795 ( .B1(n17636), .B2(n17635), .A(n16901), .ZN(n20330) );
  AOI22_X1 U20796 ( .A1(n17638), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n17637), .B2(n20330), .ZN(n17648) );
  AOI222_X1 U20797 ( .A1(n17642), .A2(n12521), .B1(n12878), .B2(n17641), .C1(
        n17640), .C2(n17639), .ZN(n17647) );
  NAND2_X1 U20798 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n20376), .ZN(n17646) );
  NAND3_X1 U20799 ( .A1(n17644), .A2(n17663), .A3(n17643), .ZN(n17645) );
  NAND4_X1 U20800 ( .A1(n17648), .A2(n17647), .A3(n17646), .A4(n17645), .ZN(
        P2_U3038) );
  OAI21_X1 U20801 ( .B1(n17650), .B2(n17649), .A(n17635), .ZN(n20472) );
  OAI22_X1 U20802 ( .A1(n20472), .A2(n17671), .B1(n17672), .B2(n20342), .ZN(
        n17654) );
  OAI22_X1 U20803 ( .A1(n17652), .A2(n17669), .B1(n17651), .B2(n17681), .ZN(
        n17653) );
  AOI211_X1 U20804 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n20376), .A(n17654), .B(
        n17653), .ZN(n17655) );
  OAI221_X1 U20805 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17658), .C1(
        n17657), .C2(n17656), .A(n17655), .ZN(P2_U3039) );
  AOI22_X1 U20806 ( .A1(n13907), .A2(n12878), .B1(n20376), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n17659) );
  OAI21_X1 U20807 ( .B1(n21185), .B2(n17671), .A(n17659), .ZN(n17660) );
  AOI21_X1 U20808 ( .B1(n17661), .B2(n12521), .A(n17660), .ZN(n17666) );
  AOI22_X1 U20809 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17664), .B1(
        n17663), .B2(n17662), .ZN(n17665) );
  OAI211_X1 U20810 ( .C1(n17667), .C2(n17681), .A(n17666), .B(n17665), .ZN(
        P2_U3043) );
  OAI22_X1 U20811 ( .A1(n17670), .A2(n13684), .B1(n17669), .B2(n17668), .ZN(
        n17674) );
  OAI22_X1 U20812 ( .A1(n20403), .A2(n17672), .B1(n17671), .B2(n20400), .ZN(
        n17673) );
  OR2_X1 U20813 ( .A1(n17674), .A2(n17673), .ZN(n17677) );
  NOR2_X1 U20814 ( .A1(n17675), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17676) );
  NOR2_X1 U20815 ( .A1(n17677), .A2(n17676), .ZN(n17679) );
  OAI211_X1 U20816 ( .C1(n17681), .C2(n17680), .A(n17679), .B(n17678), .ZN(
        P2_U3046) );
  NOR2_X1 U20817 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n17682), .ZN(n21084) );
  NAND4_X1 U20818 ( .A1(n12206), .A2(n20547), .A3(n17714), .A4(n17683), .ZN(
        n17684) );
  AND2_X1 U20819 ( .A1(n17684), .A2(n21241), .ZN(n17726) );
  AOI211_X1 U20820 ( .C1(n21226), .C2(n21084), .A(n17726), .B(n17685), .ZN(
        n17734) );
  INV_X1 U20821 ( .A(n17720), .ZN(n17689) );
  AND2_X1 U20822 ( .A1(n17720), .A2(n17686), .ZN(n17687) );
  AOI21_X1 U20823 ( .B1(n17688), .B2(n17689), .A(n17687), .ZN(n17699) );
  INV_X1 U20824 ( .A(n17699), .ZN(n17724) );
  NAND2_X1 U20825 ( .A1(n17690), .A2(n17689), .ZN(n17693) );
  NAND2_X1 U20826 ( .A1(n17720), .A2(n17691), .ZN(n17692) );
  NAND2_X1 U20827 ( .A1(n17693), .A2(n17692), .ZN(n17723) );
  INV_X1 U20828 ( .A(n17695), .ZN(n17697) );
  AOI211_X1 U20829 ( .C1(n21203), .C2(n17695), .A(n21212), .B(n17694), .ZN(
        n17696) );
  AOI211_X1 U20830 ( .C1(n17697), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17720), .B(n17696), .ZN(n17698) );
  OAI21_X1 U20831 ( .B1(n17699), .B2(n21194), .A(n17698), .ZN(n17700) );
  AOI21_X1 U20832 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17723), .A(
        n17700), .ZN(n17703) );
  OAI22_X1 U20833 ( .A1(n17723), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n20619), .B2(n17724), .ZN(n17702) );
  OAI21_X1 U20834 ( .B1(n17703), .B2(n17702), .A(n17701), .ZN(n17722) );
  NAND2_X1 U20835 ( .A1(n17705), .A2(n17704), .ZN(n17711) );
  AOI22_X1 U20836 ( .A1(n17709), .A2(n17708), .B1(n17707), .B2(n17706), .ZN(
        n17710) );
  NAND2_X1 U20837 ( .A1(n17711), .A2(n17710), .ZN(n21218) );
  NAND2_X1 U20838 ( .A1(n20547), .A2(n17712), .ZN(n17718) );
  OAI21_X1 U20839 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n17713), .ZN(n17717) );
  NAND2_X1 U20840 ( .A1(n17715), .A2(n17714), .ZN(n17716) );
  OAI211_X1 U20841 ( .C1(n15199), .C2(n17718), .A(n17717), .B(n17716), .ZN(
        n17719) );
  AOI211_X1 U20842 ( .C1(n17720), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n21218), .B(n17719), .ZN(n17721) );
  OAI211_X1 U20843 ( .C1(n17724), .C2(n17723), .A(n17722), .B(n17721), .ZN(
        n17728) );
  AOI22_X1 U20844 ( .A1(n21241), .A2(n17728), .B1(n17725), .B2(n17736), .ZN(
        n17733) );
  INV_X1 U20845 ( .A(n17726), .ZN(n17727) );
  NOR2_X1 U20846 ( .A1(n17728), .A2(n17727), .ZN(n17737) );
  NOR2_X1 U20847 ( .A1(n17737), .A2(n20541), .ZN(n21083) );
  OAI21_X1 U20848 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n17730), .A(n17729), 
        .ZN(n17731) );
  OAI21_X1 U20849 ( .B1(n21083), .B2(n21236), .A(n17731), .ZN(n17732) );
  NAND3_X1 U20850 ( .A1(n17734), .A2(n17733), .A3(n17732), .ZN(P2_U3176) );
  AOI211_X1 U20851 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n17737), .A(n17736), 
        .B(n17735), .ZN(n17738) );
  INV_X1 U20852 ( .A(n17738), .ZN(P2_U3593) );
  AOI22_X1 U20853 ( .A1(n19062), .A2(n17761), .B1(n19061), .B2(n17756), .ZN(
        n17752) );
  XOR2_X1 U20854 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n9845), .Z(n17924) );
  NAND2_X1 U20855 ( .A1(n17740), .A2(n19018), .ZN(n18925) );
  OAI221_X1 U20856 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17745), .C1(
        n10128), .C2(n17744), .A(n17743), .ZN(n17746) );
  AOI211_X1 U20857 ( .C1(n19071), .C2(n17924), .A(n17747), .B(n17746), .ZN(
        n17750) );
  NAND2_X1 U20858 ( .A1(n19128), .A2(n17748), .ZN(n17749) );
  OAI211_X1 U20859 ( .C1(n17752), .C2(n17751), .A(n17750), .B(n17749), .ZN(
        P3_U2800) );
  OAI21_X1 U20860 ( .B1(n19652), .B2(n17753), .A(n17936), .ZN(n17754) );
  AOI22_X1 U20861 ( .A1(n9790), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n17755), 
        .B2(n17754), .ZN(n17766) );
  NAND2_X1 U20862 ( .A1(n19061), .A2(n17756), .ZN(n17757) );
  AOI21_X1 U20863 ( .B1(n17758), .B2(n17792), .A(n17757), .ZN(n17759) );
  AOI21_X1 U20864 ( .B1(n19128), .B2(n17760), .A(n17759), .ZN(n17765) );
  OAI211_X1 U20865 ( .C1(n17794), .C2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n19062), .B(n17761), .ZN(n17764) );
  AOI21_X1 U20866 ( .B1(n17936), .B2(n13532), .A(n9845), .ZN(n17935) );
  OAI21_X1 U20867 ( .B1(n17762), .B2(n19071), .A(n17935), .ZN(n17763) );
  NAND4_X1 U20868 ( .A1(n17766), .A2(n17765), .A3(n17764), .A4(n17763), .ZN(
        P3_U2801) );
  OAI22_X1 U20869 ( .A1(n17769), .A2(n20165), .B1(n17768), .B2(n17767), .ZN(
        n17770) );
  AOI211_X1 U20870 ( .C1(n17773), .C2(n17772), .A(n17771), .B(n17770), .ZN(
        n17777) );
  AOI22_X1 U20871 ( .A1(n19443), .A2(n17775), .B1(n19374), .B2(n17774), .ZN(
        n17776) );
  OAI211_X1 U20872 ( .C1(n17778), .C2(n19439), .A(n17777), .B(n17776), .ZN(
        P3_U2831) );
  INV_X1 U20873 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17785) );
  NAND2_X1 U20874 ( .A1(n17779), .A2(n17785), .ZN(n18860) );
  INV_X1 U20875 ( .A(n19511), .ZN(n19976) );
  AOI22_X1 U20876 ( .A1(n19976), .A2(n19405), .B1(n19407), .B2(n19381), .ZN(
        n19325) );
  NAND3_X1 U20877 ( .A1(n17781), .A2(n13477), .A3(n17780), .ZN(n19505) );
  AOI21_X1 U20878 ( .B1(n20016), .B2(n20181), .A(n19482), .ZN(n19508) );
  AOI22_X1 U20879 ( .A1(n19977), .A2(n19337), .B1(n19378), .B2(n19508), .ZN(
        n17782) );
  AOI211_X1 U20880 ( .C1(n19325), .C2(n17782), .A(n19326), .B(n19318), .ZN(
        n19290) );
  NAND2_X1 U20881 ( .A1(n17783), .A2(n19290), .ZN(n19282) );
  NOR2_X1 U20882 ( .A1(n19289), .A2(n19282), .ZN(n19269) );
  NAND2_X1 U20883 ( .A1(n19466), .A2(n19269), .ZN(n19262) );
  NOR2_X1 U20884 ( .A1(n17784), .A2(n18863), .ZN(n17789) );
  OAI22_X1 U20885 ( .A1(n19119), .A2(n17785), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n19008), .ZN(n18850) );
  INV_X1 U20886 ( .A(n18864), .ZN(n17788) );
  AOI22_X1 U20887 ( .A1(n17785), .A2(n17789), .B1(n18850), .B2(n17788), .ZN(
        n17786) );
  INV_X1 U20888 ( .A(n17786), .ZN(n17787) );
  AOI22_X1 U20889 ( .A1(n9790), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n19398), 
        .B2(n17787), .ZN(n17798) );
  NOR4_X1 U20890 ( .A1(n17790), .A2(n17789), .A3(n18849), .A4(n19983), .ZN(
        n17796) );
  INV_X1 U20891 ( .A(n19381), .ZN(n19406) );
  AOI211_X1 U20892 ( .C1(n19976), .C2(n17792), .A(n19525), .B(n17791), .ZN(
        n17793) );
  OAI21_X1 U20893 ( .B1(n17794), .B2(n19406), .A(n17793), .ZN(n17795) );
  OAI211_X1 U20894 ( .C1(n17796), .C2(n17795), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n19529), .ZN(n17797) );
  OAI211_X1 U20895 ( .C1(n18860), .C2(n19262), .A(n17798), .B(n17797), .ZN(
        P3_U2834) );
  NOR3_X1 U20896 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17800) );
  NOR4_X1 U20897 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17799) );
  NAND4_X1 U20898 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17800), .A3(n17799), .A4(
        U215), .ZN(U213) );
  INV_X1 U20899 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20501) );
  INV_X2 U20900 ( .A(U214), .ZN(n17844) );
  OAI222_X1 U20901 ( .A1(U212), .A2(n20501), .B1(n17849), .B2(n17802), .C1(
        U214), .C2(n17883), .ZN(U216) );
  INV_X2 U20902 ( .A(U212), .ZN(n17847) );
  AOI222_X1 U20903 ( .A1(n17847), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17845), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17844), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n17803) );
  INV_X1 U20904 ( .A(n17803), .ZN(U217) );
  AOI222_X1 U20905 ( .A1(n17844), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n17845), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n17847), .C2(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n17804) );
  INV_X1 U20906 ( .A(n17804), .ZN(U218) );
  AOI22_X1 U20907 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17847), .ZN(n17805) );
  OAI21_X1 U20908 ( .B1(n15657), .B2(n17849), .A(n17805), .ZN(U219) );
  INV_X1 U20909 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17807) );
  AOI22_X1 U20910 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17847), .ZN(n17806) );
  OAI21_X1 U20911 ( .B1(n17807), .B2(n17849), .A(n17806), .ZN(U220) );
  AOI22_X1 U20912 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17847), .ZN(n17808) );
  OAI21_X1 U20913 ( .B1(n15667), .B2(n17849), .A(n17808), .ZN(U221) );
  AOI22_X1 U20914 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17847), .ZN(n17809) );
  OAI21_X1 U20915 ( .B1(n15673), .B2(n17849), .A(n17809), .ZN(U222) );
  AOI22_X1 U20916 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17847), .ZN(n17810) );
  OAI21_X1 U20917 ( .B1(n15678), .B2(n17849), .A(n17810), .ZN(U223) );
  INV_X1 U20918 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20580) );
  AOI22_X1 U20919 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17847), .ZN(n17811) );
  OAI21_X1 U20920 ( .B1(n20580), .B2(n17849), .A(n17811), .ZN(U224) );
  AOI222_X1 U20921 ( .A1(n17844), .A2(P1_DATAO_REG_22__SCAN_IN), .B1(n17847), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .C1(BUF1_REG_22__SCAN_IN), .C2(n17845), 
        .ZN(n17812) );
  INV_X1 U20922 ( .A(n17812), .ZN(U225) );
  INV_X1 U20923 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n17813) );
  OAI222_X1 U20924 ( .A1(U214), .A2(n17813), .B1(U212), .B2(n17871), .C1(
        n20568), .C2(n17849), .ZN(U226) );
  AOI22_X1 U20925 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17847), .ZN(n17814) );
  OAI21_X1 U20926 ( .B1(n15700), .B2(n17849), .A(n17814), .ZN(U227) );
  AOI222_X1 U20927 ( .A1(n17844), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n17847), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .C1(BUF1_REG_19__SCAN_IN), .C2(n17845), 
        .ZN(n17815) );
  INV_X1 U20928 ( .A(n17815), .ZN(U228) );
  AOI22_X1 U20929 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17847), .ZN(n17816) );
  OAI21_X1 U20930 ( .B1(n15714), .B2(n17849), .A(n17816), .ZN(U229) );
  AOI22_X1 U20931 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17847), .ZN(n17817) );
  OAI21_X1 U20932 ( .B1(n20550), .B2(n17849), .A(n17817), .ZN(U230) );
  AOI22_X1 U20933 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17847), .ZN(n17818) );
  OAI21_X1 U20934 ( .B1(n17819), .B2(n17849), .A(n17818), .ZN(U231) );
  AOI22_X1 U20935 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17847), .ZN(n17820) );
  OAI21_X1 U20936 ( .B1(n14550), .B2(n17849), .A(n17820), .ZN(U232) );
  INV_X1 U20937 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n17822) );
  AOI22_X1 U20938 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17847), .ZN(n17821) );
  OAI21_X1 U20939 ( .B1(n17822), .B2(n17849), .A(n17821), .ZN(U233) );
  AOI222_X1 U20940 ( .A1(n17847), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n17845), 
        .B2(BUF1_REG_13__SCAN_IN), .C1(n17844), .C2(P1_DATAO_REG_13__SCAN_IN), 
        .ZN(n17823) );
  INV_X1 U20941 ( .A(n17823), .ZN(U234) );
  INV_X1 U20942 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U20943 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17847), .ZN(n17824) );
  OAI21_X1 U20944 ( .B1(n17825), .B2(n17849), .A(n17824), .ZN(U235) );
  INV_X1 U20945 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U20946 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17847), .ZN(n17826) );
  OAI21_X1 U20947 ( .B1(n17827), .B2(n17849), .A(n17826), .ZN(U236) );
  AOI22_X1 U20948 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17847), .ZN(n17828) );
  OAI21_X1 U20949 ( .B1(n17829), .B2(n17849), .A(n17828), .ZN(U237) );
  INV_X1 U20950 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n17831) );
  AOI22_X1 U20951 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17847), .ZN(n17830) );
  OAI21_X1 U20952 ( .B1(n17831), .B2(n17849), .A(n17830), .ZN(U238) );
  AOI22_X1 U20953 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17847), .ZN(n17832) );
  OAI21_X1 U20954 ( .B1(n17833), .B2(n17849), .A(n17832), .ZN(U239) );
  INV_X1 U20955 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n17835) );
  AOI22_X1 U20956 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n17847), .ZN(n17834) );
  OAI21_X1 U20957 ( .B1(n17835), .B2(n17849), .A(n17834), .ZN(U240) );
  AOI22_X1 U20958 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17847), .ZN(n17836) );
  OAI21_X1 U20959 ( .B1(n17837), .B2(n17849), .A(n17836), .ZN(U241) );
  INV_X1 U20960 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n17839) );
  AOI22_X1 U20961 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17847), .ZN(n17838) );
  OAI21_X1 U20962 ( .B1(n17839), .B2(n17849), .A(n17838), .ZN(U242) );
  AOI222_X1 U20963 ( .A1(n17844), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n17847), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .C1(BUF1_REG_4__SCAN_IN), .C2(n17845), 
        .ZN(n17840) );
  INV_X1 U20964 ( .A(n17840), .ZN(U243) );
  INV_X1 U20965 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n20535) );
  AOI22_X1 U20966 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17845), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17844), .ZN(n17841) );
  OAI21_X1 U20967 ( .B1(n20535), .B2(U212), .A(n17841), .ZN(U244) );
  AOI22_X1 U20968 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17847), .ZN(n17842) );
  OAI21_X1 U20969 ( .B1(n17843), .B2(n17849), .A(n17842), .ZN(U245) );
  INV_X1 U20970 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n17852) );
  AOI22_X1 U20971 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17845), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17844), .ZN(n17846) );
  OAI21_X1 U20972 ( .B1(n17852), .B2(U212), .A(n17846), .ZN(U246) );
  AOI22_X1 U20973 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n17844), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n17847), .ZN(n17848) );
  OAI21_X1 U20974 ( .B1(n17850), .B2(n17849), .A(n17848), .ZN(U247) );
  INV_X1 U20975 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17851) );
  AOI22_X1 U20976 ( .A1(n17881), .A2(n17851), .B1(n19547), .B2(U215), .ZN(U251) );
  INV_X1 U20977 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n19556) );
  AOI22_X1 U20978 ( .A1(n17875), .A2(n17852), .B1(n19556), .B2(U215), .ZN(U252) );
  INV_X1 U20979 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17853) );
  AOI22_X1 U20980 ( .A1(n17881), .A2(n17853), .B1(n19560), .B2(U215), .ZN(U253) );
  INV_X1 U20981 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19563) );
  AOI22_X1 U20982 ( .A1(n17881), .A2(n20535), .B1(n19563), .B2(U215), .ZN(U254) );
  INV_X1 U20983 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19567) );
  AOI22_X1 U20984 ( .A1(n17881), .A2(n20531), .B1(n19567), .B2(U215), .ZN(U255) );
  INV_X1 U20985 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17854) );
  INV_X1 U20986 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19574) );
  AOI22_X1 U20987 ( .A1(n17881), .A2(n17854), .B1(n19574), .B2(U215), .ZN(U256) );
  INV_X1 U20988 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17855) );
  AOI22_X1 U20989 ( .A1(n17881), .A2(n17855), .B1(n19577), .B2(U215), .ZN(U257) );
  OAI22_X1 U20990 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n17875), .ZN(n17856) );
  INV_X1 U20991 ( .A(n17856), .ZN(U258) );
  INV_X1 U20992 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n17857) );
  INV_X1 U20993 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18828) );
  AOI22_X1 U20994 ( .A1(n17881), .A2(n17857), .B1(n18828), .B2(U215), .ZN(U259) );
  INV_X1 U20995 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17858) );
  AOI22_X1 U20996 ( .A1(n17881), .A2(n17858), .B1(n13804), .B2(U215), .ZN(U260) );
  INV_X1 U20997 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17859) );
  INV_X1 U20998 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18831) );
  AOI22_X1 U20999 ( .A1(n17875), .A2(n17859), .B1(n18831), .B2(U215), .ZN(U261) );
  OAI22_X1 U21000 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n17881), .ZN(n17860) );
  INV_X1 U21001 ( .A(n17860), .ZN(U262) );
  INV_X1 U21002 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17861) );
  INV_X1 U21003 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18836) );
  AOI22_X1 U21004 ( .A1(n17881), .A2(n17861), .B1(n18836), .B2(U215), .ZN(U263) );
  OAI22_X1 U21005 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17881), .ZN(n17862) );
  INV_X1 U21006 ( .A(n17862), .ZN(U264) );
  INV_X1 U21007 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n17863) );
  AOI22_X1 U21008 ( .A1(n17881), .A2(n17863), .B1(n18843), .B2(U215), .ZN(U265) );
  OAI22_X1 U21009 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17875), .ZN(n17864) );
  INV_X1 U21010 ( .A(n17864), .ZN(U266) );
  INV_X1 U21011 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n17865) );
  AOI22_X1 U21012 ( .A1(n17881), .A2(n17865), .B1(n19548), .B2(U215), .ZN(U267) );
  INV_X1 U21013 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n17866) );
  INV_X1 U21014 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n20549) );
  AOI22_X1 U21015 ( .A1(n17881), .A2(n17866), .B1(n20549), .B2(U215), .ZN(U268) );
  INV_X1 U21016 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n17867) );
  INV_X1 U21017 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n20555) );
  AOI22_X1 U21018 ( .A1(n17875), .A2(n17867), .B1(n20555), .B2(U215), .ZN(U269) );
  INV_X1 U21019 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n17868) );
  AOI22_X1 U21020 ( .A1(n17881), .A2(n17869), .B1(n17868), .B2(U215), .ZN(U270) );
  INV_X1 U21021 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n17870) );
  INV_X1 U21022 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n20562) );
  AOI22_X1 U21023 ( .A1(n17875), .A2(n17870), .B1(n20562), .B2(U215), .ZN(U271) );
  INV_X1 U21024 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n20567) );
  AOI22_X1 U21025 ( .A1(n17881), .A2(n17871), .B1(n20567), .B2(U215), .ZN(U272) );
  INV_X1 U21026 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19578) );
  AOI22_X1 U21027 ( .A1(n17875), .A2(n20504), .B1(n19578), .B2(U215), .ZN(U273) );
  INV_X1 U21028 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n17872) );
  INV_X1 U21029 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n20578) );
  AOI22_X1 U21030 ( .A1(n17875), .A2(n17872), .B1(n20578), .B2(U215), .ZN(U274) );
  OAI22_X1 U21031 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17875), .ZN(n17873) );
  INV_X1 U21032 ( .A(n17873), .ZN(U275) );
  OAI22_X1 U21033 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17881), .ZN(n17874) );
  INV_X1 U21034 ( .A(n17874), .ZN(U276) );
  OAI22_X1 U21035 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17875), .ZN(n17876) );
  INV_X1 U21036 ( .A(n17876), .ZN(U277) );
  OAI22_X1 U21037 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17881), .ZN(n17877) );
  INV_X1 U21038 ( .A(n17877), .ZN(U278) );
  INV_X1 U21039 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n17878) );
  INV_X1 U21040 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18600) );
  AOI22_X1 U21041 ( .A1(n17881), .A2(n17878), .B1(n18600), .B2(U215), .ZN(U279) );
  INV_X1 U21042 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n19573) );
  AOI22_X1 U21043 ( .A1(n17881), .A2(n17879), .B1(n19573), .B2(U215), .ZN(U280) );
  INV_X1 U21044 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18587) );
  AOI22_X1 U21045 ( .A1(n17881), .A2(n17880), .B1(n18587), .B2(U215), .ZN(U281) );
  OAI22_X1 U21046 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n17881), .ZN(n17882) );
  INV_X1 U21047 ( .A(n17882), .ZN(U282) );
  INV_X1 U21048 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18731) );
  AOI222_X1 U21049 ( .A1(n18731), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(n20501), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17883), .C2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n17884) );
  INV_X2 U21050 ( .A(n17886), .ZN(n17885) );
  INV_X1 U21051 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20093) );
  INV_X1 U21052 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n21129) );
  AOI22_X1 U21053 ( .A1(n17885), .A2(n20093), .B1(n21129), .B2(n17886), .ZN(
        U347) );
  INV_X1 U21054 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20091) );
  INV_X1 U21055 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n21127) );
  AOI22_X1 U21056 ( .A1(n17885), .A2(n20091), .B1(n21127), .B2(n17886), .ZN(
        U348) );
  INV_X1 U21057 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20088) );
  INV_X1 U21058 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n21125) );
  AOI22_X1 U21059 ( .A1(n17885), .A2(n20088), .B1(n21125), .B2(n17886), .ZN(
        U349) );
  INV_X1 U21060 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20087) );
  INV_X1 U21061 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n21124) );
  AOI22_X1 U21062 ( .A1(n17885), .A2(n20087), .B1(n21124), .B2(n17886), .ZN(
        U350) );
  INV_X1 U21063 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20085) );
  INV_X1 U21064 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n21122) );
  AOI22_X1 U21065 ( .A1(n17885), .A2(n20085), .B1(n21122), .B2(n17886), .ZN(
        U351) );
  INV_X1 U21066 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20083) );
  INV_X1 U21067 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n21120) );
  AOI22_X1 U21068 ( .A1(n17885), .A2(n20083), .B1(n21120), .B2(n17886), .ZN(
        U352) );
  INV_X1 U21069 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20081) );
  INV_X1 U21070 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n21119) );
  AOI22_X1 U21071 ( .A1(n17885), .A2(n20081), .B1(n21119), .B2(n17886), .ZN(
        U353) );
  INV_X1 U21072 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n20079) );
  AOI22_X1 U21073 ( .A1(n17885), .A2(n20079), .B1(n21117), .B2(n17886), .ZN(
        U354) );
  INV_X1 U21074 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20136) );
  INV_X1 U21075 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n21162) );
  AOI22_X1 U21076 ( .A1(n17885), .A2(n20136), .B1(n21162), .B2(n17886), .ZN(
        U355) );
  INV_X1 U21077 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20133) );
  INV_X1 U21078 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n21160) );
  AOI22_X1 U21079 ( .A1(n17885), .A2(n20133), .B1(n21160), .B2(n17886), .ZN(
        U356) );
  INV_X1 U21080 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20130) );
  INV_X1 U21081 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n21158) );
  AOI22_X1 U21082 ( .A1(n17885), .A2(n20130), .B1(n21158), .B2(n17886), .ZN(
        U357) );
  INV_X1 U21083 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20127) );
  INV_X1 U21084 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n21155) );
  AOI22_X1 U21085 ( .A1(n17885), .A2(n20127), .B1(n21155), .B2(n17886), .ZN(
        U358) );
  INV_X1 U21086 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20125) );
  INV_X1 U21087 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n21154) );
  AOI22_X1 U21088 ( .A1(n17885), .A2(n20125), .B1(n21154), .B2(n17886), .ZN(
        U359) );
  INV_X1 U21089 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20123) );
  AOI22_X1 U21090 ( .A1(n17885), .A2(n20123), .B1(n21152), .B2(n17886), .ZN(
        U360) );
  INV_X1 U21091 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20121) );
  INV_X1 U21092 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n21150) );
  AOI22_X1 U21093 ( .A1(n17885), .A2(n20121), .B1(n21150), .B2(n17886), .ZN(
        U361) );
  INV_X1 U21094 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20119) );
  INV_X1 U21095 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n21149) );
  AOI22_X1 U21096 ( .A1(n17885), .A2(n20119), .B1(n21149), .B2(n17886), .ZN(
        U362) );
  INV_X1 U21097 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20117) );
  INV_X1 U21098 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n21147) );
  AOI22_X1 U21099 ( .A1(n17885), .A2(n20117), .B1(n21147), .B2(n17886), .ZN(
        U363) );
  INV_X1 U21100 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20115) );
  INV_X1 U21101 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n21146) );
  AOI22_X1 U21102 ( .A1(n17885), .A2(n20115), .B1(n21146), .B2(n17886), .ZN(
        U364) );
  INV_X1 U21103 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n20077) );
  INV_X1 U21104 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n21115) );
  AOI22_X1 U21105 ( .A1(n17885), .A2(n20077), .B1(n21115), .B2(n17886), .ZN(
        U365) );
  INV_X1 U21106 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20113) );
  INV_X1 U21107 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n21144) );
  AOI22_X1 U21108 ( .A1(n17885), .A2(n20113), .B1(n21144), .B2(n17886), .ZN(
        U366) );
  INV_X1 U21109 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20111) );
  INV_X1 U21110 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n21142) );
  AOI22_X1 U21111 ( .A1(n17885), .A2(n20111), .B1(n21142), .B2(n17886), .ZN(
        U367) );
  INV_X1 U21112 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20109) );
  INV_X1 U21113 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n21140) );
  AOI22_X1 U21114 ( .A1(n17885), .A2(n20109), .B1(n21140), .B2(n17886), .ZN(
        U368) );
  INV_X1 U21115 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20107) );
  INV_X1 U21116 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n21138) );
  AOI22_X1 U21117 ( .A1(n17885), .A2(n20107), .B1(n21138), .B2(n17886), .ZN(
        U369) );
  INV_X1 U21118 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20105) );
  INV_X1 U21119 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n21136) );
  AOI22_X1 U21120 ( .A1(n17885), .A2(n20105), .B1(n21136), .B2(n17886), .ZN(
        U370) );
  INV_X1 U21121 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20103) );
  INV_X1 U21122 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n21135) );
  AOI22_X1 U21123 ( .A1(n17885), .A2(n20103), .B1(n21135), .B2(n17886), .ZN(
        U371) );
  INV_X1 U21124 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20100) );
  INV_X1 U21125 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n21134) );
  AOI22_X1 U21126 ( .A1(n17885), .A2(n20100), .B1(n21134), .B2(n17886), .ZN(
        U372) );
  INV_X1 U21127 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20099) );
  INV_X1 U21128 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n21133) );
  AOI22_X1 U21129 ( .A1(n17885), .A2(n20099), .B1(n21133), .B2(n17886), .ZN(
        U373) );
  INV_X1 U21130 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20097) );
  INV_X1 U21131 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n21132) );
  AOI22_X1 U21132 ( .A1(n17885), .A2(n20097), .B1(n21132), .B2(n17886), .ZN(
        U374) );
  INV_X1 U21133 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n21131) );
  AOI22_X1 U21134 ( .A1(n17885), .A2(n20094), .B1(n21131), .B2(n17886), .ZN(
        U375) );
  INV_X1 U21135 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20075) );
  INV_X1 U21136 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n21113) );
  AOI22_X1 U21137 ( .A1(n17885), .A2(n20075), .B1(n21113), .B2(n17886), .ZN(
        U376) );
  INV_X1 U21138 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17887) );
  INV_X1 U21139 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n20060) );
  NOR2_X1 U21140 ( .A1(n20060), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n20062) );
  OAI22_X1 U21141 ( .A1(n20071), .A2(n20062), .B1(n20060), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n20147) );
  OAI21_X1 U21142 ( .B1(n20071), .B2(n17887), .A(n20147), .ZN(P3_U2633) );
  NAND2_X1 U21143 ( .A1(n20047), .A2(n20153), .ZN(n17889) );
  OAI21_X1 U21144 ( .B1(n17893), .B2(n18796), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17888) );
  OAI21_X1 U21145 ( .B1(n17889), .B2(n20049), .A(n17888), .ZN(P3_U2634) );
  AOI21_X1 U21146 ( .B1(n20071), .B2(n20074), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17890) );
  AOI22_X1 U21147 ( .A1(n20129), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17890), 
        .B2(n20195), .ZN(P3_U2635) );
  INV_X1 U21148 ( .A(n20147), .ZN(n20150) );
  OAI21_X1 U21149 ( .B1(n20058), .B2(BS16), .A(n20150), .ZN(n20148) );
  OAI21_X1 U21150 ( .B1(n20150), .B2(n20204), .A(n20148), .ZN(P3_U2636) );
  NOR3_X1 U21151 ( .A1(n17893), .A2(n17892), .A3(n17891), .ZN(n19984) );
  NOR2_X1 U21152 ( .A1(n19984), .A2(n20202), .ZN(n20197) );
  OAI21_X1 U21153 ( .B1(n20197), .B2(n19540), .A(n17894), .ZN(P3_U2637) );
  NOR4_X1 U21154 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n17898) );
  NOR4_X1 U21155 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17897) );
  NOR4_X1 U21156 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17896) );
  NOR4_X1 U21157 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17895) );
  NAND4_X1 U21158 ( .A1(n17898), .A2(n17897), .A3(n17896), .A4(n17895), .ZN(
        n17904) );
  NOR4_X1 U21159 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n17902) );
  AOI211_X1 U21160 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n17901) );
  NOR4_X1 U21161 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n17900) );
  NOR4_X1 U21162 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n17899) );
  NAND4_X1 U21163 ( .A1(n17902), .A2(n17901), .A3(n17900), .A4(n17899), .ZN(
        n17903) );
  NOR2_X1 U21164 ( .A1(n17904), .A2(n17903), .ZN(n20190) );
  INV_X1 U21165 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20143) );
  NOR3_X1 U21166 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17906) );
  OAI21_X1 U21167 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17906), .A(n20190), .ZN(
        n17905) );
  OAI21_X1 U21168 ( .B1(n20190), .B2(n20143), .A(n17905), .ZN(P3_U2638) );
  INV_X1 U21169 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20186) );
  INV_X1 U21170 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20149) );
  AOI21_X1 U21171 ( .B1(n20186), .B2(n20149), .A(n17906), .ZN(n17907) );
  INV_X1 U21172 ( .A(n20190), .ZN(n20193) );
  AOI22_X1 U21173 ( .A1(n20190), .A2(n17907), .B1(n20140), .B2(n20193), .ZN(
        P3_U2639) );
  INV_X1 U21174 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20137) );
  NAND4_X1 U21175 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17952), .ZN(n17916) );
  NOR3_X1 U21176 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20137), .A3(n17916), 
        .ZN(n17909) );
  AOI21_X1 U21177 ( .B1(n18248), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17909), .ZN(
        n17921) );
  INV_X1 U21178 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17959) );
  NAND2_X1 U21179 ( .A1(n17960), .A2(n17959), .ZN(n17958) );
  NOR2_X1 U21180 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17958), .ZN(n17942) );
  INV_X1 U21181 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n18318) );
  NAND2_X1 U21182 ( .A1(n17942), .A2(n18318), .ZN(n17923) );
  NOR2_X1 U21183 ( .A1(n18269), .A2(n17923), .ZN(n17930) );
  INV_X1 U21184 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n18311) );
  INV_X1 U21185 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18866) );
  NOR2_X1 U21186 ( .A1(n17912), .A2(n18866), .ZN(n17911) );
  OAI21_X1 U21187 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17911), .A(
        n13532), .ZN(n18855) );
  INV_X1 U21188 ( .A(n18855), .ZN(n17945) );
  AOI21_X1 U21189 ( .B1(n17912), .B2(n18866), .A(n17911), .ZN(n18861) );
  NOR2_X1 U21190 ( .A1(n17913), .A2(n18164), .ZN(n17954) );
  NOR2_X1 U21191 ( .A1(n18861), .A2(n17954), .ZN(n17953) );
  NOR2_X1 U21192 ( .A1(n17953), .A2(n13603), .ZN(n17944) );
  NOR2_X1 U21193 ( .A1(n17945), .A2(n17944), .ZN(n17943) );
  NOR2_X1 U21194 ( .A1(n17943), .A2(n13603), .ZN(n17934) );
  NAND2_X1 U21195 ( .A1(n18224), .A2(n18225), .ZN(n18261) );
  NOR3_X1 U21196 ( .A1(n17924), .A2(n17926), .A3(n18261), .ZN(n17919) );
  NAND3_X1 U21197 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n17915) );
  INV_X1 U21198 ( .A(n17914), .ZN(n17957) );
  AOI21_X1 U21199 ( .B1(n18243), .B2(n17915), .A(n17957), .ZN(n17937) );
  NOR2_X1 U21200 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17916), .ZN(n17928) );
  INV_X1 U21201 ( .A(n17928), .ZN(n17917) );
  AOI21_X1 U21202 ( .B1(n17937), .B2(n17917), .A(n20135), .ZN(n17918) );
  OAI211_X1 U21203 ( .C1(n17922), .C2(n18260), .A(n17921), .B(n17920), .ZN(
        P3_U2640) );
  NAND2_X1 U21204 ( .A1(n18259), .A2(n17923), .ZN(n17940) );
  OAI22_X1 U21205 ( .A1(n17937), .A2(n20137), .B1(n10128), .B2(n18260), .ZN(
        n17927) );
  OAI21_X1 U21206 ( .B1(n18248), .B2(n17930), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17931) );
  OAI211_X1 U21207 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17940), .A(n17932), .B(
        n17931), .ZN(P3_U2641) );
  NOR2_X1 U21208 ( .A1(n17942), .A2(n18318), .ZN(n17941) );
  INV_X1 U21209 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20132) );
  OAI22_X1 U21210 ( .A1(n17937), .A2(n20132), .B1(n17936), .B2(n18260), .ZN(
        n17938) );
  NAND4_X1 U21211 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17952), .A4(n20132), .ZN(n17939) );
  INV_X1 U21212 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17951) );
  AOI22_X1 U21213 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n17957), .B1(n18248), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17950) );
  INV_X1 U21214 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20126) );
  INV_X1 U21215 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20131) );
  AOI22_X1 U21216 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .B1(n20126), .B2(n20131), .ZN(n17948) );
  AOI211_X1 U21217 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17958), .A(n17942), .B(
        n18269), .ZN(n17947) );
  AOI211_X1 U21218 ( .C1(n17945), .C2(n17944), .A(n17943), .B(n20053), .ZN(
        n17946) );
  AOI211_X1 U21219 ( .C1(n17952), .C2(n17948), .A(n17947), .B(n17946), .ZN(
        n17949) );
  OAI211_X1 U21220 ( .C1(n17951), .C2(n18260), .A(n17950), .B(n17949), .ZN(
        P3_U2643) );
  INV_X1 U21221 ( .A(n17952), .ZN(n17963) );
  AOI211_X1 U21222 ( .C1(n18861), .C2(n17954), .A(n17953), .B(n20053), .ZN(
        n17956) );
  OAI22_X1 U21223 ( .A1(n18866), .A2(n18260), .B1(n18270), .B2(n17959), .ZN(
        n17955) );
  AOI211_X1 U21224 ( .C1(n17957), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17956), 
        .B(n17955), .ZN(n17962) );
  OAI211_X1 U21225 ( .C1(n17960), .C2(n17959), .A(n18259), .B(n17958), .ZN(
        n17961) );
  OAI211_X1 U21226 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17963), .A(n17962), 
        .B(n17961), .ZN(P3_U2644) );
  AOI21_X1 U21227 ( .B1(n18259), .B2(n17965), .A(n18248), .ZN(n17964) );
  INV_X1 U21228 ( .A(n17964), .ZN(n17969) );
  NOR2_X1 U21229 ( .A1(n17965), .A2(n18269), .ZN(n17977) );
  AOI211_X1 U21230 ( .C1(n18893), .C2(n17967), .A(n17966), .B(n20053), .ZN(
        n17968) );
  AOI221_X1 U21231 ( .B1(n17969), .B2(P3_EBX_REG_25__SCAN_IN), .C1(n17977), 
        .C2(n18281), .A(n17968), .ZN(n17974) );
  AOI21_X1 U21232 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17976), .A(n18263), 
        .ZN(n17971) );
  OAI22_X1 U21233 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17972), .B1(n17971), 
        .B2(n17970), .ZN(n17973) );
  OAI211_X1 U21234 ( .C1(n18260), .C2(n18891), .A(n17974), .B(n17973), .ZN(
        P3_U2646) );
  INV_X1 U21235 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18902) );
  NOR2_X1 U21236 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18263), .ZN(n17975) );
  AOI22_X1 U21237 ( .A1(n18248), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17976), 
        .B2(n17975), .ZN(n17984) );
  OAI21_X1 U21238 ( .B1(n17976), .B2(n18263), .A(n18273), .ZN(n17985) );
  INV_X1 U21239 ( .A(n17977), .ZN(n17978) );
  AOI21_X1 U21240 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17992), .A(n17978), .ZN(
        n17982) );
  AOI211_X1 U21241 ( .C1(n18905), .C2(n17980), .A(n17979), .B(n20053), .ZN(
        n17981) );
  AOI211_X1 U21242 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n17985), .A(n17982), 
        .B(n17981), .ZN(n17983) );
  OAI211_X1 U21243 ( .C1(n18902), .C2(n18260), .A(n17984), .B(n17983), .ZN(
        P3_U2647) );
  INV_X1 U21244 ( .A(n17985), .ZN(n17995) );
  AOI211_X1 U21245 ( .C1(n18916), .C2(n17987), .A(n17986), .B(n20053), .ZN(
        n17991) );
  NAND2_X1 U21246 ( .A1(n18061), .A2(n20118), .ZN(n17988) );
  OAI22_X1 U21247 ( .A1(n18888), .A2(n18260), .B1(n17989), .B2(n17988), .ZN(
        n17990) );
  AOI211_X1 U21248 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n18248), .A(n17991), .B(
        n17990), .ZN(n17994) );
  OAI211_X1 U21249 ( .C1(n17996), .C2(n18278), .A(n18259), .B(n17992), .ZN(
        n17993) );
  OAI211_X1 U21250 ( .C1(n17995), .C2(n20118), .A(n17994), .B(n17993), .ZN(
        P3_U2648) );
  AOI22_X1 U21251 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18200), .B1(
        n18248), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n18007) );
  NOR2_X1 U21252 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n18076), .ZN(n18001) );
  AOI211_X1 U21253 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n18015), .A(n17996), .B(
        n18269), .ZN(n18000) );
  AOI211_X1 U21254 ( .C1(n18938), .C2(n17998), .A(n17997), .B(n20053), .ZN(
        n17999) );
  AOI211_X1 U21255 ( .C1(n18002), .C2(n18001), .A(n18000), .B(n17999), .ZN(
        n18006) );
  NOR3_X1 U21256 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n18004), .A3(n18076), 
        .ZN(n18010) );
  INV_X1 U21257 ( .A(n18273), .ZN(n18258) );
  AOI21_X1 U21258 ( .B1(n18243), .B2(n18003), .A(n18258), .ZN(n18091) );
  INV_X1 U21259 ( .A(n18091), .ZN(n18079) );
  AOI21_X1 U21260 ( .B1(n18004), .B2(n18271), .A(n18079), .ZN(n18027) );
  INV_X1 U21261 ( .A(n18027), .ZN(n18014) );
  OAI21_X1 U21262 ( .B1(n18010), .B2(n18014), .A(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n18005) );
  NAND3_X1 U21263 ( .A1(n18007), .A2(n18006), .A3(n18005), .ZN(P3_U2649) );
  AOI211_X1 U21264 ( .C1(n18954), .C2(n18009), .A(n18008), .B(n20053), .ZN(
        n18013) );
  INV_X1 U21265 ( .A(n18010), .ZN(n18011) );
  OAI21_X1 U21266 ( .B1(n18368), .B2(n18270), .A(n18011), .ZN(n18012) );
  AOI211_X1 U21267 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n18014), .A(n18013), 
        .B(n18012), .ZN(n18017) );
  OAI211_X1 U21268 ( .C1(n18022), .C2(n18368), .A(n18259), .B(n18015), .ZN(
        n18016) );
  OAI211_X1 U21269 ( .C1(n18260), .C2(n18945), .A(n18017), .B(n18016), .ZN(
        P3_U2650) );
  INV_X1 U21270 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20112) );
  NOR2_X1 U21271 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18076), .ZN(n18018) );
  AOI22_X1 U21272 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18200), .B1(
        n18019), .B2(n18018), .ZN(n18026) );
  AOI211_X1 U21273 ( .C1(n18965), .C2(n18021), .A(n18020), .B(n20053), .ZN(
        n18024) );
  AOI211_X1 U21274 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n18035), .A(n18022), .B(
        n18269), .ZN(n18023) );
  AOI211_X1 U21275 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n18248), .A(n18024), .B(
        n18023), .ZN(n18025) );
  OAI211_X1 U21276 ( .C1(n18027), .C2(n20112), .A(n18026), .B(n18025), .ZN(
        P3_U2651) );
  AOI22_X1 U21277 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18200), .B1(
        n18248), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n18039) );
  AOI211_X1 U21278 ( .C1(n18977), .C2(n18029), .A(n18028), .B(n20053), .ZN(
        n18034) );
  AOI21_X1 U21279 ( .B1(n18031), .B2(n18271), .A(n18079), .ZN(n18049) );
  NOR2_X1 U21280 ( .A1(n18031), .A2(n18076), .ZN(n18030) );
  NAND2_X1 U21281 ( .A1(n18030), .A2(n20108), .ZN(n18047) );
  AOI21_X1 U21282 ( .B1(n18049), .B2(n18047), .A(n20110), .ZN(n18033) );
  NOR4_X1 U21283 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n20108), .A3(n18031), 
        .A4(n18076), .ZN(n18032) );
  NOR3_X1 U21284 ( .A1(n18034), .A2(n18033), .A3(n18032), .ZN(n18038) );
  OAI211_X1 U21285 ( .C1(n18042), .C2(n18036), .A(n18259), .B(n18035), .ZN(
        n18037) );
  NAND4_X1 U21286 ( .A1(n18039), .A2(n18038), .A3(n19529), .A4(n18037), .ZN(
        P3_U2652) );
  AOI211_X1 U21287 ( .C1(n18985), .C2(n18041), .A(n18040), .B(n20053), .ZN(
        n18046) );
  AOI211_X1 U21288 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n18056), .A(n18042), .B(
        n18269), .ZN(n18045) );
  INV_X1 U21289 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n18043) );
  OAI22_X1 U21290 ( .A1(n18043), .A2(n18270), .B1(n18973), .B2(n18260), .ZN(
        n18044) );
  NOR4_X1 U21291 ( .A1(n9790), .A2(n18046), .A3(n18045), .A4(n18044), .ZN(
        n18048) );
  OAI211_X1 U21292 ( .C1(n18049), .C2(n20108), .A(n18048), .B(n18047), .ZN(
        P3_U2653) );
  INV_X1 U21293 ( .A(n18049), .ZN(n18055) );
  AOI21_X1 U21294 ( .B1(n19000), .B2(n18065), .A(n18976), .ZN(n18996) );
  AND2_X1 U21295 ( .A1(n19014), .A2(n18252), .ZN(n18067) );
  AOI21_X1 U21296 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18067), .A(
        n13603), .ZN(n18051) );
  OAI21_X1 U21297 ( .B1(n18996), .B2(n18051), .A(n18225), .ZN(n18050) );
  AOI21_X1 U21298 ( .B1(n18996), .B2(n18051), .A(n18050), .ZN(n18054) );
  INV_X1 U21299 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20106) );
  NAND4_X1 U21300 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(n18061), .A4(n20106), .ZN(n18052) );
  OAI211_X1 U21301 ( .C1(n18270), .C2(n18398), .A(n19529), .B(n18052), .ZN(
        n18053) );
  AOI211_X1 U21302 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n18055), .A(n18054), 
        .B(n18053), .ZN(n18058) );
  OAI211_X1 U21303 ( .C1(n18059), .C2(n18398), .A(n18259), .B(n18056), .ZN(
        n18057) );
  OAI211_X1 U21304 ( .C1(n18260), .C2(n19000), .A(n18058), .B(n18057), .ZN(
        P3_U2654) );
  INV_X1 U21305 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20104) );
  AOI211_X1 U21306 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18080), .A(n18059), .B(
        n18269), .ZN(n18064) );
  INV_X1 U21307 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n18397) );
  NAND2_X1 U21308 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n18060) );
  OAI211_X1 U21309 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(P3_REIP_REG_16__SCAN_IN), .A(n18061), .B(n18060), .ZN(n18062) );
  OAI211_X1 U21310 ( .C1(n18270), .C2(n18397), .A(n19529), .B(n18062), .ZN(
        n18063) );
  AOI211_X1 U21311 ( .C1(n18200), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n18064), .B(n18063), .ZN(n18071) );
  OAI21_X1 U21312 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18066), .A(
        n18065), .ZN(n19016) );
  INV_X1 U21313 ( .A(n19016), .ZN(n18069) );
  NOR2_X1 U21314 ( .A1(n18067), .A2(n18164), .ZN(n18074) );
  INV_X1 U21315 ( .A(n18074), .ZN(n18068) );
  OAI221_X1 U21316 ( .B1(n18069), .B2(n18074), .C1(n19016), .C2(n18068), .A(
        n18225), .ZN(n18070) );
  OAI211_X1 U21317 ( .C1(n18091), .C2(n20104), .A(n18071), .B(n18070), .ZN(
        P3_U2655) );
  AOI21_X1 U21318 ( .B1(n18224), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n20053), .ZN(n18266) );
  OAI21_X1 U21319 ( .B1(n18073), .B2(n18164), .A(n18266), .ZN(n18084) );
  OAI21_X1 U21320 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19012), .A(
        n18072), .ZN(n19022) );
  OAI22_X1 U21321 ( .A1(n18073), .A2(n18260), .B1(n18270), .B2(n18081), .ZN(
        n18078) );
  NAND3_X1 U21322 ( .A1(n18225), .A2(n18074), .A3(n19022), .ZN(n18075) );
  OAI211_X1 U21323 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n18076), .A(n18075), 
        .B(n19529), .ZN(n18077) );
  AOI211_X1 U21324 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n18079), .A(n18078), 
        .B(n18077), .ZN(n18083) );
  OAI211_X1 U21325 ( .C1(n18085), .C2(n18081), .A(n18259), .B(n18080), .ZN(
        n18082) );
  OAI211_X1 U21326 ( .C1(n18084), .C2(n19022), .A(n18083), .B(n18082), .ZN(
        P3_U2656) );
  AOI211_X1 U21327 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n18105), .A(n18085), .B(
        n18269), .ZN(n18094) );
  AOI21_X1 U21328 ( .B1(n18243), .B2(n18086), .A(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n18092) );
  INV_X1 U21329 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18088) );
  INV_X1 U21330 ( .A(n18087), .ZN(n19049) );
  NOR2_X1 U21331 ( .A1(n19208), .A2(n19049), .ZN(n19051) );
  NAND2_X1 U21332 ( .A1(n19053), .A2(n19051), .ZN(n18097) );
  AOI21_X1 U21333 ( .B1(n18088), .B2(n18097), .A(n19012), .ZN(n19036) );
  INV_X1 U21334 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18262) );
  NAND3_X1 U21335 ( .A1(n19053), .A2(n19051), .A3(n18262), .ZN(n18098) );
  NAND2_X1 U21336 ( .A1(n18224), .A2(n18098), .ZN(n18089) );
  XOR2_X1 U21337 ( .A(n19036), .B(n18089), .Z(n18090) );
  OAI22_X1 U21338 ( .A1(n18092), .A2(n18091), .B1(n20053), .B2(n18090), .ZN(
        n18093) );
  AOI211_X1 U21339 ( .C1(n18200), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n18094), .B(n18093), .ZN(n18095) );
  OAI211_X1 U21340 ( .C1(n18270), .C2(n10073), .A(n18095), .B(n19529), .ZN(
        P3_U2657) );
  NOR3_X1 U21341 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n18263), .A3(n18096), 
        .ZN(n18104) );
  OAI21_X1 U21342 ( .B1(n18263), .B2(n18112), .A(n18273), .ZN(n18120) );
  NOR2_X1 U21343 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18263), .ZN(n18111) );
  OAI21_X1 U21344 ( .B1(n18120), .B2(n18111), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n18102) );
  INV_X1 U21345 ( .A(n18261), .ZN(n18251) );
  INV_X1 U21346 ( .A(n19051), .ZN(n18123) );
  NOR2_X1 U21347 ( .A1(n19055), .A2(n18123), .ZN(n18113) );
  OAI21_X1 U21348 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18113), .A(
        n18097), .ZN(n19066) );
  NAND3_X1 U21349 ( .A1(n18251), .A2(n19066), .A3(n18098), .ZN(n18101) );
  INV_X1 U21350 ( .A(n19066), .ZN(n18099) );
  OAI211_X1 U21351 ( .C1(n19054), .C2(n18164), .A(n18099), .B(n18266), .ZN(
        n18100) );
  NAND4_X1 U21352 ( .A1(n19529), .A2(n18102), .A3(n18101), .A4(n18100), .ZN(
        n18103) );
  AOI211_X1 U21353 ( .C1(n18200), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n18104), .B(n18103), .ZN(n18107) );
  OAI211_X1 U21354 ( .C1(n18109), .C2(n18108), .A(n18259), .B(n18105), .ZN(
        n18106) );
  OAI211_X1 U21355 ( .C1(n18270), .C2(n18108), .A(n18107), .B(n18106), .ZN(
        P3_U2658) );
  AOI22_X1 U21356 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18200), .B1(
        n18248), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n18118) );
  AOI211_X1 U21357 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n18129), .A(n18109), .B(
        n18269), .ZN(n18110) );
  AOI211_X1 U21358 ( .C1(n18112), .C2(n18111), .A(n9790), .B(n18110), .ZN(
        n18117) );
  AOI21_X1 U21359 ( .B1(n19055), .B2(n18123), .A(n18113), .ZN(n19070) );
  OAI21_X1 U21360 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18123), .A(
        n18224), .ZN(n18114) );
  XNOR2_X1 U21361 ( .A(n19070), .B(n18114), .ZN(n18115) );
  AOI22_X1 U21362 ( .A1(n18225), .A2(n18115), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n18120), .ZN(n18116) );
  NAND3_X1 U21363 ( .A1(n18118), .A2(n18117), .A3(n18116), .ZN(P3_U2659) );
  INV_X1 U21364 ( .A(n18133), .ZN(n18119) );
  NOR2_X1 U21365 ( .A1(n18263), .A2(n18158), .ZN(n18154) );
  AOI21_X1 U21366 ( .B1(n18119), .B2(n18154), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n18127) );
  INV_X1 U21367 ( .A(n18120), .ZN(n18126) );
  NOR3_X1 U21368 ( .A1(n19208), .A2(n18121), .A3(n19148), .ZN(n18146) );
  AND2_X1 U21369 ( .A1(n18122), .A2(n18146), .ZN(n18137) );
  OAI21_X1 U21370 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18137), .A(
        n18123), .ZN(n19083) );
  AOI21_X1 U21371 ( .B1(n18137), .B2(n18262), .A(n18164), .ZN(n18124) );
  XOR2_X1 U21372 ( .A(n19083), .B(n18124), .Z(n18125) );
  OAI22_X1 U21373 ( .A1(n18127), .A2(n18126), .B1(n20053), .B2(n18125), .ZN(
        n18128) );
  AOI211_X1 U21374 ( .C1(n18248), .C2(P3_EBX_REG_11__SCAN_IN), .A(n9790), .B(
        n18128), .ZN(n18131) );
  OAI211_X1 U21375 ( .C1(n18132), .C2(n18484), .A(n18259), .B(n18129), .ZN(
        n18130) );
  OAI211_X1 U21376 ( .C1(n18260), .C2(n19035), .A(n18131), .B(n18130), .ZN(
        P3_U2660) );
  AOI21_X1 U21377 ( .B1(n18243), .B2(n18158), .A(n18258), .ZN(n18169) );
  INV_X1 U21378 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20092) );
  AOI211_X1 U21379 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n18144), .A(n18132), .B(
        n18269), .ZN(n18136) );
  OAI211_X1 U21380 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n18154), .B(n18133), .ZN(n18134) );
  OAI211_X1 U21381 ( .C1(n18510), .C2(n18270), .A(n19529), .B(n18134), .ZN(
        n18135) );
  AOI211_X1 U21382 ( .C1(n18200), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18136), .B(n18135), .ZN(n18142) );
  INV_X1 U21383 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19136) );
  INV_X1 U21384 ( .A(n18146), .ZN(n18186) );
  NOR2_X1 U21385 ( .A1(n19136), .A2(n18186), .ZN(n18171) );
  NAND3_X1 U21386 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(n18171), .ZN(n18147) );
  AOI21_X1 U21387 ( .B1(n18138), .B2(n18147), .A(n18137), .ZN(n19099) );
  OAI21_X1 U21388 ( .B1(n18147), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18224), .ZN(n18139) );
  INV_X1 U21389 ( .A(n18139), .ZN(n18149) );
  AOI21_X1 U21390 ( .B1(n19099), .B2(n18149), .A(n20053), .ZN(n18140) );
  OAI21_X1 U21391 ( .B1(n19099), .B2(n18149), .A(n18140), .ZN(n18141) );
  OAI211_X1 U21392 ( .C1(n18169), .C2(n20092), .A(n18142), .B(n18141), .ZN(
        P3_U2661) );
  INV_X1 U21393 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20090) );
  INV_X1 U21394 ( .A(n18157), .ZN(n18143) );
  AOI21_X1 U21395 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18143), .A(n18269), .ZN(
        n18145) );
  AOI22_X1 U21396 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18200), .B1(
        n18145), .B2(n18144), .ZN(n18156) );
  NAND3_X1 U21397 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(n18146), .ZN(n18163) );
  INV_X1 U21398 ( .A(n18163), .ZN(n18150) );
  OAI21_X1 U21399 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18150), .A(
        n18147), .ZN(n19106) );
  NAND2_X1 U21400 ( .A1(n18225), .A2(n13603), .ZN(n18255) );
  OAI22_X1 U21401 ( .A1(n18270), .A2(n18148), .B1(n19106), .B2(n18255), .ZN(
        n18153) );
  OAI221_X1 U21402 ( .B1(n19106), .B2(n18150), .C1(n19106), .C2(n18262), .A(
        n18149), .ZN(n18151) );
  OAI21_X1 U21403 ( .B1(n20053), .B2(n18151), .A(n19529), .ZN(n18152) );
  AOI211_X1 U21404 ( .C1(n18154), .C2(n20090), .A(n18153), .B(n18152), .ZN(
        n18155) );
  OAI211_X1 U21405 ( .C1(n18169), .C2(n20090), .A(n18156), .B(n18155), .ZN(
        P3_U2662) );
  INV_X1 U21406 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20089) );
  AOI211_X1 U21407 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n18178), .A(n18157), .B(
        n18269), .ZN(n18162) );
  INV_X1 U21408 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n18546) );
  NAND3_X1 U21409 ( .A1(n18159), .A2(n18243), .A3(n18158), .ZN(n18160) );
  OAI211_X1 U21410 ( .C1(n18270), .C2(n18546), .A(n19529), .B(n18160), .ZN(
        n18161) );
  AOI211_X1 U21411 ( .C1(n18200), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n18162), .B(n18161), .ZN(n18168) );
  OAI21_X1 U21412 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18171), .A(
        n18163), .ZN(n18165) );
  INV_X1 U21413 ( .A(n18165), .ZN(n19120) );
  AOI21_X1 U21414 ( .B1(n18262), .B2(n18171), .A(n18164), .ZN(n18166) );
  INV_X1 U21415 ( .A(n18166), .ZN(n18173) );
  OAI221_X1 U21416 ( .B1(n19120), .B2(n18166), .C1(n18165), .C2(n18173), .A(
        n18225), .ZN(n18167) );
  OAI211_X1 U21417 ( .C1(n18169), .C2(n20089), .A(n18168), .B(n18167), .ZN(
        P3_U2663) );
  AOI21_X1 U21418 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18200), .A(
        n9790), .ZN(n18182) );
  AOI21_X1 U21419 ( .B1(n18170), .B2(n18252), .A(n13603), .ZN(n18188) );
  AOI21_X1 U21420 ( .B1(n19136), .B2(n18186), .A(n18171), .ZN(n19140) );
  INV_X1 U21421 ( .A(n19140), .ZN(n18172) );
  AOI221_X1 U21422 ( .B1(n18188), .B2(n19140), .C1(n18173), .C2(n18172), .A(
        n20053), .ZN(n18176) );
  NOR3_X1 U21423 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n18263), .A3(n18174), .ZN(
        n18175) );
  AOI211_X1 U21424 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n18248), .A(n18176), .B(
        n18175), .ZN(n18181) );
  INV_X1 U21425 ( .A(n18177), .ZN(n18201) );
  NOR3_X1 U21426 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18263), .A3(n18201), .ZN(
        n18183) );
  OAI21_X1 U21427 ( .B1(n18177), .B2(n18263), .A(n18273), .ZN(n18206) );
  OAI21_X1 U21428 ( .B1(n18183), .B2(n18206), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n18180) );
  OAI211_X1 U21429 ( .C1(n18184), .C2(n18549), .A(n18259), .B(n18178), .ZN(
        n18179) );
  NAND4_X1 U21430 ( .A1(n18182), .A2(n18181), .A3(n18180), .A4(n18179), .ZN(
        P3_U2664) );
  AOI21_X1 U21431 ( .B1(n18200), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n18183), .ZN(n18192) );
  AOI211_X1 U21432 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18198), .A(n18184), .B(
        n18269), .ZN(n18185) );
  AOI211_X1 U21433 ( .C1(n18248), .C2(P3_EBX_REG_6__SCAN_IN), .A(n9790), .B(
        n18185), .ZN(n18191) );
  NOR2_X1 U21434 ( .A1(n19208), .A2(n18121), .ZN(n18195) );
  OAI21_X1 U21435 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18195), .A(
        n18186), .ZN(n19149) );
  AOI21_X1 U21436 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18255), .A(
        n19149), .ZN(n18187) );
  AOI22_X1 U21437 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18206), .B1(n18266), 
        .B2(n18187), .ZN(n18190) );
  NAND3_X1 U21438 ( .A1(n18225), .A2(n18188), .A3(n19149), .ZN(n18189) );
  NAND4_X1 U21439 ( .A1(n18192), .A2(n18191), .A3(n18190), .A4(n18189), .ZN(
        P3_U2665) );
  INV_X1 U21440 ( .A(n18193), .ZN(n18194) );
  INV_X1 U21441 ( .A(n18252), .ZN(n18215) );
  OAI21_X1 U21442 ( .B1(n18194), .B2(n18215), .A(n18224), .ZN(n18216) );
  NOR2_X1 U21443 ( .A1(n19208), .A2(n18194), .ZN(n18210) );
  INV_X1 U21444 ( .A(n18195), .ZN(n18196) );
  OAI21_X1 U21445 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18210), .A(
        n18196), .ZN(n19162) );
  XNOR2_X1 U21446 ( .A(n18216), .B(n19162), .ZN(n18209) );
  INV_X1 U21447 ( .A(n18211), .ZN(n18197) );
  AOI21_X1 U21448 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18197), .A(n18269), .ZN(
        n18199) );
  AOI22_X1 U21449 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n18200), .B1(
        n18199), .B2(n18198), .ZN(n18208) );
  NAND2_X1 U21450 ( .A1(n18243), .A2(n18201), .ZN(n18202) );
  OAI22_X1 U21451 ( .A1(n18270), .A2(n18204), .B1(n18203), .B2(n18202), .ZN(
        n18205) );
  AOI211_X1 U21452 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n18206), .A(n9790), .B(
        n18205), .ZN(n18207) );
  OAI211_X1 U21453 ( .C1(n20053), .C2(n18209), .A(n18208), .B(n18207), .ZN(
        P3_U2666) );
  NOR2_X1 U21454 ( .A1(n18732), .A2(n20216), .ZN(n18241) );
  AOI221_X1 U21455 ( .B1(n17067), .B2(n18241), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18241), .A(n9790), .ZN(
        n18222) );
  INV_X1 U21456 ( .A(n18255), .ZN(n18214) );
  NAND2_X1 U21457 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10117), .ZN(
        n18223) );
  AOI21_X1 U21458 ( .B1(n19178), .B2(n18223), .A(n18210), .ZN(n19175) );
  AOI211_X1 U21459 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18233), .A(n18211), .B(
        n18269), .ZN(n18213) );
  OAI22_X1 U21460 ( .A1(n19178), .A2(n18260), .B1(n18270), .B2(n18561), .ZN(
        n18212) );
  AOI211_X1 U21461 ( .C1(n18214), .C2(n19175), .A(n18213), .B(n18212), .ZN(
        n18221) );
  NAND2_X1 U21462 ( .A1(n10117), .A2(n19178), .ZN(n19169) );
  OAI22_X1 U21463 ( .A1(n19175), .A2(n18216), .B1(n18215), .B2(n19169), .ZN(
        n18217) );
  OAI21_X1 U21464 ( .B1(n18218), .B2(n18263), .A(n18273), .ZN(n18232) );
  AOI22_X1 U21465 ( .A1(n18225), .A2(n18217), .B1(P3_REIP_REG_4__SCAN_IN), 
        .B2(n18232), .ZN(n18220) );
  INV_X1 U21466 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20080) );
  NAND3_X1 U21467 ( .A1(n18243), .A2(n18218), .A3(n20080), .ZN(n18219) );
  NAND4_X1 U21468 ( .A1(n18222), .A2(n18221), .A3(n18220), .A4(n18219), .ZN(
        P3_U2667) );
  INV_X1 U21469 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18237) );
  OAI21_X1 U21470 ( .B1(n18263), .B2(n18242), .A(n20078), .ZN(n18231) );
  INV_X1 U21471 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19198) );
  NOR2_X1 U21472 ( .A1(n19208), .A2(n19198), .ZN(n18249) );
  OAI21_X1 U21473 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18249), .A(
        n18223), .ZN(n19186) );
  INV_X1 U21474 ( .A(n18249), .ZN(n18238) );
  OAI21_X1 U21475 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18238), .A(
        n18224), .ZN(n18227) );
  OAI21_X1 U21476 ( .B1(n19186), .B2(n18227), .A(n18225), .ZN(n18226) );
  AOI21_X1 U21477 ( .B1(n19186), .B2(n18227), .A(n18226), .ZN(n18230) );
  INV_X1 U21478 ( .A(n18241), .ZN(n18276) );
  NOR2_X1 U21479 ( .A1(n20169), .A2(n20177), .ZN(n20005) );
  INV_X1 U21480 ( .A(n20005), .ZN(n19989) );
  NOR2_X1 U21481 ( .A1(n20184), .A2(n19989), .ZN(n18228) );
  OAI21_X1 U21482 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18228), .A(
        n13389), .ZN(n20155) );
  OAI22_X1 U21483 ( .A1(n18270), .A2(n18234), .B1(n18276), .B2(n20155), .ZN(
        n18229) );
  AOI211_X1 U21484 ( .C1(n18232), .C2(n18231), .A(n18230), .B(n18229), .ZN(
        n18236) );
  OAI211_X1 U21485 ( .C1(n18239), .C2(n18234), .A(n18259), .B(n18233), .ZN(
        n18235) );
  OAI211_X1 U21486 ( .C1(n18260), .C2(n18237), .A(n18236), .B(n18235), .ZN(
        P3_U2668) );
  OAI21_X1 U21487 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18238), .ZN(n19195) );
  NOR2_X1 U21488 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18257) );
  INV_X1 U21489 ( .A(n18257), .ZN(n18240) );
  AOI211_X1 U21490 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18240), .A(n18239), .B(
        n18269), .ZN(n18247) );
  AOI22_X1 U21491 ( .A1(n20005), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20169), .B2(n20006), .ZN(n20166) );
  AOI22_X1 U21492 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18258), .B1(n20166), 
        .B2(n18241), .ZN(n18245) );
  OAI211_X1 U21493 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n18243), .B(n18242), .ZN(n18244) );
  OAI211_X1 U21494 ( .C1(n18260), .C2(n19198), .A(n18245), .B(n18244), .ZN(
        n18246) );
  AOI211_X1 U21495 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18248), .A(n18247), .B(
        n18246), .ZN(n18254) );
  NAND2_X1 U21496 ( .A1(n18249), .A2(n18262), .ZN(n18250) );
  OAI211_X1 U21497 ( .C1(n18252), .C2(n19195), .A(n18251), .B(n18250), .ZN(
        n18253) );
  OAI211_X1 U21498 ( .C1(n18255), .C2(n19195), .A(n18254), .B(n18253), .ZN(
        P3_U2669) );
  NAND2_X1 U21499 ( .A1(n18256), .A2(n20006), .ZN(n20170) );
  AOI21_X1 U21500 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n18257), .ZN(n18574) );
  AOI22_X1 U21501 ( .A1(n18259), .A2(n18574), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n18258), .ZN(n18268) );
  OAI21_X1 U21502 ( .B1(n18262), .B2(n18261), .A(n18260), .ZN(n18265) );
  INV_X1 U21503 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18576) );
  OAI22_X1 U21504 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18263), .B1(n18270), 
        .B2(n18576), .ZN(n18264) );
  AOI221_X1 U21505 ( .B1(n18266), .B2(n19208), .C1(n18265), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n18264), .ZN(n18267) );
  OAI211_X1 U21506 ( .C1(n20170), .C2(n18276), .A(n18268), .B(n18267), .ZN(
        P3_U2670) );
  NAND2_X1 U21507 ( .A1(n18270), .A2(n18269), .ZN(n18272) );
  AOI22_X1 U21508 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n18272), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n18271), .ZN(n18275) );
  NAND3_X1 U21509 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20154), .A3(
        n18273), .ZN(n18274) );
  OAI211_X1 U21510 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18276), .A(
        n18275), .B(n18274), .ZN(P3_U2671) );
  NOR4_X1 U21511 ( .A1(n18279), .A2(n18278), .A3(n18277), .A4(n18368), .ZN(
        n18284) );
  NAND2_X1 U21512 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n18280) );
  NOR4_X1 U21513 ( .A1(n18318), .A2(n18282), .A3(n18281), .A4(n18280), .ZN(
        n18283) );
  NAND4_X1 U21514 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18396), .A3(n18284), 
        .A4(n18283), .ZN(n18312) );
  NOR2_X1 U21515 ( .A1(n18311), .A2(n18312), .ZN(n18310) );
  NAND2_X1 U21516 ( .A1(n18570), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18286) );
  NAND2_X1 U21517 ( .A1(n18310), .A2(n19584), .ZN(n18285) );
  OAI22_X1 U21518 ( .A1(n18310), .A2(n18286), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18285), .ZN(P3_U2672) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18520), .B1(
        n9794), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18297) );
  AOI22_X1 U21520 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U21521 ( .A1(n13259), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18287) );
  OAI21_X1 U21522 ( .B1(n18288), .B2(n9787), .A(n18287), .ZN(n18294) );
  AOI22_X1 U21523 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18292) );
  AOI22_X1 U21524 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9817), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18291) );
  AOI22_X1 U21525 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18290) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n9793), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18289) );
  NAND4_X1 U21527 ( .A1(n18292), .A2(n18291), .A3(n18290), .A4(n18289), .ZN(
        n18293) );
  AOI211_X1 U21528 ( .C1(n18498), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n18294), .B(n18293), .ZN(n18295) );
  AND3_X1 U21529 ( .A1(n18297), .A2(n18296), .A3(n18295), .ZN(n18316) );
  OR3_X1 U21530 ( .A1(n18315), .A2(n18322), .A3(n18316), .ZN(n18309) );
  AOI22_X1 U21531 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n18520), .ZN(n18301) );
  AOI22_X1 U21532 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9793), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18300) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18534), .B1(
        n18503), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18299) );
  AOI22_X1 U21534 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18298) );
  NAND4_X1 U21535 ( .A1(n18301), .A2(n18300), .A3(n18299), .A4(n18298), .ZN(
        n18307) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17066), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n9817), .ZN(n18305) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17067), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n18518), .ZN(n18304) );
  AOI22_X1 U21538 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n18513), .ZN(n18303) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13311), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n18533), .ZN(n18302) );
  NAND4_X1 U21540 ( .A1(n18305), .A2(n18304), .A3(n18303), .A4(n18302), .ZN(
        n18306) );
  NOR2_X1 U21541 ( .A1(n18307), .A2(n18306), .ZN(n18308) );
  XNOR2_X1 U21542 ( .A(n18309), .B(n18308), .ZN(n18588) );
  AOI21_X1 U21543 ( .B1(n18312), .B2(n18311), .A(n18310), .ZN(n18313) );
  NAND2_X1 U21544 ( .A1(n18570), .A2(n18313), .ZN(n18314) );
  OAI21_X1 U21545 ( .B1(n18588), .B2(n18570), .A(n18314), .ZN(P3_U2673) );
  NOR2_X1 U21546 ( .A1(n18322), .A2(n18315), .ZN(n18317) );
  XOR2_X1 U21547 ( .A(n18317), .B(n18316), .Z(n18595) );
  AOI22_X1 U21548 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n18320), .B1(n18319), 
        .B2(n18318), .ZN(n18321) );
  OAI21_X1 U21549 ( .B1(n18570), .B2(n18595), .A(n18321), .ZN(P3_U2674) );
  OAI21_X1 U21550 ( .B1(n18324), .B2(n18323), .A(n18322), .ZN(n18605) );
  NAND3_X1 U21551 ( .A1(n18326), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18570), 
        .ZN(n18325) );
  OAI221_X1 U21552 ( .B1(n18326), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18570), 
        .C2(n18605), .A(n18325), .ZN(P3_U2676) );
  AOI21_X1 U21553 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18570), .A(n18334), .ZN(
        n18330) );
  OAI21_X1 U21554 ( .B1(n18329), .B2(n18328), .A(n18327), .ZN(n18609) );
  OAI22_X1 U21555 ( .A1(n18331), .A2(n18330), .B1(n18570), .B2(n18609), .ZN(
        P3_U2677) );
  AOI21_X1 U21556 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18570), .A(n18340), .ZN(
        n18333) );
  XNOR2_X1 U21557 ( .A(n18332), .B(n18336), .ZN(n18613) );
  OAI22_X1 U21558 ( .A1(n18334), .A2(n18333), .B1(n18570), .B2(n18613), .ZN(
        P3_U2678) );
  INV_X1 U21559 ( .A(n18335), .ZN(n18345) );
  AOI21_X1 U21560 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18570), .A(n18345), .ZN(
        n18339) );
  OAI21_X1 U21561 ( .B1(n18338), .B2(n18337), .A(n18336), .ZN(n18618) );
  OAI22_X1 U21562 ( .A1(n18340), .A2(n18339), .B1(n18570), .B2(n18618), .ZN(
        P3_U2679) );
  AOI21_X1 U21563 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18570), .A(n18341), .ZN(
        n18344) );
  XNOR2_X1 U21564 ( .A(n18343), .B(n18342), .ZN(n18623) );
  OAI22_X1 U21565 ( .A1(n18345), .A2(n18344), .B1(n18570), .B2(n18623), .ZN(
        P3_U2680) );
  AOI22_X1 U21566 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18349) );
  AOI22_X1 U21567 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18503), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18348) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n17066), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18347) );
  AOI22_X1 U21569 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18346) );
  NAND4_X1 U21570 ( .A1(n18349), .A2(n18348), .A3(n18347), .A4(n18346), .ZN(
        n18355) );
  AOI22_X1 U21571 ( .A1(n13259), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18353) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18455), .B1(
        P3_INSTQUEUE_REG_10__6__SCAN_IN), .B2(n18518), .ZN(n18352) );
  AOI22_X1 U21573 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18351) );
  AOI22_X1 U21574 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18350) );
  NAND4_X1 U21575 ( .A1(n18353), .A2(n18352), .A3(n18351), .A4(n18350), .ZN(
        n18354) );
  NOR2_X1 U21576 ( .A1(n18355), .A2(n18354), .ZN(n18627) );
  NAND3_X1 U21577 ( .A1(n18357), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n18570), 
        .ZN(n18356) );
  OAI221_X1 U21578 ( .B1(n18357), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n18570), 
        .C2(n18627), .A(n18356), .ZN(P3_U2681) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n17067), .B1(
        n18503), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18361) );
  AOI22_X1 U21580 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9817), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18360) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n13259), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18359) );
  AOI22_X1 U21582 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18358) );
  NAND4_X1 U21583 ( .A1(n18361), .A2(n18360), .A3(n18359), .A4(n18358), .ZN(
        n18367) );
  AOI22_X1 U21584 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18365) );
  AOI22_X1 U21585 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18364) );
  AOI22_X1 U21586 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18363) );
  AOI22_X1 U21587 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18362) );
  NAND4_X1 U21588 ( .A1(n18365), .A2(n18364), .A3(n18363), .A4(n18362), .ZN(
        n18366) );
  NOR2_X1 U21589 ( .A1(n18367), .A2(n18366), .ZN(n18633) );
  AOI21_X1 U21590 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18396), .A(n18579), .ZN(
        n18381) );
  AOI22_X1 U21591 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18381), .B1(n18369), 
        .B2(n18368), .ZN(n18370) );
  OAI21_X1 U21592 ( .B1(n18633), .B2(n18570), .A(n18370), .ZN(P3_U2682) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9795), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18374) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18539), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U21595 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18372) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18534), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18371) );
  NAND4_X1 U21597 ( .A1(n18374), .A2(n18373), .A3(n18372), .A4(n18371), .ZN(
        n18380) );
  AOI22_X1 U21598 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18378) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18518), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18377) );
  AOI22_X1 U21600 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18376) );
  AOI22_X1 U21601 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9794), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18375) );
  NAND4_X1 U21602 ( .A1(n18378), .A2(n18377), .A3(n18376), .A4(n18375), .ZN(
        n18379) );
  NOR2_X1 U21603 ( .A1(n18380), .A2(n18379), .ZN(n18640) );
  OAI21_X1 U21604 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18382), .A(n18381), .ZN(
        n18383) );
  OAI21_X1 U21605 ( .B1(n18640), .B2(n18570), .A(n18383), .ZN(P3_U2683) );
  INV_X1 U21606 ( .A(n18384), .ZN(n18410) );
  OAI21_X1 U21607 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18410), .A(n18570), .ZN(
        n18395) );
  AOI22_X1 U21608 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18388) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n17066), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18387) );
  AOI22_X1 U21610 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18386) );
  AOI22_X1 U21611 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18385) );
  NAND4_X1 U21612 ( .A1(n18388), .A2(n18387), .A3(n18386), .A4(n18385), .ZN(
        n18394) );
  AOI22_X1 U21613 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18392) );
  AOI22_X1 U21614 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18391) );
  AOI22_X1 U21615 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9794), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18390) );
  AOI22_X1 U21616 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18389) );
  NAND4_X1 U21617 ( .A1(n18392), .A2(n18391), .A3(n18390), .A4(n18389), .ZN(
        n18393) );
  NOR2_X1 U21618 ( .A1(n18394), .A2(n18393), .ZN(n18645) );
  OAI22_X1 U21619 ( .A1(n18396), .A2(n18395), .B1(n18645), .B2(n18570), .ZN(
        P3_U2684) );
  NAND2_X1 U21620 ( .A1(n19584), .A2(n18424), .ZN(n18437) );
  NOR3_X1 U21621 ( .A1(n18398), .A2(n18397), .A3(n18437), .ZN(n18423) );
  AOI21_X1 U21622 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n18570), .A(n18423), .ZN(
        n18409) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n9793), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18402) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n17067), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18401) );
  AOI22_X1 U21625 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18400) );
  AOI22_X1 U21626 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18399) );
  NAND4_X1 U21627 ( .A1(n18402), .A2(n18401), .A3(n18400), .A4(n18399), .ZN(
        n18408) );
  AOI22_X1 U21628 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18406) );
  AOI22_X1 U21629 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18405) );
  AOI22_X1 U21630 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18404) );
  AOI22_X1 U21631 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18403) );
  NAND4_X1 U21632 ( .A1(n18406), .A2(n18405), .A3(n18404), .A4(n18403), .ZN(
        n18407) );
  NOR2_X1 U21633 ( .A1(n18408), .A2(n18407), .ZN(n18651) );
  OAI22_X1 U21634 ( .A1(n18410), .A2(n18409), .B1(n18651), .B2(n18570), .ZN(
        P3_U2685) );
  INV_X1 U21635 ( .A(n18437), .ZN(n18411) );
  AOI22_X1 U21636 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18570), .B1(
        P3_EBX_REG_16__SCAN_IN), .B2(n18411), .ZN(n18422) );
  AOI22_X1 U21637 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18415) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9795), .B1(
        n18473), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18414) );
  AOI22_X1 U21639 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18413) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18472), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18412) );
  NAND4_X1 U21641 ( .A1(n18415), .A2(n18414), .A3(n18413), .A4(n18412), .ZN(
        n18421) );
  AOI22_X1 U21642 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18419) );
  AOI22_X1 U21643 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18418) );
  AOI22_X1 U21644 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18417) );
  AOI22_X1 U21645 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18416) );
  NAND4_X1 U21646 ( .A1(n18419), .A2(n18418), .A3(n18417), .A4(n18416), .ZN(
        n18420) );
  NOR2_X1 U21647 ( .A1(n18421), .A2(n18420), .ZN(n18657) );
  OAI22_X1 U21648 ( .A1(n18423), .A2(n18422), .B1(n18657), .B2(n18570), .ZN(
        P3_U2686) );
  NOR2_X1 U21649 ( .A1(n18579), .A2(n18424), .ZN(n18449) );
  AOI22_X1 U21650 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18435) );
  AOI22_X1 U21651 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9794), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18434) );
  AOI22_X1 U21652 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18425) );
  OAI21_X1 U21653 ( .B1(n9850), .B2(n18426), .A(n18425), .ZN(n18432) );
  AOI22_X1 U21654 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18430) );
  AOI22_X1 U21655 ( .A1(n18520), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18429) );
  AOI22_X1 U21656 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18428) );
  AOI22_X1 U21657 ( .A1(n18473), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18427) );
  NAND4_X1 U21658 ( .A1(n18430), .A2(n18429), .A3(n18428), .A4(n18427), .ZN(
        n18431) );
  AOI211_X1 U21659 ( .C1(n18498), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n18432), .B(n18431), .ZN(n18433) );
  NAND3_X1 U21660 ( .A1(n18435), .A2(n18434), .A3(n18433), .ZN(n18658) );
  AOI22_X1 U21661 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18449), .B1(n18579), 
        .B2(n18658), .ZN(n18436) );
  OAI21_X1 U21662 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18437), .A(n18436), .ZN(
        P3_U2687) );
  AOI22_X1 U21663 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n18518), .ZN(n18441) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n9817), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n18455), .ZN(n18440) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n9794), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18439) );
  AOI22_X1 U21666 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18438) );
  NAND4_X1 U21667 ( .A1(n18441), .A2(n18440), .A3(n18439), .A4(n18438), .ZN(
        n18447) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18503), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n18539), .ZN(n18445) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17067), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17066), .ZN(n18444) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18472), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18443) );
  AOI22_X1 U21671 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18442) );
  NAND4_X1 U21672 ( .A1(n18445), .A2(n18444), .A3(n18443), .A4(n18442), .ZN(
        n18446) );
  NOR2_X1 U21673 ( .A1(n18447), .A2(n18446), .ZN(n18667) );
  INV_X1 U21674 ( .A(n18448), .ZN(n18450) );
  OAI21_X1 U21675 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n18450), .A(n18449), .ZN(
        n18451) );
  OAI21_X1 U21676 ( .B1(n18667), .B2(n18570), .A(n18451), .ZN(P3_U2688) );
  NAND2_X1 U21677 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18481), .ZN(n18467) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n9794), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18464) );
  AOI22_X1 U21679 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18463) );
  AOI22_X1 U21680 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18452) );
  OAI21_X1 U21681 ( .B1(n18454), .B2(n18453), .A(n18452), .ZN(n18461) );
  AOI22_X1 U21682 ( .A1(n13259), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18459) );
  AOI22_X1 U21683 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18458) );
  AOI22_X1 U21684 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18457) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18455), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18456) );
  NAND4_X1 U21686 ( .A1(n18459), .A2(n18458), .A3(n18457), .A4(n18456), .ZN(
        n18460) );
  AOI211_X1 U21687 ( .C1(n18498), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n18461), .B(n18460), .ZN(n18462) );
  NAND3_X1 U21688 ( .A1(n18464), .A2(n18463), .A3(n18462), .ZN(n18672) );
  AOI22_X1 U21689 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18465), .B1(n18579), 
        .B2(n18672), .ZN(n18466) );
  OAI21_X1 U21690 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n18467), .A(n18466), .ZN(
        P3_U2689) );
  AOI22_X1 U21691 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18471) );
  AOI22_X1 U21692 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18470) );
  AOI22_X1 U21693 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18469) );
  AOI22_X1 U21694 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18468) );
  NAND4_X1 U21695 ( .A1(n18471), .A2(n18470), .A3(n18469), .A4(n18468), .ZN(
        n18479) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18533), .B1(
        n18519), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18477) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13311), .B1(
        n18472), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18476) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n17067), .B1(
        n18473), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18475) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18520), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18474) );
  NAND4_X1 U21700 ( .A1(n18477), .A2(n18476), .A3(n18475), .A4(n18474), .ZN(
        n18478) );
  NOR2_X1 U21701 ( .A1(n18479), .A2(n18478), .ZN(n18681) );
  OAI21_X1 U21702 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n18482), .A(n18570), .ZN(
        n18480) );
  OAI22_X1 U21703 ( .A1(n18681), .A2(n18570), .B1(n18481), .B2(n18480), .ZN(
        P3_U2691) );
  AOI21_X1 U21704 ( .B1(n18484), .B2(n18483), .A(n18482), .ZN(n18497) );
  AOI22_X1 U21705 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18496) );
  AOI22_X1 U21706 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18495) );
  AOI22_X1 U21707 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18485) );
  OAI21_X1 U21708 ( .B1(n18487), .B2(n18486), .A(n18485), .ZN(n18493) );
  AOI22_X1 U21709 ( .A1(n17067), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18491) );
  AOI22_X1 U21710 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18490) );
  AOI22_X1 U21711 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18489) );
  AOI22_X1 U21712 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18488) );
  NAND4_X1 U21713 ( .A1(n18491), .A2(n18490), .A3(n18489), .A4(n18488), .ZN(
        n18492) );
  AOI211_X1 U21714 ( .C1(n18472), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n18493), .B(n18492), .ZN(n18494) );
  NAND3_X1 U21715 ( .A1(n18496), .A2(n18495), .A3(n18494), .ZN(n18684) );
  MUX2_X1 U21716 ( .A(n18497), .B(n18684), .S(n18579), .Z(P3_U2692) );
  AOI22_X1 U21717 ( .A1(n18473), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18502) );
  AOI22_X1 U21718 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18501) );
  AOI22_X1 U21719 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18500) );
  AOI22_X1 U21720 ( .A1(n18534), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18499) );
  NAND4_X1 U21721 ( .A1(n18502), .A2(n18501), .A3(n18500), .A4(n18499), .ZN(
        n18509) );
  AOI22_X1 U21722 ( .A1(n13311), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18507) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18503), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18506) );
  AOI22_X1 U21724 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9794), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18505) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18518), .B1(
        n18472), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18504) );
  NAND4_X1 U21726 ( .A1(n18507), .A2(n18506), .A3(n18505), .A4(n18504), .ZN(
        n18508) );
  NOR2_X1 U21727 ( .A1(n18509), .A2(n18508), .ZN(n18687) );
  NOR2_X1 U21728 ( .A1(n18579), .A2(n18511), .ZN(n18529) );
  OAI222_X1 U21729 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n19584), .B1(
        P3_EBX_REG_10__SCAN_IN), .B2(n18511), .C1(n18529), .C2(n18510), .ZN(
        n18512) );
  OAI21_X1 U21730 ( .B1(n18687), .B2(n18570), .A(n18512), .ZN(P3_U2693) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13311), .B1(
        n18533), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18517) );
  AOI22_X1 U21732 ( .A1(n18539), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18516) );
  AOI22_X1 U21733 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18515) );
  AOI22_X1 U21734 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18514) );
  NAND4_X1 U21735 ( .A1(n18517), .A2(n18516), .A3(n18515), .A4(n18514), .ZN(
        n18527) );
  AOI22_X1 U21736 ( .A1(n18503), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18518), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18525) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18519), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18524) );
  AOI22_X1 U21738 ( .A1(n9817), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18523) );
  AOI22_X1 U21739 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18520), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18522) );
  NAND4_X1 U21740 ( .A1(n18525), .A2(n18524), .A3(n18523), .A4(n18522), .ZN(
        n18526) );
  NOR2_X1 U21741 ( .A1(n18527), .A2(n18526), .ZN(n18691) );
  INV_X1 U21742 ( .A(n18528), .ZN(n18530) );
  OAI21_X1 U21743 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18530), .A(n18529), .ZN(
        n18531) );
  OAI21_X1 U21744 ( .B1(n18691), .B2(n18570), .A(n18531), .ZN(P3_U2694) );
  AOI22_X1 U21745 ( .A1(n18520), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18532), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18538) );
  AOI22_X1 U21746 ( .A1(n13258), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18537) );
  AOI22_X1 U21747 ( .A1(n18533), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9817), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18536) );
  AOI22_X1 U21748 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18534), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18535) );
  NAND4_X1 U21749 ( .A1(n18538), .A2(n18537), .A3(n18536), .A4(n18535), .ZN(
        n18545) );
  AOI22_X1 U21750 ( .A1(n18519), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13394), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18543) );
  AOI22_X1 U21751 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18542) );
  AOI22_X1 U21752 ( .A1(n9794), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13311), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18541) );
  AOI22_X1 U21753 ( .A1(n18472), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18513), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18540) );
  NAND4_X1 U21754 ( .A1(n18543), .A2(n18542), .A3(n18541), .A4(n18540), .ZN(
        n18544) );
  NOR2_X1 U21755 ( .A1(n18545), .A2(n18544), .ZN(n18697) );
  NOR2_X1 U21756 ( .A1(n18579), .A2(n18547), .ZN(n18551) );
  OAI222_X1 U21757 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n19584), .B1(
        P3_EBX_REG_8__SCAN_IN), .B2(n18547), .C1(n18551), .C2(n18546), .ZN(
        n18548) );
  OAI21_X1 U21758 ( .B1(n18697), .B2(n18570), .A(n18548), .ZN(P3_U2695) );
  INV_X1 U21759 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18553) );
  NOR3_X1 U21760 ( .A1(n18624), .A2(n18557), .A3(n18554), .ZN(n18550) );
  AOI22_X1 U21761 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n18551), .B1(n18550), .B2(
        n18549), .ZN(n18552) );
  OAI21_X1 U21762 ( .B1(n18553), .B2(n18570), .A(n18552), .ZN(P3_U2696) );
  NAND2_X1 U21763 ( .A1(n18570), .A2(n18554), .ZN(n18559) );
  NOR2_X1 U21764 ( .A1(n18624), .A2(n18554), .ZN(n18555) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18579), .B1(
        n18555), .B2(n18557), .ZN(n18556) );
  OAI21_X1 U21766 ( .B1(n18557), .B2(n18559), .A(n18556), .ZN(P3_U2697) );
  NOR2_X1 U21767 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n18565), .ZN(n18560) );
  INV_X1 U21768 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18558) );
  OAI22_X1 U21769 ( .A1(n18560), .A2(n18559), .B1(n18558), .B2(n18570), .ZN(
        P3_U2698) );
  AOI21_X1 U21770 ( .B1(n18561), .B2(n18566), .A(n18579), .ZN(n18562) );
  INV_X1 U21771 ( .A(n18562), .ZN(n18564) );
  INV_X1 U21772 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18563) );
  OAI22_X1 U21773 ( .A1(n18565), .A2(n18564), .B1(n18563), .B2(n18570), .ZN(
        P3_U2699) );
  INV_X1 U21774 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18568) );
  OAI21_X1 U21775 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18573), .A(n18566), .ZN(
        n18567) );
  AOI22_X1 U21776 ( .A1(n18579), .A2(n18568), .B1(n18567), .B2(n18570), .ZN(
        P3_U2700) );
  OAI21_X1 U21777 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n18569), .A(n18570), .ZN(
        n18572) );
  INV_X1 U21778 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18571) );
  OAI22_X1 U21779 ( .A1(n18573), .A2(n18572), .B1(n18571), .B2(n18570), .ZN(
        P3_U2701) );
  OAI221_X1 U21780 ( .B1(n19584), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .C1(
        n18624), .C2(n18574), .A(n18577), .ZN(n18575) );
  OAI21_X1 U21781 ( .B1(n18577), .B2(n18576), .A(n18575), .ZN(P3_U2702) );
  NAND2_X1 U21782 ( .A1(n19584), .A2(n18577), .ZN(n18581) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18579), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18578), .ZN(n18580) );
  OAI21_X1 U21784 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18581), .A(n18580), .ZN(
        P3_U2703) );
  INV_X1 U21785 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18738) );
  INV_X1 U21786 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18742) );
  INV_X1 U21787 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18762) );
  INV_X1 U21788 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18784) );
  INV_X1 U21789 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18787) );
  NAND4_X1 U21790 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n18582) );
  NOR3_X1 U21791 ( .A1(n18784), .A2(n18787), .A3(n18582), .ZN(n18670) );
  INV_X1 U21792 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18775) );
  NAND2_X1 U21793 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n18671) );
  NAND4_X1 U21794 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n18583)
         );
  NAND4_X1 U21795 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n18625)
         );
  NAND2_X1 U21796 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18601), .ZN(n18597) );
  INV_X1 U21797 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18734) );
  OR2_X1 U21798 ( .A1(n18591), .A2(n18734), .ZN(n18586) );
  NOR2_X2 U21799 ( .A1(n19579), .A2(n18726), .ZN(n18659) );
  AOI22_X1 U21800 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18659), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18584), .ZN(n18585) );
  OAI21_X1 U21801 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n18586), .A(n18585), .ZN(
        P3_U2704) );
  NOR2_X2 U21802 ( .A1(n19571), .A2(n18726), .ZN(n18652) );
  INV_X1 U21803 ( .A(n18659), .ZN(n18632) );
  OAI22_X1 U21804 ( .A1(n18588), .A2(n18717), .B1(n18587), .B2(n18632), .ZN(
        n18589) );
  AOI21_X1 U21805 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18652), .A(n18589), .ZN(
        n18590) );
  OAI221_X1 U21806 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18591), .C1(n18734), 
        .C2(n9916), .A(n18590), .ZN(P3_U2705) );
  AOI22_X1 U21807 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18659), .ZN(n18594) );
  OAI211_X1 U21808 ( .C1(n18592), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18726), .B(
        n18591), .ZN(n18593) );
  OAI211_X1 U21809 ( .C1(n18717), .C2(n18595), .A(n18594), .B(n18593), .ZN(
        P3_U2706) );
  AOI22_X1 U21810 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18652), .B1(n18596), .B2(
        n18722), .ZN(n18599) );
  OAI211_X1 U21811 ( .C1(n18601), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18726), .B(
        n18597), .ZN(n18598) );
  OAI211_X1 U21812 ( .C1(n18632), .C2(n18600), .A(n18599), .B(n18598), .ZN(
        P3_U2707) );
  AOI22_X1 U21813 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18659), .ZN(n18604) );
  AOI211_X1 U21814 ( .C1(n18738), .C2(n18606), .A(n18601), .B(n18646), .ZN(
        n18602) );
  INV_X1 U21815 ( .A(n18602), .ZN(n18603) );
  OAI211_X1 U21816 ( .C1(n18717), .C2(n18605), .A(n18604), .B(n18603), .ZN(
        P3_U2708) );
  AOI22_X1 U21817 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18659), .ZN(n18608) );
  OAI211_X1 U21818 ( .C1(n9898), .C2(P3_EAX_REG_26__SCAN_IN), .A(n18726), .B(
        n18606), .ZN(n18607) );
  OAI211_X1 U21819 ( .C1(n18717), .C2(n18609), .A(n18608), .B(n18607), .ZN(
        P3_U2709) );
  AOI22_X1 U21820 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18659), .ZN(n18612) );
  AOI211_X1 U21821 ( .C1(n18742), .C2(n18614), .A(n9898), .B(n18646), .ZN(
        n18610) );
  INV_X1 U21822 ( .A(n18610), .ZN(n18611) );
  OAI211_X1 U21823 ( .C1(n18717), .C2(n18613), .A(n18612), .B(n18611), .ZN(
        P3_U2710) );
  AOI22_X1 U21824 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18659), .ZN(n18617) );
  OAI211_X1 U21825 ( .C1(n18615), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18726), .B(
        n18614), .ZN(n18616) );
  OAI211_X1 U21826 ( .C1(n18717), .C2(n18618), .A(n18617), .B(n18616), .ZN(
        P3_U2711) );
  AOI22_X1 U21827 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18659), .ZN(n18622) );
  OAI211_X1 U21828 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18620), .A(n18726), .B(
        n18619), .ZN(n18621) );
  OAI211_X1 U21829 ( .C1(n18717), .C2(n18623), .A(n18622), .B(n18621), .ZN(
        P3_U2712) );
  INV_X1 U21830 ( .A(n18652), .ZN(n18663) );
  NOR2_X1 U21831 ( .A1(n18625), .A2(n18653), .ZN(n18630) );
  NAND2_X1 U21832 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n18626) );
  NAND2_X1 U21833 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18641), .ZN(n18637) );
  NAND2_X1 U21834 ( .A1(n18726), .A2(n18637), .ZN(n18636) );
  OAI21_X1 U21835 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18668), .A(n18636), .ZN(
        n18629) );
  OAI22_X1 U21836 ( .A1(n18627), .A2(n18717), .B1(n19578), .B2(n18632), .ZN(
        n18628) );
  AOI221_X1 U21837 ( .B1(n18630), .B2(n18746), .C1(n18629), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n18628), .ZN(n18631) );
  OAI21_X1 U21838 ( .B1(n19577), .B2(n18663), .A(n18631), .ZN(P3_U2713) );
  OAI22_X1 U21839 ( .A1(n18633), .A2(n18717), .B1(n20567), .B2(n18632), .ZN(
        n18634) );
  AOI21_X1 U21840 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n18652), .A(n18634), .ZN(
        n18635) );
  OAI221_X1 U21841 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18637), .C1(n18748), 
        .C2(n18636), .A(n18635), .ZN(P3_U2714) );
  AOI22_X1 U21842 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18659), .ZN(n18639) );
  OAI211_X1 U21843 ( .C1(n18641), .C2(P3_EAX_REG_20__SCAN_IN), .A(n18726), .B(
        n18637), .ZN(n18638) );
  OAI211_X1 U21844 ( .C1(n18640), .C2(n18717), .A(n18639), .B(n18638), .ZN(
        P3_U2715) );
  AOI22_X1 U21845 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18659), .ZN(n18644) );
  INV_X1 U21846 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18754) );
  NOR2_X1 U21847 ( .A1(n18754), .A2(n18653), .ZN(n18647) );
  INV_X1 U21848 ( .A(n18641), .ZN(n18642) );
  OAI211_X1 U21849 ( .C1(n18647), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18726), .B(
        n18642), .ZN(n18643) );
  OAI211_X1 U21850 ( .C1(n18645), .C2(n18717), .A(n18644), .B(n18643), .ZN(
        P3_U2716) );
  AOI22_X1 U21851 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18659), .ZN(n18650) );
  AOI211_X1 U21852 ( .C1(n18754), .C2(n18653), .A(n18647), .B(n18646), .ZN(
        n18648) );
  INV_X1 U21853 ( .A(n18648), .ZN(n18649) );
  OAI211_X1 U21854 ( .C1(n18651), .C2(n18717), .A(n18650), .B(n18649), .ZN(
        P3_U2717) );
  AOI22_X1 U21855 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18652), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18659), .ZN(n18656) );
  OAI211_X1 U21856 ( .C1(n18654), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18726), .B(
        n18653), .ZN(n18655) );
  OAI211_X1 U21857 ( .C1(n18657), .C2(n18717), .A(n18656), .B(n18655), .ZN(
        P3_U2718) );
  AOI22_X1 U21858 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n18659), .B1(n18722), .B2(
        n18658), .ZN(n18662) );
  OAI211_X1 U21859 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18664), .A(n18726), .B(
        n18660), .ZN(n18661) );
  OAI211_X1 U21860 ( .C1(n18663), .C2(n19547), .A(n18662), .B(n18661), .ZN(
        P3_U2719) );
  AOI21_X1 U21861 ( .B1(n18762), .B2(n18673), .A(n18664), .ZN(n18665) );
  AOI22_X1 U21862 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18723), .B1(n18665), .B2(
        n18726), .ZN(n18666) );
  OAI21_X1 U21863 ( .B1(n18667), .B2(n18717), .A(n18666), .ZN(P3_U2720) );
  NAND2_X1 U21864 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n18669) );
  NAND2_X1 U21865 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18693), .ZN(n18686) );
  NOR2_X1 U21866 ( .A1(n18671), .A2(n18686), .ZN(n18683) );
  NAND2_X1 U21867 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18683), .ZN(n18676) );
  AOI22_X1 U21868 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18723), .B1(n18722), .B2(
        n18672), .ZN(n18675) );
  NAND3_X1 U21869 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18726), .A3(n18673), 
        .ZN(n18674) );
  OAI211_X1 U21870 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n18676), .A(n18675), .B(
        n18674), .ZN(P3_U2721) );
  INV_X1 U21871 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n18838) );
  INV_X1 U21872 ( .A(n18676), .ZN(n18679) );
  AOI21_X1 U21873 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18726), .A(n18683), .ZN(
        n18678) );
  OAI222_X1 U21874 ( .A1(n18720), .A2(n18838), .B1(n18679), .B2(n18678), .C1(
        n18717), .C2(n18677), .ZN(P3_U2722) );
  INV_X1 U21875 ( .A(n18686), .ZN(n18680) );
  AOI22_X1 U21876 ( .A1(n18680), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n18726), .ZN(n18682) );
  OAI222_X1 U21877 ( .A1(n18720), .A2(n18836), .B1(n18683), .B2(n18682), .C1(
        n18717), .C2(n18681), .ZN(P3_U2723) );
  INV_X1 U21878 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18834) );
  NAND2_X1 U21879 ( .A1(n18726), .A2(n18686), .ZN(n18689) );
  AOI22_X1 U21880 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18723), .B1(n18722), .B2(
        n18684), .ZN(n18685) );
  OAI221_X1 U21881 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18686), .C1(n18834), 
        .C2(n18689), .A(n18685), .ZN(P3_U2724) );
  NOR2_X1 U21882 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18693), .ZN(n18688) );
  OAI222_X1 U21883 ( .A1(n18720), .A2(n18831), .B1(n18689), .B2(n18688), .C1(
        n18717), .C2(n18687), .ZN(P3_U2725) );
  AOI21_X1 U21884 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18726), .A(n18690), .ZN(
        n18692) );
  OAI222_X1 U21885 ( .A1(n18720), .A2(n13804), .B1(n18693), .B2(n18692), .C1(
        n18717), .C2(n18691), .ZN(P3_U2726) );
  AOI22_X1 U21886 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18723), .B1(n18701), .B2(
        n18775), .ZN(n18696) );
  NAND3_X1 U21887 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18726), .A3(n18694), .ZN(
        n18695) );
  OAI211_X1 U21888 ( .C1(n18697), .C2(n18717), .A(n18696), .B(n18695), .ZN(
        P3_U2727) );
  INV_X1 U21889 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18778) );
  INV_X1 U21890 ( .A(n18715), .ZN(n18725) );
  NOR3_X1 U21891 ( .A1(n18784), .A2(n18787), .A3(n18725), .ZN(n18714) );
  AND2_X1 U21892 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18714), .ZN(n18711) );
  NAND2_X1 U21893 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18711), .ZN(n18702) );
  NOR2_X1 U21894 ( .A1(n18778), .A2(n18702), .ZN(n18704) );
  OAI21_X1 U21895 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18704), .A(n18726), .ZN(
        n18700) );
  AOI22_X1 U21896 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18723), .B1(n18722), .B2(
        n18698), .ZN(n18699) );
  OAI21_X1 U21897 ( .B1(n18701), .B2(n18700), .A(n18699), .ZN(P3_U2728) );
  INV_X1 U21898 ( .A(n18702), .ZN(n18708) );
  AOI21_X1 U21899 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18726), .A(n18708), .ZN(
        n18705) );
  OAI222_X1 U21900 ( .A1(n18720), .A2(n19577), .B1(n18705), .B2(n18704), .C1(
        n18717), .C2(n18703), .ZN(P3_U2729) );
  AOI21_X1 U21901 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18726), .A(n18711), .ZN(
        n18707) );
  OAI222_X1 U21902 ( .A1(n19574), .A2(n18720), .B1(n18708), .B2(n18707), .C1(
        n18717), .C2(n18706), .ZN(P3_U2730) );
  AOI21_X1 U21903 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18726), .A(n18714), .ZN(
        n18710) );
  OAI222_X1 U21904 ( .A1(n19567), .A2(n18720), .B1(n18711), .B2(n18710), .C1(
        n18717), .C2(n18709), .ZN(P3_U2731) );
  AOI22_X1 U21905 ( .A1(n18715), .A2(P3_EAX_REG_2__SCAN_IN), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(n18726), .ZN(n18713) );
  OAI222_X1 U21906 ( .A1(n19563), .A2(n18720), .B1(n18714), .B2(n18713), .C1(
        n18717), .C2(n18712), .ZN(P3_U2732) );
  NOR2_X1 U21907 ( .A1(n18787), .A2(n18725), .ZN(n18719) );
  AOI21_X1 U21908 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18726), .A(n18715), .ZN(
        n18718) );
  OAI222_X1 U21909 ( .A1(n19560), .A2(n18720), .B1(n18719), .B2(n18718), .C1(
        n18717), .C2(n18716), .ZN(P3_U2733) );
  AOI22_X1 U21910 ( .A1(n18723), .A2(BUF2_REG_1__SCAN_IN), .B1(n18722), .B2(
        n18721), .ZN(n18729) );
  AND2_X1 U21911 ( .A1(n18724), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n18727) );
  OAI211_X1 U21912 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n18727), .A(n18726), .B(
        n18725), .ZN(n18728) );
  NAND2_X1 U21913 ( .A1(n18729), .A2(n18728), .ZN(P3_U2734) );
  OR2_X1 U21914 ( .A1(n20164), .A2(n19011), .ZN(n20199) );
  NOR2_X1 U21915 ( .A1(n18759), .A2(n18731), .ZN(P3_U2736) );
  NAND2_X1 U21916 ( .A1(n18772), .A2(n18732), .ZN(n18756) );
  INV_X2 U21917 ( .A(n20199), .ZN(n18790) );
  AOI22_X1 U21918 ( .A1(n18790), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18733) );
  OAI21_X1 U21919 ( .B1(n18734), .B2(n18756), .A(n18733), .ZN(P3_U2737) );
  AOI22_X1 U21920 ( .A1(n18790), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18735) );
  OAI21_X1 U21921 ( .B1(n10017), .B2(n18756), .A(n18735), .ZN(P3_U2738) );
  INV_X1 U21922 ( .A(n18756), .ZN(n18757) );
  AOI22_X1 U21923 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18757), .B1(n18790), 
        .B2(P3_UWORD_REG_12__SCAN_IN), .ZN(n18736) );
  OAI21_X1 U21924 ( .B1(n18737), .B2(n18759), .A(n18736), .ZN(P3_U2739) );
  INV_X1 U21925 ( .A(P3_UWORD_REG_11__SCAN_IN), .ZN(n18812) );
  OAI222_X1 U21926 ( .A1(n18812), .A2(n20199), .B1(n18759), .B2(n18739), .C1(
        n18738), .C2(n18756), .ZN(P3_U2740) );
  AOI22_X1 U21927 ( .A1(n18790), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18740) );
  OAI21_X1 U21928 ( .B1(n10020), .B2(n18756), .A(n18740), .ZN(P3_U2741) );
  AOI22_X1 U21929 ( .A1(n18790), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18741) );
  OAI21_X1 U21930 ( .B1(n18742), .B2(n18756), .A(n18741), .ZN(P3_U2742) );
  AOI22_X1 U21931 ( .A1(n18790), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18743) );
  OAI21_X1 U21932 ( .B1(n10019), .B2(n18756), .A(n18743), .ZN(P3_U2743) );
  INV_X1 U21933 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18806) );
  AOI22_X1 U21934 ( .A1(n18790), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18744) );
  OAI21_X1 U21935 ( .B1(n18806), .B2(n18756), .A(n18744), .ZN(P3_U2744) );
  AOI22_X1 U21936 ( .A1(n18790), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18745) );
  OAI21_X1 U21937 ( .B1(n18746), .B2(n18756), .A(n18745), .ZN(P3_U2745) );
  AOI22_X1 U21938 ( .A1(P3_UWORD_REG_5__SCAN_IN), .A2(n18790), .B1(n18789), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18747) );
  OAI21_X1 U21939 ( .B1(n18748), .B2(n18756), .A(n18747), .ZN(P3_U2746) );
  INV_X1 U21940 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18750) );
  AOI22_X1 U21941 ( .A1(n18790), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18749) );
  OAI21_X1 U21942 ( .B1(n18750), .B2(n18756), .A(n18749), .ZN(P3_U2747) );
  AOI22_X1 U21943 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18757), .B1(n18790), 
        .B2(P3_UWORD_REG_3__SCAN_IN), .ZN(n18751) );
  OAI21_X1 U21944 ( .B1(n18752), .B2(n18759), .A(n18751), .ZN(P3_U2748) );
  AOI22_X1 U21945 ( .A1(n18790), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18753) );
  OAI21_X1 U21946 ( .B1(n18754), .B2(n18756), .A(n18753), .ZN(P3_U2749) );
  AOI22_X1 U21947 ( .A1(n18790), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18755) );
  OAI21_X1 U21948 ( .B1(n18799), .B2(n18756), .A(n18755), .ZN(P3_U2750) );
  AOI22_X1 U21949 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18757), .B1(n18790), 
        .B2(P3_UWORD_REG_0__SCAN_IN), .ZN(n18758) );
  OAI21_X1 U21950 ( .B1(n18760), .B2(n18759), .A(n18758), .ZN(P3_U2751) );
  AOI22_X1 U21951 ( .A1(P3_LWORD_REG_15__SCAN_IN), .A2(n18790), .B1(n18789), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18761) );
  OAI21_X1 U21952 ( .B1(n18762), .B2(n18792), .A(n18761), .ZN(P3_U2752) );
  INV_X1 U21953 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18764) );
  AOI22_X1 U21954 ( .A1(n18790), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18763) );
  OAI21_X1 U21955 ( .B1(n18764), .B2(n18792), .A(n18763), .ZN(P3_U2753) );
  AOI22_X1 U21956 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18772), .B1(n18789), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18765) );
  OAI21_X1 U21957 ( .B1(n18766), .B2(n20199), .A(n18765), .ZN(P3_U2754) );
  INV_X1 U21958 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18768) );
  AOI22_X1 U21959 ( .A1(n18790), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18767) );
  OAI21_X1 U21960 ( .B1(n18768), .B2(n18792), .A(n18767), .ZN(P3_U2755) );
  AOI22_X1 U21961 ( .A1(n18790), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18769) );
  OAI21_X1 U21962 ( .B1(n18834), .B2(n18792), .A(n18769), .ZN(P3_U2756) );
  INV_X1 U21963 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18771) );
  AOI22_X1 U21964 ( .A1(n18790), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18785), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18770) );
  OAI21_X1 U21965 ( .B1(n18771), .B2(n18792), .A(n18770), .ZN(P3_U2757) );
  AOI222_X1 U21966 ( .A1(P3_LWORD_REG_9__SCAN_IN), .A2(n18790), .B1(n18789), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .C1(P3_EAX_REG_9__SCAN_IN), .C2(n18772), 
        .ZN(n18773) );
  INV_X1 U21967 ( .A(n18773), .ZN(P3_U2758) );
  AOI22_X1 U21968 ( .A1(n18790), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18785), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18774) );
  OAI21_X1 U21969 ( .B1(n18775), .B2(n18792), .A(n18774), .ZN(P3_U2759) );
  INV_X1 U21970 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18826) );
  AOI22_X1 U21971 ( .A1(n18790), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18785), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18776) );
  OAI21_X1 U21972 ( .B1(n18826), .B2(n18792), .A(n18776), .ZN(P3_U2760) );
  AOI22_X1 U21973 ( .A1(n18790), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18785), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18777) );
  OAI21_X1 U21974 ( .B1(n18778), .B2(n18792), .A(n18777), .ZN(P3_U2761) );
  INV_X1 U21975 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18780) );
  AOI22_X1 U21976 ( .A1(n18790), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18785), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18779) );
  OAI21_X1 U21977 ( .B1(n18780), .B2(n18792), .A(n18779), .ZN(P3_U2762) );
  INV_X1 U21978 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18782) );
  AOI22_X1 U21979 ( .A1(n18790), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18785), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18781) );
  OAI21_X1 U21980 ( .B1(n18782), .B2(n18792), .A(n18781), .ZN(P3_U2763) );
  AOI22_X1 U21981 ( .A1(n18790), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18785), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18783) );
  OAI21_X1 U21982 ( .B1(n18784), .B2(n18792), .A(n18783), .ZN(P3_U2764) );
  AOI22_X1 U21983 ( .A1(n18790), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18785), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18786) );
  OAI21_X1 U21984 ( .B1(n18787), .B2(n18792), .A(n18786), .ZN(P3_U2765) );
  INV_X1 U21985 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18819) );
  AOI22_X1 U21986 ( .A1(n18790), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18788) );
  OAI21_X1 U21987 ( .B1(n18819), .B2(n18792), .A(n18788), .ZN(P3_U2766) );
  AOI22_X1 U21988 ( .A1(n18790), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18789), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18791) );
  OAI21_X1 U21989 ( .B1(n18793), .B2(n18792), .A(n18791), .ZN(P3_U2767) );
  AOI211_X1 U21990 ( .C1(n10001), .C2(n19555), .A(n18794), .B(n18796), .ZN(
        n18813) );
  NAND2_X1 U21991 ( .A1(n18813), .A2(n19555), .ZN(n18808) );
  INV_X1 U21992 ( .A(n18795), .ZN(n20039) );
  INV_X2 U21993 ( .A(n18813), .ZN(n18839) );
  AOI22_X1 U21994 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18839), .ZN(n18797) );
  OAI21_X1 U21995 ( .B1(n19547), .B2(n18808), .A(n18797), .ZN(P3_U2768) );
  INV_X1 U21996 ( .A(n18808), .ZN(n18844) );
  AOI22_X1 U21997 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18844), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18839), .ZN(n18798) );
  OAI21_X1 U21998 ( .B1(n18799), .B2(n18833), .A(n18798), .ZN(P3_U2769) );
  INV_X2 U21999 ( .A(n18833), .ZN(n18840) );
  AOI22_X1 U22000 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18839), .ZN(n18800) );
  OAI21_X1 U22001 ( .B1(n19560), .B2(n18808), .A(n18800), .ZN(P3_U2770) );
  AOI22_X1 U22002 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18839), .ZN(n18801) );
  OAI21_X1 U22003 ( .B1(n19563), .B2(n18808), .A(n18801), .ZN(P3_U2771) );
  AOI22_X1 U22004 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18839), .ZN(n18802) );
  OAI21_X1 U22005 ( .B1(n19567), .B2(n18808), .A(n18802), .ZN(P3_U2772) );
  AOI22_X1 U22006 ( .A1(P3_UWORD_REG_5__SCAN_IN), .A2(n18839), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n18840), .ZN(n18803) );
  OAI21_X1 U22007 ( .B1(n19574), .B2(n18808), .A(n18803), .ZN(P3_U2773) );
  AOI22_X1 U22008 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18839), .ZN(n18804) );
  OAI21_X1 U22009 ( .B1(n19577), .B2(n18808), .A(n18804), .ZN(P3_U2774) );
  AOI22_X1 U22010 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18844), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18839), .ZN(n18805) );
  OAI21_X1 U22011 ( .B1(n18806), .B2(n18833), .A(n18805), .ZN(P3_U2775) );
  AOI22_X1 U22012 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18839), .ZN(n18807) );
  OAI21_X1 U22013 ( .B1(n18828), .B2(n18808), .A(n18807), .ZN(P3_U2776) );
  AOI22_X1 U22014 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18839), .ZN(n18809) );
  OAI21_X1 U22015 ( .B1(n13804), .B2(n18842), .A(n18809), .ZN(P3_U2777) );
  AOI22_X1 U22016 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18839), .ZN(n18810) );
  OAI21_X1 U22017 ( .B1(n18831), .B2(n18842), .A(n18810), .ZN(P3_U2778) );
  AOI22_X1 U22018 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18844), .B1(
        P3_EAX_REG_27__SCAN_IN), .B2(n18840), .ZN(n18811) );
  OAI21_X1 U22019 ( .B1(n18813), .B2(n18812), .A(n18811), .ZN(P3_U2779) );
  AOI22_X1 U22020 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18839), .ZN(n18814) );
  OAI21_X1 U22021 ( .B1(n18836), .B2(n18842), .A(n18814), .ZN(P3_U2780) );
  AOI22_X1 U22022 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18839), .ZN(n18815) );
  OAI21_X1 U22023 ( .B1(n18838), .B2(n18842), .A(n18815), .ZN(P3_U2781) );
  AOI22_X1 U22024 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18840), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18839), .ZN(n18816) );
  OAI21_X1 U22025 ( .B1(n18843), .B2(n18842), .A(n18816), .ZN(P3_U2782) );
  AOI22_X1 U22026 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18839), .ZN(n18817) );
  OAI21_X1 U22027 ( .B1(n19547), .B2(n18842), .A(n18817), .ZN(P3_U2783) );
  AOI22_X1 U22028 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18844), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18839), .ZN(n18818) );
  OAI21_X1 U22029 ( .B1(n18819), .B2(n18833), .A(n18818), .ZN(P3_U2784) );
  AOI22_X1 U22030 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18839), .ZN(n18820) );
  OAI21_X1 U22031 ( .B1(n19560), .B2(n18842), .A(n18820), .ZN(P3_U2785) );
  AOI22_X1 U22032 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18839), .ZN(n18821) );
  OAI21_X1 U22033 ( .B1(n19563), .B2(n18842), .A(n18821), .ZN(P3_U2786) );
  AOI22_X1 U22034 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18839), .ZN(n18822) );
  OAI21_X1 U22035 ( .B1(n19567), .B2(n18842), .A(n18822), .ZN(P3_U2787) );
  AOI22_X1 U22036 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18839), .ZN(n18823) );
  OAI21_X1 U22037 ( .B1(n19574), .B2(n18842), .A(n18823), .ZN(P3_U2788) );
  AOI22_X1 U22038 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18839), .ZN(n18824) );
  OAI21_X1 U22039 ( .B1(n19577), .B2(n18842), .A(n18824), .ZN(P3_U2789) );
  AOI22_X1 U22040 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18844), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18839), .ZN(n18825) );
  OAI21_X1 U22041 ( .B1(n18826), .B2(n18833), .A(n18825), .ZN(P3_U2790) );
  AOI22_X1 U22042 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18839), .ZN(n18827) );
  OAI21_X1 U22043 ( .B1(n18828), .B2(n18842), .A(n18827), .ZN(P3_U2791) );
  AOI22_X1 U22044 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18839), .ZN(n18829) );
  OAI21_X1 U22045 ( .B1(n13804), .B2(n18842), .A(n18829), .ZN(P3_U2792) );
  AOI22_X1 U22046 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18839), .ZN(n18830) );
  OAI21_X1 U22047 ( .B1(n18831), .B2(n18842), .A(n18830), .ZN(P3_U2793) );
  AOI22_X1 U22048 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18844), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18839), .ZN(n18832) );
  OAI21_X1 U22049 ( .B1(n18834), .B2(n18833), .A(n18832), .ZN(P3_U2794) );
  AOI22_X1 U22050 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18839), .ZN(n18835) );
  OAI21_X1 U22051 ( .B1(n18836), .B2(n18842), .A(n18835), .ZN(P3_U2795) );
  AOI22_X1 U22052 ( .A1(P3_LWORD_REG_13__SCAN_IN), .A2(n18839), .B1(
        P3_EAX_REG_13__SCAN_IN), .B2(n18840), .ZN(n18837) );
  OAI21_X1 U22053 ( .B1(n18838), .B2(n18842), .A(n18837), .ZN(P3_U2796) );
  AOI22_X1 U22054 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18840), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18839), .ZN(n18841) );
  OAI21_X1 U22055 ( .B1(n18843), .B2(n18842), .A(n18841), .ZN(P3_U2797) );
  AOI222_X1 U22056 ( .A1(n18844), .A2(BUF2_REG_15__SCAN_IN), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18839), .C1(P3_EAX_REG_15__SCAN_IN), 
        .C2(n18840), .ZN(n18845) );
  INV_X1 U22057 ( .A(n18845), .ZN(P3_U2798) );
  OAI21_X1 U22058 ( .B1(n18846), .B2(n19121), .A(n19212), .ZN(n18847) );
  AOI21_X1 U22059 ( .B1(n19048), .B2(n18848), .A(n18847), .ZN(n18876) );
  OAI21_X1 U22060 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18964), .A(
        n18876), .ZN(n18862) );
  NAND2_X1 U22061 ( .A1(n9790), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n18854) );
  NAND3_X1 U22062 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18851) );
  NAND2_X1 U22063 ( .A1(n18887), .A2(n19052), .ZN(n18903) );
  NOR2_X1 U22064 ( .A1(n18851), .A2(n18903), .ZN(n18867) );
  OAI211_X1 U22065 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n18867), .B(n18852), .ZN(n18853) );
  OAI211_X1 U22066 ( .C1(n19067), .C2(n18855), .A(n18854), .B(n18853), .ZN(
        n18856) );
  NAND2_X1 U22067 ( .A1(n19126), .A2(n19218), .ZN(n18960) );
  AOI22_X1 U22068 ( .A1(n19062), .A2(n19226), .B1(n19061), .B2(n18857), .ZN(
        n18883) );
  NAND2_X1 U22069 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18883), .ZN(
        n18868) );
  NAND3_X1 U22070 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18960), .A3(
        n18868), .ZN(n18858) );
  OAI211_X1 U22071 ( .C1(n18925), .C2(n18860), .A(n18859), .B(n18858), .ZN(
        P3_U2802) );
  AOI22_X1 U22072 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18862), .B1(
        n19071), .B2(n18861), .ZN(n18872) );
  NAND2_X1 U22073 ( .A1(n18864), .A2(n18863), .ZN(n18865) );
  XNOR2_X1 U22074 ( .A(n19119), .B(n18865), .ZN(n19229) );
  AOI22_X1 U22075 ( .A1(n19128), .A2(n19229), .B1(n18867), .B2(n18866), .ZN(
        n18871) );
  NOR2_X1 U22076 ( .A1(n19219), .A2(n18925), .ZN(n18869) );
  OAI21_X1 U22077 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18869), .A(
        n18868), .ZN(n18870) );
  NAND2_X1 U22078 ( .A1(n9790), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n19230) );
  NAND4_X1 U22079 ( .A1(n18872), .A2(n18871), .A3(n18870), .A4(n19230), .ZN(
        P3_U2803) );
  NOR2_X1 U22080 ( .A1(n18873), .A2(n19652), .ZN(n18918) );
  AOI21_X1 U22081 ( .B1(n18874), .B2(n18918), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18875) );
  OAI22_X1 U22082 ( .A1(n18876), .A2(n18875), .B1(n19529), .B2(n20124), .ZN(
        n18880) );
  AOI21_X1 U22083 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18878), .A(
        n18877), .ZN(n19233) );
  NAND3_X1 U22084 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19244), .A3(
        n10202), .ZN(n19239) );
  OAI22_X1 U22085 ( .A1(n19233), .A2(n19101), .B1(n18925), .B2(n19239), .ZN(
        n18879) );
  AOI211_X1 U22086 ( .C1(n18881), .C2(n19174), .A(n18880), .B(n18879), .ZN(
        n18882) );
  OAI21_X1 U22087 ( .B1(n18883), .B2(n10202), .A(n18882), .ZN(P3_U2804) );
  NAND2_X1 U22088 ( .A1(n19347), .A2(n18900), .ZN(n19256) );
  NOR2_X1 U22089 ( .A1(n19256), .A2(n18912), .ZN(n18884) );
  XNOR2_X1 U22090 ( .A(n18884), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n19254) );
  INV_X1 U22091 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20122) );
  NOR2_X1 U22092 ( .A1(n19529), .A2(n20122), .ZN(n19248) );
  INV_X1 U22093 ( .A(n18964), .ZN(n18934) );
  AOI21_X1 U22094 ( .B1(n19048), .B2(n18885), .A(n19163), .ZN(n18886) );
  OAI21_X1 U22095 ( .B1(n18887), .B2(n19652), .A(n18886), .ZN(n18917) );
  AOI21_X1 U22096 ( .B1(n18934), .B2(n18888), .A(n18917), .ZN(n18901) );
  OAI21_X1 U22097 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18889), .ZN(n18890) );
  OAI22_X1 U22098 ( .A1(n18901), .A2(n18891), .B1(n18903), .B2(n18890), .ZN(
        n18892) );
  AOI211_X1 U22099 ( .C1(n18893), .C2(n19071), .A(n19248), .B(n18892), .ZN(
        n18899) );
  NAND3_X1 U22100 ( .A1(n19350), .A2(n18900), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18894) );
  XNOR2_X1 U22101 ( .A(n18894), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n19250) );
  AOI21_X1 U22102 ( .B1(n9797), .B2(n19119), .A(n18895), .ZN(n18897) );
  XNOR2_X1 U22103 ( .A(n18897), .B(n19240), .ZN(n19249) );
  AOI22_X1 U22104 ( .A1(n19062), .A2(n19250), .B1(n19128), .B2(n19249), .ZN(
        n18898) );
  OAI211_X1 U22105 ( .C1(n19218), .C2(n19254), .A(n18899), .B(n18898), .ZN(
        P3_U2805) );
  NAND2_X1 U22106 ( .A1(n19350), .A2(n18900), .ZN(n19255) );
  AOI22_X1 U22107 ( .A1(n19062), .A2(n19255), .B1(n19061), .B2(n19256), .ZN(
        n18923) );
  NAND2_X1 U22108 ( .A1(n9790), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n19266) );
  OAI221_X1 U22109 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18903), .C1(
        n18902), .C2(n18901), .A(n19266), .ZN(n18904) );
  AOI21_X1 U22110 ( .B1(n19071), .B2(n18905), .A(n18904), .ZN(n18911) );
  AOI21_X1 U22111 ( .B1(n18907), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n18906), .ZN(n18908) );
  INV_X1 U22112 ( .A(n18908), .ZN(n19265) );
  INV_X1 U22113 ( .A(n18925), .ZN(n18909) );
  NOR2_X1 U22114 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18924), .ZN(
        n19263) );
  AOI22_X1 U22115 ( .A1(n19128), .A2(n19265), .B1(n18909), .B2(n19263), .ZN(
        n18910) );
  OAI211_X1 U22116 ( .C1(n18923), .C2(n18912), .A(n18911), .B(n18910), .ZN(
        P3_U2806) );
  AOI22_X1 U22117 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19119), .B1(
        n18913), .B2(n18928), .ZN(n18914) );
  NAND2_X1 U22118 ( .A1(n18957), .A2(n18914), .ZN(n18915) );
  XNOR2_X1 U22119 ( .A(n18915), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n19270) );
  OAI21_X1 U22120 ( .B1(n19071), .B2(n18934), .A(n18916), .ZN(n18920) );
  OAI21_X1 U22121 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18918), .A(
        n18917), .ZN(n18919) );
  OAI211_X1 U22122 ( .C1(n20118), .C2(n19529), .A(n18920), .B(n18919), .ZN(
        n18921) );
  AOI21_X1 U22123 ( .B1(n19128), .B2(n19270), .A(n18921), .ZN(n18922) );
  OAI221_X1 U22124 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18925), 
        .C1(n18924), .C2(n18923), .A(n18922), .ZN(P3_U2807) );
  NAND2_X1 U22125 ( .A1(n18926), .A2(n19018), .ZN(n18943) );
  INV_X1 U22126 ( .A(n18926), .ZN(n19278) );
  OAI22_X1 U22127 ( .A1(n19350), .A2(n19126), .B1(n19347), .B2(n19218), .ZN(
        n19019) );
  AOI21_X1 U22128 ( .B1(n19278), .B2(n18960), .A(n19019), .ZN(n18956) );
  INV_X1 U22129 ( .A(n18957), .ZN(n18927) );
  AOI221_X1 U22130 ( .B1(n18929), .B2(n18928), .C1(n18947), .C2(n18928), .A(
        n18927), .ZN(n18930) );
  XNOR2_X1 U22131 ( .A(n18930), .B(n19289), .ZN(n19285) );
  AOI21_X1 U22132 ( .B1(n19048), .B2(n18931), .A(n19163), .ZN(n18932) );
  OAI21_X1 U22133 ( .B1(n18935), .B2(n19121), .A(n18932), .ZN(n18963) );
  AOI21_X1 U22134 ( .B1(n18934), .B2(n18933), .A(n18963), .ZN(n18944) );
  NAND2_X1 U22135 ( .A1(n18935), .A2(n19052), .ZN(n18946) );
  AOI21_X1 U22136 ( .B1(n18945), .B2(n18940), .A(n18946), .ZN(n18937) );
  AOI22_X1 U22137 ( .A1(n18938), .A2(n19071), .B1(n18937), .B2(n18936), .ZN(
        n18939) );
  NAND2_X1 U22138 ( .A1(n9790), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n19287) );
  OAI211_X1 U22139 ( .C1(n18944), .C2(n18940), .A(n18939), .B(n19287), .ZN(
        n18941) );
  AOI21_X1 U22140 ( .B1(n19128), .B2(n19285), .A(n18941), .ZN(n18942) );
  OAI221_X1 U22141 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18943), 
        .C1(n19289), .C2(n18956), .A(n18942), .ZN(P3_U2808) );
  NAND2_X1 U22142 ( .A1(n9790), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n19300) );
  OAI221_X1 U22143 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18946), .C1(
        n18945), .C2(n18944), .A(n19300), .ZN(n18953) );
  INV_X1 U22144 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19274) );
  NOR3_X1 U22145 ( .A1(n19119), .A2(n19274), .A3(n18947), .ZN(n18970) );
  AOI22_X1 U22146 ( .A1(n19280), .A2(n18970), .B1(n18992), .B2(n18949), .ZN(
        n18950) );
  XOR2_X1 U22147 ( .A(n18950), .B(n19296), .Z(n19299) );
  INV_X1 U22148 ( .A(n19299), .ZN(n18951) );
  NAND2_X1 U22149 ( .A1(n19280), .A2(n19296), .ZN(n19302) );
  NOR2_X1 U22150 ( .A1(n19318), .A2(n19274), .ZN(n19292) );
  NAND2_X1 U22151 ( .A1(n19018), .A2(n19292), .ZN(n18984) );
  OAI22_X1 U22152 ( .A1(n18951), .A2(n19101), .B1(n19302), .B2(n18984), .ZN(
        n18952) );
  AOI211_X1 U22153 ( .C1(n19071), .C2(n18954), .A(n18953), .B(n18952), .ZN(
        n18955) );
  OAI21_X1 U22154 ( .B1(n18956), .B2(n19296), .A(n18955), .ZN(P3_U2809) );
  OAI221_X1 U22155 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18991), 
        .C1(n18983), .C2(n18970), .A(n18957), .ZN(n18958) );
  XNOR2_X1 U22156 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18958), .ZN(
        n19303) );
  NAND3_X1 U22157 ( .A1(n18959), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n19306) );
  AOI21_X1 U22158 ( .B1(n18960), .B2(n19306), .A(n19019), .ZN(n18982) );
  NAND2_X1 U22159 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18961), .ZN(
        n19311) );
  OAI22_X1 U22160 ( .A1(n18982), .A2(n18961), .B1(n19311), .B2(n18984), .ZN(
        n18962) );
  AOI21_X1 U22161 ( .B1(n19128), .B2(n19303), .A(n18962), .ZN(n18969) );
  NAND2_X1 U22162 ( .A1(n9790), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18968) );
  OAI221_X1 U22163 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10350), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19922), .A(n18963), .ZN(
        n18967) );
  OAI21_X1 U22164 ( .B1(n19071), .B2(n18934), .A(n18965), .ZN(n18966) );
  NAND4_X1 U22165 ( .A1(n18969), .A2(n18968), .A3(n18967), .A4(n18966), .ZN(
        P3_U2810) );
  AOI21_X1 U22166 ( .B1(n18991), .B2(n18992), .A(n18970), .ZN(n18971) );
  XNOR2_X1 U22167 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n18971), .ZN(
        n19312) );
  NAND2_X1 U22168 ( .A1(n18974), .A2(n19052), .ZN(n18987) );
  AOI221_X1 U22169 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n18973), .C2(n18972), .A(
        n18987), .ZN(n18980) );
  INV_X1 U22170 ( .A(n18974), .ZN(n18975) );
  AOI21_X1 U22171 ( .B1(n19165), .B2(n18975), .A(n19163), .ZN(n18999) );
  OAI21_X1 U22172 ( .B1(n18976), .B2(n19011), .A(n18999), .ZN(n18990) );
  AOI22_X1 U22173 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18990), .B1(
        n19071), .B2(n18977), .ZN(n18978) );
  OAI21_X1 U22174 ( .B1(n19529), .B2(n20110), .A(n18978), .ZN(n18979) );
  AOI211_X1 U22175 ( .C1(n19128), .C2(n19312), .A(n18980), .B(n18979), .ZN(
        n18981) );
  OAI221_X1 U22176 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18984), 
        .C1(n18983), .C2(n18982), .A(n18981), .ZN(P3_U2811) );
  AOI21_X1 U22177 ( .B1(n19018), .B2(n19318), .A(n19019), .ZN(n19006) );
  NOR2_X1 U22178 ( .A1(n19529), .A2(n20108), .ZN(n18989) );
  INV_X1 U22179 ( .A(n18985), .ZN(n18986) );
  OAI22_X1 U22180 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18987), .B1(
        n18986), .B2(n19067), .ZN(n18988) );
  AOI211_X1 U22181 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18990), .A(
        n18989), .B(n18988), .ZN(n18995) );
  AOI21_X1 U22182 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n19008), .A(
        n18991), .ZN(n18993) );
  XOR2_X1 U22183 ( .A(n18993), .B(n18992), .Z(n19328) );
  NOR2_X1 U22184 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n19318), .ZN(
        n19327) );
  AOI22_X1 U22185 ( .A1(n19128), .A2(n19328), .B1(n19018), .B2(n19327), .ZN(
        n18994) );
  OAI211_X1 U22186 ( .C1(n19006), .C2(n19274), .A(n18995), .B(n18994), .ZN(
        P3_U2812) );
  AOI21_X1 U22187 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19018), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19005) );
  AOI22_X1 U22188 ( .A1(n9790), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18996), 
        .B2(n19174), .ZN(n19004) );
  OAI21_X1 U22189 ( .B1(n18998), .B2(n19333), .A(n18997), .ZN(n19331) );
  AOI221_X1 U22190 ( .B1(n19001), .B2(n19000), .C1(n19652), .C2(n19000), .A(
        n18999), .ZN(n19002) );
  AOI21_X1 U22191 ( .B1(n19128), .B2(n19331), .A(n19002), .ZN(n19003) );
  OAI211_X1 U22192 ( .C1(n19006), .C2(n19005), .A(n19004), .B(n19003), .ZN(
        P3_U2813) );
  NAND2_X1 U22193 ( .A1(n19008), .A2(n19116), .ZN(n19080) );
  OAI22_X1 U22194 ( .A1(n19008), .A2(n19007), .B1(n19080), .B2(n19326), .ZN(
        n19009) );
  XNOR2_X1 U22195 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n19009), .ZN(
        n19346) );
  INV_X1 U22196 ( .A(n19052), .ZN(n19010) );
  NOR3_X1 U22197 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19010), .A3(
        n13599), .ZN(n19024) );
  AOI21_X1 U22198 ( .B1(n19165), .B2(n13599), .A(n19163), .ZN(n19047) );
  OAI21_X1 U22199 ( .B1(n19012), .B2(n19011), .A(n19047), .ZN(n19025) );
  NAND2_X1 U22200 ( .A1(n9790), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n19344) );
  INV_X1 U22201 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n19013) );
  NAND3_X1 U22202 ( .A1(n19014), .A2(n19013), .A3(n19052), .ZN(n19015) );
  OAI211_X1 U22203 ( .C1(n19067), .C2(n19016), .A(n19344), .B(n19015), .ZN(
        n19017) );
  AOI221_X1 U22204 ( .B1(n19024), .B2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(
        n19025), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n19017), .ZN(
        n19021) );
  AOI22_X1 U22205 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19019), .B1(
        n19018), .B2(n19341), .ZN(n19020) );
  OAI211_X1 U22206 ( .C1(n19346), .C2(n19101), .A(n19021), .B(n19020), .ZN(
        P3_U2814) );
  AND2_X1 U22207 ( .A1(n19352), .A2(n19351), .ZN(n19033) );
  OR2_X1 U22208 ( .A1(n19126), .A2(n19350), .ZN(n19032) );
  NAND2_X1 U22209 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n9790), .ZN(n19358) );
  OAI21_X1 U22210 ( .B1(n19067), .B2(n19022), .A(n19358), .ZN(n19023) );
  AOI211_X1 U22211 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19025), .A(
        n19024), .B(n19023), .ZN(n19031) );
  NAND2_X1 U22212 ( .A1(n19026), .A2(n19119), .ZN(n19068) );
  NOR2_X1 U22213 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19068), .ZN(
        n19040) );
  NOR3_X1 U22214 ( .A1(n19392), .A2(n19078), .A3(n19080), .ZN(n19041) );
  NAND2_X1 U22215 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19385), .ZN(
        n19060) );
  OAI221_X1 U22216 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n19040), 
        .C1(n19369), .C2(n19041), .A(n19060), .ZN(n19027) );
  XNOR2_X1 U22217 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n19027), .ZN(
        n19357) );
  NOR2_X1 U22218 ( .A1(n19347), .A2(n19218), .ZN(n19029) );
  NAND2_X1 U22219 ( .A1(n19351), .A2(n19028), .ZN(n19355) );
  AOI22_X1 U22220 ( .A1(n19128), .A2(n19357), .B1(n19029), .B2(n19355), .ZN(
        n19030) );
  OAI211_X1 U22221 ( .C1(n19033), .C2(n19032), .A(n19031), .B(n19030), .ZN(
        P3_U2815) );
  NOR3_X1 U22222 ( .A1(n19034), .A2(n19035), .A3(n19652), .ZN(n19085) );
  AOI21_X1 U22223 ( .B1(n19053), .B2(n19085), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n19046) );
  AOI22_X1 U22224 ( .A1(n9790), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n19036), 
        .B2(n19174), .ZN(n19045) );
  AOI21_X1 U22225 ( .B1(n19369), .B2(n19038), .A(n19037), .ZN(n19373) );
  OAI21_X1 U22226 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n19039), .A(
        n19352), .ZN(n19371) );
  OAI21_X1 U22227 ( .B1(n19041), .B2(n19040), .A(n19060), .ZN(n19042) );
  XNOR2_X1 U22228 ( .A(n19042), .B(n19369), .ZN(n19370) );
  OAI22_X1 U22229 ( .A1(n19126), .A2(n19371), .B1(n19101), .B2(n19370), .ZN(
        n19043) );
  AOI21_X1 U22230 ( .B1(n19061), .B2(n19373), .A(n19043), .ZN(n19044) );
  OAI211_X1 U22231 ( .C1(n19047), .C2(n19046), .A(n19045), .B(n19044), .ZN(
        P3_U2816) );
  AOI21_X1 U22232 ( .B1(n19165), .B2(n19049), .A(n19048), .ZN(n19050) );
  OAI21_X1 U22233 ( .B1(n19051), .B2(n19050), .A(n19212), .ZN(n19072) );
  NAND2_X1 U22234 ( .A1(n18087), .A2(n19052), .ZN(n19074) );
  AOI211_X1 U22235 ( .C1(n19055), .C2(n19054), .A(n19053), .B(n19074), .ZN(
        n19056) );
  NOR2_X1 U22236 ( .A1(n19529), .A2(n20098), .ZN(n19387) );
  AOI211_X1 U22237 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n19072), .A(
        n19056), .B(n19387), .ZN(n19065) );
  AOI22_X1 U22238 ( .A1(n19116), .A2(n19361), .B1(n19119), .B2(n19078), .ZN(
        n19058) );
  NOR2_X1 U22239 ( .A1(n19058), .A2(n19057), .ZN(n19059) );
  XNOR2_X1 U22240 ( .A(n19059), .B(n19385), .ZN(n19389) );
  OR2_X1 U22241 ( .A1(n19392), .A2(n19060), .ZN(n19391) );
  NAND2_X1 U22242 ( .A1(n19407), .A2(n19361), .ZN(n19380) );
  NAND2_X1 U22243 ( .A1(n19361), .A2(n19405), .ZN(n19382) );
  AOI22_X1 U22244 ( .A1(n19062), .A2(n19380), .B1(n19061), .B2(n19382), .ZN(
        n19079) );
  OAI22_X1 U22245 ( .A1(n19113), .A2(n19391), .B1(n19079), .B2(n19385), .ZN(
        n19063) );
  AOI21_X1 U22246 ( .B1(n19128), .B2(n19389), .A(n19063), .ZN(n19064) );
  OAI211_X1 U22247 ( .C1(n19067), .C2(n19066), .A(n19065), .B(n19064), .ZN(
        P3_U2817) );
  OAI21_X1 U22248 ( .B1(n19080), .B2(n19392), .A(n19068), .ZN(n19069) );
  XNOR2_X1 U22249 ( .A(n19069), .B(n19078), .ZN(n19397) );
  NOR3_X1 U22250 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19113), .A3(
        n19392), .ZN(n19076) );
  AOI22_X1 U22251 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n19070), .ZN(n19073) );
  NAND2_X1 U22252 ( .A1(n9790), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n19399) );
  OAI211_X1 U22253 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n19074), .A(
        n19073), .B(n19399), .ZN(n19075) );
  AOI211_X1 U22254 ( .C1(n19128), .C2(n19397), .A(n19076), .B(n19075), .ZN(
        n19077) );
  OAI21_X1 U22255 ( .B1(n19079), .B2(n19078), .A(n19077), .ZN(P3_U2818) );
  NAND2_X1 U22256 ( .A1(n19412), .A2(n13344), .ZN(n19417) );
  INV_X1 U22257 ( .A(n19080), .ZN(n19103) );
  NOR2_X1 U22258 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19096) );
  NOR2_X1 U22259 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19081), .ZN(
        n19104) );
  AOI22_X1 U22260 ( .A1(n19412), .A2(n19103), .B1(n19096), .B2(n19104), .ZN(
        n19082) );
  XNOR2_X1 U22261 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19082), .ZN(
        n19403) );
  NOR2_X1 U22262 ( .A1(n19529), .A2(n20095), .ZN(n19087) );
  NAND2_X1 U22263 ( .A1(n19212), .A2(n19121), .ZN(n19199) );
  NOR2_X1 U22264 ( .A1(n19034), .A2(n19652), .ZN(n19094) );
  AOI21_X1 U22265 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19199), .A(
        n19094), .ZN(n19084) );
  OAI22_X1 U22266 ( .A1(n19085), .A2(n19084), .B1(n19209), .B2(n19083), .ZN(
        n19086) );
  AOI211_X1 U22267 ( .C1(n19128), .C2(n19403), .A(n19087), .B(n19086), .ZN(
        n19089) );
  NOR2_X1 U22268 ( .A1(n19412), .A2(n19113), .ZN(n19091) );
  OAI22_X1 U22269 ( .A1(n19407), .A2(n19126), .B1(n19218), .B2(n19405), .ZN(
        n19102) );
  OAI21_X1 U22270 ( .B1(n19091), .B2(n19102), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n19088) );
  OAI211_X1 U22271 ( .C1(n19113), .C2(n19417), .A(n19089), .B(n19088), .ZN(
        P3_U2819) );
  AOI22_X1 U22272 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n19103), .B1(
        n19104), .B2(n13343), .ZN(n19090) );
  XNOR2_X1 U22273 ( .A(n19090), .B(n13342), .ZN(n19426) );
  NOR2_X1 U22274 ( .A1(n19529), .A2(n20092), .ZN(n19098) );
  AOI21_X1 U22275 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n19102), .A(
        n19091), .ZN(n19095) );
  NAND2_X1 U22276 ( .A1(n18170), .A2(n19922), .ZN(n19134) );
  NOR2_X1 U22277 ( .A1(n19092), .A2(n19134), .ZN(n19108) );
  AOI21_X1 U22278 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19199), .A(
        n19108), .ZN(n19093) );
  OAI22_X1 U22279 ( .A1(n19096), .A2(n19095), .B1(n19094), .B2(n19093), .ZN(
        n19097) );
  AOI211_X1 U22280 ( .C1(n19099), .C2(n19174), .A(n19098), .B(n19097), .ZN(
        n19100) );
  OAI21_X1 U22281 ( .B1(n19426), .B2(n19101), .A(n19100), .ZN(P3_U2820) );
  INV_X1 U22282 ( .A(n19102), .ZN(n19112) );
  NOR2_X1 U22283 ( .A1(n19104), .A2(n19103), .ZN(n19105) );
  XNOR2_X1 U22284 ( .A(n19105), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n19434) );
  NAND2_X1 U22285 ( .A1(n9790), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n19435) );
  INV_X1 U22286 ( .A(n19435), .ZN(n19110) );
  NOR2_X1 U22287 ( .A1(n19136), .A2(n19134), .ZN(n19123) );
  AOI22_X1 U22288 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19123), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19199), .ZN(n19107) );
  OAI22_X1 U22289 ( .A1(n19108), .A2(n19107), .B1(n19209), .B2(n19106), .ZN(
        n19109) );
  AOI211_X1 U22290 ( .C1(n19128), .C2(n19434), .A(n19110), .B(n19109), .ZN(
        n19111) );
  OAI221_X1 U22291 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19113), .C1(
        n13343), .C2(n19112), .A(n19111), .ZN(P3_U2821) );
  OAI21_X1 U22292 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n19115), .A(
        n19114), .ZN(n19440) );
  INV_X1 U22293 ( .A(n19116), .ZN(n19117) );
  NAND2_X1 U22294 ( .A1(n19118), .A2(n19117), .ZN(n19438) );
  XNOR2_X1 U22295 ( .A(n19119), .B(n19438), .ZN(n19442) );
  AOI22_X1 U22296 ( .A1(n9790), .A2(P3_REIP_REG_8__SCAN_IN), .B1(n19120), .B2(
        n19174), .ZN(n19125) );
  AOI21_X1 U22297 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(n19652), .ZN(n19122) );
  OAI21_X1 U22298 ( .B1(n18170), .B2(n19121), .A(n19212), .ZN(n19135) );
  OAI22_X1 U22299 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19123), .B1(
        n19122), .B2(n19135), .ZN(n19124) );
  OAI211_X1 U22300 ( .C1(n19438), .C2(n19126), .A(n19125), .B(n19124), .ZN(
        n19127) );
  AOI21_X1 U22301 ( .B1(n19128), .B2(n19442), .A(n19127), .ZN(n19129) );
  OAI21_X1 U22302 ( .B1(n19218), .B2(n19440), .A(n19129), .ZN(P3_U2822) );
  OAI21_X1 U22303 ( .B1(n19132), .B2(n19131), .A(n19130), .ZN(n19133) );
  XNOR2_X1 U22304 ( .A(n19133), .B(n19456), .ZN(n19463) );
  INV_X1 U22305 ( .A(n19134), .ZN(n19137) );
  NOR2_X1 U22306 ( .A1(n19529), .A2(n20086), .ZN(n19455) );
  AOI221_X1 U22307 ( .B1(n19137), .B2(n19136), .C1(n19135), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n19455), .ZN(n19142) );
  AOI21_X1 U22308 ( .B1(n19456), .B2(n19139), .A(n19138), .ZN(n19458) );
  AOI22_X1 U22309 ( .A1(n19205), .A2(n19458), .B1(n19140), .B2(n19174), .ZN(
        n19141) );
  OAI211_X1 U22310 ( .C1(n19218), .C2(n19463), .A(n19142), .B(n19141), .ZN(
        P3_U2823) );
  OAI21_X1 U22311 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19144), .A(
        n19143), .ZN(n19473) );
  NOR2_X1 U22312 ( .A1(n18121), .A2(n19652), .ZN(n19145) );
  AOI22_X1 U22313 ( .A1(n9790), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n19145), .B2(
        n19148), .ZN(n19152) );
  AOI21_X1 U22314 ( .B1(n9928), .B2(n19147), .A(n19146), .ZN(n19471) );
  OAI21_X1 U22315 ( .B1(n19652), .B2(n18121), .A(n19199), .ZN(n19158) );
  OAI22_X1 U22316 ( .A1(n19209), .A2(n19149), .B1(n19148), .B2(n19158), .ZN(
        n19150) );
  AOI21_X1 U22317 ( .B1(n19205), .B2(n19471), .A(n19150), .ZN(n19151) );
  OAI211_X1 U22318 ( .C1(n19218), .C2(n19473), .A(n19152), .B(n19151), .ZN(
        P3_U2824) );
  AOI21_X1 U22319 ( .B1(n19480), .B2(n19154), .A(n19153), .ZN(n19477) );
  NOR2_X1 U22320 ( .A1(n19529), .A2(n20082), .ZN(n19476) );
  AOI21_X1 U22321 ( .B1(n18193), .B2(n19212), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19159) );
  OAI21_X1 U22322 ( .B1(n19157), .B2(n19156), .A(n19155), .ZN(n19474) );
  OAI22_X1 U22323 ( .A1(n19159), .A2(n19158), .B1(n19218), .B2(n19474), .ZN(
        n19160) );
  AOI211_X1 U22324 ( .C1(n19205), .C2(n19477), .A(n19476), .B(n19160), .ZN(
        n19161) );
  OAI21_X1 U22325 ( .B1(n19209), .B2(n19162), .A(n19161), .ZN(P3_U2825) );
  AOI21_X1 U22326 ( .B1(n19165), .B2(n19164), .A(n19163), .ZN(n19184) );
  OAI21_X1 U22327 ( .B1(n19168), .B2(n19167), .A(n19166), .ZN(n19492) );
  OAI22_X1 U22328 ( .A1(n19218), .A2(n19492), .B1(n19652), .B2(n19169), .ZN(
        n19170) );
  AOI21_X1 U22329 ( .B1(n9790), .B2(P3_REIP_REG_4__SCAN_IN), .A(n19170), .ZN(
        n19177) );
  AOI21_X1 U22330 ( .B1(n19173), .B2(n19172), .A(n19171), .ZN(n19487) );
  AOI22_X1 U22331 ( .A1(n19205), .A2(n19487), .B1(n19175), .B2(n19174), .ZN(
        n19176) );
  OAI211_X1 U22332 ( .C1(n19178), .C2(n19184), .A(n19177), .B(n19176), .ZN(
        P3_U2826) );
  OAI21_X1 U22333 ( .B1(n19181), .B2(n19180), .A(n19179), .ZN(n19502) );
  AOI21_X1 U22334 ( .B1(n19496), .B2(n19183), .A(n19182), .ZN(n19500) );
  AOI21_X1 U22335 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19212), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19185) );
  OAI22_X1 U22336 ( .A1(n19209), .A2(n19186), .B1(n19185), .B2(n19184), .ZN(
        n19187) );
  AOI21_X1 U22337 ( .B1(n19205), .B2(n19500), .A(n19187), .ZN(n19188) );
  NAND2_X1 U22338 ( .A1(n9790), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19495) );
  OAI211_X1 U22339 ( .C1(n19218), .C2(n19502), .A(n19188), .B(n19495), .ZN(
        P3_U2827) );
  AOI21_X1 U22340 ( .B1(n19191), .B2(n19190), .A(n19189), .ZN(n19515) );
  INV_X1 U22341 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20076) );
  NOR2_X1 U22342 ( .A1(n19529), .A2(n20076), .ZN(n19517) );
  OAI21_X1 U22343 ( .B1(n19194), .B2(n19193), .A(n19192), .ZN(n19512) );
  OAI22_X1 U22344 ( .A1(n19209), .A2(n19195), .B1(n19218), .B2(n19512), .ZN(
        n19196) );
  AOI211_X1 U22345 ( .C1(n19205), .C2(n19515), .A(n19517), .B(n19196), .ZN(
        n19197) );
  OAI221_X1 U22346 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19652), .C1(
        n19198), .C2(n19212), .A(n19197), .ZN(P3_U2828) );
  INV_X1 U22347 ( .A(n19199), .ZN(n19207) );
  AOI21_X1 U22348 ( .B1(n19201), .B2(n19211), .A(n19200), .ZN(n19523) );
  AOI21_X1 U22349 ( .B1(n19203), .B2(n19210), .A(n19202), .ZN(n19528) );
  OAI22_X1 U22350 ( .A1(n19528), .A2(n19218), .B1(n19529), .B2(n20186), .ZN(
        n19204) );
  AOI21_X1 U22351 ( .B1(n19205), .B2(n19523), .A(n19204), .ZN(n19206) );
  OAI221_X1 U22352 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19209), .C1(
        n19208), .C2(n19207), .A(n19206), .ZN(P3_U2829) );
  NAND2_X1 U22353 ( .A1(n19211), .A2(n19210), .ZN(n19217) );
  INV_X1 U22354 ( .A(n19217), .ZN(n19537) );
  INV_X1 U22355 ( .A(n20056), .ZN(n20209) );
  OAI21_X1 U22356 ( .B1(n19213), .B2(n20209), .A(n19212), .ZN(n19214) );
  AOI22_X1 U22357 ( .A1(n9790), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19214), .ZN(n19215) );
  OAI221_X1 U22358 ( .B1(n19537), .B2(n19218), .C1(n19217), .C2(n19216), .A(
        n19215), .ZN(P3_U2830) );
  OAI22_X1 U22359 ( .A1(n19219), .A2(n19262), .B1(n19232), .B2(n19533), .ZN(
        n19228) );
  NOR2_X1 U22360 ( .A1(n19427), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19506) );
  NOR2_X1 U22361 ( .A1(n19506), .A2(n19220), .ZN(n19258) );
  AOI21_X1 U22362 ( .B1(n19244), .B2(n19258), .A(n19482), .ZN(n19241) );
  AOI22_X1 U22363 ( .A1(n19988), .A2(n19240), .B1(n20014), .B2(n19221), .ZN(
        n19222) );
  OAI211_X1 U22364 ( .C1(n19224), .C2(n19511), .A(n19223), .B(n19222), .ZN(
        n19225) );
  AOI211_X1 U22365 ( .C1(n19381), .C2(n19226), .A(n19241), .B(n19225), .ZN(
        n19234) );
  OAI211_X1 U22366 ( .C1(n20016), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n19234), .ZN(n19227) );
  AOI22_X1 U22367 ( .A1(n19443), .A2(n19229), .B1(n19228), .B2(n19227), .ZN(
        n19231) );
  OAI211_X1 U22368 ( .C1(n19497), .C2(n19232), .A(n19231), .B(n19230), .ZN(
        P3_U2835) );
  INV_X1 U22369 ( .A(n19233), .ZN(n19237) );
  NOR2_X1 U22370 ( .A1(n19529), .A2(n20124), .ZN(n19236) );
  AOI211_X1 U22371 ( .C1(n19466), .C2(n19234), .A(n9790), .B(n10202), .ZN(
        n19235) );
  AOI211_X1 U22372 ( .C1(n19443), .C2(n19237), .A(n19236), .B(n19235), .ZN(
        n19238) );
  OAI21_X1 U22373 ( .B1(n19262), .B2(n19239), .A(n19238), .ZN(P3_U2836) );
  NOR3_X1 U22374 ( .A1(n19242), .A2(n19241), .A3(n19240), .ZN(n19246) );
  AOI21_X1 U22375 ( .B1(n19244), .B2(n19243), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19245) );
  NOR3_X1 U22376 ( .A1(n19246), .A2(n19245), .A3(n19533), .ZN(n19247) );
  AOI211_X1 U22377 ( .C1(n19525), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n19248), .B(n19247), .ZN(n19253) );
  AOI22_X1 U22378 ( .A1(n19251), .A2(n19250), .B1(n19398), .B2(n19249), .ZN(
        n19252) );
  OAI211_X1 U22379 ( .C1(n19536), .C2(n19254), .A(n19253), .B(n19252), .ZN(
        P3_U2837) );
  AOI22_X1 U22380 ( .A1(n19976), .A2(n19256), .B1(n19381), .B2(n19255), .ZN(
        n19257) );
  OAI211_X1 U22381 ( .C1(n19482), .C2(n19258), .A(n19257), .B(n19497), .ZN(
        n19261) );
  OAI21_X1 U22382 ( .B1(n19259), .B2(n20009), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19260) );
  OAI21_X1 U22383 ( .B1(n19261), .B2(n19260), .A(n19529), .ZN(n19272) );
  INV_X1 U22384 ( .A(n19364), .ZN(n19448) );
  OAI21_X1 U22385 ( .B1(n19448), .B2(n19261), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n19268) );
  INV_X1 U22386 ( .A(n19262), .ZN(n19264) );
  AOI22_X1 U22387 ( .A1(n19443), .A2(n19265), .B1(n19264), .B2(n19263), .ZN(
        n19267) );
  OAI211_X1 U22388 ( .C1(n19272), .C2(n19268), .A(n19267), .B(n19266), .ZN(
        P3_U2838) );
  AOI21_X1 U22389 ( .B1(n19269), .B2(n19497), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19273) );
  AOI22_X1 U22390 ( .A1(n9790), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n19443), 
        .B2(n19270), .ZN(n19271) );
  OAI21_X1 U22391 ( .B1(n19273), .B2(n19272), .A(n19271), .ZN(P3_U2839) );
  OAI22_X1 U22392 ( .A1(n19350), .A2(n19406), .B1(n19347), .B2(n19511), .ZN(
        n19291) );
  NAND2_X1 U22393 ( .A1(n19511), .A2(n19406), .ZN(n19404) );
  INV_X1 U22394 ( .A(n19306), .ZN(n19276) );
  OAI21_X1 U22395 ( .B1(n19274), .B2(n19319), .A(n19977), .ZN(n19275) );
  OAI221_X1 U22396 ( .B1(n20016), .B2(n19277), .C1(n20016), .C2(n19276), .A(
        n19275), .ZN(n19304) );
  AOI21_X1 U22397 ( .B1(n19278), .B2(n19404), .A(n19304), .ZN(n19279) );
  OAI21_X1 U22398 ( .B1(n20016), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n19279), .ZN(n19293) );
  AOI211_X1 U22399 ( .C1(n19419), .C2(n19296), .A(n19291), .B(n19293), .ZN(
        n19284) );
  INV_X1 U22400 ( .A(n19280), .ZN(n19294) );
  AOI22_X1 U22401 ( .A1(n19977), .A2(n19294), .B1(n20014), .B2(n19281), .ZN(
        n19283) );
  OAI222_X1 U22402 ( .A1(n19289), .A2(n19284), .B1(n19289), .B2(n19283), .C1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n19282), .ZN(n19286) );
  AOI22_X1 U22403 ( .A1(n19466), .A2(n19286), .B1(n19443), .B2(n19285), .ZN(
        n19288) );
  OAI211_X1 U22404 ( .C1(n19497), .C2(n19289), .A(n19288), .B(n19287), .ZN(
        P3_U2840) );
  NAND3_X1 U22405 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n19466), .A3(
        n19290), .ZN(n19316) );
  NOR2_X1 U22406 ( .A1(n19977), .A2(n20014), .ZN(n19524) );
  INV_X1 U22407 ( .A(n19524), .ZN(n19295) );
  AOI21_X1 U22408 ( .B1(n19338), .B2(n19292), .A(n19427), .ZN(n19305) );
  AOI211_X1 U22409 ( .C1(n19295), .C2(n19294), .A(n19305), .B(n19293), .ZN(
        n19297) );
  AOI211_X1 U22410 ( .C1(n19340), .C2(n19297), .A(n9790), .B(n19296), .ZN(
        n19298) );
  AOI21_X1 U22411 ( .B1(n19443), .B2(n19299), .A(n19298), .ZN(n19301) );
  OAI211_X1 U22412 ( .C1(n19302), .C2(n19316), .A(n19301), .B(n19300), .ZN(
        P3_U2841) );
  AOI22_X1 U22413 ( .A1(n9790), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n19398), 
        .B2(n19303), .ZN(n19310) );
  AOI211_X1 U22414 ( .C1(n19306), .C2(n19404), .A(n19305), .B(n19304), .ZN(
        n19307) );
  AOI21_X1 U22415 ( .B1(n19340), .B2(n19307), .A(n9790), .ZN(n19313) );
  NOR3_X1 U22416 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19524), .A3(
        n20047), .ZN(n19308) );
  OAI21_X1 U22417 ( .B1(n19313), .B2(n19308), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19309) );
  OAI211_X1 U22418 ( .C1(n19311), .C2(n19316), .A(n19310), .B(n19309), .ZN(
        P3_U2842) );
  AOI22_X1 U22419 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19313), .B1(
        n19398), .B2(n19312), .ZN(n19315) );
  NAND2_X1 U22420 ( .A1(n9790), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n19314) );
  OAI211_X1 U22421 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n19316), .A(
        n19315), .B(n19314), .ZN(P3_U2843) );
  NOR3_X1 U22422 ( .A1(n19506), .A2(n19317), .A3(n19341), .ZN(n19321) );
  AOI22_X1 U22423 ( .A1(n19977), .A2(n19319), .B1(n19318), .B2(n19404), .ZN(
        n19320) );
  OAI211_X1 U22424 ( .C1(n19482), .C2(n19321), .A(n19340), .B(n19320), .ZN(
        n19332) );
  OAI221_X1 U22425 ( .B1(n19332), .B2(n19333), .C1(n19332), .C2(n19505), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19330) );
  AOI22_X1 U22426 ( .A1(n19977), .A2(n19504), .B1(n19483), .B2(n19508), .ZN(
        n19494) );
  INV_X1 U22427 ( .A(n19322), .ZN(n19323) );
  NOR2_X1 U22428 ( .A1(n19494), .A2(n19323), .ZN(n19464) );
  INV_X1 U22429 ( .A(n19464), .ZN(n19457) );
  NAND2_X1 U22430 ( .A1(n19325), .A2(n19365), .ZN(n19393) );
  NAND2_X1 U22431 ( .A1(n19466), .A2(n19393), .ZN(n19437) );
  NOR2_X1 U22432 ( .A1(n19326), .A2(n19437), .ZN(n19342) );
  AOI22_X1 U22433 ( .A1(n19443), .A2(n19328), .B1(n19342), .B2(n19327), .ZN(
        n19329) );
  OAI221_X1 U22434 ( .B1(n9790), .B2(n19330), .C1(n19529), .C2(n20108), .A(
        n19329), .ZN(P3_U2844) );
  AOI22_X1 U22435 ( .A1(n9790), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n19443), 
        .B2(n19331), .ZN(n19336) );
  NAND3_X1 U22436 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n19529), .A3(
        n19332), .ZN(n19335) );
  NAND3_X1 U22437 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19342), .A3(
        n19333), .ZN(n19334) );
  NAND3_X1 U22438 ( .A1(n19336), .A2(n19335), .A3(n19334), .ZN(P3_U2845) );
  INV_X1 U22439 ( .A(n19398), .ZN(n19425) );
  NOR2_X1 U22440 ( .A1(n19337), .A2(n20009), .ZN(n19409) );
  OR2_X1 U22441 ( .A1(n20016), .A2(n19378), .ZN(n19420) );
  OAI211_X1 U22442 ( .C1(n19338), .C2(n19427), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n19420), .ZN(n19339) );
  AOI211_X1 U22443 ( .C1(n19419), .C2(n19349), .A(n19409), .B(n19339), .ZN(
        n19348) );
  AOI221_X1 U22444 ( .B1(n19364), .B2(n19340), .C1(n19348), .C2(n19340), .A(
        n9790), .ZN(n19343) );
  AOI22_X1 U22445 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19343), .B1(
        n19342), .B2(n19341), .ZN(n19345) );
  OAI211_X1 U22446 ( .C1(n19346), .C2(n19425), .A(n19345), .B(n19344), .ZN(
        P3_U2846) );
  NOR2_X1 U22447 ( .A1(n19347), .A2(n19511), .ZN(n19356) );
  AOI221_X1 U22448 ( .B1(n19349), .B2(n19351), .C1(n19365), .C2(n19351), .A(
        n19348), .ZN(n19354) );
  AOI211_X1 U22449 ( .C1(n19352), .C2(n19351), .A(n19350), .B(n19406), .ZN(
        n19353) );
  AOI211_X1 U22450 ( .C1(n19356), .C2(n19355), .A(n19354), .B(n19353), .ZN(
        n19360) );
  AOI22_X1 U22451 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19525), .B1(
        n19443), .B2(n19357), .ZN(n19359) );
  OAI211_X1 U22452 ( .C1(n19360), .C2(n19533), .A(n19359), .B(n19358), .ZN(
        P3_U2847) );
  INV_X1 U22453 ( .A(n19361), .ZN(n19362) );
  AOI221_X1 U22454 ( .B1(n19362), .B2(n20014), .C1(n19429), .C2(n20014), .A(
        n19409), .ZN(n19384) );
  OAI211_X1 U22455 ( .C1(n19364), .C2(n19363), .A(n19384), .B(n19420), .ZN(
        n19368) );
  OAI21_X1 U22456 ( .B1(n19366), .B2(n19365), .A(n19369), .ZN(n19367) );
  OAI21_X1 U22457 ( .B1(n19369), .B2(n19368), .A(n19367), .ZN(n19377) );
  AOI22_X1 U22458 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19525), .B1(
        n9790), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n19376) );
  OAI22_X1 U22459 ( .A1(n19439), .A2(n19371), .B1(n19425), .B2(n19370), .ZN(
        n19372) );
  AOI21_X1 U22460 ( .B1(n19374), .B2(n19373), .A(n19372), .ZN(n19375) );
  OAI211_X1 U22461 ( .C1(n19533), .C2(n19377), .A(n19376), .B(n19375), .ZN(
        P3_U2848) );
  OAI21_X1 U22462 ( .B1(n20016), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19396) );
  AOI21_X1 U22463 ( .B1(n19412), .B2(n19378), .A(n20016), .ZN(n19379) );
  AOI21_X1 U22464 ( .B1(n19977), .B2(n19392), .A(n19379), .ZN(n19413) );
  AOI22_X1 U22465 ( .A1(n19976), .A2(n19382), .B1(n19381), .B2(n19380), .ZN(
        n19383) );
  NAND3_X1 U22466 ( .A1(n19413), .A2(n19384), .A3(n19383), .ZN(n19395) );
  AOI211_X1 U22467 ( .C1(n19419), .C2(n19396), .A(n19533), .B(n19395), .ZN(
        n19386) );
  NOR3_X1 U22468 ( .A1(n9790), .A2(n19386), .A3(n19385), .ZN(n19388) );
  AOI211_X1 U22469 ( .C1(n19389), .C2(n19443), .A(n19388), .B(n19387), .ZN(
        n19390) );
  OAI21_X1 U22470 ( .B1(n19437), .B2(n19391), .A(n19390), .ZN(P3_U2849) );
  INV_X1 U22471 ( .A(n19392), .ZN(n19394) );
  AOI21_X1 U22472 ( .B1(n19394), .B2(n19393), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19402) );
  OAI21_X1 U22473 ( .B1(n19396), .B2(n19395), .A(n19466), .ZN(n19401) );
  AOI22_X1 U22474 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19525), .B1(
        n19398), .B2(n19397), .ZN(n19400) );
  OAI211_X1 U22475 ( .C1(n19402), .C2(n19401), .A(n19400), .B(n19399), .ZN(
        P3_U2850) );
  AOI22_X1 U22476 ( .A1(n9790), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n19443), 
        .B2(n19403), .ZN(n19416) );
  INV_X1 U22477 ( .A(n19404), .ZN(n19411) );
  OAI22_X1 U22478 ( .A1(n19407), .A2(n19406), .B1(n19511), .B2(n19405), .ZN(
        n19408) );
  NOR3_X1 U22479 ( .A1(n19409), .A2(n19533), .A3(n19408), .ZN(n19432) );
  OAI21_X1 U22480 ( .B1(n13343), .B2(n19429), .A(n20014), .ZN(n19410) );
  OAI211_X1 U22481 ( .C1(n19412), .C2(n19411), .A(n19432), .B(n19410), .ZN(
        n19418) );
  OAI21_X1 U22482 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n19427), .A(
        n19413), .ZN(n19414) );
  OAI211_X1 U22483 ( .C1(n19418), .C2(n19414), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19529), .ZN(n19415) );
  OAI211_X1 U22484 ( .C1(n19417), .C2(n19437), .A(n19416), .B(n19415), .ZN(
        P3_U2851) );
  AOI21_X1 U22485 ( .B1(n13343), .B2(n19419), .A(n19418), .ZN(n19421) );
  AOI21_X1 U22486 ( .B1(n19421), .B2(n19420), .A(n13342), .ZN(n19423) );
  NOR3_X1 U22487 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n13343), .A3(
        n19437), .ZN(n19422) );
  AOI221_X1 U22488 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n9790), .C1(n19423), 
        .C2(n19529), .A(n19422), .ZN(n19424) );
  OAI21_X1 U22489 ( .B1(n19426), .B2(n19425), .A(n19424), .ZN(P3_U2852) );
  AOI21_X1 U22490 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n19427), .A(
        n19482), .ZN(n19430) );
  AOI22_X1 U22491 ( .A1(n19430), .A2(n19429), .B1(n19988), .B2(n19428), .ZN(
        n19431) );
  AOI211_X1 U22492 ( .C1(n19432), .C2(n19431), .A(n9790), .B(n13343), .ZN(
        n19433) );
  AOI21_X1 U22493 ( .B1(n19443), .B2(n19434), .A(n19433), .ZN(n19436) );
  OAI211_X1 U22494 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n19437), .A(
        n19436), .B(n19435), .ZN(P3_U2853) );
  OAI22_X1 U22495 ( .A1(n19536), .A2(n19440), .B1(n19439), .B2(n19438), .ZN(
        n19441) );
  AOI21_X1 U22496 ( .B1(n19443), .B2(n19442), .A(n19441), .ZN(n19454) );
  NAND2_X1 U22497 ( .A1(n9790), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n19453) );
  AOI21_X1 U22498 ( .B1(n19977), .B2(n19444), .A(n19506), .ZN(n19445) );
  OAI21_X1 U22499 ( .B1(n19446), .B2(n19482), .A(n19445), .ZN(n19465) );
  AOI211_X1 U22500 ( .C1(n19448), .C2(n19468), .A(n19456), .B(n19465), .ZN(
        n19447) );
  NOR2_X1 U22501 ( .A1(n19447), .A2(n19533), .ZN(n19460) );
  OAI221_X1 U22502 ( .B1(n19525), .B2(n19460), .C1(n19525), .C2(n19448), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n19452) );
  NAND4_X1 U22503 ( .A1(n19466), .A2(n19450), .A3(n19464), .A4(n19449), .ZN(
        n19451) );
  NAND4_X1 U22504 ( .A1(n19454), .A2(n19453), .A3(n19452), .A4(n19451), .ZN(
        P3_U2854) );
  AOI21_X1 U22505 ( .B1(n19525), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19455), .ZN(n19462) );
  OAI21_X1 U22506 ( .B1(n19468), .B2(n19457), .A(n19456), .ZN(n19459) );
  NOR2_X1 U22507 ( .A1(n19983), .A2(n19533), .ZN(n19532) );
  AOI22_X1 U22508 ( .A1(n19460), .A2(n19459), .B1(n19458), .B2(n19532), .ZN(
        n19461) );
  OAI211_X1 U22509 ( .C1(n19536), .C2(n19463), .A(n19462), .B(n19461), .ZN(
        P3_U2855) );
  NAND2_X1 U22510 ( .A1(n19466), .A2(n19464), .ZN(n19469) );
  AOI21_X1 U22511 ( .B1(n19466), .B2(n19465), .A(n19525), .ZN(n19479) );
  NAND2_X1 U22512 ( .A1(n9790), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n19467) );
  OAI221_X1 U22513 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19469), .C1(
        n19468), .C2(n19479), .A(n19467), .ZN(n19470) );
  AOI21_X1 U22514 ( .B1(n19532), .B2(n19471), .A(n19470), .ZN(n19472) );
  OAI21_X1 U22515 ( .B1(n19536), .B2(n19473), .A(n19472), .ZN(P3_U2856) );
  NOR2_X1 U22516 ( .A1(n19494), .A2(n19533), .ZN(n19489) );
  NAND3_X1 U22517 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n19489), .ZN(n19481) );
  NOR2_X1 U22518 ( .A1(n19536), .A2(n19474), .ZN(n19475) );
  AOI211_X1 U22519 ( .C1(n19532), .C2(n19477), .A(n19476), .B(n19475), .ZN(
        n19478) );
  OAI221_X1 U22520 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n19481), .C1(
        n19480), .C2(n19479), .A(n19478), .ZN(P3_U2857) );
  NOR2_X1 U22521 ( .A1(n19529), .A2(n20080), .ZN(n19486) );
  OAI22_X1 U22522 ( .A1(n19483), .A2(n19482), .B1(n20009), .B2(n19504), .ZN(
        n19484) );
  NOR3_X1 U22523 ( .A1(n19506), .A2(n19496), .A3(n19484), .ZN(n19493) );
  AOI221_X1 U22524 ( .B1(n19493), .B2(n19497), .C1(n19520), .C2(n19497), .A(
        n19488), .ZN(n19485) );
  AOI211_X1 U22525 ( .C1(n19487), .C2(n19532), .A(n19486), .B(n19485), .ZN(
        n19491) );
  NAND3_X1 U22526 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19489), .A3(
        n19488), .ZN(n19490) );
  OAI211_X1 U22527 ( .C1(n19492), .C2(n19536), .A(n19491), .B(n19490), .ZN(
        P3_U2858) );
  AOI211_X1 U22528 ( .C1(n19494), .C2(n19496), .A(n19493), .B(n19533), .ZN(
        n19499) );
  OAI21_X1 U22529 ( .B1(n19497), .B2(n19496), .A(n19495), .ZN(n19498) );
  AOI211_X1 U22530 ( .C1(n19500), .C2(n19532), .A(n19499), .B(n19498), .ZN(
        n19501) );
  OAI21_X1 U22531 ( .B1(n19536), .B2(n19502), .A(n19501), .ZN(P3_U2859) );
  INV_X1 U22532 ( .A(n19983), .ZN(n19516) );
  NAND2_X1 U22533 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19503) );
  AOI221_X1 U22534 ( .B1(n19507), .B2(n19504), .C1(n19503), .C2(n19504), .A(
        n20009), .ZN(n19514) );
  OAI211_X1 U22535 ( .C1(n19506), .C2(n9952), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n19505), .ZN(n19510) );
  NAND3_X1 U22536 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19508), .A3(
        n19507), .ZN(n19509) );
  OAI211_X1 U22537 ( .C1(n19512), .C2(n19511), .A(n19510), .B(n19509), .ZN(
        n19513) );
  AOI211_X1 U22538 ( .C1(n19516), .C2(n19515), .A(n19514), .B(n19513), .ZN(
        n19519) );
  AOI21_X1 U22539 ( .B1(n19525), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n19517), .ZN(n19518) );
  OAI21_X1 U22540 ( .B1(n19519), .B2(n19533), .A(n19518), .ZN(P3_U2860) );
  NOR2_X1 U22541 ( .A1(n19529), .A2(n20186), .ZN(n19522) );
  AOI211_X1 U22542 ( .C1(n20016), .C2(n20181), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n19520), .ZN(n19521) );
  AOI211_X1 U22543 ( .C1(n19523), .C2(n19532), .A(n19522), .B(n19521), .ZN(
        n19527) );
  NOR3_X1 U22544 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19524), .A3(
        n19533), .ZN(n19530) );
  OAI21_X1 U22545 ( .B1(n19525), .B2(n19530), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19526) );
  OAI211_X1 U22546 ( .C1(n19528), .C2(n19536), .A(n19527), .B(n19526), .ZN(
        P3_U2861) );
  INV_X1 U22547 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n20192) );
  NOR2_X1 U22548 ( .A1(n19529), .A2(n20192), .ZN(n19531) );
  AOI211_X1 U22549 ( .C1(n19532), .C2(n19537), .A(n19531), .B(n19530), .ZN(
        n19535) );
  OAI211_X1 U22550 ( .C1(n19988), .C2(n19533), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n19529), .ZN(n19534) );
  OAI211_X1 U22551 ( .C1(n19537), .C2(n19536), .A(n19535), .B(n19534), .ZN(
        P3_U2862) );
  AOI21_X1 U22552 ( .B1(n19540), .B2(n19539), .A(n19538), .ZN(n20041) );
  OAI21_X1 U22553 ( .B1(n20041), .B2(n19588), .A(n19546), .ZN(n19541) );
  OAI221_X1 U22554 ( .B1(n20019), .B2(n19542), .C1(n20019), .C2(n19546), .A(
        n19541), .ZN(P3_U2863) );
  NOR2_X1 U22555 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20029), .ZN(
        n19813) );
  NAND2_X1 U22556 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20029), .ZN(
        n19676) );
  INV_X1 U22557 ( .A(n19676), .ZN(n19721) );
  NOR2_X1 U22558 ( .A1(n19813), .A2(n19721), .ZN(n19544) );
  OAI22_X1 U22559 ( .A1(n19545), .A2(n20029), .B1(n19544), .B2(n19543), .ZN(
        P3_U2866) );
  NOR2_X1 U22560 ( .A1(n20030), .A2(n19546), .ZN(P3_U2867) );
  NAND2_X1 U22561 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19922), .ZN(n19890) );
  NOR3_X1 U22562 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20026), .A3(
        n20029), .ZN(n19921) );
  NAND2_X1 U22563 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19921), .ZN(
        n19963) );
  NOR2_X2 U22564 ( .A1(n19651), .A2(n19547), .ZN(n19917) );
  NOR2_X1 U22565 ( .A1(n20029), .A2(n19697), .ZN(n19920) );
  INV_X1 U22566 ( .A(n19920), .ZN(n19916) );
  NOR2_X2 U22567 ( .A1(n20019), .A2(n19916), .ZN(n19959) );
  NAND2_X1 U22568 ( .A1(n20021), .A2(n20019), .ZN(n20022) );
  NAND2_X1 U22569 ( .A1(n20026), .A2(n20029), .ZN(n19607) );
  NOR2_X2 U22570 ( .A1(n20022), .A2(n19607), .ZN(n19643) );
  NOR2_X1 U22571 ( .A1(n19959), .A2(n19643), .ZN(n19609) );
  NOR2_X1 U22572 ( .A1(n20050), .A2(n19609), .ZN(n19582) );
  NOR2_X2 U22573 ( .A1(n19652), .A2(n19548), .ZN(n19923) );
  NOR2_X2 U22574 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19916), .ZN(
        n19906) );
  AOI22_X1 U22575 ( .A1(n19917), .A2(n19582), .B1(n19923), .B2(n19906), .ZN(
        n19554) );
  INV_X1 U22576 ( .A(n19963), .ZN(n19969) );
  NOR2_X1 U22577 ( .A1(n19969), .A2(n19906), .ZN(n19882) );
  OAI21_X1 U22578 ( .B1(n20019), .B2(n20153), .A(n19886), .ZN(n19743) );
  OAI22_X1 U22579 ( .A1(n19652), .A2(n19882), .B1(n19743), .B2(n19609), .ZN(
        n19549) );
  INV_X1 U22580 ( .A(n19549), .ZN(n19585) );
  NOR2_X1 U22581 ( .A1(n19551), .A2(n19550), .ZN(n19572) );
  INV_X1 U22582 ( .A(n19572), .ZN(n19583) );
  NOR2_X1 U22583 ( .A1(n19552), .A2(n19583), .ZN(n19887) );
  AOI22_X1 U22584 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19585), .B1(
        n19887), .B2(n19643), .ZN(n19553) );
  OAI211_X1 U22585 ( .C1(n19890), .C2(n19963), .A(n19554), .B(n19553), .ZN(
        P3_U2868) );
  NAND2_X1 U22586 ( .A1(n19572), .A2(n19555), .ZN(n19932) );
  INV_X1 U22587 ( .A(n19643), .ZN(n19650) );
  NOR2_X2 U22588 ( .A1(n19652), .A2(n20549), .ZN(n19929) );
  NOR2_X2 U22589 ( .A1(n19651), .A2(n19556), .ZN(n19927) );
  AOI22_X1 U22590 ( .A1(n19929), .A2(n19906), .B1(n19927), .B2(n19582), .ZN(
        n19558) );
  AND2_X1 U22591 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19922), .ZN(n19928) );
  AOI22_X1 U22592 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19585), .B1(
        n19928), .B2(n19969), .ZN(n19557) );
  OAI211_X1 U22593 ( .C1(n19932), .C2(n19650), .A(n19558), .B(n19557), .ZN(
        P3_U2869) );
  NAND2_X1 U22594 ( .A1(n19572), .A2(n19559), .ZN(n19938) );
  NOR2_X2 U22595 ( .A1(n19651), .A2(n19560), .ZN(n19933) );
  AND2_X1 U22596 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19922), .ZN(n19934) );
  AOI22_X1 U22597 ( .A1(n19933), .A2(n19582), .B1(n19934), .B2(n19969), .ZN(
        n19562) );
  NOR2_X2 U22598 ( .A1(n19652), .A2(n20555), .ZN(n19935) );
  AOI22_X1 U22599 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19585), .B1(
        n19935), .B2(n19906), .ZN(n19561) );
  OAI211_X1 U22600 ( .C1(n19938), .C2(n19650), .A(n19562), .B(n19561), .ZN(
        P3_U2870) );
  NAND2_X1 U22601 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19922), .ZN(n19898) );
  NAND2_X1 U22602 ( .A1(n19922), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19944) );
  INV_X1 U22603 ( .A(n19944), .ZN(n19895) );
  NOR2_X2 U22604 ( .A1(n19651), .A2(n19563), .ZN(n19939) );
  AOI22_X1 U22605 ( .A1(n19895), .A2(n19906), .B1(n19939), .B2(n19582), .ZN(
        n19566) );
  NOR2_X2 U22606 ( .A1(n19564), .A2(n19583), .ZN(n19941) );
  AOI22_X1 U22607 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19585), .B1(
        n19941), .B2(n19643), .ZN(n19565) );
  OAI211_X1 U22608 ( .C1(n19898), .C2(n19963), .A(n19566), .B(n19565), .ZN(
        P3_U2871) );
  NAND2_X1 U22609 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19922), .ZN(n19902) );
  NOR2_X2 U22610 ( .A1(n19651), .A2(n19567), .ZN(n19945) );
  NOR2_X2 U22611 ( .A1(n19652), .A2(n20562), .ZN(n19947) );
  AOI22_X1 U22612 ( .A1(n19945), .A2(n19582), .B1(n19947), .B2(n19906), .ZN(
        n19570) );
  NOR2_X1 U22613 ( .A1(n19568), .A2(n19583), .ZN(n19899) );
  AOI22_X1 U22614 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19585), .B1(
        n19899), .B2(n19643), .ZN(n19569) );
  OAI211_X1 U22615 ( .C1(n19902), .C2(n19963), .A(n19570), .B(n19569), .ZN(
        P3_U2872) );
  NAND2_X1 U22616 ( .A1(n19572), .A2(n19571), .ZN(n19956) );
  NOR2_X2 U22617 ( .A1(n19573), .A2(n19652), .ZN(n19953) );
  NOR2_X2 U22618 ( .A1(n19651), .A2(n19574), .ZN(n19951) );
  AOI22_X1 U22619 ( .A1(n19953), .A2(n19969), .B1(n19951), .B2(n19582), .ZN(
        n19576) );
  NOR2_X2 U22620 ( .A1(n19652), .A2(n20567), .ZN(n19952) );
  AOI22_X1 U22621 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19585), .B1(
        n19952), .B2(n19906), .ZN(n19575) );
  OAI211_X1 U22622 ( .C1(n19956), .C2(n19650), .A(n19576), .B(n19575), .ZN(
        P3_U2873) );
  NAND2_X1 U22623 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19922), .ZN(n19852) );
  NOR2_X2 U22624 ( .A1(n19577), .A2(n19651), .ZN(n19957) );
  NOR2_X1 U22625 ( .A1(n19578), .A2(n19652), .ZN(n19849) );
  AOI22_X1 U22626 ( .A1(n19957), .A2(n19582), .B1(n19849), .B2(n19906), .ZN(
        n19581) );
  NOR2_X2 U22627 ( .A1(n19579), .A2(n19583), .ZN(n19960) );
  AOI22_X1 U22628 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19585), .B1(
        n19960), .B2(n19643), .ZN(n19580) );
  OAI211_X1 U22629 ( .C1(n19852), .C2(n19963), .A(n19581), .B(n19580), .ZN(
        P3_U2874) );
  NAND2_X1 U22630 ( .A1(n19922), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19880) );
  NOR2_X2 U22631 ( .A1(n20578), .A2(n19652), .ZN(n19970) );
  AND2_X1 U22632 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n19886), .ZN(n19966) );
  AOI22_X1 U22633 ( .A1(n19970), .A2(n19906), .B1(n19966), .B2(n19582), .ZN(
        n19587) );
  NOR2_X1 U22634 ( .A1(n19584), .A2(n19583), .ZN(n19876) );
  AOI22_X1 U22635 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19585), .B1(
        n19876), .B2(n19643), .ZN(n19586) );
  OAI211_X1 U22636 ( .C1(n19880), .C2(n19963), .A(n19587), .B(n19586), .ZN(
        P3_U2875) );
  INV_X1 U22637 ( .A(n19887), .ZN(n19926) );
  NOR2_X1 U22638 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20019), .ZN(
        n19766) );
  INV_X1 U22639 ( .A(n19607), .ZN(n19630) );
  NAND2_X1 U22640 ( .A1(n19766), .A2(n19630), .ZN(n19675) );
  INV_X1 U22641 ( .A(n19890), .ZN(n19918) );
  AOI22_X1 U22642 ( .A1(n19918), .A2(n19906), .B1(n19917), .B2(n19603), .ZN(
        n19590) );
  NOR2_X1 U22643 ( .A1(n19651), .A2(n19588), .ZN(n19919) );
  AND2_X1 U22644 ( .A1(n20021), .A2(n19919), .ZN(n19768) );
  AOI22_X1 U22645 ( .A1(n19922), .A2(n19920), .B1(n19630), .B2(n19768), .ZN(
        n19604) );
  AOI22_X1 U22646 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19604), .B1(
        n19923), .B2(n19959), .ZN(n19589) );
  OAI211_X1 U22647 ( .C1(n19926), .C2(n19675), .A(n19590), .B(n19589), .ZN(
        P3_U2876) );
  AOI22_X1 U22648 ( .A1(n19927), .A2(n19603), .B1(n19928), .B2(n19906), .ZN(
        n19592) );
  AOI22_X1 U22649 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19604), .B1(
        n19929), .B2(n19959), .ZN(n19591) );
  OAI211_X1 U22650 ( .C1(n19932), .C2(n19675), .A(n19592), .B(n19591), .ZN(
        P3_U2877) );
  AOI22_X1 U22651 ( .A1(n19935), .A2(n19959), .B1(n19933), .B2(n19603), .ZN(
        n19594) );
  AOI22_X1 U22652 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19604), .B1(
        n19934), .B2(n19906), .ZN(n19593) );
  OAI211_X1 U22653 ( .C1(n19938), .C2(n19675), .A(n19594), .B(n19593), .ZN(
        P3_U2878) );
  INV_X1 U22654 ( .A(n19906), .ZN(n19915) );
  AOI22_X1 U22655 ( .A1(n19895), .A2(n19959), .B1(n19939), .B2(n19603), .ZN(
        n19596) );
  INV_X1 U22656 ( .A(n19675), .ZN(n19666) );
  AOI22_X1 U22657 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19604), .B1(
        n19941), .B2(n19666), .ZN(n19595) );
  OAI211_X1 U22658 ( .C1(n19898), .C2(n19915), .A(n19596), .B(n19595), .ZN(
        P3_U2879) );
  INV_X1 U22659 ( .A(n19899), .ZN(n19950) );
  INV_X1 U22660 ( .A(n19902), .ZN(n19946) );
  AOI22_X1 U22661 ( .A1(n19946), .A2(n19906), .B1(n19945), .B2(n19603), .ZN(
        n19598) );
  AOI22_X1 U22662 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19604), .B1(
        n19947), .B2(n19959), .ZN(n19597) );
  OAI211_X1 U22663 ( .C1(n19950), .C2(n19675), .A(n19598), .B(n19597), .ZN(
        P3_U2880) );
  AOI22_X1 U22664 ( .A1(n19952), .A2(n19959), .B1(n19951), .B2(n19603), .ZN(
        n19600) );
  AOI22_X1 U22665 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19604), .B1(
        n19953), .B2(n19906), .ZN(n19599) );
  OAI211_X1 U22666 ( .C1(n19956), .C2(n19675), .A(n19600), .B(n19599), .ZN(
        P3_U2881) );
  AOI22_X1 U22667 ( .A1(n19957), .A2(n19603), .B1(n19849), .B2(n19959), .ZN(
        n19602) );
  AOI22_X1 U22668 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19604), .B1(
        n19960), .B2(n19666), .ZN(n19601) );
  OAI211_X1 U22669 ( .C1(n19852), .C2(n19915), .A(n19602), .B(n19601), .ZN(
        P3_U2882) );
  INV_X1 U22670 ( .A(n19876), .ZN(n19975) );
  INV_X1 U22671 ( .A(n19880), .ZN(n19967) );
  AOI22_X1 U22672 ( .A1(n19967), .A2(n19906), .B1(n19966), .B2(n19603), .ZN(
        n19606) );
  AOI22_X1 U22673 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19604), .B1(
        n19970), .B2(n19959), .ZN(n19605) );
  OAI211_X1 U22674 ( .C1(n19975), .C2(n19675), .A(n19606), .B(n19605), .ZN(
        P3_U2883) );
  NOR2_X1 U22675 ( .A1(n20021), .A2(n19607), .ZN(n19677) );
  NAND2_X1 U22676 ( .A1(n19677), .A2(n20019), .ZN(n19663) );
  NOR2_X1 U22677 ( .A1(n19666), .A2(n19693), .ZN(n19653) );
  NOR2_X1 U22678 ( .A1(n20050), .A2(n19653), .ZN(n19625) );
  AOI22_X1 U22679 ( .A1(n19918), .A2(n19959), .B1(n19917), .B2(n19625), .ZN(
        n19612) );
  INV_X1 U22680 ( .A(n19608), .ZN(n19883) );
  OAI21_X1 U22681 ( .B1(n19609), .B2(n19883), .A(n19653), .ZN(n19610) );
  OAI211_X1 U22682 ( .C1(n19693), .C2(n20153), .A(n19886), .B(n19610), .ZN(
        n19626) );
  AOI22_X1 U22683 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19626), .B1(
        n19923), .B2(n19643), .ZN(n19611) );
  OAI211_X1 U22684 ( .C1(n19926), .C2(n19663), .A(n19612), .B(n19611), .ZN(
        P3_U2884) );
  AOI22_X1 U22685 ( .A1(n19927), .A2(n19625), .B1(n19928), .B2(n19959), .ZN(
        n19614) );
  AOI22_X1 U22686 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19626), .B1(
        n19929), .B2(n19643), .ZN(n19613) );
  OAI211_X1 U22687 ( .C1(n19932), .C2(n19663), .A(n19614), .B(n19613), .ZN(
        P3_U2885) );
  AOI22_X1 U22688 ( .A1(n19935), .A2(n19643), .B1(n19933), .B2(n19625), .ZN(
        n19616) );
  AOI22_X1 U22689 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19626), .B1(
        n19934), .B2(n19959), .ZN(n19615) );
  OAI211_X1 U22690 ( .C1(n19938), .C2(n19663), .A(n19616), .B(n19615), .ZN(
        P3_U2886) );
  INV_X1 U22691 ( .A(n19898), .ZN(n19940) );
  AOI22_X1 U22692 ( .A1(n19940), .A2(n19959), .B1(n19939), .B2(n19625), .ZN(
        n19618) );
  AOI22_X1 U22693 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19626), .B1(
        n19941), .B2(n19693), .ZN(n19617) );
  OAI211_X1 U22694 ( .C1(n19944), .C2(n19650), .A(n19618), .B(n19617), .ZN(
        P3_U2887) );
  AOI22_X1 U22695 ( .A1(n19945), .A2(n19625), .B1(n19947), .B2(n19643), .ZN(
        n19620) );
  AOI22_X1 U22696 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19626), .B1(
        n19946), .B2(n19959), .ZN(n19619) );
  OAI211_X1 U22697 ( .C1(n19950), .C2(n19663), .A(n19620), .B(n19619), .ZN(
        P3_U2888) );
  AOI22_X1 U22698 ( .A1(n19952), .A2(n19643), .B1(n19951), .B2(n19625), .ZN(
        n19622) );
  AOI22_X1 U22699 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19626), .B1(
        n19953), .B2(n19959), .ZN(n19621) );
  OAI211_X1 U22700 ( .C1(n19956), .C2(n19663), .A(n19622), .B(n19621), .ZN(
        P3_U2889) );
  INV_X1 U22701 ( .A(n19959), .ZN(n19974) );
  AOI22_X1 U22702 ( .A1(n19957), .A2(n19625), .B1(n19849), .B2(n19643), .ZN(
        n19624) );
  AOI22_X1 U22703 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19626), .B1(
        n19960), .B2(n19693), .ZN(n19623) );
  OAI211_X1 U22704 ( .C1(n19852), .C2(n19974), .A(n19624), .B(n19623), .ZN(
        P3_U2890) );
  AOI22_X1 U22705 ( .A1(n19967), .A2(n19959), .B1(n19966), .B2(n19625), .ZN(
        n19628) );
  AOI22_X1 U22706 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19626), .B1(
        n19970), .B2(n19643), .ZN(n19627) );
  OAI211_X1 U22707 ( .C1(n19975), .C2(n19663), .A(n19628), .B(n19627), .ZN(
        P3_U2891) );
  NAND2_X1 U22708 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19677), .ZN(
        n19719) );
  INV_X1 U22709 ( .A(n19677), .ZN(n19629) );
  NOR2_X1 U22710 ( .A1(n20050), .A2(n19629), .ZN(n19646) );
  AOI22_X1 U22711 ( .A1(n19917), .A2(n19646), .B1(n19923), .B2(n19666), .ZN(
        n19632) );
  INV_X1 U22712 ( .A(n19719), .ZN(n19710) );
  AOI21_X1 U22713 ( .B1(n20021), .B2(n19883), .A(n19651), .ZN(n19722) );
  OAI211_X1 U22714 ( .C1(n19710), .C2(n20153), .A(n19630), .B(n19722), .ZN(
        n19647) );
  AOI22_X1 U22715 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19647), .B1(
        n19918), .B2(n19643), .ZN(n19631) );
  OAI211_X1 U22716 ( .C1(n19926), .C2(n19719), .A(n19632), .B(n19631), .ZN(
        P3_U2892) );
  AOI22_X1 U22717 ( .A1(n19927), .A2(n19646), .B1(n19928), .B2(n19643), .ZN(
        n19634) );
  AOI22_X1 U22718 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19647), .B1(
        n19929), .B2(n19666), .ZN(n19633) );
  OAI211_X1 U22719 ( .C1(n19932), .C2(n19719), .A(n19634), .B(n19633), .ZN(
        P3_U2893) );
  AOI22_X1 U22720 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19647), .B1(
        n19933), .B2(n19646), .ZN(n19636) );
  AOI22_X1 U22721 ( .A1(n19935), .A2(n19666), .B1(n19934), .B2(n19643), .ZN(
        n19635) );
  OAI211_X1 U22722 ( .C1(n19938), .C2(n19719), .A(n19636), .B(n19635), .ZN(
        P3_U2894) );
  AOI22_X1 U22723 ( .A1(n19895), .A2(n19666), .B1(n19939), .B2(n19646), .ZN(
        n19638) );
  AOI22_X1 U22724 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19647), .B1(
        n19941), .B2(n19710), .ZN(n19637) );
  OAI211_X1 U22725 ( .C1(n19898), .C2(n19650), .A(n19638), .B(n19637), .ZN(
        P3_U2895) );
  AOI22_X1 U22726 ( .A1(n19946), .A2(n19643), .B1(n19945), .B2(n19646), .ZN(
        n19640) );
  AOI22_X1 U22727 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19647), .B1(
        n19947), .B2(n19666), .ZN(n19639) );
  OAI211_X1 U22728 ( .C1(n19950), .C2(n19719), .A(n19640), .B(n19639), .ZN(
        P3_U2896) );
  AOI22_X1 U22729 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19647), .B1(
        n19951), .B2(n19646), .ZN(n19642) );
  AOI22_X1 U22730 ( .A1(n19952), .A2(n19666), .B1(n19953), .B2(n19643), .ZN(
        n19641) );
  OAI211_X1 U22731 ( .C1(n19956), .C2(n19719), .A(n19642), .B(n19641), .ZN(
        P3_U2897) );
  INV_X1 U22732 ( .A(n19849), .ZN(n19964) );
  INV_X1 U22733 ( .A(n19852), .ZN(n19958) );
  AOI22_X1 U22734 ( .A1(n19958), .A2(n19643), .B1(n19957), .B2(n19646), .ZN(
        n19645) );
  AOI22_X1 U22735 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19647), .B1(
        n19960), .B2(n19710), .ZN(n19644) );
  OAI211_X1 U22736 ( .C1(n19964), .C2(n19675), .A(n19645), .B(n19644), .ZN(
        P3_U2898) );
  AOI22_X1 U22737 ( .A1(n19970), .A2(n19666), .B1(n19966), .B2(n19646), .ZN(
        n19649) );
  AOI22_X1 U22738 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19647), .B1(
        n19876), .B2(n19710), .ZN(n19648) );
  OAI211_X1 U22739 ( .C1(n19880), .C2(n19650), .A(n19649), .B(n19648), .ZN(
        P3_U2899) );
  NOR2_X2 U22740 ( .A1(n20022), .A2(n19676), .ZN(n19735) );
  NOR2_X1 U22741 ( .A1(n19710), .A2(n19735), .ZN(n19698) );
  NOR2_X1 U22742 ( .A1(n20050), .A2(n19698), .ZN(n19671) );
  AOI22_X1 U22743 ( .A1(n19917), .A2(n19671), .B1(n19923), .B2(n19693), .ZN(
        n19656) );
  OAI22_X1 U22744 ( .A1(n19653), .A2(n19652), .B1(n19698), .B2(n19651), .ZN(
        n19654) );
  OAI21_X1 U22745 ( .B1(n19735), .B2(n20153), .A(n19654), .ZN(n19672) );
  AOI22_X1 U22746 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19672), .B1(
        n19887), .B2(n19735), .ZN(n19655) );
  OAI211_X1 U22747 ( .C1(n19890), .C2(n19675), .A(n19656), .B(n19655), .ZN(
        P3_U2900) );
  INV_X1 U22748 ( .A(n19735), .ZN(n19742) );
  AOI22_X1 U22749 ( .A1(n19927), .A2(n19671), .B1(n19928), .B2(n19666), .ZN(
        n19658) );
  AOI22_X1 U22750 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19672), .B1(
        n19929), .B2(n19693), .ZN(n19657) );
  OAI211_X1 U22751 ( .C1(n19932), .C2(n19742), .A(n19658), .B(n19657), .ZN(
        P3_U2901) );
  AOI22_X1 U22752 ( .A1(n19935), .A2(n19693), .B1(n19933), .B2(n19671), .ZN(
        n19660) );
  AOI22_X1 U22753 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19672), .B1(
        n19934), .B2(n19666), .ZN(n19659) );
  OAI211_X1 U22754 ( .C1(n19938), .C2(n19742), .A(n19660), .B(n19659), .ZN(
        P3_U2902) );
  AOI22_X1 U22755 ( .A1(n19940), .A2(n19666), .B1(n19939), .B2(n19671), .ZN(
        n19662) );
  AOI22_X1 U22756 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19672), .B1(
        n19941), .B2(n19735), .ZN(n19661) );
  OAI211_X1 U22757 ( .C1(n19944), .C2(n19663), .A(n19662), .B(n19661), .ZN(
        P3_U2903) );
  AOI22_X1 U22758 ( .A1(n19946), .A2(n19666), .B1(n19945), .B2(n19671), .ZN(
        n19665) );
  AOI22_X1 U22759 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19672), .B1(
        n19947), .B2(n19693), .ZN(n19664) );
  OAI211_X1 U22760 ( .C1(n19950), .C2(n19742), .A(n19665), .B(n19664), .ZN(
        P3_U2904) );
  AOI22_X1 U22761 ( .A1(n19952), .A2(n19693), .B1(n19951), .B2(n19671), .ZN(
        n19668) );
  AOI22_X1 U22762 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19672), .B1(
        n19953), .B2(n19666), .ZN(n19667) );
  OAI211_X1 U22763 ( .C1(n19956), .C2(n19742), .A(n19668), .B(n19667), .ZN(
        P3_U2905) );
  AOI22_X1 U22764 ( .A1(n19957), .A2(n19671), .B1(n19849), .B2(n19693), .ZN(
        n19670) );
  AOI22_X1 U22765 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19672), .B1(
        n19960), .B2(n19735), .ZN(n19669) );
  OAI211_X1 U22766 ( .C1(n19852), .C2(n19675), .A(n19670), .B(n19669), .ZN(
        P3_U2906) );
  AOI22_X1 U22767 ( .A1(n19970), .A2(n19693), .B1(n19966), .B2(n19671), .ZN(
        n19674) );
  AOI22_X1 U22768 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19672), .B1(
        n19876), .B2(n19735), .ZN(n19673) );
  OAI211_X1 U22769 ( .C1(n19880), .C2(n19675), .A(n19674), .B(n19673), .ZN(
        P3_U2907) );
  NAND2_X1 U22770 ( .A1(n19766), .A2(n19721), .ZN(n19754) );
  AOI22_X1 U22771 ( .A1(n19918), .A2(n19693), .B1(n19917), .B2(n19692), .ZN(
        n19679) );
  AOI22_X1 U22772 ( .A1(n19922), .A2(n19677), .B1(n19768), .B2(n19721), .ZN(
        n19694) );
  AOI22_X1 U22773 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19694), .B1(
        n19923), .B2(n19710), .ZN(n19678) );
  OAI211_X1 U22774 ( .C1(n19926), .C2(n19754), .A(n19679), .B(n19678), .ZN(
        P3_U2908) );
  AOI22_X1 U22775 ( .A1(n19927), .A2(n19692), .B1(n19928), .B2(n19693), .ZN(
        n19681) );
  AOI22_X1 U22776 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19694), .B1(
        n19929), .B2(n19710), .ZN(n19680) );
  OAI211_X1 U22777 ( .C1(n19932), .C2(n19754), .A(n19681), .B(n19680), .ZN(
        P3_U2909) );
  AOI22_X1 U22778 ( .A1(n19935), .A2(n19710), .B1(n19933), .B2(n19692), .ZN(
        n19683) );
  AOI22_X1 U22779 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19694), .B1(
        n19934), .B2(n19693), .ZN(n19682) );
  OAI211_X1 U22780 ( .C1(n19938), .C2(n19754), .A(n19683), .B(n19682), .ZN(
        P3_U2910) );
  AOI22_X1 U22781 ( .A1(n19940), .A2(n19693), .B1(n19939), .B2(n19692), .ZN(
        n19685) );
  INV_X1 U22782 ( .A(n19754), .ZN(n19762) );
  AOI22_X1 U22783 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19694), .B1(
        n19941), .B2(n19762), .ZN(n19684) );
  OAI211_X1 U22784 ( .C1(n19944), .C2(n19719), .A(n19685), .B(n19684), .ZN(
        P3_U2911) );
  AOI22_X1 U22785 ( .A1(n19946), .A2(n19693), .B1(n19945), .B2(n19692), .ZN(
        n19687) );
  AOI22_X1 U22786 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19694), .B1(
        n19947), .B2(n19710), .ZN(n19686) );
  OAI211_X1 U22787 ( .C1(n19950), .C2(n19754), .A(n19687), .B(n19686), .ZN(
        P3_U2912) );
  AOI22_X1 U22788 ( .A1(n19953), .A2(n19693), .B1(n19951), .B2(n19692), .ZN(
        n19689) );
  AOI22_X1 U22789 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19694), .B1(
        n19952), .B2(n19710), .ZN(n19688) );
  OAI211_X1 U22790 ( .C1(n19956), .C2(n19754), .A(n19689), .B(n19688), .ZN(
        P3_U2913) );
  AOI22_X1 U22791 ( .A1(n19958), .A2(n19693), .B1(n19957), .B2(n19692), .ZN(
        n19691) );
  AOI22_X1 U22792 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19694), .B1(
        n19960), .B2(n19762), .ZN(n19690) );
  OAI211_X1 U22793 ( .C1(n19964), .C2(n19719), .A(n19691), .B(n19690), .ZN(
        P3_U2914) );
  AOI22_X1 U22794 ( .A1(n19967), .A2(n19693), .B1(n19966), .B2(n19692), .ZN(
        n19696) );
  AOI22_X1 U22795 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19694), .B1(
        n19970), .B2(n19710), .ZN(n19695) );
  OAI211_X1 U22796 ( .C1(n19975), .C2(n19754), .A(n19696), .B(n19695), .ZN(
        P3_U2915) );
  NOR2_X1 U22797 ( .A1(n19697), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19769) );
  INV_X1 U22798 ( .A(n19769), .ZN(n19720) );
  NOR2_X2 U22799 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19720), .ZN(
        n19780) );
  NOR2_X1 U22800 ( .A1(n19762), .A2(n19780), .ZN(n19744) );
  NOR2_X1 U22801 ( .A1(n20050), .A2(n19744), .ZN(n19715) );
  AOI22_X1 U22802 ( .A1(n19917), .A2(n19715), .B1(n19923), .B2(n19735), .ZN(
        n19701) );
  OAI21_X1 U22803 ( .B1(n19698), .B2(n19883), .A(n19744), .ZN(n19699) );
  OAI211_X1 U22804 ( .C1(n19780), .C2(n20153), .A(n19886), .B(n19699), .ZN(
        n19716) );
  AOI22_X1 U22805 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19716), .B1(
        n19887), .B2(n19780), .ZN(n19700) );
  OAI211_X1 U22806 ( .C1(n19890), .C2(n19719), .A(n19701), .B(n19700), .ZN(
        P3_U2916) );
  INV_X1 U22807 ( .A(n19780), .ZN(n19789) );
  AOI22_X1 U22808 ( .A1(n19929), .A2(n19735), .B1(n19927), .B2(n19715), .ZN(
        n19703) );
  AOI22_X1 U22809 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19716), .B1(
        n19928), .B2(n19710), .ZN(n19702) );
  OAI211_X1 U22810 ( .C1(n19932), .C2(n19789), .A(n19703), .B(n19702), .ZN(
        P3_U2917) );
  AOI22_X1 U22811 ( .A1(n19935), .A2(n19735), .B1(n19933), .B2(n19715), .ZN(
        n19705) );
  AOI22_X1 U22812 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19716), .B1(
        n19934), .B2(n19710), .ZN(n19704) );
  OAI211_X1 U22813 ( .C1(n19938), .C2(n19789), .A(n19705), .B(n19704), .ZN(
        P3_U2918) );
  AOI22_X1 U22814 ( .A1(n19895), .A2(n19735), .B1(n19939), .B2(n19715), .ZN(
        n19707) );
  AOI22_X1 U22815 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19716), .B1(
        n19941), .B2(n19780), .ZN(n19706) );
  OAI211_X1 U22816 ( .C1(n19898), .C2(n19719), .A(n19707), .B(n19706), .ZN(
        P3_U2919) );
  AOI22_X1 U22817 ( .A1(n19946), .A2(n19710), .B1(n19945), .B2(n19715), .ZN(
        n19709) );
  AOI22_X1 U22818 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19716), .B1(
        n19947), .B2(n19735), .ZN(n19708) );
  OAI211_X1 U22819 ( .C1(n19950), .C2(n19789), .A(n19709), .B(n19708), .ZN(
        P3_U2920) );
  AOI22_X1 U22820 ( .A1(n19952), .A2(n19735), .B1(n19951), .B2(n19715), .ZN(
        n19712) );
  AOI22_X1 U22821 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19716), .B1(
        n19953), .B2(n19710), .ZN(n19711) );
  OAI211_X1 U22822 ( .C1(n19956), .C2(n19789), .A(n19712), .B(n19711), .ZN(
        P3_U2921) );
  AOI22_X1 U22823 ( .A1(n19957), .A2(n19715), .B1(n19849), .B2(n19735), .ZN(
        n19714) );
  AOI22_X1 U22824 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19716), .B1(
        n19960), .B2(n19780), .ZN(n19713) );
  OAI211_X1 U22825 ( .C1(n19852), .C2(n19719), .A(n19714), .B(n19713), .ZN(
        P3_U2922) );
  AOI22_X1 U22826 ( .A1(n19970), .A2(n19735), .B1(n19966), .B2(n19715), .ZN(
        n19718) );
  AOI22_X1 U22827 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19716), .B1(
        n19876), .B2(n19780), .ZN(n19717) );
  OAI211_X1 U22828 ( .C1(n19880), .C2(n19719), .A(n19718), .B(n19717), .ZN(
        P3_U2923) );
  NOR2_X1 U22829 ( .A1(n20050), .A2(n19720), .ZN(n19738) );
  AOI22_X1 U22830 ( .A1(n19917), .A2(n19738), .B1(n19923), .B2(n19762), .ZN(
        n19724) );
  NOR2_X2 U22831 ( .A1(n20019), .A2(n19720), .ZN(n19804) );
  OAI211_X1 U22832 ( .C1(n19804), .C2(n20153), .A(n19722), .B(n19721), .ZN(
        n19739) );
  AOI22_X1 U22833 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19739), .B1(
        n19887), .B2(n19804), .ZN(n19723) );
  OAI211_X1 U22834 ( .C1(n19890), .C2(n19742), .A(n19724), .B(n19723), .ZN(
        P3_U2924) );
  INV_X1 U22835 ( .A(n19804), .ZN(n19811) );
  AOI22_X1 U22836 ( .A1(n19927), .A2(n19738), .B1(n19928), .B2(n19735), .ZN(
        n19726) );
  AOI22_X1 U22837 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19739), .B1(
        n19929), .B2(n19762), .ZN(n19725) );
  OAI211_X1 U22838 ( .C1(n19932), .C2(n19811), .A(n19726), .B(n19725), .ZN(
        P3_U2925) );
  AOI22_X1 U22839 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19739), .B1(
        n19933), .B2(n19738), .ZN(n19728) );
  AOI22_X1 U22840 ( .A1(n19935), .A2(n19762), .B1(n19934), .B2(n19735), .ZN(
        n19727) );
  OAI211_X1 U22841 ( .C1(n19938), .C2(n19811), .A(n19728), .B(n19727), .ZN(
        P3_U2926) );
  AOI22_X1 U22842 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19739), .B1(
        n19939), .B2(n19738), .ZN(n19730) );
  AOI22_X1 U22843 ( .A1(n19941), .A2(n19804), .B1(n19895), .B2(n19762), .ZN(
        n19729) );
  OAI211_X1 U22844 ( .C1(n19898), .C2(n19742), .A(n19730), .B(n19729), .ZN(
        P3_U2927) );
  AOI22_X1 U22845 ( .A1(n19945), .A2(n19738), .B1(n19947), .B2(n19762), .ZN(
        n19732) );
  AOI22_X1 U22846 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19739), .B1(
        n19899), .B2(n19804), .ZN(n19731) );
  OAI211_X1 U22847 ( .C1(n19902), .C2(n19742), .A(n19732), .B(n19731), .ZN(
        P3_U2928) );
  AOI22_X1 U22848 ( .A1(n19953), .A2(n19735), .B1(n19951), .B2(n19738), .ZN(
        n19734) );
  AOI22_X1 U22849 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19739), .B1(
        n19952), .B2(n19762), .ZN(n19733) );
  OAI211_X1 U22850 ( .C1(n19956), .C2(n19811), .A(n19734), .B(n19733), .ZN(
        P3_U2929) );
  AOI22_X1 U22851 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19739), .B1(
        n19957), .B2(n19738), .ZN(n19737) );
  AOI22_X1 U22852 ( .A1(n19958), .A2(n19735), .B1(n19960), .B2(n19804), .ZN(
        n19736) );
  OAI211_X1 U22853 ( .C1(n19964), .C2(n19754), .A(n19737), .B(n19736), .ZN(
        P3_U2930) );
  AOI22_X1 U22854 ( .A1(n19970), .A2(n19762), .B1(n19966), .B2(n19738), .ZN(
        n19741) );
  AOI22_X1 U22855 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19739), .B1(
        n19876), .B2(n19804), .ZN(n19740) );
  OAI211_X1 U22856 ( .C1(n19880), .C2(n19742), .A(n19741), .B(n19740), .ZN(
        P3_U2931) );
  INV_X1 U22857 ( .A(n19813), .ZN(n19767) );
  NOR2_X2 U22858 ( .A1(n20022), .A2(n19767), .ZN(n19830) );
  NOR2_X1 U22859 ( .A1(n19804), .A2(n19830), .ZN(n19790) );
  NOR2_X1 U22860 ( .A1(n20050), .A2(n19790), .ZN(n19761) );
  AOI22_X1 U22861 ( .A1(n19917), .A2(n19761), .B1(n19923), .B2(n19780), .ZN(
        n19747) );
  AOI221_X1 U22862 ( .B1(n19790), .B2(n19883), .C1(n19790), .C2(n19744), .A(
        n19743), .ZN(n19745) );
  INV_X1 U22863 ( .A(n19745), .ZN(n19763) );
  AOI22_X1 U22864 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19763), .B1(
        n19887), .B2(n19830), .ZN(n19746) );
  OAI211_X1 U22865 ( .C1(n19890), .C2(n19754), .A(n19747), .B(n19746), .ZN(
        P3_U2932) );
  INV_X1 U22866 ( .A(n19830), .ZN(n19828) );
  AOI22_X1 U22867 ( .A1(n19929), .A2(n19780), .B1(n19927), .B2(n19761), .ZN(
        n19749) );
  AOI22_X1 U22868 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19763), .B1(
        n19928), .B2(n19762), .ZN(n19748) );
  OAI211_X1 U22869 ( .C1(n19932), .C2(n19828), .A(n19749), .B(n19748), .ZN(
        P3_U2933) );
  AOI22_X1 U22870 ( .A1(n19935), .A2(n19780), .B1(n19933), .B2(n19761), .ZN(
        n19751) );
  AOI22_X1 U22871 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19763), .B1(
        n19934), .B2(n19762), .ZN(n19750) );
  OAI211_X1 U22872 ( .C1(n19938), .C2(n19828), .A(n19751), .B(n19750), .ZN(
        P3_U2934) );
  AOI22_X1 U22873 ( .A1(n19895), .A2(n19780), .B1(n19939), .B2(n19761), .ZN(
        n19753) );
  AOI22_X1 U22874 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19763), .B1(
        n19941), .B2(n19830), .ZN(n19752) );
  OAI211_X1 U22875 ( .C1(n19898), .C2(n19754), .A(n19753), .B(n19752), .ZN(
        P3_U2935) );
  AOI22_X1 U22876 ( .A1(n19946), .A2(n19762), .B1(n19945), .B2(n19761), .ZN(
        n19756) );
  AOI22_X1 U22877 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19763), .B1(
        n19947), .B2(n19780), .ZN(n19755) );
  OAI211_X1 U22878 ( .C1(n19950), .C2(n19828), .A(n19756), .B(n19755), .ZN(
        P3_U2936) );
  AOI22_X1 U22879 ( .A1(n19953), .A2(n19762), .B1(n19951), .B2(n19761), .ZN(
        n19758) );
  AOI22_X1 U22880 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19763), .B1(
        n19952), .B2(n19780), .ZN(n19757) );
  OAI211_X1 U22881 ( .C1(n19956), .C2(n19828), .A(n19758), .B(n19757), .ZN(
        P3_U2937) );
  AOI22_X1 U22882 ( .A1(n19958), .A2(n19762), .B1(n19957), .B2(n19761), .ZN(
        n19760) );
  AOI22_X1 U22883 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19763), .B1(
        n19960), .B2(n19830), .ZN(n19759) );
  OAI211_X1 U22884 ( .C1(n19964), .C2(n19789), .A(n19760), .B(n19759), .ZN(
        P3_U2938) );
  AOI22_X1 U22885 ( .A1(n19967), .A2(n19762), .B1(n19966), .B2(n19761), .ZN(
        n19765) );
  AOI22_X1 U22886 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19763), .B1(
        n19970), .B2(n19780), .ZN(n19764) );
  OAI211_X1 U22887 ( .C1(n19975), .C2(n19828), .A(n19765), .B(n19764), .ZN(
        P3_U2939) );
  NAND2_X1 U22888 ( .A1(n19813), .A2(n19766), .ZN(n19857) );
  AOI22_X1 U22889 ( .A1(n19918), .A2(n19780), .B1(n19917), .B2(n19785), .ZN(
        n19771) );
  AOI22_X1 U22890 ( .A1(n19922), .A2(n19769), .B1(n19813), .B2(n19768), .ZN(
        n19786) );
  AOI22_X1 U22891 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19786), .B1(
        n19923), .B2(n19804), .ZN(n19770) );
  OAI211_X1 U22892 ( .C1(n19857), .C2(n19926), .A(n19771), .B(n19770), .ZN(
        P3_U2940) );
  AOI22_X1 U22893 ( .A1(n19927), .A2(n19785), .B1(n19928), .B2(n19780), .ZN(
        n19773) );
  AOI22_X1 U22894 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19786), .B1(
        n19929), .B2(n19804), .ZN(n19772) );
  OAI211_X1 U22895 ( .C1(n19857), .C2(n19932), .A(n19773), .B(n19772), .ZN(
        P3_U2941) );
  AOI22_X1 U22896 ( .A1(n19935), .A2(n19804), .B1(n19933), .B2(n19785), .ZN(
        n19775) );
  AOI22_X1 U22897 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19786), .B1(
        n19934), .B2(n19780), .ZN(n19774) );
  OAI211_X1 U22898 ( .C1(n19857), .C2(n19938), .A(n19775), .B(n19774), .ZN(
        P3_U2942) );
  AOI22_X1 U22899 ( .A1(n19940), .A2(n19780), .B1(n19939), .B2(n19785), .ZN(
        n19777) );
  INV_X1 U22900 ( .A(n19857), .ZN(n19846) );
  AOI22_X1 U22901 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19786), .B1(
        n19846), .B2(n19941), .ZN(n19776) );
  OAI211_X1 U22902 ( .C1(n19944), .C2(n19811), .A(n19777), .B(n19776), .ZN(
        P3_U2943) );
  AOI22_X1 U22903 ( .A1(n19946), .A2(n19780), .B1(n19945), .B2(n19785), .ZN(
        n19779) );
  AOI22_X1 U22904 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19786), .B1(
        n19947), .B2(n19804), .ZN(n19778) );
  OAI211_X1 U22905 ( .C1(n19857), .C2(n19950), .A(n19779), .B(n19778), .ZN(
        P3_U2944) );
  AOI22_X1 U22906 ( .A1(n19952), .A2(n19804), .B1(n19951), .B2(n19785), .ZN(
        n19782) );
  AOI22_X1 U22907 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19786), .B1(
        n19953), .B2(n19780), .ZN(n19781) );
  OAI211_X1 U22908 ( .C1(n19857), .C2(n19956), .A(n19782), .B(n19781), .ZN(
        P3_U2945) );
  AOI22_X1 U22909 ( .A1(n19957), .A2(n19785), .B1(n19849), .B2(n19804), .ZN(
        n19784) );
  AOI22_X1 U22910 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19786), .B1(
        n19846), .B2(n19960), .ZN(n19783) );
  OAI211_X1 U22911 ( .C1(n19852), .C2(n19789), .A(n19784), .B(n19783), .ZN(
        P3_U2946) );
  AOI22_X1 U22912 ( .A1(n19970), .A2(n19804), .B1(n19966), .B2(n19785), .ZN(
        n19788) );
  AOI22_X1 U22913 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19786), .B1(
        n19846), .B2(n19876), .ZN(n19787) );
  OAI211_X1 U22914 ( .C1(n19880), .C2(n19789), .A(n19788), .B(n19787), .ZN(
        P3_U2947) );
  NAND2_X1 U22915 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19813), .ZN(
        n19812) );
  NOR2_X2 U22916 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19812), .ZN(
        n19872) );
  INV_X1 U22917 ( .A(n19872), .ZN(n19881) );
  NOR2_X1 U22918 ( .A1(n19846), .A2(n19872), .ZN(n19834) );
  NOR2_X1 U22919 ( .A1(n20050), .A2(n19834), .ZN(n19807) );
  AOI22_X1 U22920 ( .A1(n19918), .A2(n19804), .B1(n19917), .B2(n19807), .ZN(
        n19793) );
  OAI21_X1 U22921 ( .B1(n19790), .B2(n19883), .A(n19834), .ZN(n19791) );
  OAI211_X1 U22922 ( .C1(n19872), .C2(n20153), .A(n19886), .B(n19791), .ZN(
        n19808) );
  AOI22_X1 U22923 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19808), .B1(
        n19923), .B2(n19830), .ZN(n19792) );
  OAI211_X1 U22924 ( .C1(n19881), .C2(n19926), .A(n19793), .B(n19792), .ZN(
        P3_U2948) );
  AOI22_X1 U22925 ( .A1(n19929), .A2(n19830), .B1(n19927), .B2(n19807), .ZN(
        n19795) );
  AOI22_X1 U22926 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19808), .B1(
        n19928), .B2(n19804), .ZN(n19794) );
  OAI211_X1 U22927 ( .C1(n19881), .C2(n19932), .A(n19795), .B(n19794), .ZN(
        P3_U2949) );
  AOI22_X1 U22928 ( .A1(n19933), .A2(n19807), .B1(n19934), .B2(n19804), .ZN(
        n19797) );
  AOI22_X1 U22929 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19808), .B1(
        n19935), .B2(n19830), .ZN(n19796) );
  OAI211_X1 U22930 ( .C1(n19881), .C2(n19938), .A(n19797), .B(n19796), .ZN(
        P3_U2950) );
  AOI22_X1 U22931 ( .A1(n19895), .A2(n19830), .B1(n19939), .B2(n19807), .ZN(
        n19799) );
  AOI22_X1 U22932 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19808), .B1(
        n19872), .B2(n19941), .ZN(n19798) );
  OAI211_X1 U22933 ( .C1(n19898), .C2(n19811), .A(n19799), .B(n19798), .ZN(
        P3_U2951) );
  AOI22_X1 U22934 ( .A1(n19946), .A2(n19804), .B1(n19945), .B2(n19807), .ZN(
        n19801) );
  AOI22_X1 U22935 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19808), .B1(
        n19947), .B2(n19830), .ZN(n19800) );
  OAI211_X1 U22936 ( .C1(n19881), .C2(n19950), .A(n19801), .B(n19800), .ZN(
        P3_U2952) );
  AOI22_X1 U22937 ( .A1(n19953), .A2(n19804), .B1(n19951), .B2(n19807), .ZN(
        n19803) );
  AOI22_X1 U22938 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19808), .B1(
        n19952), .B2(n19830), .ZN(n19802) );
  OAI211_X1 U22939 ( .C1(n19881), .C2(n19956), .A(n19803), .B(n19802), .ZN(
        P3_U2953) );
  AOI22_X1 U22940 ( .A1(n19958), .A2(n19804), .B1(n19957), .B2(n19807), .ZN(
        n19806) );
  AOI22_X1 U22941 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19808), .B1(
        n19872), .B2(n19960), .ZN(n19805) );
  OAI211_X1 U22942 ( .C1(n19964), .C2(n19828), .A(n19806), .B(n19805), .ZN(
        P3_U2954) );
  AOI22_X1 U22943 ( .A1(n19970), .A2(n19830), .B1(n19966), .B2(n19807), .ZN(
        n19810) );
  AOI22_X1 U22944 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19808), .B1(
        n19872), .B2(n19876), .ZN(n19809) );
  OAI211_X1 U22945 ( .C1(n19880), .C2(n19811), .A(n19810), .B(n19809), .ZN(
        P3_U2955) );
  INV_X1 U22946 ( .A(n19812), .ZN(n19859) );
  NAND2_X1 U22947 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19859), .ZN(
        n19903) );
  NOR2_X1 U22948 ( .A1(n20050), .A2(n19812), .ZN(n19829) );
  AOI22_X1 U22949 ( .A1(n19846), .A2(n19923), .B1(n19917), .B2(n19829), .ZN(
        n19815) );
  AOI22_X1 U22950 ( .A1(n19922), .A2(n19813), .B1(n19859), .B2(n19919), .ZN(
        n19831) );
  AOI22_X1 U22951 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19831), .B1(
        n19918), .B2(n19830), .ZN(n19814) );
  OAI211_X1 U22952 ( .C1(n19903), .C2(n19926), .A(n19815), .B(n19814), .ZN(
        P3_U2956) );
  AOI22_X1 U22953 ( .A1(n19927), .A2(n19829), .B1(n19928), .B2(n19830), .ZN(
        n19817) );
  AOI22_X1 U22954 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19831), .B1(
        n19846), .B2(n19929), .ZN(n19816) );
  OAI211_X1 U22955 ( .C1(n19903), .C2(n19932), .A(n19817), .B(n19816), .ZN(
        P3_U2957) );
  AOI22_X1 U22956 ( .A1(n19846), .A2(n19935), .B1(n19933), .B2(n19829), .ZN(
        n19819) );
  AOI22_X1 U22957 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19831), .B1(
        n19934), .B2(n19830), .ZN(n19818) );
  OAI211_X1 U22958 ( .C1(n19903), .C2(n19938), .A(n19819), .B(n19818), .ZN(
        P3_U2958) );
  AOI22_X1 U22959 ( .A1(n19846), .A2(n19895), .B1(n19939), .B2(n19829), .ZN(
        n19821) );
  INV_X1 U22960 ( .A(n19903), .ZN(n19911) );
  AOI22_X1 U22961 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19831), .B1(
        n19911), .B2(n19941), .ZN(n19820) );
  OAI211_X1 U22962 ( .C1(n19898), .C2(n19828), .A(n19821), .B(n19820), .ZN(
        P3_U2959) );
  AOI22_X1 U22963 ( .A1(n19846), .A2(n19947), .B1(n19945), .B2(n19829), .ZN(
        n19823) );
  AOI22_X1 U22964 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19831), .B1(
        n19911), .B2(n19899), .ZN(n19822) );
  OAI211_X1 U22965 ( .C1(n19902), .C2(n19828), .A(n19823), .B(n19822), .ZN(
        P3_U2960) );
  AOI22_X1 U22966 ( .A1(n19953), .A2(n19830), .B1(n19951), .B2(n19829), .ZN(
        n19825) );
  AOI22_X1 U22967 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19831), .B1(
        n19846), .B2(n19952), .ZN(n19824) );
  OAI211_X1 U22968 ( .C1(n19903), .C2(n19956), .A(n19825), .B(n19824), .ZN(
        P3_U2961) );
  AOI22_X1 U22969 ( .A1(n19846), .A2(n19849), .B1(n19957), .B2(n19829), .ZN(
        n19827) );
  AOI22_X1 U22970 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19831), .B1(
        n19911), .B2(n19960), .ZN(n19826) );
  OAI211_X1 U22971 ( .C1(n19852), .C2(n19828), .A(n19827), .B(n19826), .ZN(
        P3_U2962) );
  AOI22_X1 U22972 ( .A1(n19967), .A2(n19830), .B1(n19966), .B2(n19829), .ZN(
        n19833) );
  AOI22_X1 U22973 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19831), .B1(
        n19846), .B2(n19970), .ZN(n19832) );
  OAI211_X1 U22974 ( .C1(n19903), .C2(n19975), .A(n19833), .B(n19832), .ZN(
        P3_U2963) );
  NAND2_X1 U22975 ( .A1(n19921), .A2(n20019), .ZN(n19909) );
  AOI21_X1 U22976 ( .B1(n19909), .B2(n19903), .A(n20050), .ZN(n19853) );
  AOI22_X1 U22977 ( .A1(n19872), .A2(n19923), .B1(n19917), .B2(n19853), .ZN(
        n19837) );
  AOI221_X1 U22978 ( .B1(n19834), .B2(n19903), .C1(n19883), .C2(n19903), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19835) );
  OAI21_X1 U22979 ( .B1(n19968), .B2(n19835), .A(n19886), .ZN(n19854) );
  AOI22_X1 U22980 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19854), .B1(
        n19968), .B2(n19887), .ZN(n19836) );
  OAI211_X1 U22981 ( .C1(n19890), .C2(n19857), .A(n19837), .B(n19836), .ZN(
        P3_U2964) );
  AOI22_X1 U22982 ( .A1(n19846), .A2(n19928), .B1(n19853), .B2(n19927), .ZN(
        n19839) );
  AOI22_X1 U22983 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19854), .B1(
        n19872), .B2(n19929), .ZN(n19838) );
  OAI211_X1 U22984 ( .C1(n19909), .C2(n19932), .A(n19839), .B(n19838), .ZN(
        P3_U2965) );
  AOI22_X1 U22985 ( .A1(n19846), .A2(n19934), .B1(n19853), .B2(n19933), .ZN(
        n19841) );
  AOI22_X1 U22986 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19854), .B1(
        n19872), .B2(n19935), .ZN(n19840) );
  OAI211_X1 U22987 ( .C1(n19909), .C2(n19938), .A(n19841), .B(n19840), .ZN(
        P3_U2966) );
  AOI22_X1 U22988 ( .A1(n19872), .A2(n19895), .B1(n19853), .B2(n19939), .ZN(
        n19843) );
  AOI22_X1 U22989 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19854), .B1(
        n19968), .B2(n19941), .ZN(n19842) );
  OAI211_X1 U22990 ( .C1(n19857), .C2(n19898), .A(n19843), .B(n19842), .ZN(
        P3_U2967) );
  AOI22_X1 U22991 ( .A1(n19872), .A2(n19947), .B1(n19853), .B2(n19945), .ZN(
        n19845) );
  AOI22_X1 U22992 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19854), .B1(
        n19968), .B2(n19899), .ZN(n19844) );
  OAI211_X1 U22993 ( .C1(n19857), .C2(n19902), .A(n19845), .B(n19844), .ZN(
        P3_U2968) );
  AOI22_X1 U22994 ( .A1(n19846), .A2(n19953), .B1(n19853), .B2(n19951), .ZN(
        n19848) );
  AOI22_X1 U22995 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19854), .B1(
        n19872), .B2(n19952), .ZN(n19847) );
  OAI211_X1 U22996 ( .C1(n19909), .C2(n19956), .A(n19848), .B(n19847), .ZN(
        P3_U2969) );
  AOI22_X1 U22997 ( .A1(n19872), .A2(n19849), .B1(n19853), .B2(n19957), .ZN(
        n19851) );
  AOI22_X1 U22998 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19854), .B1(
        n19968), .B2(n19960), .ZN(n19850) );
  OAI211_X1 U22999 ( .C1(n19857), .C2(n19852), .A(n19851), .B(n19850), .ZN(
        P3_U2970) );
  AOI22_X1 U23000 ( .A1(n19872), .A2(n19970), .B1(n19853), .B2(n19966), .ZN(
        n19856) );
  AOI22_X1 U23001 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19854), .B1(
        n19968), .B2(n19876), .ZN(n19855) );
  OAI211_X1 U23002 ( .C1(n19857), .C2(n19880), .A(n19856), .B(n19855), .ZN(
        P3_U2971) );
  INV_X1 U23003 ( .A(n19921), .ZN(n19858) );
  NOR2_X1 U23004 ( .A1(n20050), .A2(n19858), .ZN(n19875) );
  AOI22_X1 U23005 ( .A1(n19911), .A2(n19923), .B1(n19917), .B2(n19875), .ZN(
        n19861) );
  AOI22_X1 U23006 ( .A1(n19922), .A2(n19859), .B1(n19921), .B2(n19919), .ZN(
        n19877) );
  AOI22_X1 U23007 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19877), .B1(
        n19887), .B2(n19969), .ZN(n19860) );
  OAI211_X1 U23008 ( .C1(n19890), .C2(n19881), .A(n19861), .B(n19860), .ZN(
        P3_U2972) );
  AOI22_X1 U23009 ( .A1(n19911), .A2(n19929), .B1(n19927), .B2(n19875), .ZN(
        n19863) );
  AOI22_X1 U23010 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19877), .B1(
        n19872), .B2(n19928), .ZN(n19862) );
  OAI211_X1 U23011 ( .C1(n19932), .C2(n19963), .A(n19863), .B(n19862), .ZN(
        P3_U2973) );
  AOI22_X1 U23012 ( .A1(n19911), .A2(n19935), .B1(n19933), .B2(n19875), .ZN(
        n19865) );
  AOI22_X1 U23013 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19877), .B1(
        n19872), .B2(n19934), .ZN(n19864) );
  OAI211_X1 U23014 ( .C1(n19938), .C2(n19963), .A(n19865), .B(n19864), .ZN(
        P3_U2974) );
  AOI22_X1 U23015 ( .A1(n19872), .A2(n19940), .B1(n19939), .B2(n19875), .ZN(
        n19867) );
  AOI22_X1 U23016 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19877), .B1(
        n19941), .B2(n19969), .ZN(n19866) );
  OAI211_X1 U23017 ( .C1(n19903), .C2(n19944), .A(n19867), .B(n19866), .ZN(
        P3_U2975) );
  AOI22_X1 U23018 ( .A1(n19872), .A2(n19946), .B1(n19945), .B2(n19875), .ZN(
        n19869) );
  AOI22_X1 U23019 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19877), .B1(
        n19911), .B2(n19947), .ZN(n19868) );
  OAI211_X1 U23020 ( .C1(n19950), .C2(n19963), .A(n19869), .B(n19868), .ZN(
        P3_U2976) );
  AOI22_X1 U23021 ( .A1(n19911), .A2(n19952), .B1(n19951), .B2(n19875), .ZN(
        n19871) );
  AOI22_X1 U23022 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19877), .B1(
        n19872), .B2(n19953), .ZN(n19870) );
  OAI211_X1 U23023 ( .C1(n19956), .C2(n19963), .A(n19871), .B(n19870), .ZN(
        P3_U2977) );
  AOI22_X1 U23024 ( .A1(n19872), .A2(n19958), .B1(n19957), .B2(n19875), .ZN(
        n19874) );
  AOI22_X1 U23025 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19877), .B1(
        n19960), .B2(n19969), .ZN(n19873) );
  OAI211_X1 U23026 ( .C1(n19903), .C2(n19964), .A(n19874), .B(n19873), .ZN(
        P3_U2978) );
  AOI22_X1 U23027 ( .A1(n19911), .A2(n19970), .B1(n19966), .B2(n19875), .ZN(
        n19879) );
  AOI22_X1 U23028 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19877), .B1(
        n19876), .B2(n19969), .ZN(n19878) );
  OAI211_X1 U23029 ( .C1(n19881), .C2(n19880), .A(n19879), .B(n19878), .ZN(
        P3_U2979) );
  NOR2_X1 U23030 ( .A1(n20050), .A2(n19882), .ZN(n19910) );
  AOI22_X1 U23031 ( .A1(n19968), .A2(n19923), .B1(n19917), .B2(n19910), .ZN(
        n19889) );
  NOR2_X1 U23032 ( .A1(n19968), .A2(n19911), .ZN(n19884) );
  OAI21_X1 U23033 ( .B1(n19884), .B2(n19883), .A(n19882), .ZN(n19885) );
  OAI211_X1 U23034 ( .C1(n19906), .C2(n20153), .A(n19886), .B(n19885), .ZN(
        n19912) );
  AOI22_X1 U23035 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19912), .B1(
        n19887), .B2(n19906), .ZN(n19888) );
  OAI211_X1 U23036 ( .C1(n19890), .C2(n19903), .A(n19889), .B(n19888), .ZN(
        P3_U2980) );
  AOI22_X1 U23037 ( .A1(n19911), .A2(n19928), .B1(n19927), .B2(n19910), .ZN(
        n19892) );
  AOI22_X1 U23038 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19912), .B1(
        n19968), .B2(n19929), .ZN(n19891) );
  OAI211_X1 U23039 ( .C1(n19932), .C2(n19915), .A(n19892), .B(n19891), .ZN(
        P3_U2981) );
  AOI22_X1 U23040 ( .A1(n19968), .A2(n19935), .B1(n19933), .B2(n19910), .ZN(
        n19894) );
  AOI22_X1 U23041 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19912), .B1(
        n19911), .B2(n19934), .ZN(n19893) );
  OAI211_X1 U23042 ( .C1(n19938), .C2(n19915), .A(n19894), .B(n19893), .ZN(
        P3_U2982) );
  AOI22_X1 U23043 ( .A1(n19968), .A2(n19895), .B1(n19939), .B2(n19910), .ZN(
        n19897) );
  AOI22_X1 U23044 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19912), .B1(
        n19941), .B2(n19906), .ZN(n19896) );
  OAI211_X1 U23045 ( .C1(n19903), .C2(n19898), .A(n19897), .B(n19896), .ZN(
        P3_U2983) );
  AOI22_X1 U23046 ( .A1(n19968), .A2(n19947), .B1(n19945), .B2(n19910), .ZN(
        n19901) );
  AOI22_X1 U23047 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19912), .B1(
        n19899), .B2(n19906), .ZN(n19900) );
  OAI211_X1 U23048 ( .C1(n19903), .C2(n19902), .A(n19901), .B(n19900), .ZN(
        P3_U2984) );
  AOI22_X1 U23049 ( .A1(n19968), .A2(n19952), .B1(n19951), .B2(n19910), .ZN(
        n19905) );
  AOI22_X1 U23050 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19912), .B1(
        n19911), .B2(n19953), .ZN(n19904) );
  OAI211_X1 U23051 ( .C1(n19956), .C2(n19915), .A(n19905), .B(n19904), .ZN(
        P3_U2985) );
  AOI22_X1 U23052 ( .A1(n19911), .A2(n19958), .B1(n19957), .B2(n19910), .ZN(
        n19908) );
  AOI22_X1 U23053 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19912), .B1(
        n19960), .B2(n19906), .ZN(n19907) );
  OAI211_X1 U23054 ( .C1(n19909), .C2(n19964), .A(n19908), .B(n19907), .ZN(
        P3_U2986) );
  AOI22_X1 U23055 ( .A1(n19911), .A2(n19967), .B1(n19966), .B2(n19910), .ZN(
        n19914) );
  AOI22_X1 U23056 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19912), .B1(
        n19968), .B2(n19970), .ZN(n19913) );
  OAI211_X1 U23057 ( .C1(n19975), .C2(n19915), .A(n19914), .B(n19913), .ZN(
        P3_U2987) );
  NOR2_X1 U23058 ( .A1(n20050), .A2(n19916), .ZN(n19965) );
  AOI22_X1 U23059 ( .A1(n19918), .A2(n19968), .B1(n19917), .B2(n19965), .ZN(
        n19925) );
  AOI22_X1 U23060 ( .A1(n19922), .A2(n19921), .B1(n19920), .B2(n19919), .ZN(
        n19971) );
  AOI22_X1 U23061 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19971), .B1(
        n19923), .B2(n19969), .ZN(n19924) );
  OAI211_X1 U23062 ( .C1(n19926), .C2(n19974), .A(n19925), .B(n19924), .ZN(
        P3_U2988) );
  AOI22_X1 U23063 ( .A1(n19968), .A2(n19928), .B1(n19927), .B2(n19965), .ZN(
        n19931) );
  AOI22_X1 U23064 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19971), .B1(
        n19929), .B2(n19969), .ZN(n19930) );
  OAI211_X1 U23065 ( .C1(n19932), .C2(n19974), .A(n19931), .B(n19930), .ZN(
        P3_U2989) );
  AOI22_X1 U23066 ( .A1(n19968), .A2(n19934), .B1(n19933), .B2(n19965), .ZN(
        n19937) );
  AOI22_X1 U23067 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19971), .B1(
        n19935), .B2(n19969), .ZN(n19936) );
  OAI211_X1 U23068 ( .C1(n19938), .C2(n19974), .A(n19937), .B(n19936), .ZN(
        P3_U2990) );
  AOI22_X1 U23069 ( .A1(n19968), .A2(n19940), .B1(n19939), .B2(n19965), .ZN(
        n19943) );
  AOI22_X1 U23070 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19971), .B1(
        n19941), .B2(n19959), .ZN(n19942) );
  OAI211_X1 U23071 ( .C1(n19944), .C2(n19963), .A(n19943), .B(n19942), .ZN(
        P3_U2991) );
  AOI22_X1 U23072 ( .A1(n19968), .A2(n19946), .B1(n19945), .B2(n19965), .ZN(
        n19949) );
  AOI22_X1 U23073 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19971), .B1(
        n19947), .B2(n19969), .ZN(n19948) );
  OAI211_X1 U23074 ( .C1(n19950), .C2(n19974), .A(n19949), .B(n19948), .ZN(
        P3_U2992) );
  AOI22_X1 U23075 ( .A1(n19952), .A2(n19969), .B1(n19951), .B2(n19965), .ZN(
        n19955) );
  AOI22_X1 U23076 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19971), .B1(
        n19968), .B2(n19953), .ZN(n19954) );
  OAI211_X1 U23077 ( .C1(n19956), .C2(n19974), .A(n19955), .B(n19954), .ZN(
        P3_U2993) );
  AOI22_X1 U23078 ( .A1(n19968), .A2(n19958), .B1(n19957), .B2(n19965), .ZN(
        n19962) );
  AOI22_X1 U23079 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19971), .B1(
        n19960), .B2(n19959), .ZN(n19961) );
  OAI211_X1 U23080 ( .C1(n19964), .C2(n19963), .A(n19962), .B(n19961), .ZN(
        P3_U2994) );
  AOI22_X1 U23081 ( .A1(n19968), .A2(n19967), .B1(n19966), .B2(n19965), .ZN(
        n19973) );
  AOI22_X1 U23082 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19971), .B1(
        n19970), .B2(n19969), .ZN(n19972) );
  OAI211_X1 U23083 ( .C1(n19975), .C2(n19974), .A(n19973), .B(n19972), .ZN(
        P3_U2995) );
  NOR2_X1 U23084 ( .A1(n19977), .A2(n19976), .ZN(n19979) );
  OAI222_X1 U23085 ( .A1(n19983), .A2(n19982), .B1(n19981), .B2(n19980), .C1(
        n19979), .C2(n19978), .ZN(n20198) );
  OAI21_X1 U23086 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19984), .ZN(n19985) );
  OAI211_X1 U23087 ( .C1(n20013), .C2(n19987), .A(n19986), .B(n19985), .ZN(
        n20035) );
  AND2_X1 U23088 ( .A1(n20169), .A2(n20006), .ZN(n19999) );
  NOR2_X1 U23089 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19988), .ZN(
        n20017) );
  OAI22_X1 U23090 ( .A1(n20009), .A2(n19999), .B1(n19989), .B2(n20017), .ZN(
        n19990) );
  AND2_X1 U23091 ( .A1(n20160), .A2(n19990), .ZN(n20157) );
  AOI22_X1 U23092 ( .A1(n19993), .A2(n19992), .B1(n13477), .B2(n19991), .ZN(
        n19998) );
  NAND2_X1 U23093 ( .A1(n19994), .A2(n19998), .ZN(n20007) );
  NOR2_X1 U23094 ( .A1(n19996), .A2(n19995), .ZN(n19997) );
  AOI21_X1 U23095 ( .B1(n19998), .B2(n19997), .A(n20005), .ZN(n20000) );
  AOI211_X1 U23096 ( .C1(n20184), .C2(n20007), .A(n20000), .B(n19999), .ZN(
        n20158) );
  AOI21_X1 U23097 ( .B1(n20158), .B2(n20013), .A(n20160), .ZN(n20001) );
  AOI21_X1 U23098 ( .B1(n20013), .B2(n20157), .A(n20001), .ZN(n20033) );
  NAND2_X1 U23099 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20014), .ZN(
        n20002) );
  AOI211_X1 U23100 ( .C1(n20003), .C2(n20002), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n20177), .ZN(n20012) );
  AOI211_X1 U23101 ( .C1(n20169), .C2(n20177), .A(n20005), .B(n20004), .ZN(
        n20011) );
  OAI221_X1 U23102 ( .B1(n20007), .B2(n20177), .C1(n20007), .C2(n10008), .A(
        n20006), .ZN(n20008) );
  OAI22_X1 U23103 ( .A1(n20166), .A2(n20009), .B1(n20169), .B2(n20008), .ZN(
        n20010) );
  NOR3_X1 U23104 ( .A1(n20012), .A2(n20011), .A3(n20010), .ZN(n20163) );
  AOI22_X1 U23105 ( .A1(n20024), .A2(n20169), .B1(n20163), .B2(n20013), .ZN(
        n20028) );
  NOR2_X1 U23106 ( .A1(n20015), .A2(n20014), .ZN(n20018) );
  AOI22_X1 U23107 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20016), .B1(
        n20018), .B2(n20184), .ZN(n20179) );
  OAI22_X1 U23108 ( .A1(n20018), .A2(n20170), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20017), .ZN(n20175) );
  OR3_X1 U23109 ( .A1(n20179), .A2(n20021), .A3(n20019), .ZN(n20020) );
  AOI22_X1 U23110 ( .A1(n20179), .A2(n20021), .B1(n20175), .B2(n20020), .ZN(
        n20023) );
  OAI21_X1 U23111 ( .B1(n20024), .B2(n20023), .A(n20022), .ZN(n20027) );
  AND2_X1 U23112 ( .A1(n20028), .A2(n20027), .ZN(n20025) );
  OAI221_X1 U23113 ( .B1(n20028), .B2(n20027), .C1(n20026), .C2(n20025), .A(
        n20030), .ZN(n20032) );
  AOI21_X1 U23114 ( .B1(n20030), .B2(n20029), .A(n20028), .ZN(n20031) );
  AOI222_X1 U23115 ( .A1(n20033), .A2(n20032), .B1(n20033), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n20032), .C2(n20031), .ZN(
        n20034) );
  NOR4_X1 U23116 ( .A1(n20036), .A2(n20198), .A3(n20035), .A4(n20034), .ZN(
        n20046) );
  AOI22_X1 U23117 ( .A1(n20178), .A2(n20209), .B1(n10001), .B2(n18790), .ZN(
        n20037) );
  INV_X1 U23118 ( .A(n20037), .ZN(n20043) );
  OAI211_X1 U23119 ( .C1(n20040), .C2(n20039), .A(n20038), .B(n20046), .ZN(
        n20152) );
  OAI21_X1 U23120 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n20206), .A(n20152), 
        .ZN(n20048) );
  NOR2_X1 U23121 ( .A1(n20041), .A2(n20048), .ZN(n20042) );
  MUX2_X1 U23122 ( .A(n20043), .B(n20042), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n20045) );
  OAI211_X1 U23123 ( .C1(n20046), .C2(n20202), .A(n20045), .B(n20044), .ZN(
        P3_U2996) );
  NAND2_X1 U23124 ( .A1(n10001), .A2(n18790), .ZN(n20052) );
  NAND4_X1 U23125 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n10001), .A4(n20047), .ZN(n20054) );
  OR3_X1 U23126 ( .A1(n20050), .A2(n20049), .A3(n20048), .ZN(n20051) );
  NAND4_X1 U23127 ( .A1(n20053), .A2(n20052), .A3(n20054), .A4(n20051), .ZN(
        P3_U2997) );
  AND4_X1 U23128 ( .A1(n20056), .A2(n20055), .A3(n20054), .A4(n20151), .ZN(
        P3_U2998) );
  AND2_X1 U23129 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n20147), .ZN(
        P3_U2999) );
  AND2_X1 U23130 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n20147), .ZN(
        P3_U3000) );
  AND2_X1 U23131 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n20057), .ZN(
        P3_U3001) );
  AND2_X1 U23132 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n20057), .ZN(
        P3_U3002) );
  AND2_X1 U23133 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n20057), .ZN(
        P3_U3003) );
  AND2_X1 U23134 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n20057), .ZN(
        P3_U3004) );
  AND2_X1 U23135 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n20057), .ZN(
        P3_U3005) );
  AND2_X1 U23136 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n20057), .ZN(
        P3_U3006) );
  AND2_X1 U23137 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n20057), .ZN(
        P3_U3007) );
  AND2_X1 U23138 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n20057), .ZN(
        P3_U3008) );
  AND2_X1 U23139 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n20057), .ZN(
        P3_U3009) );
  AND2_X1 U23140 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n20057), .ZN(
        P3_U3010) );
  AND2_X1 U23141 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n20057), .ZN(
        P3_U3011) );
  AND2_X1 U23142 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n20057), .ZN(
        P3_U3012) );
  AND2_X1 U23143 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n20057), .ZN(
        P3_U3013) );
  AND2_X1 U23144 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n20057), .ZN(
        P3_U3014) );
  AND2_X1 U23145 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n20057), .ZN(
        P3_U3015) );
  AND2_X1 U23146 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n20057), .ZN(
        P3_U3016) );
  AND2_X1 U23147 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n20057), .ZN(
        P3_U3017) );
  AND2_X1 U23148 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n20057), .ZN(
        P3_U3018) );
  AND2_X1 U23149 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n20057), .ZN(
        P3_U3019) );
  AND2_X1 U23150 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n20057), .ZN(
        P3_U3020) );
  AND2_X1 U23151 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n20057), .ZN(P3_U3021) );
  AND2_X1 U23152 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n20147), .ZN(P3_U3022) );
  AND2_X1 U23153 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n20147), .ZN(P3_U3023) );
  AND2_X1 U23154 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n20147), .ZN(P3_U3024) );
  AND2_X1 U23155 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n20147), .ZN(P3_U3025) );
  AND2_X1 U23156 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n20147), .ZN(P3_U3026) );
  AND2_X1 U23157 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n20057), .ZN(P3_U3027) );
  AND2_X1 U23158 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n20147), .ZN(P3_U3028) );
  NOR2_X1 U23159 ( .A1(n20206), .A2(n20060), .ZN(n20065) );
  OAI21_X1 U23160 ( .B1(n20058), .B2(n21444), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n20059) );
  AOI22_X1 U23161 ( .A1(n20065), .A2(n20074), .B1(n20195), .B2(n20059), .ZN(
        n20061) );
  NAND3_X1 U23162 ( .A1(NA), .A2(n20071), .A3(n20060), .ZN(n20066) );
  OAI211_X1 U23163 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n20061), .B(n20066), .ZN(P3_U3029) );
  NOR2_X1 U23164 ( .A1(n20074), .A2(n21444), .ZN(n20069) );
  INV_X1 U23165 ( .A(n20069), .ZN(n20063) );
  AOI22_X1 U23166 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n20063), .B1(HOLD), 
        .B2(n20062), .ZN(n20064) );
  INV_X1 U23167 ( .A(n20065), .ZN(n20067) );
  OAI211_X1 U23168 ( .C1(n20064), .C2(n20071), .A(n20067), .B(n20203), .ZN(
        P3_U3030) );
  AOI21_X1 U23169 ( .B1(n20071), .B2(n20066), .A(n20065), .ZN(n20072) );
  OAI22_X1 U23170 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n20067), .ZN(n20068) );
  OAI22_X1 U23171 ( .A1(n20069), .A2(n20068), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n20070) );
  OAI22_X1 U23172 ( .A1(n20072), .A2(n20074), .B1(n20071), .B2(n20070), .ZN(
        P3_U3031) );
  NAND2_X1 U23173 ( .A1(n20129), .A2(n20074), .ZN(n20128) );
  CLKBUF_X1 U23174 ( .A(n20128), .Z(n20134) );
  OAI222_X1 U23175 ( .A1(n20186), .A2(n20138), .B1(n20075), .B2(n20129), .C1(
        n20076), .C2(n20134), .ZN(P3_U3032) );
  OAI222_X1 U23176 ( .A1(n20134), .A2(n20078), .B1(n20077), .B2(n20129), .C1(
        n20076), .C2(n20138), .ZN(P3_U3033) );
  OAI222_X1 U23177 ( .A1(n20134), .A2(n20080), .B1(n20079), .B2(n20129), .C1(
        n20078), .C2(n20138), .ZN(P3_U3034) );
  OAI222_X1 U23178 ( .A1(n20134), .A2(n20082), .B1(n20081), .B2(n20129), .C1(
        n20080), .C2(n20138), .ZN(P3_U3035) );
  INV_X1 U23179 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20084) );
  OAI222_X1 U23180 ( .A1(n20134), .A2(n20084), .B1(n20083), .B2(n20129), .C1(
        n20082), .C2(n20138), .ZN(P3_U3036) );
  OAI222_X1 U23181 ( .A1(n20134), .A2(n20086), .B1(n20085), .B2(n20129), .C1(
        n20084), .C2(n20138), .ZN(P3_U3037) );
  OAI222_X1 U23182 ( .A1(n20134), .A2(n20089), .B1(n20087), .B2(n20129), .C1(
        n20086), .C2(n20138), .ZN(P3_U3038) );
  OAI222_X1 U23183 ( .A1(n20089), .A2(n20138), .B1(n20088), .B2(n20129), .C1(
        n20090), .C2(n20134), .ZN(P3_U3039) );
  OAI222_X1 U23184 ( .A1(n20134), .A2(n20092), .B1(n20091), .B2(n20129), .C1(
        n20090), .C2(n20138), .ZN(P3_U3040) );
  OAI222_X1 U23185 ( .A1(n20134), .A2(n20095), .B1(n20093), .B2(n20129), .C1(
        n20092), .C2(n20138), .ZN(P3_U3041) );
  INV_X1 U23186 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20096) );
  OAI222_X1 U23187 ( .A1(n20095), .A2(n20138), .B1(n20094), .B2(n20129), .C1(
        n20096), .C2(n20134), .ZN(P3_U3042) );
  OAI222_X1 U23188 ( .A1(n20134), .A2(n20098), .B1(n20097), .B2(n20129), .C1(
        n20096), .C2(n20138), .ZN(P3_U3043) );
  INV_X1 U23189 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20101) );
  OAI222_X1 U23190 ( .A1(n20134), .A2(n20101), .B1(n20099), .B2(n20129), .C1(
        n20098), .C2(n20138), .ZN(P3_U3044) );
  INV_X1 U23191 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20102) );
  OAI222_X1 U23192 ( .A1(n20138), .A2(n20101), .B1(n20100), .B2(n20129), .C1(
        n20102), .C2(n20134), .ZN(P3_U3045) );
  OAI222_X1 U23193 ( .A1(n20128), .A2(n20104), .B1(n20103), .B2(n20129), .C1(
        n20102), .C2(n20138), .ZN(P3_U3046) );
  OAI222_X1 U23194 ( .A1(n20128), .A2(n20106), .B1(n20105), .B2(n20129), .C1(
        n20104), .C2(n20138), .ZN(P3_U3047) );
  OAI222_X1 U23195 ( .A1(n20128), .A2(n20108), .B1(n20107), .B2(n20129), .C1(
        n20106), .C2(n20138), .ZN(P3_U3048) );
  OAI222_X1 U23196 ( .A1(n20128), .A2(n20110), .B1(n20109), .B2(n20129), .C1(
        n20108), .C2(n20138), .ZN(P3_U3049) );
  OAI222_X1 U23197 ( .A1(n20128), .A2(n20112), .B1(n20111), .B2(n20129), .C1(
        n20110), .C2(n20138), .ZN(P3_U3050) );
  OAI222_X1 U23198 ( .A1(n20128), .A2(n20114), .B1(n20113), .B2(n20129), .C1(
        n20112), .C2(n20138), .ZN(P3_U3051) );
  INV_X1 U23199 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20116) );
  OAI222_X1 U23200 ( .A1(n20128), .A2(n20116), .B1(n20115), .B2(n20129), .C1(
        n20114), .C2(n20138), .ZN(P3_U3052) );
  OAI222_X1 U23201 ( .A1(n20134), .A2(n20118), .B1(n20117), .B2(n20129), .C1(
        n20116), .C2(n20138), .ZN(P3_U3053) );
  INV_X1 U23202 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20120) );
  OAI222_X1 U23203 ( .A1(n20134), .A2(n20120), .B1(n20119), .B2(n20129), .C1(
        n20118), .C2(n20138), .ZN(P3_U3054) );
  OAI222_X1 U23204 ( .A1(n20128), .A2(n20122), .B1(n20121), .B2(n20129), .C1(
        n20120), .C2(n20138), .ZN(P3_U3055) );
  OAI222_X1 U23205 ( .A1(n20134), .A2(n20124), .B1(n20123), .B2(n20129), .C1(
        n20122), .C2(n20138), .ZN(P3_U3056) );
  OAI222_X1 U23206 ( .A1(n20134), .A2(n20126), .B1(n20125), .B2(n20129), .C1(
        n20124), .C2(n20138), .ZN(P3_U3057) );
  OAI222_X1 U23207 ( .A1(n20128), .A2(n20131), .B1(n20127), .B2(n20129), .C1(
        n20126), .C2(n20138), .ZN(P3_U3058) );
  OAI222_X1 U23208 ( .A1(n20131), .A2(n20138), .B1(n20130), .B2(n20129), .C1(
        n20132), .C2(n20134), .ZN(P3_U3059) );
  OAI222_X1 U23209 ( .A1(n20134), .A2(n20137), .B1(n20133), .B2(n20129), .C1(
        n20132), .C2(n20138), .ZN(P3_U3060) );
  OAI222_X1 U23210 ( .A1(n20138), .A2(n20137), .B1(n20136), .B2(n20129), .C1(
        n20135), .C2(n20134), .ZN(P3_U3061) );
  INV_X1 U23211 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n20139) );
  AOI22_X1 U23212 ( .A1(n20129), .A2(n20140), .B1(n20139), .B2(n20195), .ZN(
        P3_U3274) );
  INV_X1 U23213 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20188) );
  INV_X1 U23214 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n20141) );
  AOI22_X1 U23215 ( .A1(n20129), .A2(n20188), .B1(n20141), .B2(n20195), .ZN(
        P3_U3275) );
  INV_X1 U23216 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n20142) );
  AOI22_X1 U23217 ( .A1(n20129), .A2(n20143), .B1(n20142), .B2(n20195), .ZN(
        P3_U3276) );
  INV_X1 U23218 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20194) );
  INV_X1 U23219 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n20144) );
  AOI22_X1 U23220 ( .A1(n20129), .A2(n20194), .B1(n20144), .B2(n20195), .ZN(
        P3_U3277) );
  INV_X1 U23221 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20146) );
  INV_X1 U23222 ( .A(n20148), .ZN(n20145) );
  AOI21_X1 U23223 ( .B1(n20147), .B2(n20146), .A(n20145), .ZN(P3_U3280) );
  OAI21_X1 U23224 ( .B1(n20150), .B2(n20149), .A(n20148), .ZN(P3_U3281) );
  OAI221_X1 U23225 ( .B1(n20153), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n20153), 
        .C2(n20152), .A(n20151), .ZN(P3_U3282) );
  INV_X1 U23226 ( .A(n20154), .ZN(n20180) );
  INV_X1 U23227 ( .A(n20155), .ZN(n20156) );
  AOI22_X1 U23228 ( .A1(n20180), .A2(n20157), .B1(n20178), .B2(n20156), .ZN(
        n20162) );
  INV_X1 U23229 ( .A(n20158), .ZN(n20159) );
  AOI21_X1 U23230 ( .B1(n20180), .B2(n20159), .A(n20185), .ZN(n20161) );
  OAI22_X1 U23231 ( .A1(n20185), .A2(n20162), .B1(n20161), .B2(n20160), .ZN(
        P3_U3285) );
  INV_X1 U23232 ( .A(n20163), .ZN(n20167) );
  NOR2_X1 U23233 ( .A1(n20164), .A2(n20181), .ZN(n20172) );
  AOI22_X1 U23234 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n9952), .B2(n20165), .ZN(
        n20171) );
  AOI222_X1 U23235 ( .A1(n20167), .A2(n20180), .B1(n20172), .B2(n20171), .C1(
        n20178), .C2(n20166), .ZN(n20168) );
  AOI22_X1 U23236 ( .A1(n20185), .A2(n20169), .B1(n20168), .B2(n20182), .ZN(
        P3_U3288) );
  INV_X1 U23237 ( .A(n20170), .ZN(n20174) );
  INV_X1 U23238 ( .A(n20171), .ZN(n20173) );
  AOI222_X1 U23239 ( .A1(n20175), .A2(n20180), .B1(n20178), .B2(n20174), .C1(
        n20173), .C2(n20172), .ZN(n20176) );
  AOI22_X1 U23240 ( .A1(n20185), .A2(n20177), .B1(n20176), .B2(n20182), .ZN(
        P3_U3289) );
  AOI222_X1 U23241 ( .A1(n20181), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n20180), 
        .B2(n20179), .C1(n20184), .C2(n20178), .ZN(n20183) );
  AOI22_X1 U23242 ( .A1(n20185), .A2(n20184), .B1(n20183), .B2(n20182), .ZN(
        P3_U3290) );
  AOI21_X1 U23243 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20187) );
  AOI22_X1 U23244 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n20187), .B2(n20186), .ZN(n20189) );
  AOI22_X1 U23245 ( .A1(n20190), .A2(n20189), .B1(n20188), .B2(n20193), .ZN(
        P3_U3292) );
  NOR2_X1 U23246 ( .A1(n20193), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n20191) );
  AOI22_X1 U23247 ( .A1(n20194), .A2(n20193), .B1(n20192), .B2(n20191), .ZN(
        P3_U3293) );
  INV_X1 U23248 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n20196) );
  AOI22_X1 U23249 ( .A1(n20129), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n20196), 
        .B2(n20195), .ZN(P3_U3294) );
  MUX2_X1 U23250 ( .A(P3_MORE_REG_SCAN_IN), .B(n20198), .S(n20197), .Z(
        P3_U3295) );
  OAI21_X1 U23251 ( .B1(n10001), .B2(n20199), .A(n20216), .ZN(n20200) );
  AOI21_X1 U23252 ( .B1(n20202), .B2(n20201), .A(n20200), .ZN(n20213) );
  AOI21_X1 U23253 ( .B1(n20205), .B2(n20204), .A(n20203), .ZN(n20207) );
  OAI211_X1 U23254 ( .C1(n20208), .C2(n20207), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n20206), .ZN(n20210) );
  AOI21_X1 U23255 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20210), .A(n20209), 
        .ZN(n20212) );
  NAND2_X1 U23256 ( .A1(n20213), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20211) );
  OAI21_X1 U23257 ( .B1(n20213), .B2(n20212), .A(n20211), .ZN(P3_U3296) );
  MUX2_X1 U23258 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20129), .Z(P3_U3297) );
  OAI21_X1 U23259 ( .B1(n20217), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n20216), 
        .ZN(n20214) );
  OAI21_X1 U23260 ( .B1(n20216), .B2(n20215), .A(n20214), .ZN(P3_U3298) );
  NOR2_X1 U23261 ( .A1(n20217), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n20219)
         );
  OAI21_X1 U23262 ( .B1(n20220), .B2(n20219), .A(n20218), .ZN(P3_U3299) );
  INV_X1 U23263 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n20221) );
  INV_X1 U23264 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21112) );
  AND2_X1 U23265 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21112), .ZN(n21102) );
  NOR2_X1 U23266 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n21094) );
  AOI21_X1 U23267 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21102), .A(n21094), 
        .ZN(n21090) );
  INV_X1 U23268 ( .A(n21090), .ZN(n21175) );
  INV_X1 U23269 ( .A(n21175), .ZN(n21092) );
  OAI21_X1 U23270 ( .B1(n21099), .B2(n20221), .A(n21092), .ZN(P2_U2815) );
  AOI22_X1 U23271 ( .A1(n21082), .A2(n21084), .B1(n21239), .B2(
        P2_CODEFETCH_REG_SCAN_IN), .ZN(n20222) );
  INV_X1 U23272 ( .A(n20222), .ZN(P2_U2816) );
  INV_X1 U23273 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n20223) );
  AOI22_X1 U23274 ( .A1(n21244), .A2(n20223), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n21245), .ZN(n20224) );
  OAI21_X1 U23275 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21106), .A(n20224), 
        .ZN(P2_U2817) );
  OAI21_X1 U23276 ( .B1(n21095), .B2(BS16), .A(n21175), .ZN(n21173) );
  OAI21_X1 U23277 ( .B1(n21175), .B2(n12132), .A(n21173), .ZN(P2_U2818) );
  INV_X1 U23278 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21171) );
  NOR4_X1 U23279 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20234) );
  NOR4_X1 U23280 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20233) );
  AOI211_X1 U23281 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_5__SCAN_IN), .B(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20225) );
  NAND3_X1 U23282 ( .A1(n20225), .A2(n21091), .A3(n21089), .ZN(n20231) );
  NOR4_X1 U23283 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20229) );
  NOR4_X1 U23284 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20228) );
  NOR4_X1 U23285 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20227) );
  NOR4_X1 U23286 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20226) );
  NAND4_X1 U23287 ( .A1(n20229), .A2(n20228), .A3(n20227), .A4(n20226), .ZN(
        n20230) );
  NOR4_X1 U23288 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(n20231), .A4(n20230), .ZN(n20232) );
  NAND3_X1 U23289 ( .A1(n20234), .A2(n20233), .A3(n20232), .ZN(n20237) );
  NOR2_X1 U23290 ( .A1(n20237), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n20235) );
  AOI22_X1 U23291 ( .A1(n21171), .A2(n20237), .B1(n20395), .B2(n20235), .ZN(
        P2_U2820) );
  INV_X1 U23292 ( .A(n20237), .ZN(n20243) );
  INV_X1 U23293 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21169) );
  NOR2_X1 U23294 ( .A1(P2_DATAWIDTH_REG_1__SCAN_IN), .A2(n20237), .ZN(n20238)
         );
  INV_X1 U23295 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20236) );
  NAND3_X1 U23296 ( .A1(n20238), .A2(n20395), .A3(n20236), .ZN(n20242) );
  OAI221_X1 U23297 ( .B1(n20243), .B2(n21169), .C1(n20237), .C2(n21114), .A(
        n20242), .ZN(P2_U2821) );
  NAND2_X1 U23298 ( .A1(n20238), .A2(n21114), .ZN(n20241) );
  OAI21_X1 U23299 ( .B1(n20395), .B2(n21114), .A(n20243), .ZN(n20239) );
  OAI21_X1 U23300 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n20243), .A(n20239), 
        .ZN(n20240) );
  OAI221_X1 U23301 ( .B1(n20241), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n20241), .C2(P2_REIP_REG_0__SCAN_IN), .A(n20240), .ZN(P2_U2822) );
  INV_X1 U23302 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21165) );
  OAI211_X1 U23303 ( .C1(n20243), .C2(n21165), .A(n20242), .B(n20241), .ZN(
        P2_U2823) );
  AOI22_X1 U23304 ( .A1(n20244), .A2(n20328), .B1(P2_REIP_REG_20__SCAN_IN), 
        .B2(n20406), .ZN(n20252) );
  AOI22_X1 U23305 ( .A1(n20359), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20412), .ZN(n20251) );
  AOI22_X1 U23306 ( .A1(n10332), .A2(n20378), .B1(n20385), .B2(n20245), .ZN(
        n20250) );
  AOI21_X1 U23307 ( .B1(n20247), .B2(n9935), .A(n20246), .ZN(n20248) );
  NAND2_X1 U23308 ( .A1(n20370), .A2(n20248), .ZN(n20249) );
  NAND4_X1 U23309 ( .A1(n20252), .A2(n20251), .A3(n20250), .A4(n20249), .ZN(
        P2_U2835) );
  NOR2_X1 U23310 ( .A1(n12815), .A2(n20253), .ZN(n20254) );
  XNOR2_X1 U23311 ( .A(n20255), .B(n20254), .ZN(n20262) );
  OAI21_X1 U23312 ( .B1(n20396), .B2(n11920), .A(n20324), .ZN(n20259) );
  INV_X1 U23313 ( .A(n20256), .ZN(n20257) );
  OAI22_X1 U23314 ( .A1(n20257), .A2(n20399), .B1(n10149), .B2(n20380), .ZN(
        n20258) );
  AOI211_X1 U23315 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n20406), .A(n20259), 
        .B(n20258), .ZN(n20261) );
  AOI22_X1 U23316 ( .A1(n20446), .A2(n20378), .B1(n20385), .B2(n20418), .ZN(
        n20260) );
  OAI211_X1 U23317 ( .C1(n21086), .C2(n20262), .A(n20261), .B(n20260), .ZN(
        P2_U2839) );
  XNOR2_X1 U23318 ( .A(n20264), .B(n20263), .ZN(n20272) );
  AOI22_X1 U23319 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20412), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n20406), .ZN(n20265) );
  OAI211_X1 U23320 ( .C1(n20396), .C2(n20266), .A(n20265), .B(n20347), .ZN(
        n20267) );
  AOI21_X1 U23321 ( .B1(n20268), .B2(n20328), .A(n20267), .ZN(n20271) );
  AOI22_X1 U23322 ( .A1(n20452), .A2(n20378), .B1(n20385), .B2(n20269), .ZN(
        n20270) );
  OAI211_X1 U23323 ( .C1(n21086), .C2(n20272), .A(n20271), .B(n20270), .ZN(
        P2_U2841) );
  NOR2_X1 U23324 ( .A1(n12815), .A2(n20273), .ZN(n20275) );
  XOR2_X1 U23325 ( .A(n20275), .B(n20274), .Z(n20285) );
  INV_X1 U23326 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n20425) );
  INV_X1 U23327 ( .A(n20276), .ZN(n20278) );
  OAI211_X1 U23328 ( .C1(n20425), .C2(n20278), .A(n20277), .B(n20328), .ZN(
        n20281) );
  OR2_X1 U23329 ( .A1(n20396), .A2(n20425), .ZN(n20280) );
  NAND2_X1 U23330 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20412), .ZN(
        n20279) );
  NAND4_X1 U23331 ( .A1(n20281), .A2(n20324), .A3(n20280), .A4(n20279), .ZN(
        n20282) );
  AOI21_X1 U23332 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n20406), .A(n20282), 
        .ZN(n20284) );
  AOI22_X1 U23333 ( .A1(n20458), .A2(n20378), .B1(n20385), .B2(n10334), .ZN(
        n20283) );
  OAI211_X1 U23334 ( .C1(n21086), .C2(n20285), .A(n20284), .B(n20283), .ZN(
        P2_U2843) );
  OAI21_X1 U23335 ( .B1(n20396), .B2(n20286), .A(n20347), .ZN(n20290) );
  OAI22_X1 U23336 ( .A1(n20288), .A2(n20399), .B1(n20287), .B2(n20380), .ZN(
        n20289) );
  AOI211_X1 U23337 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n20406), .A(n20290), 
        .B(n20289), .ZN(n20297) );
  NAND2_X1 U23338 ( .A1(n15196), .A2(n20291), .ZN(n20292) );
  XNOR2_X1 U23339 ( .A(n20293), .B(n20292), .ZN(n20295) );
  AOI22_X1 U23340 ( .A1(n20295), .A2(n20370), .B1(n20385), .B2(n20294), .ZN(
        n20296) );
  OAI211_X1 U23341 ( .C1(n20462), .C2(n20401), .A(n20297), .B(n20296), .ZN(
        P2_U2844) );
  NAND2_X1 U23342 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20412), .ZN(
        n20298) );
  OAI211_X1 U23343 ( .C1(n20396), .C2(n20433), .A(n20347), .B(n20298), .ZN(
        n20299) );
  AOI21_X1 U23344 ( .B1(n20300), .B2(n20328), .A(n20299), .ZN(n20301) );
  INV_X1 U23345 ( .A(n20301), .ZN(n20302) );
  AOI21_X1 U23346 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n20406), .A(n20302), 
        .ZN(n20308) );
  NOR2_X1 U23347 ( .A1(n12815), .A2(n20303), .ZN(n20305) );
  XNOR2_X1 U23348 ( .A(n20305), .B(n20304), .ZN(n20306) );
  AOI22_X1 U23349 ( .A1(n20306), .A2(n20370), .B1(n20385), .B2(n20431), .ZN(
        n20307) );
  OAI211_X1 U23350 ( .C1(n20401), .C2(n20465), .A(n20308), .B(n20307), .ZN(
        P2_U2845) );
  OAI21_X1 U23351 ( .B1(n20396), .B2(n10232), .A(n20347), .ZN(n20312) );
  OAI22_X1 U23352 ( .A1(n20310), .A2(n20399), .B1(n20309), .B2(n20380), .ZN(
        n20311) );
  AOI211_X1 U23353 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n20406), .A(n20312), .B(
        n20311), .ZN(n20319) );
  NAND2_X1 U23354 ( .A1(n15196), .A2(n20313), .ZN(n20314) );
  XNOR2_X1 U23355 ( .A(n20315), .B(n20314), .ZN(n20317) );
  AOI22_X1 U23356 ( .A1(n20317), .A2(n20370), .B1(n20385), .B2(n20316), .ZN(
        n20318) );
  OAI211_X1 U23357 ( .C1(n20401), .C2(n20467), .A(n20319), .B(n20318), .ZN(
        P2_U2846) );
  NOR2_X1 U23358 ( .A1(n12815), .A2(n20320), .ZN(n20322) );
  XOR2_X1 U23359 ( .A(n20322), .B(n20321), .Z(n20335) );
  INV_X1 U23360 ( .A(n20323), .ZN(n20329) );
  INV_X1 U23361 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n20326) );
  AOI22_X1 U23362 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20412), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n20406), .ZN(n20325) );
  OAI211_X1 U23363 ( .C1(n20396), .C2(n20326), .A(n20325), .B(n20324), .ZN(
        n20327) );
  AOI21_X1 U23364 ( .B1(n20329), .B2(n20328), .A(n20327), .ZN(n20334) );
  INV_X1 U23365 ( .A(n20330), .ZN(n20471) );
  OAI22_X1 U23366 ( .A1(n20402), .A2(n20331), .B1(n20401), .B2(n20471), .ZN(
        n20332) );
  INV_X1 U23367 ( .A(n20332), .ZN(n20333) );
  OAI211_X1 U23368 ( .C1(n21086), .C2(n20335), .A(n20334), .B(n20333), .ZN(
        P2_U2847) );
  NAND2_X1 U23369 ( .A1(n15196), .A2(n20336), .ZN(n20338) );
  XOR2_X1 U23370 ( .A(n20338), .B(n20337), .Z(n20346) );
  OAI21_X1 U23371 ( .B1(n20396), .B2(n11874), .A(n20347), .ZN(n20339) );
  AOI21_X1 U23372 ( .B1(n20406), .B2(P2_REIP_REG_7__SCAN_IN), .A(n20339), .ZN(
        n20340) );
  OAI21_X1 U23373 ( .B1(n20341), .B2(n20399), .A(n20340), .ZN(n20344) );
  OAI22_X1 U23374 ( .A1(n20472), .A2(n20401), .B1(n20402), .B2(n20342), .ZN(
        n20343) );
  AOI211_X1 U23375 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n20412), .A(
        n20344), .B(n20343), .ZN(n20345) );
  OAI21_X1 U23376 ( .B1(n20346), .B2(n21086), .A(n20345), .ZN(P2_U2848) );
  OAI21_X1 U23377 ( .B1(n20396), .B2(n20348), .A(n20347), .ZN(n20351) );
  OAI22_X1 U23378 ( .A1(n20374), .A2(n21121), .B1(n20399), .B2(n20349), .ZN(
        n20350) );
  AOI211_X1 U23379 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n20412), .A(
        n20351), .B(n20350), .ZN(n20358) );
  NOR2_X1 U23380 ( .A1(n12815), .A2(n20352), .ZN(n20354) );
  XNOR2_X1 U23381 ( .A(n20354), .B(n20353), .ZN(n20356) );
  AOI22_X1 U23382 ( .A1(n20356), .A2(n20370), .B1(n20385), .B2(n20355), .ZN(
        n20357) );
  OAI211_X1 U23383 ( .C1(n20401), .C2(n20474), .A(n20358), .B(n20357), .ZN(
        P2_U2849) );
  NAND2_X1 U23384 ( .A1(n20406), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n20361) );
  AOI21_X1 U23385 ( .B1(n20359), .B2(P2_EBX_REG_5__SCAN_IN), .A(n20376), .ZN(
        n20360) );
  OAI211_X1 U23386 ( .C1(n20362), .C2(n20399), .A(n20361), .B(n20360), .ZN(
        n20363) );
  INV_X1 U23387 ( .A(n20363), .ZN(n20372) );
  NAND2_X1 U23388 ( .A1(n15196), .A2(n20364), .ZN(n20365) );
  XNOR2_X1 U23389 ( .A(n20366), .B(n20365), .ZN(n20369) );
  OAI22_X1 U23390 ( .A1(n20482), .A2(n20401), .B1(n20402), .B2(n20367), .ZN(
        n20368) );
  AOI21_X1 U23391 ( .B1(n20370), .B2(n20369), .A(n20368), .ZN(n20371) );
  OAI211_X1 U23392 ( .C1(n20373), .C2(n20380), .A(n20372), .B(n20371), .ZN(
        P2_U2850) );
  OAI22_X1 U23393 ( .A1(n20374), .A2(n12303), .B1(n12041), .B2(n20396), .ZN(
        n20375) );
  AOI211_X1 U23394 ( .C1(n20378), .C2(n20377), .A(n20376), .B(n20375), .ZN(
        n20394) );
  OAI22_X1 U23395 ( .A1(n20399), .A2(n20381), .B1(n20380), .B2(n20379), .ZN(
        n20382) );
  INV_X1 U23396 ( .A(n20382), .ZN(n20393) );
  INV_X1 U23397 ( .A(n20383), .ZN(n20478) );
  INV_X1 U23398 ( .A(n20384), .ZN(n20408) );
  AOI22_X1 U23399 ( .A1(n20478), .A2(n20408), .B1(n20385), .B2(n20434), .ZN(
        n20392) );
  INV_X1 U23400 ( .A(n20386), .ZN(n20390) );
  NOR2_X1 U23401 ( .A1(n12815), .A2(n20387), .ZN(n20389) );
  AOI21_X1 U23402 ( .B1(n20390), .B2(n20389), .A(n21086), .ZN(n20388) );
  OAI21_X1 U23403 ( .B1(n20390), .B2(n20389), .A(n20388), .ZN(n20391) );
  NAND4_X1 U23404 ( .A1(n20394), .A2(n20393), .A3(n20392), .A4(n20391), .ZN(
        P2_U2851) );
  OAI22_X1 U23405 ( .A1(n20399), .A2(n20398), .B1(n20397), .B2(n20396), .ZN(
        n20405) );
  OAI22_X1 U23406 ( .A1(n20403), .A2(n20402), .B1(n20401), .B2(n20400), .ZN(
        n20404) );
  AOI211_X1 U23407 ( .C1(n20406), .C2(P2_REIP_REG_0__SCAN_IN), .A(n20405), .B(
        n20404), .ZN(n20415) );
  AOI22_X1 U23408 ( .A1(n20410), .A2(n20409), .B1(n20408), .B2(n20407), .ZN(
        n20414) );
  OAI21_X1 U23409 ( .B1(n20412), .B2(n20411), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20413) );
  NAND3_X1 U23410 ( .A1(n20415), .A2(n20414), .A3(n20413), .ZN(P2_U2855) );
  AOI21_X1 U23411 ( .B1(n20417), .B2(n20416), .A(n15211), .ZN(n20445) );
  AOI22_X1 U23412 ( .A1(n20445), .A2(n20435), .B1(n13216), .B2(n20418), .ZN(
        n20419) );
  OAI21_X1 U23413 ( .B1(n20437), .B2(n11920), .A(n20419), .ZN(P2_U2871) );
  AOI21_X1 U23414 ( .B1(n9925), .B2(n20421), .A(n20420), .ZN(n20422) );
  NOR3_X1 U23415 ( .A1(n20422), .A2(n14509), .A3(n20428), .ZN(n20423) );
  AOI21_X1 U23416 ( .B1(n10334), .B2(n13216), .A(n20423), .ZN(n20424) );
  OAI21_X1 U23417 ( .B1(n20437), .B2(n20425), .A(n20424), .ZN(P2_U2875) );
  AOI21_X1 U23418 ( .B1(n13970), .B2(n20427), .A(n20426), .ZN(n20429) );
  NOR3_X1 U23419 ( .A1(n20429), .A2(n9925), .A3(n20428), .ZN(n20430) );
  AOI21_X1 U23420 ( .B1(n20431), .B2(n13216), .A(n20430), .ZN(n20432) );
  OAI21_X1 U23421 ( .B1(n20437), .B2(n20433), .A(n20432), .ZN(P2_U2877) );
  AOI22_X1 U23422 ( .A1(n20478), .A2(n20435), .B1(n13216), .B2(n20434), .ZN(
        n20436) );
  OAI21_X1 U23423 ( .B1(n20437), .B2(n12041), .A(n20436), .ZN(P2_U2883) );
  INV_X1 U23424 ( .A(n16369), .ZN(n20438) );
  AOI22_X1 U23425 ( .A1(n20438), .A2(n20492), .B1(n20444), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n20440) );
  AOI22_X1 U23426 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n20491), .B1(n20443), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n20439) );
  NAND2_X1 U23427 ( .A1(n20440), .A2(n20439), .ZN(P2_U2888) );
  AOI22_X1 U23428 ( .A1(n20442), .A2(n20441), .B1(n20491), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n20449) );
  AOI22_X1 U23429 ( .A1(n20444), .A2(BUF2_REG_16__SCAN_IN), .B1(n20443), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n20448) );
  AOI22_X1 U23430 ( .A1(n20446), .A2(n20492), .B1(n20477), .B2(n20445), .ZN(
        n20447) );
  NAND3_X1 U23431 ( .A1(n20449), .A2(n20448), .A3(n20447), .ZN(P2_U2903) );
  OAI222_X1 U23432 ( .A1(n20451), .A2(n20483), .B1(n13921), .B2(n20475), .C1(
        n20450), .C2(n20500), .ZN(P2_U2904) );
  INV_X1 U23433 ( .A(n20452), .ZN(n20454) );
  INV_X1 U23434 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20511) );
  OAI222_X1 U23435 ( .A1(n20454), .A2(n20483), .B1(n20511), .B2(n20475), .C1(
        n20500), .C2(n20453), .ZN(P2_U2905) );
  INV_X1 U23436 ( .A(n20455), .ZN(n20457) );
  INV_X1 U23437 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20513) );
  OAI222_X1 U23438 ( .A1(n20457), .A2(n20483), .B1(n20513), .B2(n20475), .C1(
        n20500), .C2(n20456), .ZN(P2_U2906) );
  INV_X1 U23439 ( .A(n20458), .ZN(n20460) );
  INV_X1 U23440 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20515) );
  OAI222_X1 U23441 ( .A1(n20460), .A2(n20483), .B1(n20515), .B2(n20475), .C1(
        n20500), .C2(n20459), .ZN(P2_U2907) );
  INV_X1 U23442 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20517) );
  OAI222_X1 U23443 ( .A1(n20462), .A2(n20483), .B1(n20517), .B2(n20475), .C1(
        n20500), .C2(n20461), .ZN(P2_U2908) );
  AOI22_X1 U23444 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n20491), .B1(n20463), 
        .B2(n20468), .ZN(n20464) );
  OAI21_X1 U23445 ( .B1(n20483), .B2(n20465), .A(n20464), .ZN(P2_U2909) );
  OAI222_X1 U23446 ( .A1(n20467), .A2(n20483), .B1(n20521), .B2(n20475), .C1(
        n20500), .C2(n20466), .ZN(P2_U2910) );
  AOI22_X1 U23447 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n20491), .B1(n20469), .B2(
        n20468), .ZN(n20470) );
  OAI21_X1 U23448 ( .B1(n20483), .B2(n20471), .A(n20470), .ZN(P2_U2911) );
  OAI222_X1 U23449 ( .A1(n20472), .A2(n20483), .B1(n20525), .B2(n20475), .C1(
        n20500), .C2(n20576), .ZN(P2_U2912) );
  INV_X1 U23450 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20527) );
  OAI222_X1 U23451 ( .A1(n20474), .A2(n20483), .B1(n20527), .B2(n20475), .C1(
        n20500), .C2(n20473), .ZN(P2_U2913) );
  INV_X1 U23452 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n20529) );
  OAI22_X1 U23453 ( .A1(n20529), .A2(n20475), .B1(n20566), .B2(n20500), .ZN(
        n20476) );
  INV_X1 U23454 ( .A(n20476), .ZN(n20481) );
  NAND3_X1 U23455 ( .A1(n20479), .A2(n20478), .A3(n20477), .ZN(n20480) );
  OAI211_X1 U23456 ( .C1(n20483), .C2(n20482), .A(n20481), .B(n20480), .ZN(
        P2_U2914) );
  AOI22_X1 U23457 ( .A1(n20484), .A2(n20492), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20491), .ZN(n20490) );
  AOI21_X1 U23458 ( .B1(n20487), .B2(n20486), .A(n20485), .ZN(n20488) );
  OR2_X1 U23459 ( .A1(n20488), .A2(n20496), .ZN(n20489) );
  OAI211_X1 U23460 ( .C1(n20558), .C2(n20500), .A(n20490), .B(n20489), .ZN(
        P2_U2916) );
  AOI22_X1 U23461 ( .A1(n20492), .A2(n21201), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n20491), .ZN(n20499) );
  AOI21_X1 U23462 ( .B1(n20495), .B2(n20494), .A(n20493), .ZN(n20497) );
  OR2_X1 U23463 ( .A1(n20497), .A2(n20496), .ZN(n20498) );
  OAI211_X1 U23464 ( .C1(n20548), .C2(n20500), .A(n20499), .B(n20498), .ZN(
        P2_U2918) );
  NOR2_X1 U23465 ( .A1(n20534), .A2(n20501), .ZN(P2_U2920) );
  INV_X1 U23466 ( .A(n20502), .ZN(n20505) );
  AOI22_X1 U23467 ( .A1(n20505), .A2(P2_EAX_REG_22__SCAN_IN), .B1(
        P2_UWORD_REG_6__SCAN_IN), .B2(n20541), .ZN(n20503) );
  OAI21_X1 U23468 ( .B1(n20504), .B2(n20534), .A(n20503), .ZN(P2_U2929) );
  AOI22_X1 U23469 ( .A1(n20540), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(n20505), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n20506) );
  OAI21_X1 U23470 ( .B1(n20508), .B2(n20507), .A(n20506), .ZN(P2_U2931) );
  AOI22_X1 U23471 ( .A1(n20541), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n20509) );
  OAI21_X1 U23472 ( .B1(n13921), .B2(n20543), .A(n20509), .ZN(P2_U2936) );
  AOI22_X1 U23473 ( .A1(n20541), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n20510) );
  OAI21_X1 U23474 ( .B1(n20511), .B2(n20543), .A(n20510), .ZN(P2_U2937) );
  AOI22_X1 U23475 ( .A1(n20541), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n20512) );
  OAI21_X1 U23476 ( .B1(n20513), .B2(n20543), .A(n20512), .ZN(P2_U2938) );
  AOI22_X1 U23477 ( .A1(n20541), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n20514) );
  OAI21_X1 U23478 ( .B1(n20515), .B2(n20543), .A(n20514), .ZN(P2_U2939) );
  AOI22_X1 U23479 ( .A1(n20541), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n20516) );
  OAI21_X1 U23480 ( .B1(n20517), .B2(n20543), .A(n20516), .ZN(P2_U2940) );
  AOI22_X1 U23481 ( .A1(n20541), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n20518) );
  OAI21_X1 U23482 ( .B1(n20519), .B2(n20543), .A(n20518), .ZN(P2_U2941) );
  AOI22_X1 U23483 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n20541), .B1(n20540), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n20520) );
  OAI21_X1 U23484 ( .B1(n20521), .B2(n20543), .A(n20520), .ZN(P2_U2942) );
  AOI22_X1 U23485 ( .A1(n20541), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n20522) );
  OAI21_X1 U23486 ( .B1(n20523), .B2(n20543), .A(n20522), .ZN(P2_U2943) );
  AOI22_X1 U23487 ( .A1(n20541), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n20524) );
  OAI21_X1 U23488 ( .B1(n20525), .B2(n20543), .A(n20524), .ZN(P2_U2944) );
  AOI22_X1 U23489 ( .A1(n20541), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n20526) );
  OAI21_X1 U23490 ( .B1(n20527), .B2(n20543), .A(n20526), .ZN(P2_U2945) );
  AOI22_X1 U23491 ( .A1(n20541), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n20528) );
  OAI21_X1 U23492 ( .B1(n20529), .B2(n20543), .A(n20528), .ZN(P2_U2946) );
  AOI22_X1 U23493 ( .A1(P2_EAX_REG_4__SCAN_IN), .A2(n20532), .B1(n20541), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n20530) );
  OAI21_X1 U23494 ( .B1(n20531), .B2(n20534), .A(n20530), .ZN(P2_U2947) );
  AOI22_X1 U23495 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n20532), .B1(n20541), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n20533) );
  OAI21_X1 U23496 ( .B1(n20535), .B2(n20534), .A(n20533), .ZN(P2_U2948) );
  INV_X1 U23497 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20537) );
  AOI22_X1 U23498 ( .A1(n20541), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n20536) );
  OAI21_X1 U23499 ( .B1(n20537), .B2(n20543), .A(n20536), .ZN(P2_U2949) );
  AOI22_X1 U23500 ( .A1(n20541), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n20538) );
  OAI21_X1 U23501 ( .B1(n20539), .B2(n20543), .A(n20538), .ZN(P2_U2950) );
  AOI22_X1 U23502 ( .A1(n20541), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n20540), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n20542) );
  OAI21_X1 U23503 ( .B1(n13916), .B2(n20543), .A(n20542), .ZN(P2_U2951) );
  AOI22_X1 U23504 ( .A1(n20944), .A2(n21075), .B1(n21020), .B2(n20575), .ZN(
        n20545) );
  AOI22_X1 U23505 ( .A1(n21021), .A2(n20581), .B1(n20607), .B2(n21030), .ZN(
        n20544) );
  OAI211_X1 U23506 ( .C1(n20585), .C2(n20546), .A(n20545), .B(n20544), .ZN(
        P2_U3048) );
  AOI22_X1 U23507 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20572), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20571), .ZN(n21039) );
  INV_X1 U23508 ( .A(n21039), .ZN(n20985) );
  NOR2_X2 U23509 ( .A1(n20574), .A2(n20547), .ZN(n21034) );
  AOI22_X1 U23510 ( .A1(n20985), .A2(n21075), .B1(n20575), .B2(n21034), .ZN(
        n20552) );
  NOR2_X2 U23511 ( .A1(n20548), .A2(n20977), .ZN(n21035) );
  OAI22_X2 U23512 ( .A1(n20550), .A2(n20579), .B1(n20549), .B2(n20577), .ZN(
        n21036) );
  AOI22_X1 U23513 ( .A1(n21035), .A2(n20581), .B1(n20607), .B2(n21036), .ZN(
        n20551) );
  OAI211_X1 U23514 ( .C1(n20585), .C2(n12919), .A(n20552), .B(n20551), .ZN(
        P2_U3049) );
  AOI22_X1 U23515 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20572), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20571), .ZN(n21045) );
  INV_X1 U23516 ( .A(n21045), .ZN(n20989) );
  NOR2_X2 U23517 ( .A1(n20574), .A2(n11482), .ZN(n21040) );
  AOI22_X1 U23518 ( .A1(n20989), .A2(n21075), .B1(n20575), .B2(n21040), .ZN(
        n20557) );
  INV_X1 U23519 ( .A(n20553), .ZN(n20554) );
  NOR2_X2 U23520 ( .A1(n20554), .A2(n20977), .ZN(n21041) );
  AOI22_X1 U23521 ( .A1(n21041), .A2(n20581), .B1(n20607), .B2(n21042), .ZN(
        n20556) );
  OAI211_X1 U23522 ( .C1(n20585), .C2(n12912), .A(n20557), .B(n20556), .ZN(
        P2_U3050) );
  AOI22_X1 U23523 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20571), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20572), .ZN(n21051) );
  INV_X1 U23524 ( .A(n21051), .ZN(n20993) );
  AOI22_X1 U23525 ( .A1(n20993), .A2(n21075), .B1(n20575), .B2(n9786), .ZN(
        n20560) );
  NOR2_X2 U23526 ( .A1(n20558), .A2(n20977), .ZN(n21047) );
  AOI22_X1 U23527 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20572), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20571), .ZN(n20996) );
  AOI22_X1 U23528 ( .A1(n21047), .A2(n20581), .B1(n20607), .B2(n21048), .ZN(
        n20559) );
  OAI211_X1 U23529 ( .C1(n20585), .C2(n12899), .A(n20560), .B(n20559), .ZN(
        P2_U3051) );
  INV_X1 U23530 ( .A(n21057), .ZN(n20954) );
  NOR2_X2 U23531 ( .A1(n20574), .A2(n12215), .ZN(n21052) );
  AOI22_X1 U23532 ( .A1(n20954), .A2(n21075), .B1(n20575), .B2(n21052), .ZN(
        n20564) );
  NOR2_X2 U23533 ( .A1(n20561), .A2(n20977), .ZN(n21053) );
  OAI22_X2 U23534 ( .A1(n15700), .A2(n20579), .B1(n20562), .B2(n20577), .ZN(
        n21054) );
  AOI22_X1 U23535 ( .A1(n21053), .A2(n20581), .B1(n20607), .B2(n21054), .ZN(
        n20563) );
  OAI211_X1 U23536 ( .C1(n20585), .C2(n12931), .A(n20564), .B(n20563), .ZN(
        P2_U3052) );
  AOI22_X1 U23537 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20572), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20571), .ZN(n21063) );
  INV_X1 U23538 ( .A(n21063), .ZN(n20958) );
  NOR2_X2 U23539 ( .A1(n20574), .A2(n20565), .ZN(n21058) );
  AOI22_X1 U23540 ( .A1(n20958), .A2(n21075), .B1(n20575), .B2(n21058), .ZN(
        n20570) );
  NOR2_X2 U23541 ( .A1(n20566), .A2(n20977), .ZN(n21059) );
  OAI22_X2 U23542 ( .A1(n20568), .A2(n20579), .B1(n20567), .B2(n20577), .ZN(
        n21060) );
  AOI22_X1 U23543 ( .A1(n21059), .A2(n20581), .B1(n20607), .B2(n21060), .ZN(
        n20569) );
  OAI211_X1 U23544 ( .C1(n20585), .C2(n13946), .A(n20570), .B(n20569), .ZN(
        P2_U3053) );
  INV_X1 U23545 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20584) );
  AOI22_X1 U23546 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20572), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20571), .ZN(n21080) );
  INV_X1 U23547 ( .A(n21080), .ZN(n21009) );
  NOR2_X2 U23548 ( .A1(n20574), .A2(n20573), .ZN(n21070) );
  AOI22_X1 U23549 ( .A1(n21009), .A2(n21075), .B1(n20575), .B2(n21070), .ZN(
        n20583) );
  NOR2_X2 U23550 ( .A1(n20576), .A2(n20977), .ZN(n21072) );
  OAI22_X2 U23551 ( .A1(n20580), .A2(n20579), .B1(n20578), .B2(n20577), .ZN(
        n21074) );
  AOI22_X1 U23552 ( .A1(n21072), .A2(n20581), .B1(n20607), .B2(n21074), .ZN(
        n20582) );
  OAI211_X1 U23553 ( .C1(n20585), .C2(n20584), .A(n20583), .B(n20582), .ZN(
        P2_U3055) );
  INV_X1 U23554 ( .A(n20607), .ZN(n20615) );
  NOR2_X1 U23555 ( .A1(n20797), .A2(n20619), .ZN(n20610) );
  INV_X1 U23556 ( .A(n20610), .ZN(n20586) );
  AND3_X1 U23557 ( .A1(n20587), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20586), 
        .ZN(n20590) );
  AOI211_X2 U23558 ( .C1(n20591), .C2(n21225), .A(n20588), .B(n20590), .ZN(
        n20611) );
  AOI22_X1 U23559 ( .A1(n20611), .A2(n21021), .B1(n21020), .B2(n20610), .ZN(
        n20596) );
  INV_X1 U23560 ( .A(n20700), .ZN(n20589) );
  NAND2_X1 U23561 ( .A1(n20589), .A2(n20810), .ZN(n20592) );
  AOI21_X1 U23562 ( .B1(n20592), .B2(n20591), .A(n20590), .ZN(n20593) );
  OAI211_X1 U23563 ( .C1(n20610), .C2(n20975), .A(n21023), .B(n20593), .ZN(
        n20612) );
  AOI22_X1 U23564 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20612), .B1(
        n20621), .B2(n21030), .ZN(n20595) );
  OAI211_X1 U23565 ( .C1(n21033), .C2(n20615), .A(n20596), .B(n20595), .ZN(
        P2_U3056) );
  AOI22_X1 U23566 ( .A1(n20611), .A2(n21035), .B1(n21034), .B2(n20610), .ZN(
        n20598) );
  AOI22_X1 U23567 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20612), .B1(
        n20621), .B2(n21036), .ZN(n20597) );
  OAI211_X1 U23568 ( .C1(n21039), .C2(n20615), .A(n20598), .B(n20597), .ZN(
        P2_U3057) );
  AOI22_X1 U23569 ( .A1(n20611), .A2(n21041), .B1(n21040), .B2(n20610), .ZN(
        n20600) );
  AOI22_X1 U23570 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20612), .B1(
        n20607), .B2(n20989), .ZN(n20599) );
  OAI211_X1 U23571 ( .C1(n20992), .C2(n20645), .A(n20600), .B(n20599), .ZN(
        P2_U3058) );
  AOI22_X1 U23572 ( .A1(n20611), .A2(n21047), .B1(n9786), .B2(n20610), .ZN(
        n20602) );
  AOI22_X1 U23573 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20612), .B1(
        n20607), .B2(n20993), .ZN(n20601) );
  OAI211_X1 U23574 ( .C1(n20996), .C2(n20645), .A(n20602), .B(n20601), .ZN(
        P2_U3059) );
  AOI22_X1 U23575 ( .A1(n20611), .A2(n21053), .B1(n21052), .B2(n20610), .ZN(
        n20604) );
  AOI22_X1 U23576 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20612), .B1(
        n20621), .B2(n21054), .ZN(n20603) );
  OAI211_X1 U23577 ( .C1(n21057), .C2(n20615), .A(n20604), .B(n20603), .ZN(
        P2_U3060) );
  AOI22_X1 U23578 ( .A1(n20611), .A2(n21059), .B1(n21058), .B2(n20610), .ZN(
        n20606) );
  AOI22_X1 U23579 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20612), .B1(
        n20621), .B2(n21060), .ZN(n20605) );
  OAI211_X1 U23580 ( .C1(n21063), .C2(n20615), .A(n20606), .B(n20605), .ZN(
        P2_U3061) );
  AOI22_X1 U23581 ( .A1(n20611), .A2(n21065), .B1(n21064), .B2(n20610), .ZN(
        n20609) );
  AOI22_X1 U23582 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20612), .B1(
        n20607), .B2(n21003), .ZN(n20608) );
  OAI211_X1 U23583 ( .C1(n21006), .C2(n20645), .A(n20609), .B(n20608), .ZN(
        P2_U3062) );
  AOI22_X1 U23584 ( .A1(n20611), .A2(n21072), .B1(n21070), .B2(n20610), .ZN(
        n20614) );
  AOI22_X1 U23585 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20612), .B1(
        n20621), .B2(n21074), .ZN(n20613) );
  OAI211_X1 U23586 ( .C1(n21080), .C2(n20615), .A(n20614), .B(n20613), .ZN(
        P2_U3063) );
  NOR2_X1 U23587 ( .A1(n20833), .A2(n20619), .ZN(n20640) );
  INV_X1 U23588 ( .A(n20640), .ZN(n20616) );
  NAND2_X1 U23589 ( .A1(n20617), .A2(n20616), .ZN(n20623) );
  INV_X1 U23590 ( .A(n20623), .ZN(n20618) );
  OAI22_X1 U23591 ( .A1(n20618), .A2(n21225), .B1(n20619), .B2(n20836), .ZN(
        n20641) );
  AOI22_X1 U23592 ( .A1(n20641), .A2(n21021), .B1(n21020), .B2(n20640), .ZN(
        n20627) );
  NOR2_X1 U23593 ( .A1(n20836), .A2(n20619), .ZN(n20620) );
  AOI221_X1 U23594 ( .B1(n20661), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20621), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n20620), .ZN(n20622) );
  NAND2_X1 U23595 ( .A1(n20622), .A2(n20975), .ZN(n20624) );
  MUX2_X1 U23596 ( .A(n20624), .B(n20623), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n20625) );
  OAI211_X1 U23597 ( .C1(n20640), .C2(n20975), .A(n21023), .B(n20625), .ZN(
        n20642) );
  AOI22_X1 U23598 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20642), .B1(
        n20661), .B2(n21030), .ZN(n20626) );
  OAI211_X1 U23599 ( .C1(n21033), .C2(n20645), .A(n20627), .B(n20626), .ZN(
        P2_U3064) );
  AOI22_X1 U23600 ( .A1(n20641), .A2(n21035), .B1(n21034), .B2(n20640), .ZN(
        n20629) );
  AOI22_X1 U23601 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20642), .B1(
        n20661), .B2(n21036), .ZN(n20628) );
  OAI211_X1 U23602 ( .C1(n21039), .C2(n20645), .A(n20629), .B(n20628), .ZN(
        P2_U3065) );
  AOI22_X1 U23603 ( .A1(n20641), .A2(n21041), .B1(n21040), .B2(n20640), .ZN(
        n20631) );
  AOI22_X1 U23604 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20642), .B1(
        n20661), .B2(n21042), .ZN(n20630) );
  OAI211_X1 U23605 ( .C1(n21045), .C2(n20645), .A(n20631), .B(n20630), .ZN(
        P2_U3066) );
  AOI22_X1 U23606 ( .A1(n20641), .A2(n21047), .B1(n9786), .B2(n20640), .ZN(
        n20633) );
  AOI22_X1 U23607 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20642), .B1(
        n20661), .B2(n21048), .ZN(n20632) );
  OAI211_X1 U23608 ( .C1(n21051), .C2(n20645), .A(n20633), .B(n20632), .ZN(
        P2_U3067) );
  AOI22_X1 U23609 ( .A1(n20641), .A2(n21053), .B1(n21052), .B2(n20640), .ZN(
        n20635) );
  AOI22_X1 U23610 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20642), .B1(
        n20661), .B2(n21054), .ZN(n20634) );
  OAI211_X1 U23611 ( .C1(n21057), .C2(n20645), .A(n20635), .B(n20634), .ZN(
        P2_U3068) );
  AOI22_X1 U23612 ( .A1(n20641), .A2(n21059), .B1(n21058), .B2(n20640), .ZN(
        n20637) );
  AOI22_X1 U23613 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20642), .B1(
        n20661), .B2(n21060), .ZN(n20636) );
  OAI211_X1 U23614 ( .C1(n21063), .C2(n20645), .A(n20637), .B(n20636), .ZN(
        P2_U3069) );
  AOI22_X1 U23615 ( .A1(n20641), .A2(n21065), .B1(n21064), .B2(n20640), .ZN(
        n20639) );
  AOI22_X1 U23616 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20642), .B1(
        n20661), .B2(n21066), .ZN(n20638) );
  OAI211_X1 U23617 ( .C1(n21069), .C2(n20645), .A(n20639), .B(n20638), .ZN(
        P2_U3070) );
  AOI22_X1 U23618 ( .A1(n20641), .A2(n21072), .B1(n21070), .B2(n20640), .ZN(
        n20644) );
  AOI22_X1 U23619 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20642), .B1(
        n20661), .B2(n21074), .ZN(n20643) );
  OAI211_X1 U23620 ( .C1(n21080), .C2(n20645), .A(n20644), .B(n20643), .ZN(
        P2_U3071) );
  AOI22_X1 U23621 ( .A1(n20985), .A2(n20661), .B1(n20660), .B2(n21034), .ZN(
        n20647) );
  AOI22_X1 U23622 ( .A1(n21035), .A2(n20662), .B1(n20690), .B2(n21036), .ZN(
        n20646) );
  OAI211_X1 U23623 ( .C1(n20666), .C2(n11619), .A(n20647), .B(n20646), .ZN(
        P2_U3073) );
  INV_X1 U23624 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n20650) );
  AOI22_X1 U23625 ( .A1(n20989), .A2(n20661), .B1(n20660), .B2(n21040), .ZN(
        n20649) );
  AOI22_X1 U23626 ( .A1(n21041), .A2(n20662), .B1(n20690), .B2(n21042), .ZN(
        n20648) );
  OAI211_X1 U23627 ( .C1(n20666), .C2(n20650), .A(n20649), .B(n20648), .ZN(
        P2_U3074) );
  AOI22_X1 U23628 ( .A1(n20993), .A2(n20661), .B1(n20660), .B2(n9786), .ZN(
        n20652) );
  AOI22_X1 U23629 ( .A1(n21047), .A2(n20662), .B1(n20690), .B2(n21048), .ZN(
        n20651) );
  OAI211_X1 U23630 ( .C1(n20666), .C2(n11567), .A(n20652), .B(n20651), .ZN(
        P2_U3075) );
  INV_X1 U23631 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n20655) );
  AOI22_X1 U23632 ( .A1(n20954), .A2(n20661), .B1(n20660), .B2(n21052), .ZN(
        n20654) );
  AOI22_X1 U23633 ( .A1(n21053), .A2(n20662), .B1(n20690), .B2(n21054), .ZN(
        n20653) );
  OAI211_X1 U23634 ( .C1(n20666), .C2(n20655), .A(n20654), .B(n20653), .ZN(
        P2_U3076) );
  AOI22_X1 U23635 ( .A1(n20958), .A2(n20661), .B1(n20660), .B2(n21058), .ZN(
        n20657) );
  AOI22_X1 U23636 ( .A1(n21059), .A2(n20662), .B1(n20690), .B2(n21060), .ZN(
        n20656) );
  OAI211_X1 U23637 ( .C1(n20666), .C2(n11707), .A(n20657), .B(n20656), .ZN(
        P2_U3077) );
  AOI22_X1 U23638 ( .A1(n21003), .A2(n20661), .B1(n21064), .B2(n20660), .ZN(
        n20659) );
  AOI22_X1 U23639 ( .A1(n21065), .A2(n20662), .B1(n20690), .B2(n21066), .ZN(
        n20658) );
  OAI211_X1 U23640 ( .C1(n20666), .C2(n11825), .A(n20659), .B(n20658), .ZN(
        P2_U3078) );
  AOI22_X1 U23641 ( .A1(n21074), .A2(n20690), .B1(n20660), .B2(n21070), .ZN(
        n20664) );
  AOI22_X1 U23642 ( .A1(n21072), .A2(n20662), .B1(n20661), .B2(n21009), .ZN(
        n20663) );
  OAI211_X1 U23643 ( .C1(n20666), .C2(n20665), .A(n20664), .B(n20663), .ZN(
        P2_U3079) );
  INV_X1 U23644 ( .A(n21177), .ZN(n20908) );
  INV_X1 U23645 ( .A(n20667), .ZN(n20668) );
  NAND2_X1 U23646 ( .A1(n20669), .A2(n20668), .ZN(n20906) );
  NOR2_X1 U23647 ( .A1(n20906), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20677) );
  INV_X1 U23648 ( .A(n20677), .ZN(n20671) );
  NOR2_X1 U23649 ( .A1(n20699), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20702) );
  INV_X1 U23650 ( .A(n20702), .ZN(n20705) );
  NOR2_X1 U23651 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20705), .ZN(
        n20693) );
  OAI21_X1 U23652 ( .B1(n11723), .B2(n20693), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20670) );
  OAI21_X1 U23653 ( .B1(n20908), .B2(n20671), .A(n20670), .ZN(n20694) );
  AOI22_X1 U23654 ( .A1(n20694), .A2(n21021), .B1(n21020), .B2(n20693), .ZN(
        n20679) );
  AOI21_X1 U23655 ( .B1(n20698), .B2(n20718), .A(n12132), .ZN(n20676) );
  OAI21_X1 U23656 ( .B1(n11723), .B2(n21225), .A(n20975), .ZN(n20674) );
  INV_X1 U23657 ( .A(n20693), .ZN(n20673) );
  NAND2_X1 U23658 ( .A1(n20674), .A2(n20673), .ZN(n20675) );
  OAI211_X1 U23659 ( .C1(n20677), .C2(n20676), .A(n20675), .B(n21023), .ZN(
        n20695) );
  AOI22_X1 U23660 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20695), .B1(
        n20724), .B2(n21030), .ZN(n20678) );
  OAI211_X1 U23661 ( .C1(n21033), .C2(n20698), .A(n20679), .B(n20678), .ZN(
        P2_U3080) );
  INV_X1 U23662 ( .A(n21036), .ZN(n20988) );
  AOI22_X1 U23663 ( .A1(n20694), .A2(n21035), .B1(n21034), .B2(n20693), .ZN(
        n20681) );
  AOI22_X1 U23664 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20695), .B1(
        n20690), .B2(n20985), .ZN(n20680) );
  OAI211_X1 U23665 ( .C1(n20988), .C2(n20718), .A(n20681), .B(n20680), .ZN(
        P2_U3081) );
  AOI22_X1 U23666 ( .A1(n20694), .A2(n21041), .B1(n21040), .B2(n20693), .ZN(
        n20683) );
  AOI22_X1 U23667 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20695), .B1(
        n20690), .B2(n20989), .ZN(n20682) );
  OAI211_X1 U23668 ( .C1(n20992), .C2(n20718), .A(n20683), .B(n20682), .ZN(
        P2_U3082) );
  AOI22_X1 U23669 ( .A1(n20694), .A2(n21047), .B1(n9786), .B2(n20693), .ZN(
        n20685) );
  AOI22_X1 U23670 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20695), .B1(
        n20724), .B2(n21048), .ZN(n20684) );
  OAI211_X1 U23671 ( .C1(n21051), .C2(n20698), .A(n20685), .B(n20684), .ZN(
        P2_U3083) );
  AOI22_X1 U23672 ( .A1(n20694), .A2(n21053), .B1(n21052), .B2(n20693), .ZN(
        n20687) );
  AOI22_X1 U23673 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20695), .B1(
        n20724), .B2(n21054), .ZN(n20686) );
  OAI211_X1 U23674 ( .C1(n21057), .C2(n20698), .A(n20687), .B(n20686), .ZN(
        P2_U3084) );
  AOI22_X1 U23675 ( .A1(n20694), .A2(n21059), .B1(n21058), .B2(n20693), .ZN(
        n20689) );
  AOI22_X1 U23676 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20695), .B1(
        n20724), .B2(n21060), .ZN(n20688) );
  OAI211_X1 U23677 ( .C1(n21063), .C2(n20698), .A(n20689), .B(n20688), .ZN(
        P2_U3085) );
  AOI22_X1 U23678 ( .A1(n20694), .A2(n21065), .B1(n21064), .B2(n20693), .ZN(
        n20692) );
  AOI22_X1 U23679 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20695), .B1(
        n20690), .B2(n21003), .ZN(n20691) );
  OAI211_X1 U23680 ( .C1(n21006), .C2(n20718), .A(n20692), .B(n20691), .ZN(
        P2_U3086) );
  AOI22_X1 U23681 ( .A1(n20694), .A2(n21072), .B1(n21070), .B2(n20693), .ZN(
        n20697) );
  AOI22_X1 U23682 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20695), .B1(
        n20724), .B2(n21074), .ZN(n20696) );
  OAI211_X1 U23683 ( .C1(n21080), .C2(n20698), .A(n20697), .B(n20696), .ZN(
        P2_U3087) );
  NOR2_X1 U23684 ( .A1(n20797), .A2(n20699), .ZN(n20723) );
  AOI22_X1 U23685 ( .A1(n21030), .A2(n20715), .B1(n21020), .B2(n20723), .ZN(
        n20708) );
  OAI21_X1 U23686 ( .B1(n20700), .B2(n20931), .A(n21177), .ZN(n20706) );
  OAI211_X1 U23687 ( .C1(n20706), .C2(n20702), .A(n21023), .B(n20701), .ZN(
        n20726) );
  OAI21_X1 U23688 ( .B1(n20703), .B2(n20723), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20704) );
  OAI21_X1 U23689 ( .B1(n20706), .B2(n20705), .A(n20704), .ZN(n20725) );
  AOI22_X1 U23690 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20726), .B1(
        n21021), .B2(n20725), .ZN(n20707) );
  OAI211_X1 U23691 ( .C1(n21033), .C2(n20718), .A(n20708), .B(n20707), .ZN(
        P2_U3088) );
  AOI22_X1 U23692 ( .A1(n20985), .A2(n20724), .B1(n20723), .B2(n21034), .ZN(
        n20710) );
  AOI22_X1 U23693 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20726), .B1(
        n21035), .B2(n20725), .ZN(n20709) );
  OAI211_X1 U23694 ( .C1(n20988), .C2(n20747), .A(n20710), .B(n20709), .ZN(
        P2_U3089) );
  AOI22_X1 U23695 ( .A1(n21042), .A2(n20715), .B1(n21040), .B2(n20723), .ZN(
        n20712) );
  AOI22_X1 U23696 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20726), .B1(
        n21041), .B2(n20725), .ZN(n20711) );
  OAI211_X1 U23697 ( .C1(n21045), .C2(n20718), .A(n20712), .B(n20711), .ZN(
        P2_U3090) );
  AOI22_X1 U23698 ( .A1(n21048), .A2(n20715), .B1(n20723), .B2(n9786), .ZN(
        n20714) );
  AOI22_X1 U23699 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20726), .B1(
        n21047), .B2(n20725), .ZN(n20713) );
  OAI211_X1 U23700 ( .C1(n21051), .C2(n20718), .A(n20714), .B(n20713), .ZN(
        P2_U3091) );
  AOI22_X1 U23701 ( .A1(n21054), .A2(n20715), .B1(n20723), .B2(n21052), .ZN(
        n20717) );
  AOI22_X1 U23702 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20726), .B1(
        n21053), .B2(n20725), .ZN(n20716) );
  OAI211_X1 U23703 ( .C1(n21057), .C2(n20718), .A(n20717), .B(n20716), .ZN(
        P2_U3092) );
  INV_X1 U23704 ( .A(n21060), .ZN(n20961) );
  AOI22_X1 U23705 ( .A1(n20958), .A2(n20724), .B1(n20723), .B2(n21058), .ZN(
        n20720) );
  AOI22_X1 U23706 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20726), .B1(
        n21059), .B2(n20725), .ZN(n20719) );
  OAI211_X1 U23707 ( .C1(n20961), .C2(n20747), .A(n20720), .B(n20719), .ZN(
        P2_U3093) );
  AOI22_X1 U23708 ( .A1(n21003), .A2(n20724), .B1(n21064), .B2(n20723), .ZN(
        n20722) );
  AOI22_X1 U23709 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20726), .B1(
        n21065), .B2(n20725), .ZN(n20721) );
  OAI211_X1 U23710 ( .C1(n21006), .C2(n20747), .A(n20722), .B(n20721), .ZN(
        P2_U3094) );
  INV_X1 U23711 ( .A(n21074), .ZN(n21014) );
  AOI22_X1 U23712 ( .A1(n21009), .A2(n20724), .B1(n20723), .B2(n21070), .ZN(
        n20728) );
  AOI22_X1 U23713 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20726), .B1(
        n21072), .B2(n20725), .ZN(n20727) );
  OAI211_X1 U23714 ( .C1(n21014), .C2(n20747), .A(n20728), .B(n20727), .ZN(
        P2_U3095) );
  AOI22_X1 U23715 ( .A1(n20743), .A2(n21035), .B1(n20742), .B2(n21034), .ZN(
        n20731) );
  AOI22_X1 U23716 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20744), .B1(
        n20764), .B2(n21036), .ZN(n20730) );
  OAI211_X1 U23717 ( .C1(n21039), .C2(n20747), .A(n20731), .B(n20730), .ZN(
        P2_U3097) );
  AOI22_X1 U23718 ( .A1(n20743), .A2(n21041), .B1(n20742), .B2(n21040), .ZN(
        n20733) );
  AOI22_X1 U23719 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20744), .B1(
        n20764), .B2(n21042), .ZN(n20732) );
  OAI211_X1 U23720 ( .C1(n21045), .C2(n20747), .A(n20733), .B(n20732), .ZN(
        P2_U3098) );
  AOI22_X1 U23721 ( .A1(n20743), .A2(n21047), .B1(n20742), .B2(n9786), .ZN(
        n20735) );
  AOI22_X1 U23722 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20744), .B1(
        n20764), .B2(n21048), .ZN(n20734) );
  OAI211_X1 U23723 ( .C1(n21051), .C2(n20747), .A(n20735), .B(n20734), .ZN(
        P2_U3099) );
  AOI22_X1 U23724 ( .A1(n20743), .A2(n21053), .B1(n20742), .B2(n21052), .ZN(
        n20737) );
  AOI22_X1 U23725 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20744), .B1(
        n20764), .B2(n21054), .ZN(n20736) );
  OAI211_X1 U23726 ( .C1(n21057), .C2(n20747), .A(n20737), .B(n20736), .ZN(
        P2_U3100) );
  AOI22_X1 U23727 ( .A1(n20743), .A2(n21059), .B1(n20742), .B2(n21058), .ZN(
        n20739) );
  AOI22_X1 U23728 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20744), .B1(
        n20764), .B2(n21060), .ZN(n20738) );
  OAI211_X1 U23729 ( .C1(n21063), .C2(n20747), .A(n20739), .B(n20738), .ZN(
        P2_U3101) );
  AOI22_X1 U23730 ( .A1(n20743), .A2(n21065), .B1(n20742), .B2(n21064), .ZN(
        n20741) );
  AOI22_X1 U23731 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20744), .B1(
        n20764), .B2(n21066), .ZN(n20740) );
  OAI211_X1 U23732 ( .C1(n21069), .C2(n20747), .A(n20741), .B(n20740), .ZN(
        P2_U3102) );
  AOI22_X1 U23733 ( .A1(n20743), .A2(n21072), .B1(n20742), .B2(n21070), .ZN(
        n20746) );
  AOI22_X1 U23734 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20744), .B1(
        n20764), .B2(n21074), .ZN(n20745) );
  OAI211_X1 U23735 ( .C1(n21080), .C2(n20747), .A(n20746), .B(n20745), .ZN(
        P2_U3103) );
  AOI22_X1 U23736 ( .A1(n20763), .A2(n21021), .B1(n21020), .B2(n20774), .ZN(
        n20749) );
  AOI22_X1 U23737 ( .A1(n20759), .A2(n21030), .B1(n20764), .B2(n20944), .ZN(
        n20748) );
  OAI211_X1 U23738 ( .C1(n20762), .C2(n20750), .A(n20749), .B(n20748), .ZN(
        P2_U3104) );
  AOI22_X1 U23739 ( .A1(n20763), .A2(n21035), .B1(n20774), .B2(n21034), .ZN(
        n20752) );
  AOI22_X1 U23740 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20765), .B1(
        n20764), .B2(n20985), .ZN(n20751) );
  OAI211_X1 U23741 ( .C1(n20988), .C2(n20796), .A(n20752), .B(n20751), .ZN(
        P2_U3105) );
  AOI22_X1 U23742 ( .A1(n20763), .A2(n21041), .B1(n20774), .B2(n21040), .ZN(
        n20754) );
  AOI22_X1 U23743 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20765), .B1(
        n20764), .B2(n20989), .ZN(n20753) );
  OAI211_X1 U23744 ( .C1(n20992), .C2(n20796), .A(n20754), .B(n20753), .ZN(
        P2_U3106) );
  AOI22_X1 U23745 ( .A1(n20763), .A2(n21047), .B1(n20774), .B2(n9786), .ZN(
        n20756) );
  AOI22_X1 U23746 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20765), .B1(
        n20764), .B2(n20993), .ZN(n20755) );
  OAI211_X1 U23747 ( .C1(n20996), .C2(n20796), .A(n20756), .B(n20755), .ZN(
        P2_U3107) );
  AOI22_X1 U23748 ( .A1(n20763), .A2(n21053), .B1(n20774), .B2(n21052), .ZN(
        n20758) );
  AOI22_X1 U23749 ( .A1(n20759), .A2(n21054), .B1(n20764), .B2(n20954), .ZN(
        n20757) );
  OAI211_X1 U23750 ( .C1(n20762), .C2(n12996), .A(n20758), .B(n20757), .ZN(
        P2_U3108) );
  AOI22_X1 U23751 ( .A1(n20763), .A2(n21059), .B1(n20774), .B2(n21058), .ZN(
        n20761) );
  AOI22_X1 U23752 ( .A1(n20759), .A2(n21060), .B1(n20764), .B2(n20958), .ZN(
        n20760) );
  OAI211_X1 U23753 ( .C1(n20762), .C2(n11708), .A(n20761), .B(n20760), .ZN(
        P2_U3109) );
  AOI22_X1 U23754 ( .A1(n20763), .A2(n21072), .B1(n20774), .B2(n21070), .ZN(
        n20767) );
  AOI22_X1 U23755 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20765), .B1(
        n20764), .B2(n21009), .ZN(n20766) );
  OAI211_X1 U23756 ( .C1(n21014), .C2(n20796), .A(n20767), .B(n20766), .ZN(
        P2_U3111) );
  NOR2_X1 U23757 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n12896), .ZN(
        n20867) );
  NAND2_X1 U23758 ( .A1(n20867), .A2(n21203), .ZN(n20805) );
  NOR2_X1 U23759 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20805), .ZN(
        n20791) );
  AOI22_X1 U23760 ( .A1(n21030), .A2(n20828), .B1(n21020), .B2(n20791), .ZN(
        n20778) );
  NAND2_X1 U23761 ( .A1(n20825), .A2(n20796), .ZN(n20769) );
  AOI21_X1 U23762 ( .B1(n20769), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20908), 
        .ZN(n20773) );
  OAI21_X1 U23763 ( .B1(n11834), .B2(n21225), .A(n20975), .ZN(n20770) );
  AOI21_X1 U23764 ( .B1(n20773), .B2(n20771), .A(n20770), .ZN(n20772) );
  OAI21_X1 U23765 ( .B1(n20791), .B2(n20772), .A(n21023), .ZN(n20793) );
  OAI21_X1 U23766 ( .B1(n20774), .B2(n20791), .A(n20773), .ZN(n20776) );
  OAI21_X1 U23767 ( .B1(n11834), .B2(n20791), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20775) );
  NAND2_X1 U23768 ( .A1(n20776), .A2(n20775), .ZN(n20792) );
  AOI22_X1 U23769 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20793), .B1(
        n21021), .B2(n20792), .ZN(n20777) );
  OAI211_X1 U23770 ( .C1(n21033), .C2(n20796), .A(n20778), .B(n20777), .ZN(
        P2_U3112) );
  AOI22_X1 U23771 ( .A1(n21036), .A2(n20828), .B1(n20791), .B2(n21034), .ZN(
        n20780) );
  AOI22_X1 U23772 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21035), .ZN(n20779) );
  OAI211_X1 U23773 ( .C1(n21039), .C2(n20796), .A(n20780), .B(n20779), .ZN(
        P2_U3113) );
  AOI22_X1 U23774 ( .A1(n21042), .A2(n20828), .B1(n21040), .B2(n20791), .ZN(
        n20782) );
  AOI22_X1 U23775 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21041), .ZN(n20781) );
  OAI211_X1 U23776 ( .C1(n21045), .C2(n20796), .A(n20782), .B(n20781), .ZN(
        P2_U3114) );
  AOI22_X1 U23777 ( .A1(n21048), .A2(n20828), .B1(n20791), .B2(n9786), .ZN(
        n20784) );
  AOI22_X1 U23778 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21047), .ZN(n20783) );
  OAI211_X1 U23779 ( .C1(n21051), .C2(n20796), .A(n20784), .B(n20783), .ZN(
        P2_U3115) );
  AOI22_X1 U23780 ( .A1(n21054), .A2(n20828), .B1(n20791), .B2(n21052), .ZN(
        n20786) );
  AOI22_X1 U23781 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21053), .ZN(n20785) );
  OAI211_X1 U23782 ( .C1(n21057), .C2(n20796), .A(n20786), .B(n20785), .ZN(
        P2_U3116) );
  AOI22_X1 U23783 ( .A1(n21060), .A2(n20828), .B1(n20791), .B2(n21058), .ZN(
        n20788) );
  AOI22_X1 U23784 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21059), .ZN(n20787) );
  OAI211_X1 U23785 ( .C1(n21063), .C2(n20796), .A(n20788), .B(n20787), .ZN(
        P2_U3117) );
  AOI22_X1 U23786 ( .A1(n21066), .A2(n20828), .B1(n21064), .B2(n20791), .ZN(
        n20790) );
  AOI22_X1 U23787 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21065), .ZN(n20789) );
  OAI211_X1 U23788 ( .C1(n21069), .C2(n20796), .A(n20790), .B(n20789), .ZN(
        P2_U3118) );
  AOI22_X1 U23789 ( .A1(n21074), .A2(n20828), .B1(n20791), .B2(n21070), .ZN(
        n20795) );
  AOI22_X1 U23790 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20793), .B1(
        n20792), .B2(n21072), .ZN(n20794) );
  OAI211_X1 U23791 ( .C1(n21080), .C2(n20796), .A(n20795), .B(n20794), .ZN(
        P2_U3119) );
  NAND2_X1 U23792 ( .A1(n20807), .A2(n20975), .ZN(n20799) );
  INV_X1 U23793 ( .A(n20867), .ZN(n20837) );
  NOR2_X1 U23794 ( .A1(n20797), .A2(n20837), .ZN(n20839) );
  INV_X1 U23795 ( .A(n20839), .ZN(n20798) );
  NAND2_X1 U23796 ( .A1(n20799), .A2(n20798), .ZN(n20803) );
  NOR2_X1 U23797 ( .A1(n20800), .A2(n12132), .ZN(n21027) );
  NAND2_X1 U23798 ( .A1(n21027), .A2(n20810), .ZN(n20801) );
  NAND2_X1 U23799 ( .A1(n20801), .A2(n20805), .ZN(n20802) );
  MUX2_X1 U23800 ( .A(n20803), .B(n20802), .S(n21177), .Z(n20804) );
  AND2_X1 U23801 ( .A1(n20804), .A2(n21023), .ZN(n20816) );
  AOI22_X1 U23802 ( .A1(n20944), .A2(n20828), .B1(n21020), .B2(n20839), .ZN(
        n20812) );
  INV_X1 U23803 ( .A(n20805), .ZN(n20806) );
  NAND2_X1 U23804 ( .A1(n20806), .A2(n21177), .ZN(n20809) );
  OAI21_X1 U23805 ( .B1(n20807), .B2(n20839), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20808) );
  NAND2_X1 U23806 ( .A1(n20809), .A2(n20808), .ZN(n20829) );
  AOI22_X1 U23807 ( .A1(n21021), .A2(n20829), .B1(n20840), .B2(n21030), .ZN(
        n20811) );
  OAI211_X1 U23808 ( .C1(n20816), .C2(n20813), .A(n20812), .B(n20811), .ZN(
        P2_U3120) );
  AOI22_X1 U23809 ( .A1(n21036), .A2(n20840), .B1(n21034), .B2(n20839), .ZN(
        n20815) );
  AOI22_X1 U23810 ( .A1(n20828), .A2(n20985), .B1(n21035), .B2(n20829), .ZN(
        n20814) );
  OAI211_X1 U23811 ( .C1(n20816), .C2(n11621), .A(n20815), .B(n20814), .ZN(
        P2_U3121) );
  AOI22_X1 U23812 ( .A1(n20989), .A2(n20828), .B1(n21040), .B2(n20839), .ZN(
        n20818) );
  AOI22_X1 U23813 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20830), .B1(
        n21041), .B2(n20829), .ZN(n20817) );
  OAI211_X1 U23814 ( .C1(n20992), .C2(n20863), .A(n20818), .B(n20817), .ZN(
        P2_U3122) );
  AOI22_X1 U23815 ( .A1(n21048), .A2(n20840), .B1(n20839), .B2(n9786), .ZN(
        n20820) );
  AOI22_X1 U23816 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20830), .B1(
        n21047), .B2(n20829), .ZN(n20819) );
  OAI211_X1 U23817 ( .C1(n21051), .C2(n20825), .A(n20820), .B(n20819), .ZN(
        P2_U3123) );
  AOI22_X1 U23818 ( .A1(n21054), .A2(n20840), .B1(n20839), .B2(n21052), .ZN(
        n20822) );
  AOI22_X1 U23819 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20830), .B1(
        n21053), .B2(n20829), .ZN(n20821) );
  OAI211_X1 U23820 ( .C1(n21057), .C2(n20825), .A(n20822), .B(n20821), .ZN(
        P2_U3124) );
  AOI22_X1 U23821 ( .A1(n21060), .A2(n20840), .B1(n20839), .B2(n21058), .ZN(
        n20824) );
  AOI22_X1 U23822 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20830), .B1(
        n21059), .B2(n20829), .ZN(n20823) );
  OAI211_X1 U23823 ( .C1(n21063), .C2(n20825), .A(n20824), .B(n20823), .ZN(
        P2_U3125) );
  AOI22_X1 U23824 ( .A1(n21003), .A2(n20828), .B1(n21064), .B2(n20839), .ZN(
        n20827) );
  AOI22_X1 U23825 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20830), .B1(
        n21065), .B2(n20829), .ZN(n20826) );
  OAI211_X1 U23826 ( .C1(n21006), .C2(n20863), .A(n20827), .B(n20826), .ZN(
        P2_U3126) );
  AOI22_X1 U23827 ( .A1(n21009), .A2(n20828), .B1(n20839), .B2(n21070), .ZN(
        n20832) );
  AOI22_X1 U23828 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20830), .B1(
        n21072), .B2(n20829), .ZN(n20831) );
  OAI211_X1 U23829 ( .C1(n21014), .C2(n20863), .A(n20832), .B(n20831), .ZN(
        P2_U3127) );
  INV_X1 U23830 ( .A(n20842), .ZN(n20834) );
  NOR2_X1 U23831 ( .A1(n20833), .A2(n20837), .ZN(n20858) );
  OAI21_X1 U23832 ( .B1(n20834), .B2(n20858), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20835) );
  OAI21_X1 U23833 ( .B1(n20837), .B2(n20836), .A(n20835), .ZN(n20859) );
  AOI22_X1 U23834 ( .A1(n20859), .A2(n21021), .B1(n21020), .B2(n20858), .ZN(
        n20845) );
  NOR2_X2 U23835 ( .A1(n20971), .A2(n20838), .ZN(n20895) );
  AOI221_X1 U23836 ( .B1(n20895), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20840), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n20839), .ZN(n20841) );
  AOI211_X1 U23837 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20842), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20841), .ZN(n20843) );
  AOI22_X1 U23838 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20860), .B1(
        n20895), .B2(n21030), .ZN(n20844) );
  OAI211_X1 U23839 ( .C1(n21033), .C2(n20863), .A(n20845), .B(n20844), .ZN(
        P2_U3128) );
  AOI22_X1 U23840 ( .A1(n20859), .A2(n21035), .B1(n21034), .B2(n20858), .ZN(
        n20847) );
  AOI22_X1 U23841 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20860), .B1(
        n20895), .B2(n21036), .ZN(n20846) );
  OAI211_X1 U23842 ( .C1(n21039), .C2(n20863), .A(n20847), .B(n20846), .ZN(
        P2_U3129) );
  AOI22_X1 U23843 ( .A1(n20859), .A2(n21041), .B1(n21040), .B2(n20858), .ZN(
        n20849) );
  AOI22_X1 U23844 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20860), .B1(
        n20895), .B2(n21042), .ZN(n20848) );
  OAI211_X1 U23845 ( .C1(n21045), .C2(n20863), .A(n20849), .B(n20848), .ZN(
        P2_U3130) );
  AOI22_X1 U23846 ( .A1(n20859), .A2(n21047), .B1(n9786), .B2(n20858), .ZN(
        n20851) );
  AOI22_X1 U23847 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20860), .B1(
        n20895), .B2(n21048), .ZN(n20850) );
  OAI211_X1 U23848 ( .C1(n21051), .C2(n20863), .A(n20851), .B(n20850), .ZN(
        P2_U3131) );
  AOI22_X1 U23849 ( .A1(n20859), .A2(n21053), .B1(n21052), .B2(n20858), .ZN(
        n20853) );
  AOI22_X1 U23850 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20860), .B1(
        n20895), .B2(n21054), .ZN(n20852) );
  OAI211_X1 U23851 ( .C1(n21057), .C2(n20863), .A(n20853), .B(n20852), .ZN(
        P2_U3132) );
  AOI22_X1 U23852 ( .A1(n20859), .A2(n21059), .B1(n21058), .B2(n20858), .ZN(
        n20855) );
  AOI22_X1 U23853 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20860), .B1(
        n20895), .B2(n21060), .ZN(n20854) );
  OAI211_X1 U23854 ( .C1(n21063), .C2(n20863), .A(n20855), .B(n20854), .ZN(
        P2_U3133) );
  AOI22_X1 U23855 ( .A1(n20859), .A2(n21065), .B1(n21064), .B2(n20858), .ZN(
        n20857) );
  AOI22_X1 U23856 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20860), .B1(
        n20895), .B2(n21066), .ZN(n20856) );
  OAI211_X1 U23857 ( .C1(n21069), .C2(n20863), .A(n20857), .B(n20856), .ZN(
        P2_U3134) );
  AOI22_X1 U23858 ( .A1(n20859), .A2(n21072), .B1(n21070), .B2(n20858), .ZN(
        n20862) );
  AOI22_X1 U23859 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20860), .B1(
        n20895), .B2(n21074), .ZN(n20861) );
  OAI211_X1 U23860 ( .C1(n21080), .C2(n20863), .A(n20862), .B(n20861), .ZN(
        P2_U3135) );
  NAND2_X1 U23861 ( .A1(n21027), .A2(n21178), .ZN(n20864) );
  NAND2_X1 U23862 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20867), .ZN(
        n20875) );
  NAND2_X1 U23863 ( .A1(n20864), .A2(n20875), .ZN(n20871) );
  NAND2_X1 U23864 ( .A1(n20865), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20866) );
  NAND2_X1 U23865 ( .A1(n20866), .A2(n20975), .ZN(n20869) );
  NAND2_X1 U23866 ( .A1(n20868), .A2(n20867), .ZN(n20872) );
  AOI21_X1 U23867 ( .B1(n20869), .B2(n20872), .A(n20977), .ZN(n20870) );
  INV_X1 U23868 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20878) );
  INV_X1 U23869 ( .A(n20872), .ZN(n20893) );
  OAI21_X1 U23870 ( .B1(n20873), .B2(n20893), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20874) );
  OAI21_X1 U23871 ( .B1(n20875), .B2(n20908), .A(n20874), .ZN(n20894) );
  AOI22_X1 U23872 ( .A1(n20894), .A2(n21021), .B1(n21020), .B2(n20893), .ZN(
        n20877) );
  INV_X1 U23873 ( .A(n20930), .ZN(n20904) );
  AOI22_X1 U23874 ( .A1(n20904), .A2(n21030), .B1(n20895), .B2(n20944), .ZN(
        n20876) );
  OAI211_X1 U23875 ( .C1(n20899), .C2(n20878), .A(n20877), .B(n20876), .ZN(
        P2_U3136) );
  AOI22_X1 U23876 ( .A1(n20894), .A2(n21035), .B1(n21034), .B2(n20893), .ZN(
        n20880) );
  INV_X1 U23877 ( .A(n20899), .ZN(n20890) );
  AOI22_X1 U23878 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20890), .B1(
        n20895), .B2(n20985), .ZN(n20879) );
  OAI211_X1 U23879 ( .C1(n20988), .C2(n20930), .A(n20880), .B(n20879), .ZN(
        P2_U3137) );
  AOI22_X1 U23880 ( .A1(n20894), .A2(n21041), .B1(n21040), .B2(n20893), .ZN(
        n20882) );
  AOI22_X1 U23881 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20890), .B1(
        n20895), .B2(n20989), .ZN(n20881) );
  OAI211_X1 U23882 ( .C1(n20992), .C2(n20930), .A(n20882), .B(n20881), .ZN(
        P2_U3138) );
  AOI22_X1 U23883 ( .A1(n20894), .A2(n21047), .B1(n9786), .B2(n20893), .ZN(
        n20884) );
  AOI22_X1 U23884 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20890), .B1(
        n20895), .B2(n20993), .ZN(n20883) );
  OAI211_X1 U23885 ( .C1(n20996), .C2(n20930), .A(n20884), .B(n20883), .ZN(
        P2_U3139) );
  AOI22_X1 U23886 ( .A1(n20894), .A2(n21053), .B1(n21052), .B2(n20893), .ZN(
        n20886) );
  AOI22_X1 U23887 ( .A1(n20904), .A2(n21054), .B1(n20895), .B2(n20954), .ZN(
        n20885) );
  OAI211_X1 U23888 ( .C1(n20899), .C2(n20887), .A(n20886), .B(n20885), .ZN(
        P2_U3140) );
  AOI22_X1 U23889 ( .A1(n20894), .A2(n21059), .B1(n21058), .B2(n20893), .ZN(
        n20889) );
  AOI22_X1 U23890 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20890), .B1(
        n20895), .B2(n20958), .ZN(n20888) );
  OAI211_X1 U23891 ( .C1(n20961), .C2(n20930), .A(n20889), .B(n20888), .ZN(
        P2_U3141) );
  AOI22_X1 U23892 ( .A1(n20894), .A2(n21065), .B1(n21064), .B2(n20893), .ZN(
        n20892) );
  AOI22_X1 U23893 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20890), .B1(
        n20895), .B2(n21003), .ZN(n20891) );
  OAI211_X1 U23894 ( .C1(n21006), .C2(n20930), .A(n20892), .B(n20891), .ZN(
        P2_U3142) );
  AOI22_X1 U23895 ( .A1(n20894), .A2(n21072), .B1(n21070), .B2(n20893), .ZN(
        n20897) );
  AOI22_X1 U23896 ( .A1(n20904), .A2(n21074), .B1(n20895), .B2(n21009), .ZN(
        n20896) );
  OAI211_X1 U23897 ( .C1(n20899), .C2(n20898), .A(n20897), .B(n20896), .ZN(
        P2_U3143) );
  INV_X1 U23898 ( .A(n20900), .ZN(n20903) );
  INV_X1 U23899 ( .A(n11728), .ZN(n20901) );
  NOR3_X1 U23900 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21194), .A3(
        n12896), .ZN(n20933) );
  INV_X1 U23901 ( .A(n20933), .ZN(n20938) );
  NOR2_X1 U23902 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20938), .ZN(
        n20925) );
  OAI21_X1 U23903 ( .B1(n20901), .B2(n20925), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20902) );
  OAI21_X1 U23904 ( .B1(n20903), .B2(n20906), .A(n20902), .ZN(n20926) );
  AOI22_X1 U23905 ( .A1(n20926), .A2(n21021), .B1(n21020), .B2(n20925), .ZN(
        n20912) );
  NOR2_X2 U23906 ( .A1(n20971), .A2(n20931), .ZN(n20966) );
  OAI21_X1 U23907 ( .B1(n20966), .B2(n20904), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20905) );
  OAI21_X1 U23908 ( .B1(n20906), .B2(n12896), .A(n20905), .ZN(n20910) );
  INV_X1 U23909 ( .A(n20925), .ZN(n20907) );
  OAI211_X1 U23910 ( .C1(n11728), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20908), 
        .B(n20907), .ZN(n20909) );
  NAND3_X1 U23911 ( .A1(n20910), .A2(n21023), .A3(n20909), .ZN(n20927) );
  AOI22_X1 U23912 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20927), .B1(
        n20966), .B2(n21030), .ZN(n20911) );
  OAI211_X1 U23913 ( .C1(n21033), .C2(n20930), .A(n20912), .B(n20911), .ZN(
        P2_U3144) );
  AOI22_X1 U23914 ( .A1(n20926), .A2(n21035), .B1(n21034), .B2(n20925), .ZN(
        n20914) );
  AOI22_X1 U23915 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20927), .B1(
        n20966), .B2(n21036), .ZN(n20913) );
  OAI211_X1 U23916 ( .C1(n21039), .C2(n20930), .A(n20914), .B(n20913), .ZN(
        P2_U3145) );
  AOI22_X1 U23917 ( .A1(n20926), .A2(n21041), .B1(n21040), .B2(n20925), .ZN(
        n20916) );
  AOI22_X1 U23918 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20927), .B1(
        n20966), .B2(n21042), .ZN(n20915) );
  OAI211_X1 U23919 ( .C1(n21045), .C2(n20930), .A(n20916), .B(n20915), .ZN(
        P2_U3146) );
  AOI22_X1 U23920 ( .A1(n20926), .A2(n21047), .B1(n9786), .B2(n20925), .ZN(
        n20918) );
  AOI22_X1 U23921 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20927), .B1(
        n20966), .B2(n21048), .ZN(n20917) );
  OAI211_X1 U23922 ( .C1(n21051), .C2(n20930), .A(n20918), .B(n20917), .ZN(
        P2_U3147) );
  AOI22_X1 U23923 ( .A1(n20926), .A2(n21053), .B1(n21052), .B2(n20925), .ZN(
        n20920) );
  AOI22_X1 U23924 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20927), .B1(
        n20966), .B2(n21054), .ZN(n20919) );
  OAI211_X1 U23925 ( .C1(n21057), .C2(n20930), .A(n20920), .B(n20919), .ZN(
        P2_U3148) );
  AOI22_X1 U23926 ( .A1(n20926), .A2(n21059), .B1(n21058), .B2(n20925), .ZN(
        n20922) );
  AOI22_X1 U23927 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20927), .B1(
        n20966), .B2(n21060), .ZN(n20921) );
  OAI211_X1 U23928 ( .C1(n21063), .C2(n20930), .A(n20922), .B(n20921), .ZN(
        P2_U3149) );
  AOI22_X1 U23929 ( .A1(n20926), .A2(n21065), .B1(n21064), .B2(n20925), .ZN(
        n20924) );
  AOI22_X1 U23930 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20927), .B1(
        n20966), .B2(n21066), .ZN(n20923) );
  OAI211_X1 U23931 ( .C1(n21069), .C2(n20930), .A(n20924), .B(n20923), .ZN(
        P2_U3150) );
  AOI22_X1 U23932 ( .A1(n20926), .A2(n21072), .B1(n21070), .B2(n20925), .ZN(
        n20929) );
  AOI22_X1 U23933 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20927), .B1(
        n20966), .B2(n21074), .ZN(n20928) );
  OAI211_X1 U23934 ( .C1(n21080), .C2(n20930), .A(n20929), .B(n20928), .ZN(
        P2_U3151) );
  INV_X1 U23935 ( .A(n20931), .ZN(n20942) );
  NAND2_X1 U23936 ( .A1(n21027), .A2(n20942), .ZN(n20932) );
  NAND2_X1 U23937 ( .A1(n20932), .A2(n20938), .ZN(n20937) );
  NAND2_X1 U23938 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20933), .ZN(
        n20941) );
  AND2_X1 U23939 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20941), .ZN(n20934) );
  NAND2_X1 U23940 ( .A1(n11705), .A2(n20934), .ZN(n20940) );
  NAND2_X1 U23941 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20941), .ZN(n20935) );
  AND3_X1 U23942 ( .A1(n20940), .A2(n21023), .A3(n20935), .ZN(n20936) );
  INV_X1 U23943 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20947) );
  OAI21_X1 U23944 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20938), .A(n21225), 
        .ZN(n20939) );
  INV_X1 U23945 ( .A(n20941), .ZN(n20979) );
  AOI22_X1 U23946 ( .A1(n20965), .A2(n21021), .B1(n21020), .B2(n20979), .ZN(
        n20946) );
  AOI22_X1 U23947 ( .A1(n21008), .A2(n21030), .B1(n20966), .B2(n20944), .ZN(
        n20945) );
  OAI211_X1 U23948 ( .C1(n20964), .C2(n20947), .A(n20946), .B(n20945), .ZN(
        P2_U3152) );
  INV_X1 U23949 ( .A(n21008), .ZN(n21002) );
  AOI22_X1 U23950 ( .A1(n20965), .A2(n21035), .B1(n21034), .B2(n20979), .ZN(
        n20949) );
  INV_X1 U23951 ( .A(n20964), .ZN(n20967) );
  AOI22_X1 U23952 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20967), .B1(
        n20966), .B2(n20985), .ZN(n20948) );
  OAI211_X1 U23953 ( .C1(n20988), .C2(n21002), .A(n20949), .B(n20948), .ZN(
        P2_U3153) );
  AOI22_X1 U23954 ( .A1(n20965), .A2(n21041), .B1(n21040), .B2(n20979), .ZN(
        n20951) );
  AOI22_X1 U23955 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20967), .B1(
        n20966), .B2(n20989), .ZN(n20950) );
  OAI211_X1 U23956 ( .C1(n20992), .C2(n21002), .A(n20951), .B(n20950), .ZN(
        P2_U3154) );
  AOI22_X1 U23957 ( .A1(n20965), .A2(n21047), .B1(n9786), .B2(n20979), .ZN(
        n20953) );
  AOI22_X1 U23958 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20967), .B1(
        n20966), .B2(n20993), .ZN(n20952) );
  OAI211_X1 U23959 ( .C1(n20996), .C2(n21002), .A(n20953), .B(n20952), .ZN(
        P2_U3155) );
  AOI22_X1 U23960 ( .A1(n20965), .A2(n21053), .B1(n21052), .B2(n20979), .ZN(
        n20956) );
  AOI22_X1 U23961 ( .A1(n21008), .A2(n21054), .B1(n20966), .B2(n20954), .ZN(
        n20955) );
  OAI211_X1 U23962 ( .C1(n20964), .C2(n20957), .A(n20956), .B(n20955), .ZN(
        P2_U3156) );
  AOI22_X1 U23963 ( .A1(n20965), .A2(n21059), .B1(n21058), .B2(n20979), .ZN(
        n20960) );
  AOI22_X1 U23964 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20967), .B1(
        n20966), .B2(n20958), .ZN(n20959) );
  OAI211_X1 U23965 ( .C1(n20961), .C2(n21002), .A(n20960), .B(n20959), .ZN(
        P2_U3157) );
  AOI22_X1 U23966 ( .A1(n20965), .A2(n21065), .B1(n21064), .B2(n20979), .ZN(
        n20963) );
  AOI22_X1 U23967 ( .A1(n21008), .A2(n21066), .B1(n20966), .B2(n21003), .ZN(
        n20962) );
  OAI211_X1 U23968 ( .C1(n20964), .C2(n11844), .A(n20963), .B(n20962), .ZN(
        P2_U3158) );
  AOI22_X1 U23969 ( .A1(n20965), .A2(n21072), .B1(n21070), .B2(n20979), .ZN(
        n20969) );
  AOI22_X1 U23970 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20967), .B1(
        n20966), .B2(n21009), .ZN(n20968) );
  OAI211_X1 U23971 ( .C1(n21014), .C2(n21002), .A(n20969), .B(n20968), .ZN(
        P2_U3159) );
  NOR3_X2 U23972 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12896), .A3(
        n20972), .ZN(n21007) );
  AOI22_X1 U23973 ( .A1(n21030), .A2(n20999), .B1(n21020), .B2(n21007), .ZN(
        n20984) );
  NOR3_X1 U23974 ( .A1(n20973), .A2(n21007), .A3(n21225), .ZN(n20978) );
  NOR2_X1 U23975 ( .A1(n20999), .A2(n21008), .ZN(n20974) );
  OAI21_X1 U23976 ( .B1(n20974), .B2(n12132), .A(n21177), .ZN(n20982) );
  AOI221_X1 U23977 ( .B1(n20975), .B2(n20982), .C1(n20975), .C2(n20979), .A(
        n21007), .ZN(n20976) );
  NOR2_X1 U23978 ( .A1(n21007), .A2(n20979), .ZN(n20981) );
  OAI21_X1 U23979 ( .B1(n20973), .B2(n21007), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20980) );
  AOI22_X1 U23980 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21011), .B1(
        n21021), .B2(n21010), .ZN(n20983) );
  OAI211_X1 U23981 ( .C1(n21033), .C2(n21002), .A(n20984), .B(n20983), .ZN(
        P2_U3160) );
  AOI22_X1 U23982 ( .A1(n20985), .A2(n21008), .B1(n21034), .B2(n21007), .ZN(
        n20987) );
  AOI22_X1 U23983 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21011), .B1(
        n21035), .B2(n21010), .ZN(n20986) );
  OAI211_X1 U23984 ( .C1(n20988), .C2(n21079), .A(n20987), .B(n20986), .ZN(
        P2_U3161) );
  AOI22_X1 U23985 ( .A1(n20989), .A2(n21008), .B1(n21040), .B2(n21007), .ZN(
        n20991) );
  AOI22_X1 U23986 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21011), .B1(
        n21041), .B2(n21010), .ZN(n20990) );
  OAI211_X1 U23987 ( .C1(n20992), .C2(n21079), .A(n20991), .B(n20990), .ZN(
        P2_U3162) );
  AOI22_X1 U23988 ( .A1(n20993), .A2(n21008), .B1(n21007), .B2(n9786), .ZN(
        n20995) );
  AOI22_X1 U23989 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21011), .B1(
        n21047), .B2(n21010), .ZN(n20994) );
  OAI211_X1 U23990 ( .C1(n20996), .C2(n21079), .A(n20995), .B(n20994), .ZN(
        P2_U3163) );
  AOI22_X1 U23991 ( .A1(n21054), .A2(n20999), .B1(n21007), .B2(n21052), .ZN(
        n20998) );
  AOI22_X1 U23992 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21011), .B1(
        n21053), .B2(n21010), .ZN(n20997) );
  OAI211_X1 U23993 ( .C1(n21057), .C2(n21002), .A(n20998), .B(n20997), .ZN(
        P2_U3164) );
  AOI22_X1 U23994 ( .A1(n21060), .A2(n20999), .B1(n21007), .B2(n21058), .ZN(
        n21001) );
  AOI22_X1 U23995 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21011), .B1(
        n21059), .B2(n21010), .ZN(n21000) );
  OAI211_X1 U23996 ( .C1(n21063), .C2(n21002), .A(n21001), .B(n21000), .ZN(
        P2_U3165) );
  AOI22_X1 U23997 ( .A1(n21003), .A2(n21008), .B1(n21064), .B2(n21007), .ZN(
        n21005) );
  AOI22_X1 U23998 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21011), .B1(
        n21065), .B2(n21010), .ZN(n21004) );
  OAI211_X1 U23999 ( .C1(n21006), .C2(n21079), .A(n21005), .B(n21004), .ZN(
        P2_U3166) );
  AOI22_X1 U24000 ( .A1(n21009), .A2(n21008), .B1(n21070), .B2(n21007), .ZN(
        n21013) );
  AOI22_X1 U24001 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21011), .B1(
        n21072), .B2(n21010), .ZN(n21012) );
  OAI211_X1 U24002 ( .C1(n21014), .C2(n21079), .A(n21013), .B(n21012), .ZN(
        P2_U3167) );
  NAND2_X1 U24003 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21015), .ZN(
        n21022) );
  OR2_X1 U24004 ( .A1(n21022), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n21018) );
  NAND2_X1 U24005 ( .A1(n21019), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n21016) );
  NOR2_X1 U24006 ( .A1(n21017), .A2(n21016), .ZN(n21025) );
  AOI21_X1 U24007 ( .B1(n21225), .B2(n21018), .A(n21025), .ZN(n21073) );
  INV_X1 U24008 ( .A(n21019), .ZN(n21071) );
  AOI22_X1 U24009 ( .A1(n21073), .A2(n21021), .B1(n21071), .B2(n21020), .ZN(
        n21032) );
  INV_X1 U24010 ( .A(n21022), .ZN(n21029) );
  OAI21_X1 U24011 ( .B1(n21071), .B2(n20975), .A(n21023), .ZN(n21024) );
  NOR2_X1 U24012 ( .A1(n21025), .A2(n21024), .ZN(n21026) );
  OAI221_X1 U24013 ( .B1(n21029), .B2(n21028), .C1(n21029), .C2(n21027), .A(
        n21026), .ZN(n21076) );
  AOI22_X1 U24014 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21076), .B1(
        n21075), .B2(n21030), .ZN(n21031) );
  OAI211_X1 U24015 ( .C1(n21033), .C2(n21079), .A(n21032), .B(n21031), .ZN(
        P2_U3168) );
  AOI22_X1 U24016 ( .A1(n21073), .A2(n21035), .B1(n21071), .B2(n21034), .ZN(
        n21038) );
  AOI22_X1 U24017 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21076), .B1(
        n21075), .B2(n21036), .ZN(n21037) );
  OAI211_X1 U24018 ( .C1(n21039), .C2(n21079), .A(n21038), .B(n21037), .ZN(
        P2_U3169) );
  AOI22_X1 U24019 ( .A1(n21073), .A2(n21041), .B1(n21071), .B2(n21040), .ZN(
        n21044) );
  AOI22_X1 U24020 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21076), .B1(
        n21075), .B2(n21042), .ZN(n21043) );
  OAI211_X1 U24021 ( .C1(n21045), .C2(n21079), .A(n21044), .B(n21043), .ZN(
        P2_U3170) );
  AOI22_X1 U24022 ( .A1(n21073), .A2(n21047), .B1(n21071), .B2(n9786), .ZN(
        n21050) );
  AOI22_X1 U24023 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21076), .B1(
        n21075), .B2(n21048), .ZN(n21049) );
  OAI211_X1 U24024 ( .C1(n21051), .C2(n21079), .A(n21050), .B(n21049), .ZN(
        P2_U3171) );
  AOI22_X1 U24025 ( .A1(n21073), .A2(n21053), .B1(n21071), .B2(n21052), .ZN(
        n21056) );
  AOI22_X1 U24026 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21076), .B1(
        n21075), .B2(n21054), .ZN(n21055) );
  OAI211_X1 U24027 ( .C1(n21057), .C2(n21079), .A(n21056), .B(n21055), .ZN(
        P2_U3172) );
  AOI22_X1 U24028 ( .A1(n21073), .A2(n21059), .B1(n21071), .B2(n21058), .ZN(
        n21062) );
  AOI22_X1 U24029 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21076), .B1(
        n21075), .B2(n21060), .ZN(n21061) );
  OAI211_X1 U24030 ( .C1(n21063), .C2(n21079), .A(n21062), .B(n21061), .ZN(
        P2_U3173) );
  AOI22_X1 U24031 ( .A1(n21073), .A2(n21065), .B1(n21071), .B2(n21064), .ZN(
        n21068) );
  AOI22_X1 U24032 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21076), .B1(
        n21075), .B2(n21066), .ZN(n21067) );
  OAI211_X1 U24033 ( .C1(n21069), .C2(n21079), .A(n21068), .B(n21067), .ZN(
        P2_U3174) );
  AOI22_X1 U24034 ( .A1(n21073), .A2(n21072), .B1(n21071), .B2(n21070), .ZN(
        n21078) );
  AOI22_X1 U24035 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21076), .B1(
        n21075), .B2(n21074), .ZN(n21077) );
  OAI211_X1 U24036 ( .C1(n21080), .C2(n21079), .A(n21078), .B(n21077), .ZN(
        P2_U3175) );
  AOI21_X1 U24037 ( .B1(n21082), .B2(n21081), .A(n21241), .ZN(n21088) );
  INV_X1 U24038 ( .A(n21083), .ZN(n21087) );
  OAI211_X1 U24039 ( .C1(n21084), .C2(n21087), .A(n21226), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n21085) );
  OAI211_X1 U24040 ( .C1(n21088), .C2(n21087), .A(n21086), .B(n21085), .ZN(
        P2_U3177) );
  AND2_X1 U24041 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n21092), .ZN(
        P2_U3179) );
  AND2_X1 U24042 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n21092), .ZN(
        P2_U3180) );
  AND2_X1 U24043 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n21092), .ZN(
        P2_U3181) );
  AND2_X1 U24044 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n21092), .ZN(
        P2_U3182) );
  AND2_X1 U24045 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n21092), .ZN(
        P2_U3183) );
  AND2_X1 U24046 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n21092), .ZN(
        P2_U3184) );
  AND2_X1 U24047 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n21092), .ZN(
        P2_U3185) );
  AND2_X1 U24048 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n21092), .ZN(
        P2_U3186) );
  AND2_X1 U24049 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n21092), .ZN(
        P2_U3187) );
  AND2_X1 U24050 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n21092), .ZN(
        P2_U3188) );
  AND2_X1 U24051 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n21092), .ZN(
        P2_U3189) );
  AND2_X1 U24052 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n21092), .ZN(
        P2_U3190) );
  AND2_X1 U24053 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n21092), .ZN(
        P2_U3191) );
  AND2_X1 U24054 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n21092), .ZN(
        P2_U3192) );
  AND2_X1 U24055 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n21092), .ZN(
        P2_U3193) );
  AND2_X1 U24056 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n21090), .ZN(
        P2_U3194) );
  AND2_X1 U24057 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n21090), .ZN(
        P2_U3195) );
  AND2_X1 U24058 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n21090), .ZN(
        P2_U3196) );
  NOR2_X1 U24059 ( .A1(n21089), .A2(n21175), .ZN(P2_U3197) );
  AND2_X1 U24060 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n21090), .ZN(
        P2_U3198) );
  AND2_X1 U24061 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n21090), .ZN(
        P2_U3199) );
  AND2_X1 U24062 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n21090), .ZN(
        P2_U3200) );
  AND2_X1 U24063 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n21090), .ZN(P2_U3201) );
  AND2_X1 U24064 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n21092), .ZN(P2_U3202) );
  AND2_X1 U24065 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n21092), .ZN(P2_U3203) );
  AND2_X1 U24066 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n21092), .ZN(P2_U3204) );
  AND2_X1 U24067 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n21092), .ZN(P2_U3205) );
  NOR2_X1 U24068 ( .A1(n21091), .A2(n21175), .ZN(P2_U3206) );
  AND2_X1 U24069 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n21092), .ZN(P2_U3207) );
  NOR2_X1 U24070 ( .A1(n21093), .A2(n21175), .ZN(P2_U3208) );
  INV_X1 U24071 ( .A(NA), .ZN(n21455) );
  INV_X1 U24072 ( .A(n21094), .ZN(n21100) );
  OAI21_X1 U24073 ( .B1(n21455), .B2(n21100), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n21111) );
  NAND2_X1 U24074 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21226), .ZN(n21109) );
  NAND3_X1 U24075 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n21109), .ZN(n21097) );
  AOI211_X1 U24076 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21444), .A(
        n21244), .B(n21095), .ZN(n21096) );
  AOI21_X1 U24077 ( .B1(n21111), .B2(n21097), .A(n21096), .ZN(n21098) );
  INV_X1 U24078 ( .A(n21098), .ZN(P2_U3209) );
  NOR2_X1 U24079 ( .A1(HOLD), .A2(n21099), .ZN(n21110) );
  AOI21_X1 U24080 ( .B1(n21112), .B2(n21100), .A(n21110), .ZN(n21105) );
  INV_X1 U24081 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21104) );
  AOI21_X1 U24082 ( .B1(HOLD), .B2(n21102), .A(n21101), .ZN(n21103) );
  OAI211_X1 U24083 ( .C1(n21105), .C2(n21104), .A(n21103), .B(n21109), .ZN(
        P2_U3210) );
  OAI22_X1 U24084 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n21106), .B1(NA), 
        .B2(n21109), .ZN(n21107) );
  OAI211_X1 U24085 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n21107), .ZN(n21108) );
  OAI221_X1 U24086 ( .B1(n21111), .B2(n21110), .C1(n21111), .C2(n21109), .A(
        n21108), .ZN(P2_U3211) );
  OAI222_X1 U24087 ( .A1(n21161), .A2(n21114), .B1(n21113), .B2(n21244), .C1(
        n21116), .C2(n21163), .ZN(P2_U3212) );
  OAI222_X1 U24088 ( .A1(n21161), .A2(n21116), .B1(n21115), .B2(n21244), .C1(
        n21118), .C2(n21163), .ZN(P2_U3213) );
  OAI222_X1 U24089 ( .A1(n21161), .A2(n21118), .B1(n21117), .B2(n21244), .C1(
        n12303), .C2(n21163), .ZN(P2_U3214) );
  OAI222_X1 U24090 ( .A1(n21163), .A2(n15235), .B1(n21119), .B2(n21244), .C1(
        n12303), .C2(n21161), .ZN(P2_U3215) );
  OAI222_X1 U24091 ( .A1(n21163), .A2(n21121), .B1(n21120), .B2(n21244), .C1(
        n15235), .C2(n21161), .ZN(P2_U3216) );
  OAI222_X1 U24092 ( .A1(n21163), .A2(n21123), .B1(n21122), .B2(n21244), .C1(
        n21121), .C2(n21161), .ZN(P2_U3217) );
  OAI222_X1 U24093 ( .A1(n21163), .A2(n12320), .B1(n21124), .B2(n21244), .C1(
        n21123), .C2(n21161), .ZN(P2_U3218) );
  OAI222_X1 U24094 ( .A1(n21163), .A2(n21126), .B1(n21125), .B2(n21244), .C1(
        n12320), .C2(n21161), .ZN(P2_U3219) );
  OAI222_X1 U24095 ( .A1(n21163), .A2(n21128), .B1(n21127), .B2(n21244), .C1(
        n21126), .C2(n21161), .ZN(P2_U3220) );
  OAI222_X1 U24096 ( .A1(n21163), .A2(n21130), .B1(n21129), .B2(n21244), .C1(
        n21128), .C2(n21161), .ZN(P2_U3221) );
  OAI222_X1 U24097 ( .A1(n21163), .A2(n12077), .B1(n21131), .B2(n21244), .C1(
        n21130), .C2(n21161), .ZN(P2_U3222) );
  OAI222_X1 U24098 ( .A1(n21163), .A2(n15036), .B1(n21132), .B2(n21244), .C1(
        n12077), .C2(n21161), .ZN(P2_U3223) );
  OAI222_X1 U24099 ( .A1(n21163), .A2(n12083), .B1(n21133), .B2(n21244), .C1(
        n15036), .C2(n21161), .ZN(P2_U3224) );
  OAI222_X1 U24100 ( .A1(n21163), .A2(n12438), .B1(n21134), .B2(n21244), .C1(
        n12083), .C2(n21161), .ZN(P2_U3225) );
  OAI222_X1 U24101 ( .A1(n21163), .A2(n12455), .B1(n21135), .B2(n21244), .C1(
        n12438), .C2(n21161), .ZN(P2_U3226) );
  OAI222_X1 U24102 ( .A1(n21163), .A2(n21137), .B1(n21136), .B2(n21244), .C1(
        n12455), .C2(n21161), .ZN(P2_U3227) );
  OAI222_X1 U24103 ( .A1(n21163), .A2(n21139), .B1(n21138), .B2(n21244), .C1(
        n21137), .C2(n21161), .ZN(P2_U3228) );
  OAI222_X1 U24104 ( .A1(n21163), .A2(n21141), .B1(n21140), .B2(n21244), .C1(
        n21139), .C2(n21161), .ZN(P2_U3229) );
  OAI222_X1 U24105 ( .A1(n21163), .A2(n21143), .B1(n21142), .B2(n21244), .C1(
        n21141), .C2(n21161), .ZN(P2_U3230) );
  OAI222_X1 U24106 ( .A1(n21163), .A2(n21145), .B1(n21144), .B2(n21244), .C1(
        n21143), .C2(n21161), .ZN(P2_U3231) );
  OAI222_X1 U24107 ( .A1(n21163), .A2(n17121), .B1(n21146), .B2(n21244), .C1(
        n21145), .C2(n21161), .ZN(P2_U3232) );
  OAI222_X1 U24108 ( .A1(n21163), .A2(n21148), .B1(n21147), .B2(n21244), .C1(
        n17121), .C2(n21161), .ZN(P2_U3233) );
  OAI222_X1 U24109 ( .A1(n21163), .A2(n12471), .B1(n21149), .B2(n21244), .C1(
        n21148), .C2(n21161), .ZN(P2_U3234) );
  OAI222_X1 U24110 ( .A1(n21163), .A2(n21151), .B1(n21150), .B2(n21244), .C1(
        n12471), .C2(n21161), .ZN(P2_U3235) );
  OAI222_X1 U24111 ( .A1(n21163), .A2(n21153), .B1(n21152), .B2(n21244), .C1(
        n21151), .C2(n21161), .ZN(P2_U3236) );
  OAI222_X1 U24112 ( .A1(n21163), .A2(n21156), .B1(n21154), .B2(n21244), .C1(
        n21153), .C2(n21161), .ZN(P2_U3237) );
  OAI222_X1 U24113 ( .A1(n21161), .A2(n21156), .B1(n21155), .B2(n21244), .C1(
        n21157), .C2(n21163), .ZN(P2_U3238) );
  OAI222_X1 U24114 ( .A1(n21163), .A2(n21159), .B1(n21158), .B2(n21244), .C1(
        n21157), .C2(n21161), .ZN(P2_U3239) );
  OAI222_X1 U24115 ( .A1(n21163), .A2(n12860), .B1(n21160), .B2(n21244), .C1(
        n21159), .C2(n21161), .ZN(P2_U3240) );
  OAI222_X1 U24116 ( .A1(n21163), .A2(n12527), .B1(n21162), .B2(n21244), .C1(
        n12860), .C2(n21161), .ZN(P2_U3241) );
  INV_X1 U24117 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n21164) );
  AOI22_X1 U24118 ( .A1(n21244), .A2(n21165), .B1(n21164), .B2(n21245), .ZN(
        P2_U3585) );
  INV_X1 U24119 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21167) );
  AOI22_X1 U24120 ( .A1(n21244), .A2(n21167), .B1(n21166), .B2(n21245), .ZN(
        P2_U3586) );
  INV_X1 U24121 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n21168) );
  AOI22_X1 U24122 ( .A1(n21244), .A2(n21169), .B1(n21168), .B2(n21245), .ZN(
        P2_U3587) );
  INV_X1 U24123 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n21170) );
  AOI22_X1 U24124 ( .A1(n21244), .A2(n21171), .B1(n21170), .B2(n21245), .ZN(
        P2_U3588) );
  OAI21_X1 U24125 ( .B1(n21175), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n21173), 
        .ZN(n21172) );
  INV_X1 U24126 ( .A(n21172), .ZN(P2_U3591) );
  INV_X1 U24127 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21174) );
  OAI21_X1 U24128 ( .B1(n21175), .B2(n21174), .A(n21173), .ZN(P2_U3592) );
  NAND2_X1 U24129 ( .A1(n21176), .A2(n21177), .ZN(n21184) );
  AND2_X1 U24130 ( .A1(n21177), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n21199) );
  NAND2_X1 U24131 ( .A1(n21178), .A2(n21199), .ZN(n21188) );
  NAND3_X1 U24132 ( .A1(n21197), .A2(n21179), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n21180) );
  NAND2_X1 U24133 ( .A1(n21180), .A2(n21195), .ZN(n21189) );
  NAND2_X1 U24134 ( .A1(n21188), .A2(n21189), .ZN(n21182) );
  NAND2_X1 U24135 ( .A1(n21182), .A2(n21181), .ZN(n21183) );
  OAI211_X1 U24136 ( .C1(n21185), .C2(n20975), .A(n21184), .B(n21183), .ZN(
        n21186) );
  INV_X1 U24137 ( .A(n21186), .ZN(n21187) );
  AOI22_X1 U24138 ( .A1(n21210), .A2(n12896), .B1(n21187), .B2(n21211), .ZN(
        P2_U3602) );
  OAI21_X1 U24139 ( .B1(n21190), .B2(n21189), .A(n21188), .ZN(n21191) );
  AOI21_X1 U24140 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n21192), .A(n21191), 
        .ZN(n21193) );
  AOI22_X1 U24141 ( .A1(n21210), .A2(n21194), .B1(n21193), .B2(n21211), .ZN(
        P2_U3603) );
  INV_X1 U24142 ( .A(n21195), .ZN(n21240) );
  NOR2_X1 U24143 ( .A1(n21240), .A2(n21196), .ZN(n21198) );
  MUX2_X1 U24144 ( .A(n21199), .B(n21198), .S(n21197), .Z(n21200) );
  AOI21_X1 U24145 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n21201), .A(n21200), 
        .ZN(n21202) );
  AOI22_X1 U24146 ( .A1(n21210), .A2(n21203), .B1(n21202), .B2(n21211), .ZN(
        P2_U3604) );
  INV_X1 U24147 ( .A(n21204), .ZN(n21206) );
  OAI22_X1 U24148 ( .A1(n21207), .A2(n21240), .B1(n21206), .B2(n21205), .ZN(
        n21208) );
  AOI21_X1 U24149 ( .B1(n21212), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n21208), 
        .ZN(n21209) );
  OAI22_X1 U24150 ( .A1(n21212), .A2(n21211), .B1(n21210), .B2(n21209), .ZN(
        P2_U3605) );
  AOI22_X1 U24151 ( .A1(n21244), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n21213), 
        .B2(n21245), .ZN(P2_U3608) );
  INV_X1 U24152 ( .A(n21214), .ZN(n21215) );
  AOI21_X1 U24153 ( .B1(n21217), .B2(n21216), .A(n21215), .ZN(n21219) );
  AOI211_X1 U24154 ( .C1(n21221), .C2(n21220), .A(n21219), .B(n21218), .ZN(
        n21222) );
  INV_X1 U24155 ( .A(n21222), .ZN(n21224) );
  MUX2_X1 U24156 ( .A(P2_MORE_REG_SCAN_IN), .B(n21224), .S(n21223), .Z(
        P2_U3609) );
  NOR2_X1 U24157 ( .A1(n21226), .A2(n21225), .ZN(n21235) );
  OAI21_X1 U24158 ( .B1(n21229), .B2(n12132), .A(n21227), .ZN(n21232) );
  INV_X1 U24159 ( .A(n21228), .ZN(n21230) );
  NAND2_X1 U24160 ( .A1(n21230), .A2(n21229), .ZN(n21231) );
  MUX2_X1 U24161 ( .A(n21232), .B(n21231), .S(n9829), .Z(n21233) );
  OAI21_X1 U24162 ( .B1(n21235), .B2(n21234), .A(n21233), .ZN(n21243) );
  NAND3_X1 U24163 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n21237), .A3(n21236), 
        .ZN(n21238) );
  OAI211_X1 U24164 ( .C1(n21241), .C2(n21240), .A(n21239), .B(n21238), .ZN(
        n21242) );
  MUX2_X1 U24165 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n21243), .S(n21242), 
        .Z(P2_U3610) );
  OAI22_X1 U24166 ( .A1(n21245), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n21244), .ZN(n21246) );
  INV_X1 U24167 ( .A(n21246), .ZN(P2_U3611) );
  INV_X1 U24168 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21445) );
  NOR2_X1 U24169 ( .A1(n21445), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21453) );
  NOR2_X1 U24170 ( .A1(n21453), .A2(n12634), .ZN(n21253) );
  INV_X1 U24171 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21247) );
  INV_X2 U24172 ( .A(n21549), .ZN(n21552) );
  AOI21_X1 U24173 ( .B1(n21253), .B2(n21247), .A(n21552), .ZN(P1_U2802) );
  NAND2_X1 U24174 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21523), .ZN(n21251) );
  OAI21_X1 U24175 ( .B1(n21249), .B2(n21248), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n21250) );
  OAI21_X1 U24176 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21251), .A(n21250), 
        .ZN(P1_U2803) );
  NOR2_X1 U24177 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21448) );
  OAI21_X1 U24178 ( .B1(n21448), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21549), .ZN(
        n21252) );
  OAI21_X1 U24179 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21549), .A(n21252), 
        .ZN(P1_U2804) );
  NOR2_X1 U24180 ( .A1(n21253), .A2(n21552), .ZN(n21520) );
  OAI21_X1 U24181 ( .B1(BS16), .B2(n21448), .A(n21520), .ZN(n21518) );
  OAI21_X1 U24182 ( .B1(n21520), .B2(n21254), .A(n21518), .ZN(P1_U2805) );
  OAI21_X1 U24183 ( .B1(n21256), .B2(n21255), .A(n17312), .ZN(P1_U2806) );
  NOR4_X1 U24184 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n21260) );
  NOR4_X1 U24185 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21259) );
  NOR4_X1 U24186 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21258) );
  NOR4_X1 U24187 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n21257) );
  NAND4_X1 U24188 ( .A1(n21260), .A2(n21259), .A3(n21258), .A4(n21257), .ZN(
        n21266) );
  NOR4_X1 U24189 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n21264) );
  AOI211_X1 U24190 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_14__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21263) );
  NOR4_X1 U24191 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21262) );
  NOR4_X1 U24192 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n21261) );
  NAND4_X1 U24193 ( .A1(n21264), .A2(n21263), .A3(n21262), .A4(n21261), .ZN(
        n21265) );
  NOR2_X1 U24194 ( .A1(n21266), .A2(n21265), .ZN(n21532) );
  INV_X1 U24195 ( .A(n21532), .ZN(n21535) );
  OR2_X1 U24196 ( .A1(n21535), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n21531) );
  NOR3_X1 U24197 ( .A1(P1_DATAWIDTH_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(n21531), .ZN(n21268) );
  AOI21_X1 U24198 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n21532), .A(n21268), .ZN(
        n21267) );
  OAI21_X1 U24199 ( .B1(n21532), .B2(n21516), .A(n21267), .ZN(P1_U2807) );
  NAND2_X1 U24200 ( .A1(n21532), .A2(n21534), .ZN(n21270) );
  AOI21_X1 U24201 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n21535), .A(n21268), 
        .ZN(n21269) );
  OAI21_X1 U24202 ( .B1(P1_DATAWIDTH_REG_1__SCAN_IN), .B2(n21270), .A(n21269), 
        .ZN(P1_U2808) );
  NAND2_X1 U24203 ( .A1(n21317), .A2(n21271), .ZN(n21290) );
  AOI22_X1 U24204 ( .A1(n21345), .A2(n21272), .B1(n21343), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n21274) );
  OAI211_X1 U24205 ( .C1(n21349), .C2(n21275), .A(n21274), .B(n21273), .ZN(
        n21280) );
  OAI22_X1 U24206 ( .A1(n21278), .A2(n21277), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n21276), .ZN(n21279) );
  AOI211_X1 U24207 ( .C1(n21281), .C2(n21339), .A(n21280), .B(n21279), .ZN(
        n21282) );
  OAI21_X1 U24208 ( .B1(n21474), .B2(n21290), .A(n21282), .ZN(P1_U2831) );
  NAND2_X1 U24209 ( .A1(n21298), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n21291) );
  INV_X1 U24210 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21365) );
  NOR2_X1 U24211 ( .A1(n21349), .A2(n21283), .ZN(n21284) );
  AOI211_X1 U24212 ( .C1(n21285), .C2(n21339), .A(n21330), .B(n21284), .ZN(
        n21287) );
  NAND2_X1 U24213 ( .A1(n21345), .A2(n21362), .ZN(n21286) );
  OAI211_X1 U24214 ( .C1(n21365), .C2(n21308), .A(n21287), .B(n21286), .ZN(
        n21288) );
  AOI21_X1 U24215 ( .B1(n21363), .B2(n21312), .A(n21288), .ZN(n21289) );
  OAI221_X1 U24216 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n21291), .C1(n15125), 
        .C2(n21290), .A(n21289), .ZN(P1_U2832) );
  NOR3_X1 U24217 ( .A1(n21303), .A2(n21292), .A3(n21470), .ZN(n21293) );
  AOI21_X1 U24218 ( .B1(n21343), .B2(P1_EBX_REG_7__SCAN_IN), .A(n21293), .ZN(
        n21294) );
  OAI21_X1 U24219 ( .B1(n21296), .B2(n21295), .A(n21294), .ZN(n21297) );
  AOI211_X1 U24220 ( .C1(n21331), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n21330), .B(n21297), .ZN(n21301) );
  AOI22_X1 U24221 ( .A1(n21299), .A2(n21312), .B1(n21470), .B2(n21298), .ZN(
        n21300) );
  OAI211_X1 U24222 ( .C1(n21302), .C2(n21348), .A(n21301), .B(n21300), .ZN(
        P1_U2833) );
  INV_X1 U24223 ( .A(n21303), .ZN(n21304) );
  NAND3_X1 U24224 ( .A1(n21304), .A2(P1_REIP_REG_6__SCAN_IN), .A3(n21317), 
        .ZN(n21307) );
  INV_X1 U24225 ( .A(n21305), .ZN(n21366) );
  NAND2_X1 U24226 ( .A1(n21345), .A2(n21366), .ZN(n21306) );
  OAI211_X1 U24227 ( .C1(n21369), .C2(n21308), .A(n21307), .B(n21306), .ZN(
        n21309) );
  AOI211_X1 U24228 ( .C1(n21331), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n21330), .B(n21309), .ZN(n21314) );
  INV_X1 U24229 ( .A(n21310), .ZN(n21367) );
  AOI22_X1 U24230 ( .A1(n21367), .A2(n21312), .B1(n21311), .B2(n21339), .ZN(
        n21313) );
  OAI211_X1 U24231 ( .C1(P1_REIP_REG_6__SCAN_IN), .C2(n21315), .A(n21314), .B(
        n21313), .ZN(P1_U2834) );
  NAND2_X1 U24232 ( .A1(n21317), .A2(n21316), .ZN(n21327) );
  AOI22_X1 U24233 ( .A1(n21345), .A2(n21318), .B1(n21343), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n21319) );
  OAI21_X1 U24234 ( .B1(n21467), .B2(n21327), .A(n21319), .ZN(n21320) );
  AOI211_X1 U24235 ( .C1(n21331), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n21330), .B(n21320), .ZN(n21324) );
  AOI22_X1 U24236 ( .A1(n21322), .A2(n21357), .B1(n21321), .B2(n21467), .ZN(
        n21323) );
  OAI211_X1 U24237 ( .C1(n21325), .C2(n21348), .A(n21324), .B(n21323), .ZN(
        P1_U2835) );
  NOR2_X1 U24238 ( .A1(n21463), .A2(n21326), .ZN(n21329) );
  INV_X1 U24239 ( .A(n21327), .ZN(n21328) );
  MUX2_X1 U24240 ( .A(n21329), .B(n21328), .S(P1_REIP_REG_4__SCAN_IN), .Z(
        n21338) );
  NAND2_X1 U24241 ( .A1(n21345), .A2(n21370), .ZN(n21336) );
  NAND2_X1 U24242 ( .A1(n21343), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n21335) );
  AOI21_X1 U24243 ( .B1(n21331), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21330), .ZN(n21334) );
  OR2_X1 U24244 ( .A1(n21346), .A2(n21332), .ZN(n21333) );
  NAND4_X1 U24245 ( .A1(n21336), .A2(n21335), .A3(n21334), .A4(n21333), .ZN(
        n21337) );
  NOR2_X1 U24246 ( .A1(n21338), .A2(n21337), .ZN(n21342) );
  AOI22_X1 U24247 ( .A1(n21371), .A2(n21357), .B1(n21340), .B2(n21339), .ZN(
        n21341) );
  NAND2_X1 U24248 ( .A1(n21342), .A2(n21341), .ZN(P1_U2836) );
  AOI22_X1 U24249 ( .A1(n21345), .A2(n21344), .B1(n21343), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n21360) );
  INV_X1 U24250 ( .A(n21346), .ZN(n21352) );
  INV_X1 U24251 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21350) );
  OAI22_X1 U24252 ( .A1(n21350), .A2(n21349), .B1(n21348), .B2(n21347), .ZN(
        n21351) );
  AOI21_X1 U24253 ( .B1(n21353), .B2(n21352), .A(n21351), .ZN(n21354) );
  OAI21_X1 U24254 ( .B1(n21355), .B2(P1_REIP_REG_2__SCAN_IN), .A(n21354), .ZN(
        n21356) );
  AOI21_X1 U24255 ( .B1(n21358), .B2(n21357), .A(n21356), .ZN(n21359) );
  OAI211_X1 U24256 ( .C1(n21461), .C2(n21361), .A(n21360), .B(n21359), .ZN(
        P1_U2838) );
  AOI22_X1 U24257 ( .A1(n21363), .A2(n21377), .B1(n21376), .B2(n21362), .ZN(
        n21364) );
  OAI21_X1 U24258 ( .B1(n21381), .B2(n21365), .A(n21364), .ZN(P1_U2864) );
  AOI22_X1 U24259 ( .A1(n21367), .A2(n21377), .B1(n21376), .B2(n21366), .ZN(
        n21368) );
  OAI21_X1 U24260 ( .B1(n21381), .B2(n21369), .A(n21368), .ZN(P1_U2866) );
  INV_X1 U24261 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21373) );
  AOI22_X1 U24262 ( .A1(n21371), .A2(n21377), .B1(n21376), .B2(n21370), .ZN(
        n21372) );
  OAI21_X1 U24263 ( .B1(n21381), .B2(n21373), .A(n21372), .ZN(P1_U2868) );
  INV_X1 U24264 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21380) );
  INV_X1 U24265 ( .A(n21374), .ZN(n21375) );
  AOI22_X1 U24266 ( .A1(n21378), .A2(n21377), .B1(n21376), .B2(n21375), .ZN(
        n21379) );
  OAI21_X1 U24267 ( .B1(n21381), .B2(n21380), .A(n21379), .ZN(P1_U2871) );
  AOI22_X1 U24268 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n21392), .B1(n21407), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n21382) );
  OAI21_X1 U24269 ( .B1(n21540), .B2(n21383), .A(n21382), .ZN(P1_U2921) );
  INV_X1 U24270 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21385) );
  AOI22_X1 U24271 ( .A1(n21410), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n21384) );
  OAI21_X1 U24272 ( .B1(n21385), .B2(n21414), .A(n21384), .ZN(P1_U2922) );
  AOI22_X1 U24273 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n21407), .B1(n21410), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n21386) );
  OAI21_X1 U24274 ( .B1(n21387), .B2(n21414), .A(n21386), .ZN(P1_U2923) );
  INV_X1 U24275 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n21389) );
  AOI22_X1 U24276 ( .A1(n21410), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n21388) );
  OAI21_X1 U24277 ( .B1(n21389), .B2(n21414), .A(n21388), .ZN(P1_U2924) );
  AOI22_X1 U24278 ( .A1(n21410), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n21390) );
  OAI21_X1 U24279 ( .B1(n21391), .B2(n21414), .A(n21390), .ZN(P1_U2925) );
  AOI22_X1 U24280 ( .A1(P1_EAX_REG_10__SCAN_IN), .A2(n21392), .B1(n21407), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n21393) );
  OAI21_X1 U24281 ( .B1(n21394), .B2(n21540), .A(n21393), .ZN(P1_U2926) );
  AOI22_X1 U24282 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21410), .B1(n21407), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n21395) );
  OAI21_X1 U24283 ( .B1(n21396), .B2(n21414), .A(n21395), .ZN(P1_U2927) );
  AOI22_X1 U24284 ( .A1(n21410), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n21397) );
  OAI21_X1 U24285 ( .B1(n21398), .B2(n21414), .A(n21397), .ZN(P1_U2928) );
  AOI22_X1 U24286 ( .A1(n21410), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n21399) );
  OAI21_X1 U24287 ( .B1(n10733), .B2(n21414), .A(n21399), .ZN(P1_U2929) );
  AOI22_X1 U24288 ( .A1(n21410), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n21400) );
  OAI21_X1 U24289 ( .B1(n21401), .B2(n21414), .A(n21400), .ZN(P1_U2930) );
  AOI22_X1 U24290 ( .A1(n21410), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n21402) );
  OAI21_X1 U24291 ( .B1(n10705), .B2(n21414), .A(n21402), .ZN(P1_U2931) );
  AOI22_X1 U24292 ( .A1(n21410), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n21403) );
  OAI21_X1 U24293 ( .B1(n21404), .B2(n21414), .A(n21403), .ZN(P1_U2932) );
  AOI22_X1 U24294 ( .A1(n21410), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n21405) );
  OAI21_X1 U24295 ( .B1(n21406), .B2(n21414), .A(n21405), .ZN(P1_U2933) );
  AOI22_X1 U24296 ( .A1(n21410), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n21408) );
  OAI21_X1 U24297 ( .B1(n21409), .B2(n21414), .A(n21408), .ZN(P1_U2934) );
  AOI22_X1 U24298 ( .A1(n21410), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n21411) );
  OAI21_X1 U24299 ( .B1(n21412), .B2(n21414), .A(n21411), .ZN(P1_U2935) );
  AOI22_X1 U24300 ( .A1(n21410), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n21407), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n21413) );
  OAI21_X1 U24301 ( .B1(n21415), .B2(n21414), .A(n21413), .ZN(P1_U2936) );
  AOI22_X1 U24302 ( .A1(n21420), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n21419), .ZN(n21418) );
  NAND2_X1 U24303 ( .A1(n21422), .A2(n21416), .ZN(n21417) );
  NAND2_X1 U24304 ( .A1(n21418), .A2(n21417), .ZN(P1_U2964) );
  AOI22_X1 U24305 ( .A1(n21420), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n21419), .ZN(n21424) );
  NAND2_X1 U24306 ( .A1(n21422), .A2(n21421), .ZN(n21423) );
  NAND2_X1 U24307 ( .A1(n21424), .A2(n21423), .ZN(P1_U2966) );
  INV_X1 U24308 ( .A(n21425), .ZN(n21426) );
  AOI22_X1 U24309 ( .A1(n21429), .A2(n21428), .B1(n21427), .B2(n21426), .ZN(
        n21435) );
  OAI22_X1 U24310 ( .A1(n21432), .A2(n21431), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21430), .ZN(n21433) );
  NAND3_X1 U24311 ( .A1(n21435), .A2(n21434), .A3(n21433), .ZN(P1_U3031) );
  NOR2_X1 U24312 ( .A1(n21437), .A2(n21436), .ZN(P1_U3032) );
  NOR2_X1 U24313 ( .A1(n21439), .A2(n21438), .ZN(n21442) );
  OAI21_X1 U24314 ( .B1(n21442), .B2(n21441), .A(n21440), .ZN(P1_U3163) );
  AND2_X1 U24315 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21443), .ZN(
        P1_U3164) );
  AND2_X1 U24316 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21443), .ZN(
        P1_U3165) );
  AND2_X1 U24317 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21443), .ZN(
        P1_U3166) );
  AND2_X1 U24318 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21443), .ZN(
        P1_U3167) );
  AND2_X1 U24319 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21443), .ZN(
        P1_U3168) );
  AND2_X1 U24320 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21443), .ZN(
        P1_U3169) );
  AND2_X1 U24321 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21443), .ZN(
        P1_U3170) );
  AND2_X1 U24322 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21443), .ZN(
        P1_U3171) );
  AND2_X1 U24323 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21443), .ZN(
        P1_U3172) );
  AND2_X1 U24324 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21443), .ZN(
        P1_U3173) );
  AND2_X1 U24325 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21443), .ZN(
        P1_U3174) );
  AND2_X1 U24326 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21443), .ZN(
        P1_U3175) );
  AND2_X1 U24327 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21443), .ZN(
        P1_U3176) );
  AND2_X1 U24328 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21443), .ZN(
        P1_U3177) );
  AND2_X1 U24329 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21443), .ZN(
        P1_U3178) );
  AND2_X1 U24330 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21443), .ZN(
        P1_U3179) );
  AND2_X1 U24331 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21443), .ZN(
        P1_U3180) );
  AND2_X1 U24332 ( .A1(n21443), .A2(P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(
        P1_U3181) );
  AND2_X1 U24333 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21443), .ZN(
        P1_U3182) );
  AND2_X1 U24334 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21443), .ZN(
        P1_U3183) );
  AND2_X1 U24335 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21443), .ZN(
        P1_U3184) );
  AND2_X1 U24336 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21443), .ZN(
        P1_U3185) );
  AND2_X1 U24337 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21443), .ZN(P1_U3186) );
  AND2_X1 U24338 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21443), .ZN(P1_U3187) );
  AND2_X1 U24339 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21443), .ZN(P1_U3188) );
  AND2_X1 U24340 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21443), .ZN(P1_U3189) );
  AND2_X1 U24341 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21443), .ZN(P1_U3190) );
  AND2_X1 U24342 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21443), .ZN(P1_U3191) );
  AND2_X1 U24343 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21443), .ZN(P1_U3192) );
  AND2_X1 U24344 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21443), .ZN(P1_U3193) );
  NOR2_X1 U24345 ( .A1(n21445), .A2(n21444), .ZN(n21447) );
  AOI211_X1 U24346 ( .C1(NA), .C2(n12634), .A(n21447), .B(n21446), .ZN(n21450)
         );
  AOI21_X1 U24347 ( .B1(n21541), .B2(n21453), .A(n21448), .ZN(n21449) );
  OAI221_X1 U24348 ( .B1(n21552), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .C1(
        n21552), .C2(n21450), .A(n21449), .ZN(P1_U3194) );
  AOI21_X1 U24349 ( .B1(n21451), .B2(n21455), .A(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21459) );
  AOI221_X1 U24350 ( .B1(NA), .B2(n21453), .C1(n21452), .C2(n21453), .A(n12634), .ZN(n21454) );
  OAI211_X1 U24351 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21547), .A(HOLD), .B(
        n21454), .ZN(n21457) );
  OAI211_X1 U24352 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21455), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n12634), .ZN(n21456) );
  OAI211_X1 U24353 ( .C1(n21459), .C2(n21458), .A(n21457), .B(n21456), .ZN(
        P1_U3196) );
  NAND2_X1 U24354 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21552), .ZN(n21508) );
  INV_X1 U24355 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21460) );
  NAND2_X1 U24356 ( .A1(n21552), .A2(n10503), .ZN(n21512) );
  OAI222_X1 U24357 ( .A1(n21508), .A2(n21534), .B1(n21460), .B2(n21552), .C1(
        n21461), .C2(n21512), .ZN(P1_U3197) );
  INV_X1 U24358 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n21462) );
  OAI222_X1 U24359 ( .A1(n21512), .A2(n21463), .B1(n21462), .B2(n21552), .C1(
        n21461), .C2(n21508), .ZN(P1_U3198) );
  OAI222_X1 U24360 ( .A1(n21512), .A2(n14375), .B1(n21464), .B2(n21552), .C1(
        n21463), .C2(n21508), .ZN(P1_U3199) );
  INV_X1 U24361 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21465) );
  OAI222_X1 U24362 ( .A1(n21508), .A2(n14375), .B1(n21465), .B2(n21552), .C1(
        n21467), .C2(n21512), .ZN(P1_U3200) );
  OAI222_X1 U24363 ( .A1(n21508), .A2(n21467), .B1(n21466), .B2(n21552), .C1(
        n21468), .C2(n21512), .ZN(P1_U3201) );
  INV_X1 U24364 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21469) );
  OAI222_X1 U24365 ( .A1(n21512), .A2(n21470), .B1(n21469), .B2(n21552), .C1(
        n21468), .C2(n21508), .ZN(P1_U3202) );
  OAI222_X1 U24366 ( .A1(n21512), .A2(n15125), .B1(n21471), .B2(n21552), .C1(
        n21470), .C2(n21508), .ZN(P1_U3203) );
  INV_X1 U24367 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21472) );
  OAI222_X1 U24368 ( .A1(n21512), .A2(n21474), .B1(n21472), .B2(n21552), .C1(
        n15125), .C2(n21508), .ZN(P1_U3204) );
  INV_X1 U24369 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21476) );
  OAI222_X1 U24370 ( .A1(n21508), .A2(n21474), .B1(n21473), .B2(n21552), .C1(
        n21476), .C2(n21512), .ZN(P1_U3205) );
  INV_X1 U24371 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21475) );
  OAI222_X1 U24372 ( .A1(n21508), .A2(n21476), .B1(n21475), .B2(n21552), .C1(
        n16171), .C2(n21512), .ZN(P1_U3206) );
  INV_X1 U24373 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n21477) );
  OAI222_X1 U24374 ( .A1(n21508), .A2(n16171), .B1(n21477), .B2(n21552), .C1(
        n21479), .C2(n21512), .ZN(P1_U3207) );
  OAI222_X1 U24375 ( .A1(n21508), .A2(n21479), .B1(n21478), .B2(n21552), .C1(
        n21481), .C2(n21512), .ZN(P1_U3208) );
  INV_X1 U24376 ( .A(n21512), .ZN(n21506) );
  AOI22_X1 U24377 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n21549), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21506), .ZN(n21480) );
  OAI21_X1 U24378 ( .B1(n21481), .B2(n21508), .A(n21480), .ZN(P1_U3209) );
  INV_X1 U24379 ( .A(n21508), .ZN(n21510) );
  AOI22_X1 U24380 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n21549), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21510), .ZN(n21482) );
  OAI21_X1 U24381 ( .B1(n21484), .B2(n21512), .A(n21482), .ZN(P1_U3210) );
  AOI22_X1 U24382 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n21549), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21506), .ZN(n21483) );
  OAI21_X1 U24383 ( .B1(n21484), .B2(n21508), .A(n21483), .ZN(P1_U3211) );
  AOI22_X1 U24384 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21549), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21510), .ZN(n21485) );
  OAI21_X1 U24385 ( .B1(n21486), .B2(n21512), .A(n21485), .ZN(P1_U3212) );
  OAI222_X1 U24386 ( .A1(n21512), .A2(n16150), .B1(n21487), .B2(n21552), .C1(
        n21486), .C2(n21508), .ZN(P1_U3213) );
  INV_X1 U24387 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21488) );
  OAI222_X1 U24388 ( .A1(n21508), .A2(n16150), .B1(n21488), .B2(n21552), .C1(
        n21490), .C2(n21512), .ZN(P1_U3214) );
  AOI22_X1 U24389 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21549), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21506), .ZN(n21489) );
  OAI21_X1 U24390 ( .B1(n21490), .B2(n21508), .A(n21489), .ZN(P1_U3215) );
  INV_X1 U24391 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21492) );
  AOI22_X1 U24392 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n21549), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21510), .ZN(n21491) );
  OAI21_X1 U24393 ( .B1(n21492), .B2(n21512), .A(n21491), .ZN(P1_U3216) );
  AOI222_X1 U24394 ( .A1(n21510), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21549), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n21506), .ZN(n21493) );
  INV_X1 U24395 ( .A(n21493), .ZN(P1_U3217) );
  AOI222_X1 U24396 ( .A1(n21510), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n21549), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n21506), .ZN(n21494) );
  INV_X1 U24397 ( .A(n21494), .ZN(P1_U3218) );
  OAI222_X1 U24398 ( .A1(n21512), .A2(n21497), .B1(n21496), .B2(n21552), .C1(
        n21495), .C2(n21508), .ZN(P1_U3219) );
  AOI222_X1 U24399 ( .A1(n21510), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21549), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21506), .ZN(n21498) );
  INV_X1 U24400 ( .A(n21498), .ZN(P1_U3220) );
  AOI222_X1 U24401 ( .A1(n21510), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21549), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n21506), .ZN(n21499) );
  INV_X1 U24402 ( .A(n21499), .ZN(P1_U3221) );
  INV_X1 U24403 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21500) );
  OAI222_X1 U24404 ( .A1(n21508), .A2(n21501), .B1(n21500), .B2(n21552), .C1(
        n21503), .C2(n21512), .ZN(P1_U3222) );
  INV_X1 U24405 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21502) );
  OAI222_X1 U24406 ( .A1(n21508), .A2(n21503), .B1(n21502), .B2(n21552), .C1(
        n21505), .C2(n21512), .ZN(P1_U3223) );
  INV_X1 U24407 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21504) );
  OAI222_X1 U24408 ( .A1(n21508), .A2(n21505), .B1(n21504), .B2(n21552), .C1(
        n21509), .C2(n21512), .ZN(P1_U3224) );
  AOI22_X1 U24409 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(n21549), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21506), .ZN(n21507) );
  OAI21_X1 U24410 ( .B1(n21509), .B2(n21508), .A(n21507), .ZN(P1_U3225) );
  AOI22_X1 U24411 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(n21549), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21510), .ZN(n21511) );
  OAI21_X1 U24412 ( .B1(n21513), .B2(n21512), .A(n21511), .ZN(P1_U3226) );
  MUX2_X1 U24413 ( .A(P1_BE_N_REG_3__SCAN_IN), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .S(n21552), .Z(P1_U3458) );
  INV_X1 U24414 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21530) );
  INV_X1 U24415 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21514) );
  AOI22_X1 U24416 ( .A1(n21552), .A2(n21530), .B1(n21514), .B2(n21549), .ZN(
        P1_U3459) );
  INV_X1 U24417 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21515) );
  AOI22_X1 U24418 ( .A1(n21552), .A2(n21516), .B1(n21515), .B2(n21549), .ZN(
        P1_U3460) );
  MUX2_X1 U24419 ( .A(P1_BE_N_REG_0__SCAN_IN), .B(P1_BYTEENABLE_REG_0__SCAN_IN), .S(n21552), .Z(P1_U3461) );
  OAI21_X1 U24420 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21520), .A(n21518), 
        .ZN(n21517) );
  INV_X1 U24421 ( .A(n21517), .ZN(P1_U3464) );
  INV_X1 U24422 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21519) );
  OAI21_X1 U24423 ( .B1(n21520), .B2(n21519), .A(n21518), .ZN(P1_U3465) );
  AOI22_X1 U24424 ( .A1(n21524), .A2(n21523), .B1(n21522), .B2(n21521), .ZN(
        n21525) );
  INV_X1 U24425 ( .A(n21525), .ZN(n21527) );
  MUX2_X1 U24426 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21527), .S(
        n21526), .Z(P1_U3469) );
  AOI21_X1 U24427 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21528) );
  AOI221_X1 U24428 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .C1(n21534), .C2(n21528), .A(n21535), .ZN(n21529) );
  AOI21_X1 U24429 ( .B1(n21535), .B2(n21530), .A(n21529), .ZN(P1_U3481) );
  OAI21_X1 U24430 ( .B1(n21532), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21531), 
        .ZN(n21533) );
  OAI21_X1 U24431 ( .B1(n21535), .B2(n21534), .A(n21533), .ZN(P1_U3482) );
  AOI22_X1 U24432 ( .A1(n21552), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21536), 
        .B2(n21549), .ZN(P1_U3483) );
  INV_X1 U24433 ( .A(n21537), .ZN(n21538) );
  OAI211_X1 U24434 ( .C1(n21541), .C2(n21540), .A(n21539), .B(n21538), .ZN(
        n21548) );
  OAI211_X1 U24435 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21543), .A(n21542), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21544) );
  NAND3_X1 U24436 ( .A1(n21548), .A2(n21545), .A3(n21544), .ZN(n21546) );
  OAI21_X1 U24437 ( .B1(n21548), .B2(n21547), .A(n21546), .ZN(P1_U3485) );
  INV_X1 U24438 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21550) );
  AOI22_X1 U24439 ( .A1(n21552), .A2(n21551), .B1(n21550), .B2(n21549), .ZN(
        P1_U3486) );
  NOR2_X2 U11324 ( .A1(n13225), .A2(n20006), .ZN(n13394) );
  CLKBUF_X3 U11289 ( .A(n13310), .Z(n18472) );
  AOI22_X1 U11231 ( .A1(n11498), .A2(n11497), .B1(n11496), .B2(n11495), .ZN(
        n11499) );
  NOR2_X1 U11239 ( .A1(n10492), .A2(n10491), .ZN(n12783) );
  AND2_X1 U11249 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10368) );
  CLKBUF_X3 U11255 ( .A(n11607), .Z(n9791) );
  NOR2_X1 U11258 ( .A1(n10708), .A2(n10707), .ZN(n10728) );
  NAND2_X1 U11260 ( .A1(n10513), .A2(n10512), .ZN(n10596) );
  CLKBUF_X3 U11266 ( .A(n10800), .Z(n11134) );
  CLKBUF_X2 U11316 ( .A(n12732), .Z(n12759) );
  CLKBUF_X3 U11318 ( .A(n11444), .Z(n13778) );
  NAND2_X1 U11326 ( .A1(n16433), .A2(n13125), .ZN(n13143) );
  NAND2_X1 U11348 ( .A1(n12274), .A2(n20547), .ZN(n12435) );
  CLKBUF_X1 U11378 ( .A(n14029), .Z(n9830) );
  CLKBUF_X1 U11506 ( .A(n13077), .Z(n17469) );
  CLKBUF_X1 U11573 ( .A(n16419), .Z(n16420) );
  INV_X1 U11641 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n17682) );
  INV_X2 U11722 ( .A(n19212), .ZN(n19163) );
  CLKBUF_X1 U12474 ( .A(n17875), .Z(n17881) );
  OR2_X1 U12793 ( .A1(n20574), .A2(n11481), .ZN(n21553) );
endmodule

