

module b22_C_AntiSAT_k_256_7 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6638, n6639, n6640, n6641, n6642, n6643, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713;

  INV_X1 U7386 ( .A(n7910), .ZN(n12602) );
  BUF_X2 U7387 ( .A(n12497), .Z(n6643) );
  INV_X1 U7388 ( .A(n7754), .ZN(n9727) );
  INV_X1 U7389 ( .A(n8199), .ZN(n12601) );
  INV_X1 U7390 ( .A(n9029), .ZN(n9483) );
  NAND2_X1 U7391 ( .A1(n9020), .A2(n7039), .ZN(n15183) );
  INV_X4 U7392 ( .A(n9370), .ZN(n9501) );
  CLKBUF_X1 U7393 ( .A(n14101), .Z(n6638) );
  OAI21_X1 U7394 ( .B1(n10353), .B2(n11306), .A(n14507), .ZN(n14101) );
  INV_X1 U7396 ( .A(n8227), .ZN(n12746) );
  AND2_X1 U7397 ( .A1(n7216), .A2(n6753), .ZN(n10448) );
  INV_X1 U7398 ( .A(n10126), .ZN(n8052) );
  NAND2_X1 U7399 ( .A1(n8957), .A2(n8958), .ZN(n9248) );
  INV_X1 U7400 ( .A(n12262), .ZN(n12275) );
  BUF_X1 U7401 ( .A(n7723), .Z(n10126) );
  INV_X1 U7402 ( .A(n7489), .ZN(n9502) );
  INV_X1 U7403 ( .A(n8943), .ZN(n7615) );
  INV_X1 U7404 ( .A(n8317), .ZN(n8407) );
  AND2_X1 U7405 ( .A1(n6649), .A2(n14081), .ZN(n7203) );
  XNOR2_X1 U7406 ( .A(n12847), .B(n12845), .ZN(n13004) );
  MUX2_X1 U7407 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7693), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n7694) );
  NAND2_X1 U7408 ( .A1(n8217), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8219) );
  INV_X1 U7409 ( .A(n9829), .ZN(n9828) );
  INV_X1 U7410 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7780) );
  AOI211_X1 U7411 ( .C1(n9564), .C2(n15150), .A(n9510), .B(n9563), .ZN(n9568)
         );
  INV_X1 U7412 ( .A(n8443), .ZN(n8453) );
  XNOR2_X1 U7413 ( .A(n7762), .B(n7780), .ZN(n10213) );
  AND4_X1 U7414 ( .A1(n8399), .A2(n8398), .A3(n8397), .A4(n8487), .ZN(n6639)
         );
  AND4_X1 U7415 ( .A1(n6670), .A2(n6669), .A3(n6668), .A4(n6667), .ZN(n6640)
         );
  AND2_X1 U7416 ( .A1(n8950), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7417 ( .A1(n7761), .A2(n6756), .ZN(n8045) );
  NAND2_X2 U7418 ( .A1(n8378), .A2(n8380), .ZN(n9367) );
  INV_X1 U7420 ( .A(n8741), .ZN(n12497) );
  INV_X1 U7421 ( .A(n7767), .ZN(n8205) );
  NAND2_X2 U7422 ( .A1(n8428), .A2(n8427), .ZN(n14158) );
  AND3_X1 U7423 ( .A1(n8426), .A2(n8425), .A3(n8424), .ZN(n8427) );
  BUF_X4 U7425 ( .A(n6733), .Z(n6645) );
  BUF_X2 U7426 ( .A(n6654), .Z(n6733) );
  OR2_X1 U7427 ( .A1(n7686), .A2(n11963), .ZN(n7749) );
  XNOR2_X2 U7429 ( .A(n7698), .B(P3_IR_REG_1__SCAN_IN), .ZN(n7221) );
  NAND3_X2 U7430 ( .A1(n8998), .A2(n8997), .A3(n6750), .ZN(n15129) );
  NOR2_X2 U7431 ( .A1(n12570), .A2(n11995), .ZN(n11997) );
  AND2_X1 U7432 ( .A1(n7686), .A2(n11963), .ZN(n7750) );
  XNOR2_X2 U7433 ( .A(n7682), .B(n7681), .ZN(n11963) );
  OAI21_X2 U7434 ( .B1(n12028), .B2(n12027), .A(n12026), .ZN(n13470) );
  NAND3_X2 U7435 ( .A1(n7453), .A2(n7457), .A3(n7454), .ZN(n12026) );
  INV_X1 U7436 ( .A(n9006), .ZN(n6646) );
  NOR2_X4 U7437 ( .A1(n15151), .A2(n9704), .ZN(n9006) );
  NAND2_X1 U7438 ( .A1(n7694), .A2(n6752), .ZN(n6647) );
  NAND2_X1 U7439 ( .A1(n7694), .A2(n6752), .ZN(n6648) );
  NAND2_X1 U7440 ( .A1(n7694), .A2(n6752), .ZN(n12105) );
  OR2_X2 U7441 ( .A1(n13470), .A2(n13469), .ZN(n13471) );
  XNOR2_X2 U7442 ( .A(n13881), .B(n13585), .ZN(n13748) );
  AND2_X1 U7443 ( .A1(n13666), .A2(n13667), .ZN(n6725) );
  AND2_X1 U7444 ( .A1(n8409), .A2(n8408), .ZN(n12467) );
  OAI22_X1 U7445 ( .A1(n14439), .A2(n14442), .B1(n14632), .B2(n14138), .ZN(
        n14431) );
  OR2_X1 U7446 ( .A1(n13571), .A2(n7139), .ZN(n7137) );
  AND2_X1 U7447 ( .A1(n7185), .A2(n6650), .ZN(n6694) );
  OR2_X1 U7448 ( .A1(n8722), .A2(n8721), .ZN(n8724) );
  OAI21_X1 U7449 ( .B1(n11162), .B2(n11168), .A(n9606), .ZN(n11175) );
  INV_X1 U7450 ( .A(n11623), .ZN(n6649) );
  NAND2_X1 U7451 ( .A1(n11045), .A2(n12340), .ZN(n11362) );
  NAND2_X1 U7452 ( .A1(n9122), .A2(n9121), .ZN(n11099) );
  NAND2_X1 U7453 ( .A1(n6906), .A2(n8519), .ZN(n12342) );
  NOR2_X1 U7454 ( .A1(n10753), .A2(n12331), .ZN(n10879) );
  NAND2_X2 U7455 ( .A1(n7734), .A2(n7655), .ZN(n15243) );
  OR2_X1 U7456 ( .A1(n7768), .A2(n10673), .ZN(n7687) );
  NAND2_X1 U7457 ( .A1(n12299), .A2(n12298), .ZN(n12304) );
  CLKBUF_X2 U7458 ( .A(n7749), .Z(n7767) );
  NAND3_X1 U7459 ( .A1(n8985), .A2(n7466), .A3(n8986), .ZN(n15143) );
  INV_X2 U7460 ( .A(n9506), .ZN(n9262) );
  INV_X2 U7461 ( .A(n8979), .ZN(n9120) );
  NAND2_X1 U7462 ( .A1(n9884), .A2(n8407), .ZN(n8741) );
  NAND2_X1 U7463 ( .A1(n8419), .A2(n14655), .ZN(n8781) );
  OAI21_X1 U7464 ( .B1(n9300), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8961) );
  AND2_X1 U7465 ( .A1(n8419), .A2(n8414), .ZN(n8437) );
  NAND2_X1 U7466 ( .A1(n8710), .A2(n8874), .ZN(n14301) );
  XNOR2_X1 U7467 ( .A(n6675), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8419) );
  INV_X4 U7469 ( .A(n8407), .ZN(n9829) );
  NOR2_X1 U7470 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6670) );
  OR2_X1 U7471 ( .A1(n7571), .A2(n7301), .ZN(n7300) );
  NAND2_X1 U7472 ( .A1(n6689), .A2(n7438), .ZN(n12511) );
  NAND2_X1 U7473 ( .A1(n6692), .A2(n6690), .ZN(n6689) );
  NAND2_X1 U7474 ( .A1(n8873), .A2(n14338), .ZN(n6683) );
  OAI211_X1 U7475 ( .C1(n14985), .C2(n7231), .A(n6661), .B(n7645), .ZN(
        P1_U3525) );
  AOI22_X1 U7476 ( .A1(n12466), .A2(n12465), .B1(n12464), .B2(n12463), .ZN(
        n12471) );
  NAND2_X1 U7477 ( .A1(n13665), .A2(n9631), .ZN(n9633) );
  NAND2_X1 U7478 ( .A1(n13679), .A2(n6725), .ZN(n13665) );
  AOI21_X1 U7479 ( .B1(n13683), .B2(n15131), .A(n13682), .ZN(n13859) );
  NAND2_X1 U7480 ( .A1(n12461), .A2(n12462), .ZN(n12466) );
  NAND2_X1 U7481 ( .A1(n7124), .A2(n14921), .ZN(n6664) );
  NAND2_X1 U7482 ( .A1(n7124), .A2(n6663), .ZN(n6662) );
  XNOR2_X1 U7483 ( .A(n9750), .B(n12472), .ZN(n14327) );
  AND2_X1 U7484 ( .A1(n14345), .A2(n7244), .ZN(n9747) );
  OAI21_X1 U7485 ( .B1(n6714), .B2(n6699), .A(n7182), .ZN(n12461) );
  NOR2_X1 U7486 ( .A1(n7439), .A2(n6691), .ZN(n6690) );
  OAI21_X1 U7487 ( .B1(n8822), .B2(n7243), .A(n7241), .ZN(n9750) );
  NAND2_X1 U7488 ( .A1(n8822), .A2(n14339), .ZN(n14345) );
  INV_X1 U7489 ( .A(n7244), .ZN(n7243) );
  INV_X1 U7490 ( .A(n14343), .ZN(n8822) );
  INV_X1 U7491 ( .A(n7128), .ZN(n6663) );
  NAND2_X1 U7492 ( .A1(n13681), .A2(n13680), .ZN(n13679) );
  AOI21_X1 U7493 ( .B1(n7244), .B2(n7242), .A(n6806), .ZN(n7241) );
  OAI21_X1 U7494 ( .B1(n12000), .B2(n7456), .A(n12007), .ZN(n7455) );
  NAND2_X1 U7495 ( .A1(n7225), .A2(n7226), .ZN(n14343) );
  AND2_X1 U7496 ( .A1(n6715), .A2(n12456), .ZN(n6714) );
  OAI21_X1 U7497 ( .B1(n12457), .B2(n12458), .A(n6824), .ZN(n6699) );
  OR2_X1 U7498 ( .A1(n12512), .A2(n12547), .ZN(n7178) );
  XNOR2_X1 U7499 ( .A(n14332), .B(n14131), .ZN(n12542) );
  INV_X1 U7500 ( .A(n9701), .ZN(n13851) );
  NAND2_X1 U7501 ( .A1(n12891), .A2(n12840), .ZN(n12998) );
  INV_X1 U7502 ( .A(n6679), .ZN(n14368) );
  NOR2_X1 U7503 ( .A1(n12477), .A2(n12476), .ZN(n6691) );
  INV_X1 U7504 ( .A(n12467), .ZN(n14332) );
  AOI21_X1 U7505 ( .B1(n14362), .B2(n14361), .A(n8866), .ZN(n14340) );
  NAND2_X1 U7506 ( .A1(n14411), .A2(n7237), .ZN(n14394) );
  NAND2_X1 U7507 ( .A1(n6711), .A2(n12448), .ZN(n12452) );
  XNOR2_X1 U7508 ( .A(n8396), .B(n8395), .ZN(n11967) );
  AND2_X1 U7509 ( .A1(n14433), .A2(n8762), .ZN(n14409) );
  NAND2_X1 U7510 ( .A1(n14433), .A2(n6677), .ZN(n14411) );
  AND2_X1 U7511 ( .A1(n9436), .A2(n9435), .ZN(n13678) );
  NAND2_X1 U7512 ( .A1(n8813), .A2(n8812), .ZN(n14351) );
  NAND2_X1 U7513 ( .A1(n12445), .A2(n7436), .ZN(n6713) );
  NAND2_X1 U7514 ( .A1(n13330), .A2(n8037), .ZN(n13331) );
  XNOR2_X1 U7515 ( .A(n12065), .B(n12102), .ZN(n13136) );
  XNOR2_X1 U7516 ( .A(n8811), .B(SI_27_), .ZN(n11965) );
  NAND2_X1 U7517 ( .A1(n12443), .A2(n6693), .ZN(n12445) );
  AND2_X1 U7518 ( .A1(n7435), .A2(n12449), .ZN(n6712) );
  NAND2_X1 U7519 ( .A1(n7201), .A2(n7200), .ZN(n14396) );
  NOR2_X1 U7520 ( .A1(n14410), .A2(n6678), .ZN(n6677) );
  XNOR2_X1 U7521 ( .A(n9446), .B(n9447), .ZN(n8811) );
  NAND2_X1 U7522 ( .A1(n7169), .A2(n7167), .ZN(n9446) );
  NAND2_X1 U7523 ( .A1(n6695), .A2(n6694), .ZN(n6693) );
  NAND2_X1 U7524 ( .A1(n9384), .A2(n9383), .ZN(n13876) );
  OR2_X1 U7525 ( .A1(n12437), .A2(n7187), .ZN(n6695) );
  NAND2_X1 U7526 ( .A1(n8767), .A2(n8766), .ZN(n14553) );
  NAND2_X1 U7527 ( .A1(n7230), .A2(n7229), .ZN(n14471) );
  NAND2_X1 U7528 ( .A1(n14487), .A2(n6832), .ZN(n7230) );
  NAND2_X1 U7529 ( .A1(n9372), .A2(n9371), .ZN(n13881) );
  INV_X1 U7530 ( .A(n8762), .ZN(n6678) );
  NAND2_X1 U7531 ( .A1(n6877), .A2(n14091), .ZN(n14414) );
  NAND2_X1 U7532 ( .A1(n6701), .A2(n6700), .ZN(n6709) );
  NAND2_X1 U7533 ( .A1(n7179), .A2(n14490), .ZN(n6708) );
  NAND2_X1 U7534 ( .A1(n6702), .A2(n12403), .ZN(n6701) );
  NAND2_X1 U7535 ( .A1(n11915), .A2(n8674), .ZN(n14501) );
  NAND2_X1 U7536 ( .A1(n11512), .A2(n11511), .ZN(n11688) );
  NAND2_X1 U7537 ( .A1(n6718), .A2(n12401), .ZN(n6702) );
  OAI21_X1 U7538 ( .B1(n11796), .B2(n7579), .A(n6729), .ZN(n13805) );
  INV_X1 U7539 ( .A(n12442), .ZN(n6650) );
  NOR2_X1 U7540 ( .A1(n6710), .A2(n8637), .ZN(n6700) );
  NAND2_X1 U7541 ( .A1(n12415), .A2(n14490), .ZN(n6710) );
  INV_X1 U7542 ( .A(n12384), .ZN(n6684) );
  NAND2_X1 U7543 ( .A1(n9614), .A2(n9613), .ZN(n11794) );
  NAND2_X1 U7544 ( .A1(n6687), .A2(n6685), .ZN(n12384) );
  NAND2_X1 U7545 ( .A1(n8726), .A2(n8725), .ZN(n14570) );
  NAND2_X1 U7546 ( .A1(n11074), .A2(n7864), .ZN(n11153) );
  NAND2_X1 U7547 ( .A1(n6686), .A2(n12381), .ZN(n6685) );
  NAND2_X1 U7548 ( .A1(n6688), .A2(n12378), .ZN(n6687) );
  OAI21_X1 U7549 ( .B1(n11291), .B2(n7527), .A(n7523), .ZN(n11700) );
  INV_X1 U7550 ( .A(n12415), .ZN(n6651) );
  AOI21_X1 U7551 ( .B1(n11311), .B2(n8598), .A(n7246), .ZN(n11522) );
  NAND2_X1 U7552 ( .A1(n8714), .A2(n8713), .ZN(n14637) );
  INV_X1 U7553 ( .A(n7203), .ZN(n11669) );
  NAND2_X1 U7554 ( .A1(n7203), .A2(n7202), .ZN(n11837) );
  NAND2_X1 U7555 ( .A1(n11476), .A2(n8559), .ZN(n11311) );
  OAI21_X1 U7556 ( .B1(n6717), .B2(n6716), .A(n7188), .ZN(n12379) );
  NAND2_X1 U7557 ( .A1(n11477), .A2(n11481), .ZN(n11476) );
  AOI21_X1 U7558 ( .B1(n6755), .B2(n12371), .A(n12370), .ZN(n6716) );
  OAI21_X1 U7559 ( .B1(n6755), .B2(n12371), .A(n6828), .ZN(n6717) );
  NAND2_X1 U7560 ( .A1(n7205), .A2(n7204), .ZN(n11623) );
  NAND2_X1 U7561 ( .A1(n6728), .A2(n9605), .ZN(n11162) );
  NAND2_X1 U7562 ( .A1(n7575), .A2(n6826), .ZN(n6728) );
  OAI21_X1 U7563 ( .B1(n11275), .B2(n11274), .A(n11273), .ZN(n11276) );
  NAND2_X1 U7564 ( .A1(n8368), .A2(n8367), .ZN(n8369) );
  NAND2_X1 U7565 ( .A1(n11474), .A2(n12373), .ZN(n11605) );
  NAND2_X1 U7566 ( .A1(n11044), .A2(n12522), .ZN(n11043) );
  NAND2_X1 U7567 ( .A1(n10878), .A2(n10881), .ZN(n10877) );
  NAND2_X1 U7568 ( .A1(n6705), .A2(n6703), .ZN(n12334) );
  NAND2_X1 U7569 ( .A1(n8591), .A2(n8590), .ZN(n12382) );
  OAI21_X1 U7570 ( .B1(n10721), .B2(n7508), .A(n7506), .ZN(n11140) );
  NAND2_X1 U7571 ( .A1(n6727), .A2(n7592), .ZN(n10820) );
  NAND2_X1 U7572 ( .A1(n10694), .A2(n10695), .ZN(n11114) );
  AOI21_X1 U7573 ( .B1(n10881), .B2(n6672), .A(n8510), .ZN(n6671) );
  XNOR2_X1 U7574 ( .A(n11214), .B(n7313), .ZN(n10965) );
  INV_X1 U7575 ( .A(n11362), .ZN(n6652) );
  NAND2_X1 U7576 ( .A1(n6706), .A2(n12330), .ZN(n6705) );
  AND2_X1 U7577 ( .A1(n12882), .A2(n10693), .ZN(n10694) );
  NAND2_X1 U7578 ( .A1(n10608), .A2(n7590), .ZN(n6727) );
  NAND2_X1 U7579 ( .A1(n10751), .A2(n8498), .ZN(n10878) );
  AND2_X1 U7580 ( .A1(n12348), .A2(n12344), .ZN(n8510) );
  NAND2_X1 U7581 ( .A1(n9102), .A2(n9101), .ZN(n15117) );
  NAND2_X1 U7582 ( .A1(n10752), .A2(n8497), .ZN(n10751) );
  NAND2_X1 U7583 ( .A1(n10857), .A2(n9596), .ZN(n10608) );
  INV_X1 U7584 ( .A(n8498), .ZN(n6672) );
  INV_X2 U7585 ( .A(n14929), .ZN(n6653) );
  OAI21_X2 U7586 ( .B1(n9849), .B2(n9370), .A(n9085), .ZN(n10654) );
  NAND2_X1 U7587 ( .A1(n10859), .A2(n10858), .ZN(n10857) );
  NAND2_X1 U7588 ( .A1(n8501), .A2(n8512), .ZN(n9849) );
  NOR2_X2 U7589 ( .A1(n10319), .A2(n10318), .ZN(n13017) );
  OR2_X1 U7590 ( .A1(n11337), .A2(n12327), .ZN(n10753) );
  NAND2_X1 U7591 ( .A1(n6887), .A2(n8322), .ZN(n8500) );
  AND2_X2 U7592 ( .A1(n10348), .A2(n12502), .ZN(n12262) );
  NAND2_X1 U7593 ( .A1(n7709), .A2(n10244), .ZN(n12625) );
  INV_X1 U7594 ( .A(n11340), .ZN(n14975) );
  OAI22_X1 U7595 ( .A1(n14917), .A2(n14915), .B1(n14158), .B2(n10710), .ZN(
        n14893) );
  NAND2_X1 U7596 ( .A1(n14904), .A2(n11340), .ZN(n11337) );
  AND2_X1 U7597 ( .A1(n12306), .A2(n12305), .ZN(n14917) );
  NAND4_X2 U7598 ( .A1(n7758), .A2(n7757), .A3(n7756), .A4(n7755), .ZN(n12956)
         );
  NAND2_X1 U7599 ( .A1(n12311), .A2(n8451), .ZN(n14890) );
  AND2_X1 U7600 ( .A1(n8464), .A2(n6657), .ZN(n11340) );
  AND2_X1 U7601 ( .A1(n9591), .A2(n9544), .ZN(n15138) );
  INV_X1 U7602 ( .A(n14158), .ZN(n8436) );
  XNOR2_X1 U7603 ( .A(n12047), .B(n15129), .ZN(n10065) );
  OR2_X1 U7604 ( .A1(n14158), .A2(n14964), .ZN(n12305) );
  INV_X4 U7605 ( .A(n12304), .ZN(n12491) );
  NOR2_X1 U7606 ( .A1(n14907), .A2(n14969), .ZN(n14904) );
  OR2_X1 U7607 ( .A1(n14157), .A2(n14969), .ZN(n12311) );
  NAND4_X2 U7608 ( .A1(n8447), .A2(n8446), .A3(n8445), .A4(n8444), .ZN(n14157)
         );
  NAND2_X1 U7609 ( .A1(n14964), .A2(n14908), .ZN(n14907) );
  OAI211_X1 U7610 ( .C1(n8199), .C2(n9830), .A(n7701), .B(n7700), .ZN(n10307)
         );
  INV_X1 U7611 ( .A(n8837), .ZN(n8838) );
  INV_X1 U7612 ( .A(n14964), .ZN(n10710) );
  NAND4_X1 U7613 ( .A1(n8457), .A2(n8456), .A3(n8455), .A4(n8454), .ZN(n14156)
         );
  AND3_X2 U7614 ( .A1(n8435), .A2(n8434), .A3(n8433), .ZN(n14964) );
  AOI21_X1 U7615 ( .B1(n8712), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n6658), .ZN(
        n6657) );
  OR2_X1 U7616 ( .A1(n6660), .A2(n6659), .ZN(n14969) );
  NAND2_X1 U7617 ( .A1(n8443), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8447) );
  NAND4_X1 U7618 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), .ZN(n13605)
         );
  INV_X2 U7619 ( .A(n9794), .ZN(n15134) );
  OR2_X1 U7620 ( .A1(n10126), .A2(n7213), .ZN(n7742) );
  NAND2_X2 U7621 ( .A1(n7723), .A2(n9828), .ZN(n8199) );
  NAND2_X1 U7622 ( .A1(n7723), .A2(n9829), .ZN(n7910) );
  AOI21_X1 U7623 ( .B1(n7419), .B2(n7417), .A(n7416), .ZN(n7415) );
  NAND2_X1 U7624 ( .A1(n7686), .A2(n7685), .ZN(n7768) );
  INV_X1 U7625 ( .A(n9505), .ZN(n9487) );
  INV_X1 U7626 ( .A(n6749), .ZN(n12212) );
  OAI22_X1 U7627 ( .A1(n8741), .A2(n9871), .B1(n9884), .B2(n14180), .ZN(n6659)
         );
  NOR2_X1 U7628 ( .A1(n12495), .A2(n9824), .ZN(n6660) );
  AND2_X1 U7629 ( .A1(n8711), .A2(n14195), .ZN(n6658) );
  AND2_X1 U7630 ( .A1(n8887), .A2(n8886), .ZN(n11633) );
  INV_X1 U7631 ( .A(n8453), .ZN(n12478) );
  NAND2_X2 U7632 ( .A1(n9884), .A2(n9829), .ZN(n12495) );
  OR2_X1 U7633 ( .A1(n8883), .A2(n8882), .ZN(n8887) );
  CLKBUF_X1 U7634 ( .A(n9511), .Z(n13638) );
  INV_X1 U7635 ( .A(n8781), .ZN(n6654) );
  AND2_X1 U7636 ( .A1(n12561), .A2(n8414), .ZN(n8443) );
  NAND2_X1 U7637 ( .A1(n9510), .A2(n10906), .ZN(n9793) );
  NAND2_X1 U7638 ( .A1(n13463), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7679) );
  BUF_X2 U7639 ( .A(n8972), .Z(n11135) );
  XNOR2_X1 U7640 ( .A(n8829), .B(P1_IR_REG_21__SCAN_IN), .ZN(n12489) );
  INV_X1 U7641 ( .A(n8414), .ZN(n14655) );
  XNOR2_X1 U7642 ( .A(n8827), .B(P1_IR_REG_22__SCAN_IN), .ZN(n12297) );
  NAND2_X1 U7643 ( .A1(n8941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8937) );
  XNOR2_X1 U7644 ( .A(n8413), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U7645 ( .A1(n6726), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8827) );
  INV_X2 U7646 ( .A(n13465), .ZN(n12584) );
  INV_X2 U7647 ( .A(n10995), .ZN(n6655) );
  INV_X2 U7648 ( .A(n11471), .ZN(n6656) );
  NAND2_X1 U7649 ( .A1(n6886), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7123) );
  NAND2_X1 U7650 ( .A1(n8955), .A2(n7027), .ZN(n13957) );
  AND2_X1 U7651 ( .A1(n8969), .A2(n8968), .ZN(n9565) );
  NAND2_X1 U7652 ( .A1(n6697), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6675) );
  OR2_X1 U7653 ( .A1(n8969), .A2(n13945), .ZN(n8967) );
  NAND2_X2 U7654 ( .A1(n9829), .A2(P2_U3088), .ZN(n13955) );
  AOI21_X1 U7655 ( .B1(n8956), .B2(n6783), .A(n7028), .ZN(n7027) );
  NOR2_X2 U7656 ( .A1(n8211), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U7657 ( .A1(n7536), .A2(n7538), .ZN(n8412) );
  NAND2_X1 U7658 ( .A1(n7538), .A2(n6676), .ZN(n6697) );
  AND2_X1 U7659 ( .A1(n8966), .A2(n8964), .ZN(n8969) );
  AND2_X2 U7660 ( .A1(n8647), .A2(n7651), .ZN(n7538) );
  NOR2_X1 U7661 ( .A1(n8404), .A2(n6673), .ZN(n6676) );
  AND3_X1 U7662 ( .A1(n8932), .A2(n8957), .A3(n7494), .ZN(n8953) );
  NOR2_X1 U7663 ( .A1(n8404), .A2(n7535), .ZN(n7536) );
  NOR2_X1 U7664 ( .A1(n8404), .A2(n7252), .ZN(n7251) );
  NAND2_X1 U7665 ( .A1(n6674), .A2(n6696), .ZN(n6673) );
  NAND4_X1 U7666 ( .A1(n8875), .A2(n15475), .A3(n8878), .A4(n8403), .ZN(n8404)
         );
  AND2_X2 U7667 ( .A1(n7464), .A2(n9001), .ZN(n8957) );
  CLKBUF_X1 U7668 ( .A(n9001), .Z(n9017) );
  INV_X1 U7669 ( .A(n7535), .ZN(n6674) );
  AND3_X1 U7670 ( .A1(n6666), .A2(n6665), .A3(n8826), .ZN(n8875) );
  AND2_X1 U7671 ( .A1(n7668), .A2(n8006), .ZN(n8046) );
  AND2_X1 U7672 ( .A1(n8951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8952) );
  AND3_X1 U7673 ( .A1(n8930), .A2(n8929), .A3(n8928), .ZN(n8958) );
  AND2_X1 U7674 ( .A1(n8981), .A2(n8931), .ZN(n9001) );
  AND3_X1 U7675 ( .A1(n7672), .A2(n7671), .A3(n7670), .ZN(n7983) );
  AND3_X1 U7676 ( .A1(n7067), .A2(n7066), .A3(n7065), .ZN(n7464) );
  INV_X1 U7677 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8826) );
  INV_X1 U7678 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6696) );
  NOR2_X1 U7679 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6666) );
  NOR2_X1 U7680 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n6665) );
  NOR2_X1 U7681 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n8399) );
  INV_X1 U7682 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8398) );
  INV_X1 U7683 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8448) );
  INV_X1 U7684 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n15674) );
  INV_X1 U7685 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6667) );
  NOR2_X1 U7686 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7065) );
  INV_X1 U7687 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8678) );
  NOR2_X1 U7688 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7066) );
  INV_X4 U7689 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7690 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6668) );
  NOR2_X1 U7691 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7067) );
  INV_X4 U7692 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7693 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8610) );
  NOR2_X1 U7694 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6669) );
  INV_X1 U7695 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8662) );
  NOR2_X1 U7696 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n8930) );
  NOR2_X1 U7697 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8929) );
  NOR2_X1 U7698 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8928) );
  NOR2_X1 U7699 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n7024) );
  INV_X1 U7700 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6681) );
  INV_X4 U7701 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR3_X1 U7702 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .A3(
        P3_IR_REG_9__SCAN_IN), .ZN(n7673) );
  NOR2_X1 U7703 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8981) );
  NOR2_X1 U7704 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7539) );
  NOR2_X1 U7705 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7589) );
  NAND3_X1 U7706 ( .A1(n6664), .A2(n6662), .A3(n14987), .ZN(n6661) );
  OR2_X2 U7707 ( .A1(n11837), .A2(n14647), .ZN(n11917) );
  NOR2_X2 U7708 ( .A1(n14414), .A2(n14553), .ZN(n7201) );
  NOR2_X2 U7709 ( .A1(n14511), .A2(n7196), .ZN(n6877) );
  NOR2_X2 U7710 ( .A1(n11605), .A2(n12377), .ZN(n7205) );
  NOR2_X2 U7711 ( .A1(n11475), .A2(n12368), .ZN(n11474) );
  AND2_X2 U7712 ( .A1(n10879), .A2(n12348), .ZN(n11045) );
  OAI21_X1 U7713 ( .B1(n12520), .B2(n10751), .A(n6671), .ZN(n11044) );
  NAND2_X1 U7714 ( .A1(n14394), .A2(n8787), .ZN(n6679) );
  NAND2_X1 U7715 ( .A1(n6683), .A2(n14987), .ZN(n8925) );
  NAND2_X1 U7716 ( .A1(n6682), .A2(n6680), .ZN(P1_U3556) );
  OR2_X1 U7717 ( .A1(n14994), .A2(n6681), .ZN(n6680) );
  NAND2_X1 U7718 ( .A1(n6683), .A2(n14994), .ZN(n6682) );
  OAI21_X2 U7719 ( .B1(n14501), .B2(n8688), .A(n8687), .ZN(n14487) );
  NAND2_X1 U7720 ( .A1(n9755), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6698) );
  AND2_X2 U7721 ( .A1(n12561), .A2(n14655), .ZN(n9755) );
  NAND2_X1 U7722 ( .A1(n6684), .A2(n12386), .ZN(n6719) );
  INV_X1 U7723 ( .A(n12379), .ZN(n6686) );
  NAND2_X1 U7724 ( .A1(n12379), .A2(n12380), .ZN(n6688) );
  NAND3_X1 U7725 ( .A1(n7177), .A2(n7178), .A3(n12511), .ZN(n6722) );
  NAND3_X1 U7726 ( .A1(n12469), .A2(n12472), .A3(n12473), .ZN(n6692) );
  NAND4_X1 U7727 ( .A1(n8439), .A2(n8440), .A3(n8438), .A4(n6698), .ZN(n8837)
         );
  NAND2_X1 U7728 ( .A1(n6704), .A2(n12328), .ZN(n6703) );
  NAND2_X1 U7729 ( .A1(n6707), .A2(n12329), .ZN(n6704) );
  INV_X1 U7730 ( .A(n6707), .ZN(n6706) );
  NAND2_X1 U7731 ( .A1(n12325), .A2(n12326), .ZN(n6707) );
  NAND3_X1 U7732 ( .A1(n6709), .A2(n12433), .A3(n6708), .ZN(n12437) );
  NAND2_X1 U7733 ( .A1(n6713), .A2(n6712), .ZN(n6711) );
  NAND2_X1 U7734 ( .A1(n12457), .A2(n12458), .ZN(n6715) );
  NAND2_X1 U7735 ( .A1(n6720), .A2(n6719), .ZN(n6718) );
  NAND2_X1 U7736 ( .A1(n6721), .A2(n12383), .ZN(n6720) );
  NAND2_X1 U7737 ( .A1(n12384), .A2(n12385), .ZN(n6721) );
  OAI211_X1 U7738 ( .C1(n12511), .C2(n6723), .A(n9883), .B(n6722), .ZN(n6724)
         );
  NAND2_X1 U7739 ( .A1(n7177), .A2(n6834), .ZN(n6723) );
  NAND2_X1 U7740 ( .A1(n6724), .A2(n7175), .ZN(P1_U3242) );
  OAI21_X2 U7741 ( .B1(n13687), .B2(n9629), .A(n9628), .ZN(n13681) );
  NOR2_X1 U7742 ( .A1(n6726), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n8908) );
  NAND2_X1 U7743 ( .A1(n8828), .A2(n8826), .ZN(n6726) );
  INV_X1 U7744 ( .A(n11175), .ZN(n9608) );
  NAND2_X2 U7745 ( .A1(n9828), .A2(n8979), .ZN(n7489) );
  NAND2_X2 U7746 ( .A1(n9585), .A2(n13957), .ZN(n8979) );
  OAI21_X2 U7747 ( .B1(n6641), .B2(n8952), .A(n8954), .ZN(n9585) );
  OR2_X1 U7748 ( .A1(n7581), .A2(n9619), .ZN(n6729) );
  NAND2_X2 U7749 ( .A1(n6730), .A2(n9615), .ZN(n11796) );
  INV_X1 U7750 ( .A(n11794), .ZN(n6730) );
  NAND3_X1 U7751 ( .A1(n15138), .A2(n10065), .A3(n15126), .ZN(n7610) );
  NAND2_X2 U7752 ( .A1(n6731), .A2(n9005), .ZN(n12047) );
  INV_X1 U7753 ( .A(n9004), .ZN(n6731) );
  XNOR2_X1 U7754 ( .A(n8406), .B(n8405), .ZN(n14169) );
  NAND2_X1 U7755 ( .A1(n8893), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8406) );
  AOI21_X2 U7756 ( .B1(n8605), .B2(n8347), .A(n8346), .ZN(n8640) );
  BUF_X4 U7757 ( .A(n7768), .Z(n6732) );
  AOI21_X2 U7758 ( .B1(n8270), .B2(n11423), .A(n11559), .ZN(n11950) );
  INV_X2 U7759 ( .A(n8437), .ZN(n8868) );
  NAND2_X4 U7760 ( .A1(n7615), .A2(n13951), .ZN(n9029) );
  CLKBUF_X1 U7761 ( .A(n14169), .Z(n6734) );
  OAI21_X2 U7762 ( .B1(n14455), .B2(n14454), .A(n8736), .ZN(n14439) );
  INV_X1 U7763 ( .A(n9006), .ZN(n6735) );
  OR2_X1 U7764 ( .A1(n11414), .A2(n12509), .ZN(n6736) );
  OR2_X1 U7765 ( .A1(n9701), .A2(n13473), .ZN(n9631) );
  NOR2_X1 U7766 ( .A1(n8575), .A2(n7420), .ZN(n7419) );
  INV_X1 U7767 ( .A(n7422), .ZN(n7420) );
  OR2_X1 U7768 ( .A1(n9742), .A2(n12909), .ZN(n12763) );
  NOR2_X1 U7769 ( .A1(n8045), .A2(n7667), .ZN(n7676) );
  AND2_X1 U7770 ( .A1(n12526), .A2(n8850), .ZN(n7268) );
  NAND2_X1 U7771 ( .A1(n9492), .A2(n9491), .ZN(n9456) );
  AND2_X1 U7772 ( .A1(n8356), .A2(n8355), .ZN(n8661) );
  AND2_X1 U7773 ( .A1(n8604), .A2(n8607), .ZN(n8347) );
  INV_X1 U7774 ( .A(n8606), .ZN(n8346) );
  NAND2_X1 U7775 ( .A1(n7414), .A2(n7412), .ZN(n8605) );
  AOI21_X1 U7776 ( .B1(n7415), .B2(n7418), .A(n7413), .ZN(n7412) );
  NAND2_X1 U7777 ( .A1(n7152), .A2(n7154), .ZN(n7414) );
  INV_X1 U7778 ( .A(n8587), .ZN(n7413) );
  AOI22_X1 U7779 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n15483), .B1(n14735), 
        .B2(n14734), .ZN(n14741) );
  INV_X1 U7780 ( .A(n6732), .ZN(n8209) );
  AOI21_X1 U7781 ( .B1(n7561), .B2(n7558), .A(n6795), .ZN(n7557) );
  INV_X1 U7782 ( .A(n6758), .ZN(n7558) );
  INV_X1 U7783 ( .A(n13587), .ZN(n13513) );
  NAND2_X1 U7784 ( .A1(n7170), .A2(n9479), .ZN(n9701) );
  NAND2_X1 U7785 ( .A1(n11967), .A2(n9501), .ZN(n7170) );
  OAI21_X1 U7786 ( .B1(n13695), .B2(n7469), .A(n7470), .ZN(n13657) );
  INV_X1 U7787 ( .A(n7471), .ZN(n7470) );
  NAND2_X1 U7788 ( .A1(n9630), .A2(n9700), .ZN(n7469) );
  OAI21_X1 U7789 ( .B1(n13680), .B2(n6737), .A(n6796), .ZN(n7471) );
  AOI22_X1 U7790 ( .A1(n13700), .A2(n13703), .B1(n12011), .B2(n13866), .ZN(
        n13687) );
  NAND2_X1 U7791 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  NAND2_X1 U7792 ( .A1(n12305), .A2(n12304), .ZN(n12308) );
  AND3_X1 U7793 ( .A1(n9496), .A2(n7151), .A3(n9540), .ZN(n9497) );
  AND2_X1 U7794 ( .A1(n9521), .A2(n9495), .ZN(n7151) );
  NOR2_X1 U7795 ( .A1(n13918), .A2(n13911), .ZN(n7077) );
  NAND2_X1 U7796 ( .A1(n7168), .A2(SI_26_), .ZN(n7167) );
  NAND2_X1 U7797 ( .A1(n8393), .A2(n8392), .ZN(n7169) );
  NAND3_X1 U7798 ( .A1(n7398), .A2(n7396), .A3(n7155), .ZN(n7154) );
  AND2_X1 U7799 ( .A1(n8336), .A2(n8332), .ZN(n7155) );
  NAND2_X1 U7800 ( .A1(n6888), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7393) );
  INV_X1 U7801 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7695) );
  NAND2_X1 U7802 ( .A1(n7142), .A2(n7696), .ZN(n7395) );
  INV_X1 U7803 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7696) );
  INV_X1 U7804 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7143) );
  OAI21_X1 U7805 ( .B1(n14693), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14664), .ZN(
        n14665) );
  AND2_X2 U7806 ( .A1(n10303), .A2(n10302), .ZN(n12849) );
  AND2_X1 U7807 ( .A1(n7306), .A2(n7305), .ZN(n10458) );
  NAND2_X1 U7808 ( .A1(n7057), .A2(n7056), .ZN(n7315) );
  AOI21_X1 U7809 ( .B1(n11569), .B2(n7058), .A(n12074), .ZN(n7056) );
  NAND2_X1 U7810 ( .A1(n13218), .A2(n8170), .ZN(n7550) );
  OR2_X1 U7811 ( .A1(n8117), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U7812 ( .A1(n7543), .A2(n7541), .ZN(n7540) );
  INV_X1 U7813 ( .A(n7973), .ZN(n7541) );
  OR2_X1 U7814 ( .A1(n14789), .A2(n13055), .ZN(n12681) );
  OR2_X1 U7815 ( .A1(n7789), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U7816 ( .A1(n6931), .A2(n6929), .ZN(n7939) );
  AOI21_X1 U7817 ( .B1(n6835), .B2(n7903), .A(n6930), .ZN(n6929) );
  INV_X1 U7818 ( .A(n7921), .ZN(n6930) );
  NOR2_X1 U7819 ( .A1(n9861), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U7820 ( .A1(n9848), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U7821 ( .A1(n13876), .A2(n13480), .ZN(n7606) );
  AND2_X1 U7822 ( .A1(n13911), .A2(n13591), .ZN(n9689) );
  NAND2_X1 U7823 ( .A1(n9617), .A2(n13591), .ZN(n7587) );
  NAND2_X1 U7824 ( .A1(n11102), .A2(n11091), .ZN(n9602) );
  AND2_X1 U7825 ( .A1(n8933), .A2(n8951), .ZN(n7494) );
  INV_X1 U7826 ( .A(n11547), .ZN(n7528) );
  AND2_X1 U7827 ( .A1(n10348), .A2(n10343), .ZN(n11281) );
  NOR2_X1 U7828 ( .A1(n14269), .A2(n6965), .ZN(n14283) );
  AND2_X1 U7829 ( .A1(n14270), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6965) );
  NAND2_X1 U7830 ( .A1(n14637), .A2(n14096), .ZN(n12431) );
  OR2_X1 U7831 ( .A1(n14832), .A2(n12157), .ZN(n12397) );
  OR2_X1 U7832 ( .A1(n14637), .A2(n14583), .ZN(n7199) );
  NAND2_X1 U7833 ( .A1(n9456), .A2(n6866), .ZN(n9500) );
  INV_X1 U7834 ( .A(n9498), .ZN(n7144) );
  INV_X1 U7835 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8878) );
  OAI21_X1 U7836 ( .B1(n8689), .B2(n8364), .A(n6881), .ZN(n8368) );
  INV_X1 U7837 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8402) );
  XNOR2_X1 U7838 ( .A(n8365), .B(SI_19_), .ZN(n8706) );
  NAND2_X1 U7839 ( .A1(n8340), .A2(n8339), .ZN(n8575) );
  AND2_X1 U7840 ( .A1(n7154), .A2(n7153), .ZN(n8560) );
  NAND2_X2 U7841 ( .A1(n7393), .A2(n7395), .ZN(n8317) );
  XNOR2_X1 U7842 ( .A(n14667), .B(n6958), .ZN(n14698) );
  INV_X1 U7843 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6958) );
  AOI22_X1 U7844 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14221), .B1(n14703), .B2(
        n14670), .ZN(n14671) );
  INV_X2 U7845 ( .A(n12849), .ZN(n12903) );
  INV_X1 U7846 ( .A(n12848), .ZN(n7354) );
  OR2_X1 U7847 ( .A1(n7897), .A2(n7896), .ZN(n7932) );
  NAND2_X1 U7848 ( .A1(n7375), .A2(n6853), .ZN(n12761) );
  NAND2_X1 U7849 ( .A1(n7376), .A2(n12760), .ZN(n7375) );
  NAND2_X1 U7850 ( .A1(n6934), .A2(n12797), .ZN(n7376) );
  NAND2_X1 U7851 ( .A1(n7377), .A2(n6935), .ZN(n6934) );
  NOR2_X1 U7852 ( .A1(n10464), .A2(n10500), .ZN(n10499) );
  OR2_X1 U7853 ( .A1(n10483), .A2(n10482), .ZN(n7220) );
  NAND2_X1 U7854 ( .A1(n6997), .A2(n7001), .ZN(n6996) );
  INV_X1 U7855 ( .A(n6999), .ZN(n6997) );
  AOI21_X1 U7856 ( .B1(n10957), .B2(n10958), .A(n7000), .ZN(n6999) );
  INV_X1 U7857 ( .A(n11230), .ZN(n7000) );
  NOR2_X1 U7858 ( .A1(n13139), .A2(n13404), .ZN(n13138) );
  INV_X1 U7859 ( .A(n7557), .ZN(n7556) );
  AND2_X1 U7860 ( .A1(n13247), .A2(n7555), .ZN(n7554) );
  NAND2_X1 U7861 ( .A1(n7557), .A2(n7559), .ZN(n7555) );
  OR2_X1 U7862 ( .A1(n13375), .A2(n13273), .ZN(n12730) );
  NAND2_X1 U7863 ( .A1(n13331), .A2(n7548), .ZN(n13317) );
  NOR2_X1 U7864 ( .A1(n13325), .A2(n7549), .ZN(n7548) );
  INV_X1 U7865 ( .A(n8038), .ZN(n7549) );
  OR2_X1 U7866 ( .A1(n13340), .A2(n13315), .ZN(n12702) );
  INV_X1 U7867 ( .A(n12800), .ZN(n12613) );
  OR2_X1 U7868 ( .A1(n11077), .A2(n8234), .ZN(n11192) );
  NAND2_X1 U7869 ( .A1(n11252), .A2(n7551), .ZN(n11074) );
  NOR2_X1 U7870 ( .A1(n7552), .A2(n12774), .ZN(n7551) );
  INV_X1 U7871 ( .A(n7845), .ZN(n7552) );
  INV_X1 U7872 ( .A(n7910), .ZN(n7836) );
  XNOR2_X1 U7873 ( .A(n8212), .B(n7363), .ZN(n12617) );
  OR2_X1 U7874 ( .A1(n7904), .A2(n7903), .ZN(n6932) );
  INV_X1 U7875 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7663) );
  INV_X1 U7876 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7662) );
  OAI21_X1 U7877 ( .B1(n7817), .B2(n7816), .A(n7818), .ZN(n7834) );
  INV_X1 U7878 ( .A(n7815), .ZN(n7816) );
  AND2_X1 U7879 ( .A1(n7539), .A2(n10404), .ZN(n7726) );
  XNOR2_X1 U7880 ( .A(n11505), .B(n11494), .ZN(n11509) );
  XNOR2_X1 U7881 ( .A(n11997), .B(n11998), .ZN(n13479) );
  AND2_X1 U7882 ( .A1(n7138), .A2(n6831), .ZN(n7136) );
  AND2_X1 U7883 ( .A1(n9423), .A2(n9422), .ZN(n13526) );
  AND2_X1 U7884 ( .A1(n9283), .A2(n9282), .ZN(n13568) );
  NAND2_X1 U7885 ( .A1(n13675), .A2(n6745), .ZN(n7071) );
  XNOR2_X1 U7886 ( .A(n13845), .B(n13578), .ZN(n9702) );
  NAND2_X1 U7887 ( .A1(n9631), .A2(n9559), .ZN(n13656) );
  AND2_X1 U7888 ( .A1(n13691), .A2(n13678), .ZN(n13675) );
  OAI22_X1 U7889 ( .A1(n9699), .A2(n9698), .B1(n13582), .B2(n13866), .ZN(
        n13695) );
  OAI21_X1 U7890 ( .B1(n7598), .B2(n13743), .A(n7595), .ZN(n13700) );
  AOI21_X1 U7891 ( .B1(n7596), .B2(n7597), .A(n6805), .ZN(n7595) );
  INV_X1 U7892 ( .A(n7602), .ZN(n7596) );
  NAND2_X1 U7893 ( .A1(n13771), .A2(n7481), .ZN(n7480) );
  AOI21_X1 U7894 ( .B1(n7481), .B2(n13760), .A(n9694), .ZN(n7479) );
  AND2_X1 U7895 ( .A1(n13881), .A2(n13585), .ZN(n9694) );
  OR2_X1 U7896 ( .A1(n13771), .A2(n13760), .ZN(n7483) );
  NOR2_X1 U7897 ( .A1(n7044), .A2(n9692), .ZN(n7043) );
  INV_X1 U7898 ( .A(n9691), .ZN(n7044) );
  AND2_X1 U7899 ( .A1(n13896), .A2(n13569), .ZN(n9621) );
  NAND2_X1 U7900 ( .A1(n13799), .A2(n13588), .ZN(n9622) );
  OR2_X1 U7901 ( .A1(n13811), .A2(n13896), .ZN(n13794) );
  OR2_X1 U7902 ( .A1(n13918), .A2(n11691), .ZN(n9616) );
  NAND2_X1 U7903 ( .A1(n11266), .A2(n9684), .ZN(n7475) );
  NOR2_X1 U7904 ( .A1(n6775), .A2(n7037), .ZN(n7036) );
  INV_X1 U7905 ( .A(n9669), .ZN(n7037) );
  NOR2_X1 U7906 ( .A1(n10718), .A2(n10719), .ZN(n7512) );
  NAND2_X1 U7907 ( .A1(n14064), .A2(n14063), .ZN(n7516) );
  AND4_X1 U7908 ( .A1(n8658), .A2(n8657), .A3(n8656), .A4(n8655), .ZN(n11666)
         );
  NAND2_X1 U7909 ( .A1(n11633), .A2(n8907), .ZN(n10348) );
  NOR2_X1 U7910 ( .A1(n11875), .A2(n11720), .ZN(n8907) );
  AOI21_X1 U7911 ( .B1(n6740), .B2(n7228), .A(n6793), .ZN(n7226) );
  INV_X1 U7912 ( .A(n8797), .ZN(n7228) );
  NAND2_X1 U7913 ( .A1(n14379), .A2(n8865), .ZN(n14362) );
  AND2_X1 U7914 ( .A1(n7432), .A2(n8703), .ZN(n7229) );
  INV_X1 U7915 ( .A(n7260), .ZN(n7259) );
  OAI21_X1 U7916 ( .B1(n11834), .B2(n7261), .A(n8854), .ZN(n7260) );
  NAND2_X1 U7917 ( .A1(n11663), .A2(n7120), .ZN(n7122) );
  NOR2_X1 U7918 ( .A1(n7261), .A2(n7121), .ZN(n7120) );
  INV_X1 U7919 ( .A(n12397), .ZN(n7121) );
  NOR2_X2 U7920 ( .A1(n11917), .A2(n14039), .ZN(n14510) );
  AOI21_X1 U7921 ( .B1(n7113), .B2(n7112), .A(n6791), .ZN(n7111) );
  OAI21_X1 U7922 ( .B1(n14340), .B2(n14339), .A(n8867), .ZN(n9752) );
  NAND2_X1 U7923 ( .A1(n14351), .A2(n8821), .ZN(n8867) );
  NAND2_X1 U7924 ( .A1(n8377), .A2(SI_22_), .ZN(n8380) );
  NAND2_X1 U7925 ( .A1(n8738), .A2(n8737), .ZN(n8740) );
  OR2_X1 U7926 ( .A1(n8692), .A2(n8691), .ZN(n8705) );
  NAND2_X1 U7927 ( .A1(n7405), .A2(n8352), .ZN(n8660) );
  NAND2_X1 U7928 ( .A1(n8640), .A2(n7409), .ZN(n7405) );
  NAND2_X1 U7929 ( .A1(n8500), .A2(n7399), .ZN(n7401) );
  XNOR2_X1 U7930 ( .A(n8516), .B(n8515), .ZN(n9858) );
  NAND2_X1 U7931 ( .A1(n8512), .A2(n8511), .ZN(n8516) );
  NAND2_X1 U7932 ( .A1(n14707), .A2(n14706), .ZN(n14709) );
  AND2_X1 U7933 ( .A1(n6948), .A2(n6951), .ZN(n14744) );
  NAND2_X1 U7934 ( .A1(n14741), .A2(n14740), .ZN(n6948) );
  NOR2_X1 U7935 ( .A1(n6836), .A2(n14756), .ZN(n7088) );
  NOR2_X1 U7936 ( .A1(n9735), .A2(n9734), .ZN(n9736) );
  AND2_X1 U7937 ( .A1(n13205), .A2(n13206), .ZN(n13357) );
  NAND2_X1 U7938 ( .A1(n7574), .A2(n7573), .ZN(n7572) );
  NAND2_X1 U7939 ( .A1(n13353), .A2(n13359), .ZN(n7574) );
  NAND2_X1 U7940 ( .A1(n8256), .A2(n8230), .ZN(n7571) );
  NOR2_X1 U7941 ( .A1(n14863), .A2(n14748), .ZN(n14780) );
  NOR2_X1 U7942 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n14862), .ZN(n14748) );
  NAND2_X1 U7943 ( .A1(n9217), .A2(n9219), .ZN(n7623) );
  NAND2_X1 U7944 ( .A1(n12386), .A2(n12383), .ZN(n7173) );
  NAND2_X1 U7945 ( .A1(n12429), .A2(n12428), .ZN(n7181) );
  AOI21_X1 U7946 ( .B1(n6801), .B2(n12435), .A(n7186), .ZN(n7185) );
  NOR2_X1 U7947 ( .A1(n12436), .A2(n12438), .ZN(n7186) );
  NAND2_X1 U7948 ( .A1(n7432), .A2(n12434), .ZN(n12436) );
  NOR2_X1 U7949 ( .A1(n12439), .A2(n12435), .ZN(n7187) );
  NAND2_X1 U7950 ( .A1(n9334), .A2(n7633), .ZN(n7632) );
  OAI21_X1 U7951 ( .B1(n12445), .B2(n7437), .A(n6800), .ZN(n12451) );
  INV_X1 U7952 ( .A(n7435), .ZN(n7437) );
  NAND2_X1 U7953 ( .A1(n7636), .A2(n9373), .ZN(n7635) );
  NAND2_X1 U7954 ( .A1(n12460), .A2(n12459), .ZN(n7182) );
  OR2_X1 U7955 ( .A1(n12488), .A2(n12489), .ZN(n12299) );
  NAND2_X1 U7956 ( .A1(n9405), .A2(n9403), .ZN(n7638) );
  NAND2_X1 U7957 ( .A1(n12489), .A2(n12498), .ZN(n12502) );
  INV_X1 U7958 ( .A(n8763), .ZN(n8381) );
  AND2_X1 U7959 ( .A1(n7415), .A2(n7153), .ZN(n7152) );
  INV_X1 U7960 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15605) );
  NAND2_X1 U7961 ( .A1(n7214), .A2(n7213), .ZN(n7212) );
  INV_X1 U7962 ( .A(n6757), .ZN(n6976) );
  NAND2_X1 U7963 ( .A1(n7330), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7329) );
  AND2_X1 U7964 ( .A1(n7220), .A2(n7219), .ZN(n11214) );
  NAND2_X1 U7965 ( .A1(n10963), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7219) );
  NAND2_X1 U7966 ( .A1(n7059), .A2(n6851), .ZN(n11566) );
  NAND2_X1 U7967 ( .A1(n7317), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7316) );
  NAND2_X1 U7968 ( .A1(n12076), .A2(n7317), .ZN(n7314) );
  OR2_X1 U7969 ( .A1(n13088), .A2(n12097), .ZN(n12098) );
  NAND2_X1 U7970 ( .A1(n7324), .A2(n7323), .ZN(n7322) );
  NAND2_X1 U7971 ( .A1(n12088), .A2(n7326), .ZN(n7323) );
  NAND2_X1 U7972 ( .A1(n13161), .A2(n7325), .ZN(n7324) );
  NOR2_X1 U7973 ( .A1(n13275), .A2(n13049), .ZN(n7562) );
  OR2_X1 U7974 ( .A1(n13275), .A2(n13285), .ZN(n12725) );
  OR2_X1 U7975 ( .A1(n13323), .A2(n13027), .ZN(n12714) );
  NOR2_X1 U7976 ( .A1(n7999), .A2(n7544), .ZN(n7543) );
  INV_X1 U7977 ( .A(n7974), .ZN(n7544) );
  NAND2_X1 U7978 ( .A1(n12633), .A2(n12629), .ZN(n15246) );
  OAI21_X1 U7979 ( .B1(n8101), .B2(n7390), .A(n7388), .ZN(n8125) );
  INV_X1 U7980 ( .A(n7391), .ZN(n7390) );
  AOI21_X1 U7981 ( .B1(n7389), .B2(n7391), .A(n6862), .ZN(n7388) );
  NOR2_X1 U7982 ( .A1(n8122), .A2(n7392), .ZN(n7391) );
  AND2_X1 U7983 ( .A1(n7669), .A2(n8046), .ZN(n8049) );
  INV_X1 U7984 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7669) );
  INV_X1 U7985 ( .A(n7386), .ZN(n7385) );
  OAI21_X1 U7986 ( .B1(n7980), .B2(n7387), .A(n8018), .ZN(n7386) );
  INV_X1 U7987 ( .A(n8000), .ZN(n7387) );
  INV_X1 U7988 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8006) );
  NOR2_X1 U7989 ( .A1(n6840), .A2(n6918), .ZN(n6917) );
  INV_X1 U7990 ( .A(n7855), .ZN(n6918) );
  OAI21_X1 U7991 ( .B1(n6840), .B2(n6916), .A(n7872), .ZN(n6915) );
  NAND2_X1 U7992 ( .A1(n7853), .A2(n7855), .ZN(n6916) );
  NAND2_X1 U7993 ( .A1(n6917), .A2(n6912), .ZN(n6911) );
  XNOR2_X1 U7994 ( .A(n15117), .B(n12033), .ZN(n10533) );
  INV_X1 U7995 ( .A(n10928), .ZN(n11494) );
  INV_X1 U7996 ( .A(n10516), .ZN(n10928) );
  INV_X1 U7997 ( .A(n11494), .ZN(n12029) );
  AND2_X1 U7998 ( .A1(n9497), .A2(n9532), .ZN(n7619) );
  NAND2_X1 U7999 ( .A1(n7147), .A2(n9532), .ZN(n7146) );
  NAND2_X1 U8000 ( .A1(n9524), .A2(n7148), .ZN(n7147) );
  NAND2_X1 U8001 ( .A1(n7617), .A2(n9497), .ZN(n7150) );
  NOR2_X1 U8002 ( .A1(n7622), .A2(n9441), .ZN(n7617) );
  OR2_X1 U8003 ( .A1(n7080), .A2(n13866), .ZN(n7079) );
  NOR2_X1 U8004 ( .A1(n7604), .A2(n7603), .ZN(n7602) );
  INV_X1 U8005 ( .A(n7606), .ZN(n7604) );
  INV_X1 U8006 ( .A(n13748), .ZN(n7603) );
  INV_X1 U8007 ( .A(n13907), .ZN(n7076) );
  INV_X1 U8008 ( .A(n9685), .ZN(n7474) );
  NOR2_X1 U8009 ( .A1(n9612), .A2(n7614), .ZN(n7613) );
  INV_X1 U8010 ( .A(n9679), .ZN(n7487) );
  NAND2_X1 U8011 ( .A1(n7577), .A2(n9676), .ZN(n7576) );
  NOR2_X1 U8012 ( .A1(n10987), .A2(n15213), .ZN(n10988) );
  OR2_X1 U8013 ( .A1(n13881), .A2(n13765), .ZN(n13754) );
  INV_X1 U8014 ( .A(n8962), .ZN(n7465) );
  INV_X1 U8015 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8968) );
  INV_X1 U8016 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8960) );
  OR2_X1 U8017 ( .A1(n10723), .A2(n7512), .ZN(n7507) );
  NOR2_X1 U8018 ( .A1(n11538), .A2(n7532), .ZN(n7531) );
  INV_X1 U8019 ( .A(n11290), .ZN(n7532) );
  OR2_X1 U8020 ( .A1(n14616), .A2(n12274), .ZN(n12257) );
  INV_X1 U8021 ( .A(n12162), .ZN(n7521) );
  INV_X1 U8022 ( .A(n7644), .ZN(n7518) );
  INV_X1 U8023 ( .A(n7519), .ZN(n6901) );
  AOI21_X1 U8024 ( .B1(n12162), .B2(n7520), .A(n6789), .ZN(n7519) );
  INV_X1 U8025 ( .A(n14072), .ZN(n7520) );
  OAI21_X1 U8026 ( .B1(n12471), .B2(n12470), .A(n12468), .ZN(n12469) );
  OR2_X1 U8027 ( .A1(n14632), .A2(n14066), .ZN(n14421) );
  OR2_X1 U8028 ( .A1(n14637), .A2(n14096), .ZN(n7433) );
  OR2_X1 U8029 ( .A1(n7268), .A2(n7115), .ZN(n7113) );
  NOR2_X1 U8030 ( .A1(n7258), .A2(n8847), .ZN(n7256) );
  INV_X1 U8031 ( .A(n8847), .ZN(n7255) );
  INV_X1 U8032 ( .A(n14152), .ZN(n12341) );
  OAI21_X1 U8033 ( .B1(n9446), .B2(n9445), .A(n9453), .ZN(n9492) );
  OAI21_X1 U8034 ( .B1(n8789), .B2(n8788), .A(n8391), .ZN(n8800) );
  NAND2_X1 U8035 ( .A1(n8388), .A2(n8387), .ZN(n8789) );
  NAND2_X1 U8036 ( .A1(n7164), .A2(n7160), .ZN(n8388) );
  AND2_X1 U8037 ( .A1(n7163), .A2(n7161), .ZN(n7160) );
  NOR2_X1 U8038 ( .A1(n8386), .A2(n7162), .ZN(n7161) );
  AND2_X1 U8039 ( .A1(n8387), .A2(n8385), .ZN(n8775) );
  NAND2_X1 U8040 ( .A1(n8740), .A2(n8376), .ZN(n8377) );
  INV_X1 U8041 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U8042 ( .A1(n8370), .A2(SI_20_), .ZN(n8372) );
  NAND2_X1 U8043 ( .A1(n7404), .A2(n7402), .ZN(n8675) );
  AOI21_X1 U8044 ( .B1(n7406), .B2(n7408), .A(n7403), .ZN(n7402) );
  INV_X1 U8045 ( .A(n8356), .ZN(n7403) );
  AND2_X1 U8046 ( .A1(n8513), .A2(n8499), .ZN(n7399) );
  NAND2_X1 U8047 ( .A1(n8308), .A2(SI_2_), .ZN(n6891) );
  NAND2_X1 U8048 ( .A1(n7129), .A2(n7394), .ZN(n8302) );
  NAND2_X1 U8049 ( .A1(n8317), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7129) );
  XNOR2_X1 U8050 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14685) );
  OAI21_X1 U8051 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n15605), .A(n14660), .ZN(
        n14683) );
  NAND2_X1 U8052 ( .A1(n14685), .A2(n14686), .ZN(n14660) );
  NAND2_X1 U8053 ( .A1(n6959), .A2(n14666), .ZN(n14667) );
  NAND2_X1 U8054 ( .A1(n14682), .A2(n14205), .ZN(n6959) );
  NOR2_X1 U8055 ( .A1(n7338), .A2(n13049), .ZN(n7336) );
  INV_X1 U8056 ( .A(n7339), .ZN(n7338) );
  NOR2_X1 U8057 ( .A1(n7344), .A2(n12854), .ZN(n7339) );
  INV_X1 U8058 ( .A(n7345), .ZN(n7344) );
  AND2_X1 U8059 ( .A1(n7349), .A2(n7346), .ZN(n7345) );
  INV_X1 U8060 ( .A(n13036), .ZN(n7346) );
  NOR2_X1 U8061 ( .A1(n12858), .A2(n13233), .ZN(n7343) );
  AND2_X1 U8062 ( .A1(n12870), .A2(n11742), .ZN(n7365) );
  OR2_X1 U8063 ( .A1(n7910), .A2(n7697), .ZN(n7701) );
  INV_X1 U8064 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10212) );
  NAND2_X1 U8065 ( .A1(n7991), .A2(n7990), .ZN(n8010) );
  INV_X1 U8066 ( .A(n7992), .ZN(n7991) );
  INV_X1 U8067 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15587) );
  NAND2_X1 U8068 ( .A1(n11739), .A2(n7366), .ZN(n12982) );
  NOR2_X1 U8069 ( .A1(n12985), .A2(n7367), .ZN(n7366) );
  INV_X1 U8070 ( .A(n11738), .ZN(n7367) );
  NAND2_X1 U8071 ( .A1(n7931), .A2(n7930), .ZN(n7950) );
  INV_X1 U8072 ( .A(n7932), .ZN(n7931) );
  OAI21_X1 U8073 ( .B1(n12998), .B2(n7357), .A(n7355), .ZN(n12847) );
  AOI21_X1 U8074 ( .B1(n7358), .B2(n7356), .A(n6847), .ZN(n7355) );
  INV_X1 U8075 ( .A(n7358), .ZN(n7357) );
  NAND2_X1 U8076 ( .A1(n7334), .A2(n10426), .ZN(n10427) );
  AND2_X1 U8077 ( .A1(n10311), .A2(n10308), .ZN(n7334) );
  NAND2_X1 U8078 ( .A1(n11114), .A2(n11113), .ZN(n12953) );
  NAND2_X1 U8079 ( .A1(n7350), .A2(n6842), .ZN(n7349) );
  INV_X1 U8080 ( .A(n12934), .ZN(n7350) );
  NAND2_X1 U8081 ( .A1(n7348), .A2(n7347), .ZN(n7353) );
  OR2_X1 U8082 ( .A1(n13458), .A2(n8286), .ZN(n10319) );
  AND4_X1 U8083 ( .A1(n7775), .A2(n7774), .A3(n7773), .A4(n7772), .ZN(n11117)
         );
  NAND2_X1 U8084 ( .A1(n10142), .A2(n10141), .ZN(n10412) );
  OR2_X1 U8085 ( .A1(n10130), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10142) );
  NAND2_X1 U8086 ( .A1(n10130), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U8087 ( .A1(n6976), .A2(n6814), .ZN(n6974) );
  OR2_X1 U8088 ( .A1(n10210), .A2(n10216), .ZN(n7333) );
  NAND2_X1 U8089 ( .A1(n6753), .A2(n7217), .ZN(n10218) );
  OAI22_X1 U8090 ( .A1(n10201), .A2(n10200), .B1(n10213), .B2(n10199), .ZN(
        n10204) );
  NAND2_X1 U8091 ( .A1(n7333), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7332) );
  NOR2_X1 U8092 ( .A1(n10499), .A2(n10480), .ZN(n10483) );
  OR2_X1 U8093 ( .A1(n10491), .A2(n10458), .ZN(n7055) );
  NAND2_X1 U8094 ( .A1(n10460), .A2(n6837), .ZN(n7051) );
  NAND2_X1 U8095 ( .A1(n7053), .A2(n6837), .ZN(n7052) );
  OR2_X1 U8096 ( .A1(n10950), .A2(n10952), .ZN(n7312) );
  NAND2_X1 U8097 ( .A1(n7061), .A2(n7060), .ZN(n7059) );
  INV_X1 U8098 ( .A(n11211), .ZN(n7060) );
  NAND2_X1 U8099 ( .A1(n10959), .A2(n6841), .ZN(n6995) );
  AND2_X1 U8100 ( .A1(n7209), .A2(n7208), .ZN(n11560) );
  NAND2_X1 U8101 ( .A1(n11464), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7208) );
  INV_X1 U8102 ( .A(n11453), .ZN(n7209) );
  NAND2_X1 U8103 ( .A1(n6991), .A2(n6990), .ZN(n11576) );
  NAND2_X1 U8104 ( .A1(n6994), .A2(n6992), .ZN(n6990) );
  NAND2_X1 U8105 ( .A1(n10959), .A2(n6854), .ZN(n6991) );
  NOR2_X1 U8106 ( .A1(n12056), .A2(n7207), .ZN(n12057) );
  AND2_X1 U8107 ( .A1(n12073), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7207) );
  NOR2_X1 U8108 ( .A1(n13087), .A2(n6979), .ZN(n13088) );
  NAND2_X1 U8109 ( .A1(n6981), .A2(n6980), .ZN(n6979) );
  INV_X1 U8110 ( .A(n13086), .ZN(n6980) );
  INV_X1 U8111 ( .A(n13090), .ZN(n6981) );
  NAND2_X1 U8112 ( .A1(n12059), .A2(n12094), .ZN(n12061) );
  OR2_X1 U8113 ( .A1(n13115), .A2(n12064), .ZN(n12065) );
  NAND2_X1 U8114 ( .A1(n7206), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13157) );
  INV_X1 U8115 ( .A(n13136), .ZN(n7206) );
  NOR2_X1 U8116 ( .A1(n13201), .A2(n7298), .ZN(n7297) );
  INV_X1 U8117 ( .A(n8248), .ZN(n7298) );
  OR2_X1 U8118 ( .A1(n8163), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8180) );
  OR2_X1 U8119 ( .A1(n8180), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8203) );
  INV_X1 U8120 ( .A(n13233), .ZN(n13197) );
  NAND2_X1 U8121 ( .A1(n7550), .A2(n8171), .ZN(n13194) );
  NAND2_X1 U8122 ( .A1(n13228), .A2(n12792), .ZN(n8247) );
  NAND2_X1 U8123 ( .A1(n6882), .A2(n7561), .ZN(n7553) );
  NAND2_X1 U8124 ( .A1(n7563), .A2(n7560), .ZN(n13255) );
  INV_X1 U8125 ( .A(n7562), .ZN(n7560) );
  NAND2_X1 U8126 ( .A1(n7564), .A2(n6758), .ZN(n7563) );
  INV_X1 U8127 ( .A(n6882), .ZN(n7564) );
  NAND2_X1 U8128 ( .A1(n13264), .A2(n13263), .ZN(n13266) );
  AND2_X1 U8129 ( .A1(n12730), .A2(n12729), .ZN(n13263) );
  INV_X1 U8130 ( .A(n7007), .ZN(n7006) );
  AND4_X1 U8132 ( .A1(n8036), .A2(n8035), .A3(n8034), .A4(n8033), .ZN(n13315)
         );
  AND2_X1 U8133 ( .A1(n8241), .A2(n12701), .ZN(n7020) );
  AND2_X1 U8134 ( .A1(n12704), .A2(n12701), .ZN(n12789) );
  AND4_X1 U8135 ( .A1(n8015), .A2(n8014), .A3(n8013), .A4(n8012), .ZN(n12944)
         );
  AND2_X1 U8136 ( .A1(n12698), .A2(n12697), .ZN(n11848) );
  AND2_X1 U8137 ( .A1(n12691), .A2(n12696), .ZN(n12689) );
  AOI21_X1 U8138 ( .B1(n7279), .B2(n6743), .A(n7019), .ZN(n11647) );
  INV_X1 U8139 ( .A(n12680), .ZN(n7019) );
  AND4_X1 U8140 ( .A1(n7956), .A2(n7955), .A3(n7954), .A4(n7953), .ZN(n11941)
         );
  INV_X1 U8141 ( .A(n8238), .ZN(n12781) );
  AND4_X1 U8142 ( .A1(n7852), .A2(n7851), .A3(n7850), .A4(n7849), .ZN(n11740)
         );
  AND4_X1 U8143 ( .A1(n7883), .A2(n7882), .A3(n7881), .A4(n7880), .ZN(n13012)
         );
  AND4_X1 U8144 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n11744)
         );
  NAND2_X1 U8145 ( .A1(n7844), .A2(n7843), .ZN(n11252) );
  INV_X1 U8146 ( .A(n7012), .ZN(n7011) );
  OAI21_X1 U8147 ( .B1(n7274), .B2(n7843), .A(n12658), .ZN(n7012) );
  NOR2_X1 U8148 ( .A1(n12777), .A2(n12766), .ZN(n7273) );
  AOI21_X1 U8149 ( .B1(n12650), .B2(n7276), .A(n7275), .ZN(n7274) );
  INV_X1 U8150 ( .A(n12651), .ZN(n7276) );
  INV_X1 U8151 ( .A(n12653), .ZN(n7275) );
  AND3_X1 U8152 ( .A1(n7842), .A2(n7841), .A3(n7840), .ZN(n11241) );
  NAND2_X1 U8153 ( .A1(n10734), .A2(n10733), .ZN(n10736) );
  AND4_X1 U8154 ( .A1(n7831), .A2(n7830), .A3(n7829), .A4(n7828), .ZN(n11072)
         );
  AND4_X1 U8155 ( .A1(n7795), .A2(n7794), .A3(n7793), .A4(n7792), .ZN(n10918)
         );
  AND2_X1 U8156 ( .A1(n8228), .A2(n8227), .ZN(n15242) );
  NAND2_X1 U8157 ( .A1(n12617), .A2(n12618), .ZN(n15295) );
  AND2_X1 U8158 ( .A1(n10236), .A2(n13459), .ZN(n10671) );
  INV_X1 U8159 ( .A(n15242), .ZN(n13312) );
  INV_X1 U8160 ( .A(n15295), .ZN(n15302) );
  INV_X1 U8161 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U8162 ( .A1(n7567), .A2(n7565), .ZN(n8268) );
  NAND2_X1 U8163 ( .A1(n8159), .A2(n8158), .ZN(n8174) );
  NAND2_X1 U8164 ( .A1(n8261), .A2(n7677), .ZN(n8265) );
  AND2_X1 U8165 ( .A1(n7362), .A2(n8290), .ZN(n7361) );
  NOR2_X1 U8166 ( .A1(n7664), .A2(n13462), .ZN(n8258) );
  INV_X1 U8167 ( .A(n8259), .ZN(n8261) );
  OR2_X1 U8168 ( .A1(n8125), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U8169 ( .A1(n8098), .A2(n8097), .ZN(n8101) );
  NAND2_X1 U8170 ( .A1(n8101), .A2(n8100), .ZN(n8114) );
  NAND2_X1 U8171 ( .A1(n8084), .A2(n8083), .ZN(n8098) );
  NAND2_X1 U8172 ( .A1(n8067), .A2(n8066), .ZN(n8081) );
  NAND2_X1 U8173 ( .A1(n8043), .A2(n8042), .ZN(n8064) );
  NAND2_X1 U8174 ( .A1(n6907), .A2(n7978), .ZN(n7981) );
  NAND2_X1 U8175 ( .A1(n7981), .A2(n7980), .ZN(n8001) );
  NAND2_X1 U8176 ( .A1(n7939), .A2(n10079), .ZN(n7940) );
  NAND2_X1 U8177 ( .A1(n7923), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7941) );
  XNOR2_X1 U8178 ( .A(n7939), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n7923) );
  INV_X1 U8179 ( .A(n7907), .ZN(n6933) );
  NAND2_X1 U8180 ( .A1(n7888), .A2(n7887), .ZN(n7904) );
  NAND2_X1 U8181 ( .A1(n7886), .A2(n7885), .ZN(n7888) );
  AND2_X1 U8182 ( .A1(n9867), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7853) );
  OAI21_X1 U8183 ( .B1(n7834), .B2(n7833), .A(n6910), .ZN(n7854) );
  INV_X1 U8184 ( .A(n6912), .ZN(n6910) );
  NAND2_X1 U8185 ( .A1(n7799), .A2(n7798), .ZN(n7817) );
  NAND2_X1 U8186 ( .A1(n7797), .A2(n7796), .ZN(n7799) );
  XNOR2_X1 U8187 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7776) );
  NAND2_X1 U8188 ( .A1(n6807), .A2(n7737), .ZN(n6926) );
  NOR2_X1 U8189 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7292) );
  NAND2_X1 U8190 ( .A1(n7720), .A2(n7719), .ZN(n7736) );
  NOR2_X1 U8191 ( .A1(n13480), .A2(n15134), .ZN(n11996) );
  AOI21_X1 U8192 ( .B1(n7449), .B2(n13469), .A(n6803), .ZN(n7448) );
  NAND2_X1 U8193 ( .A1(n10547), .A2(n10543), .ZN(n10544) );
  AND2_X1 U8194 ( .A1(n7136), .A2(n13511), .ZN(n7135) );
  XNOR2_X1 U8195 ( .A(n11200), .B(n12033), .ZN(n12575) );
  NAND2_X1 U8196 ( .A1(n11688), .A2(n6759), .ZN(n7461) );
  INV_X1 U8197 ( .A(n11690), .ZN(n7459) );
  INV_X1 U8198 ( .A(n13564), .ZN(n7141) );
  NAND2_X1 U8199 ( .A1(n7140), .A2(n7141), .ZN(n7139) );
  INV_X1 U8200 ( .A(n7463), .ZN(n7140) );
  AND2_X1 U8201 ( .A1(n11504), .A2(n11499), .ZN(n7134) );
  INV_X1 U8202 ( .A(n15001), .ZN(n11504) );
  NAND2_X1 U8203 ( .A1(n9357), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9375) );
  INV_X1 U8204 ( .A(n9359), .ZN(n9357) );
  INV_X1 U8205 ( .A(n11086), .ZN(n11015) );
  XNOR2_X1 U8206 ( .A(n12575), .B(n11490), .ZN(n11026) );
  XNOR2_X1 U8207 ( .A(n7462), .B(n9797), .ZN(n13504) );
  INV_X1 U8208 ( .A(n12048), .ZN(n7462) );
  AND2_X1 U8209 ( .A1(n7131), .A2(n10527), .ZN(n10539) );
  INV_X1 U8210 ( .A(n10526), .ZN(n7131) );
  XNOR2_X1 U8211 ( .A(n13857), .B(n12036), .ZN(n9630) );
  NAND2_X1 U8212 ( .A1(n9505), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8996) );
  NAND2_X1 U8213 ( .A1(n9504), .A2(n9503), .ZN(n13643) );
  NAND2_X1 U8214 ( .A1(n7601), .A2(n7606), .ZN(n7600) );
  NAND2_X1 U8215 ( .A1(n9625), .A2(n7607), .ZN(n7601) );
  NAND2_X1 U8216 ( .A1(n7602), .A2(n13743), .ZN(n7599) );
  INV_X1 U8217 ( .A(n7484), .ZN(n7482) );
  NAND2_X1 U8218 ( .A1(n7485), .A2(n13558), .ZN(n7484) );
  NAND2_X1 U8219 ( .A1(n7040), .A2(n6746), .ZN(n13771) );
  NAND2_X1 U8220 ( .A1(n13808), .A2(n6780), .ZN(n7040) );
  NOR2_X1 U8221 ( .A1(n7047), .A2(n6744), .ZN(n7041) );
  NOR2_X1 U8222 ( .A1(n13794), .A2(n13891), .ZN(n13785) );
  AND2_X1 U8223 ( .A1(n13907), .A2(n13590), .ZN(n7492) );
  OR2_X1 U8224 ( .A1(n10683), .A2(n9370), .ZN(n9303) );
  NAND2_X1 U8225 ( .A1(n9618), .A2(n7584), .ZN(n7579) );
  INV_X1 U8226 ( .A(n7582), .ZN(n7581) );
  OR2_X1 U8227 ( .A1(n11819), .A2(n9689), .ZN(n7493) );
  AND2_X1 U8228 ( .A1(n9616), .A2(n7587), .ZN(n7585) );
  AOI21_X1 U8229 ( .B1(n11803), .B2(n11804), .A(n9687), .ZN(n11817) );
  AND2_X1 U8230 ( .A1(n11817), .A2(n11816), .ZN(n11819) );
  AND2_X1 U8231 ( .A1(n9610), .A2(n9609), .ZN(n7614) );
  NAND2_X1 U8232 ( .A1(n9608), .A2(n9607), .ZN(n11177) );
  AOI21_X1 U8233 ( .B1(n11173), .B2(n11174), .A(n9683), .ZN(n11266) );
  NOR2_X1 U8234 ( .A1(n11179), .A2(n14815), .ZN(n11267) );
  NAND2_X1 U8235 ( .A1(n10979), .A2(n10981), .ZN(n7488) );
  OR2_X1 U8236 ( .A1(n9866), .A2(n9370), .ZN(n9122) );
  NOR2_X1 U8237 ( .A1(n15117), .A2(n10824), .ZN(n11096) );
  AOI21_X1 U8238 ( .B1(n7593), .B2(n10639), .A(n6773), .ZN(n7592) );
  NAND2_X1 U8239 ( .A1(n7031), .A2(n7030), .ZN(n9672) );
  NAND2_X1 U8240 ( .A1(n7034), .A2(n9670), .ZN(n7030) );
  NAND2_X1 U8241 ( .A1(n10856), .A2(n7032), .ZN(n7031) );
  INV_X1 U8242 ( .A(n7036), .ZN(n7034) );
  INV_X1 U8243 ( .A(n13678), .ZN(n13857) );
  NAND2_X1 U8244 ( .A1(n9705), .A2(n10975), .ZN(n15201) );
  XNOR2_X1 U8245 ( .A(n9793), .B(n9704), .ZN(n9705) );
  NAND2_X1 U8246 ( .A1(n9825), .A2(n9501), .ZN(n7039) );
  INV_X1 U8247 ( .A(n15215), .ZN(n15196) );
  AND2_X1 U8248 ( .A1(n15166), .A2(n9789), .ZN(n11970) );
  NAND2_X1 U8249 ( .A1(n8940), .A2(n8939), .ZN(n7608) );
  NAND2_X1 U8250 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n8935), .ZN(n8939) );
  OR2_X1 U8251 ( .A1(n9098), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9118) );
  INV_X1 U8252 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9016) );
  INV_X1 U8253 ( .A(n7507), .ZN(n7511) );
  OR2_X1 U8254 ( .A1(n10721), .A2(n10720), .ZN(n7513) );
  AND2_X1 U8255 ( .A1(n13966), .A2(n7498), .ZN(n7497) );
  OR2_X1 U8256 ( .A1(n14107), .A2(n12260), .ZN(n7498) );
  AND2_X1 U8257 ( .A1(n6904), .A2(n6903), .ZN(n7530) );
  NAND2_X1 U8258 ( .A1(n11536), .A2(n6905), .ZN(n6903) );
  OR2_X1 U8259 ( .A1(n11538), .A2(n7534), .ZN(n6904) );
  AND2_X1 U8260 ( .A1(n7500), .A2(n14056), .ZN(n7499) );
  OAI22_X1 U8261 ( .A1(n10622), .A2(n10617), .B1(n12316), .B2(n12274), .ZN(
        n10718) );
  NAND2_X1 U8262 ( .A1(n14042), .A2(n12185), .ZN(n7522) );
  NOR2_X1 U8263 ( .A1(n14271), .A2(n14272), .ZN(n14285) );
  XNOR2_X1 U8264 ( .A(n14283), .B(n14282), .ZN(n14271) );
  INV_X1 U8265 ( .A(n14616), .ZN(n14358) );
  XNOR2_X1 U8266 ( .A(n14358), .B(n14133), .ZN(n14361) );
  NAND2_X1 U8267 ( .A1(n14368), .A2(n14376), .ZN(n14367) );
  AND2_X1 U8268 ( .A1(n12537), .A2(n8864), .ZN(n7116) );
  NOR2_X1 U8269 ( .A1(n8863), .A2(n7238), .ZN(n7237) );
  INV_X1 U8270 ( .A(n8774), .ZN(n7238) );
  NAND2_X1 U8271 ( .A1(n7265), .A2(n7263), .ZN(n14388) );
  NOR2_X1 U8272 ( .A1(n14385), .A2(n7264), .ZN(n7263) );
  INV_X1 U8273 ( .A(n8862), .ZN(n7264) );
  NAND2_X1 U8274 ( .A1(n7119), .A2(n7117), .ZN(n14420) );
  AND2_X1 U8275 ( .A1(n14442), .A2(n7118), .ZN(n7117) );
  NAND2_X1 U8276 ( .A1(n14456), .A2(n8858), .ZN(n7118) );
  NAND2_X1 U8277 ( .A1(n7197), .A2(n14446), .ZN(n7196) );
  INV_X1 U8278 ( .A(n7198), .ZN(n7197) );
  OR2_X1 U8279 ( .A1(n14457), .A2(n14456), .ZN(n14459) );
  NAND2_X1 U8280 ( .A1(n7122), .A2(n6786), .ZN(n14505) );
  OR2_X1 U8281 ( .A1(n14647), .A2(n11666), .ZN(n12411) );
  AOI21_X1 U8282 ( .B1(n8659), .B2(n12402), .A(n6792), .ZN(n7239) );
  NAND2_X1 U8283 ( .A1(n11663), .A2(n12397), .ZN(n11835) );
  NAND2_X1 U8284 ( .A1(n11835), .A2(n11834), .ZN(n11833) );
  AND2_X1 U8285 ( .A1(n7113), .A2(n12527), .ZN(n7114) );
  INV_X1 U8286 ( .A(n8851), .ZN(n7115) );
  INV_X1 U8287 ( .A(n11602), .ZN(n12527) );
  XNOR2_X1 U8288 ( .A(n12377), .B(n6885), .ZN(n11602) );
  AND2_X1 U8289 ( .A1(n8851), .A2(n8574), .ZN(n12526) );
  NOR2_X1 U8290 ( .A1(n11481), .A2(n7270), .ZN(n7269) );
  INV_X1 U8291 ( .A(n8849), .ZN(n7270) );
  OR2_X1 U8292 ( .A1(n11414), .A2(n12509), .ZN(n14909) );
  OR2_X1 U8293 ( .A1(n12297), .A2(n12489), .ZN(n11414) );
  NAND2_X1 U8294 ( .A1(n12486), .A2(n12485), .ZN(n14313) );
  INV_X1 U8295 ( .A(n7127), .ZN(n7125) );
  AOI21_X1 U8296 ( .B1(n10252), .B2(n8921), .A(n10253), .ZN(n11303) );
  INV_X1 U8297 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8410) );
  INV_X1 U8298 ( .A(n7651), .ZN(n7252) );
  XNOR2_X1 U8299 ( .A(n8789), .B(n8788), .ZN(n11719) );
  NAND2_X1 U8300 ( .A1(n7166), .A2(n7165), .ZN(n9369) );
  INV_X1 U8301 ( .A(n9366), .ZN(n7165) );
  INV_X1 U8302 ( .A(n8828), .ZN(n8831) );
  XNOR2_X1 U8303 ( .A(n8646), .B(n8645), .ZN(n10394) );
  NAND2_X1 U8304 ( .A1(n7411), .A2(n7415), .ZN(n8588) );
  OR2_X1 U8305 ( .A1(n8560), .A2(n7418), .ZN(n7411) );
  NAND2_X1 U8306 ( .A1(n7421), .A2(n7422), .ZN(n8576) );
  NAND2_X1 U8307 ( .A1(n8560), .A2(n7423), .ZN(n7421) );
  OR2_X1 U8308 ( .A1(n8327), .A2(n8328), .ZN(n7400) );
  AND2_X1 U8309 ( .A1(n8511), .A2(n8514), .ZN(n8328) );
  NAND2_X1 U8310 ( .A1(n8481), .A2(n8321), .ZN(n6887) );
  NAND2_X1 U8311 ( .A1(n8499), .A2(n8500), .ZN(n8512) );
  NAND2_X1 U8312 ( .A1(n8301), .A2(n7697), .ZN(n8303) );
  INV_X1 U8313 ( .A(n8302), .ZN(n8301) );
  NAND2_X1 U8314 ( .A1(n8302), .A2(SI_1_), .ZN(n8305) );
  AND2_X1 U8315 ( .A1(n7250), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14686) );
  INV_X1 U8316 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7250) );
  INV_X1 U8317 ( .A(n7081), .ZN(n14705) );
  NAND2_X1 U8318 ( .A1(n6957), .A2(n14672), .ZN(n14681) );
  NAND2_X1 U8319 ( .A1(n14710), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6957) );
  AOI21_X1 U8320 ( .B1(n14729), .B2(n14728), .A(n14847), .ZN(n14732) );
  OAI21_X1 U8321 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14678), .A(n14677), .ZN(
        n14735) );
  XNOR2_X1 U8322 ( .A(n14751), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n14752) );
  NAND2_X1 U8323 ( .A1(n8179), .A2(n8178), .ZN(n13358) );
  INV_X1 U8324 ( .A(n13053), .ZN(n12824) );
  XNOR2_X1 U8325 ( .A(n7348), .B(n12850), .ZN(n12973) );
  NAND2_X1 U8326 ( .A1(n11243), .A2(n11242), .ZN(n11739) );
  AND2_X1 U8327 ( .A1(n8137), .A2(n8136), .ZN(n13256) );
  NAND2_X1 U8328 ( .A1(n8009), .A2(n8008), .ZN(n12968) );
  AND3_X1 U8329 ( .A1(n7863), .A2(n7862), .A3(n7861), .ZN(n12988) );
  AND3_X1 U8330 ( .A1(n8121), .A2(n8120), .A3(n8119), .ZN(n13273) );
  NAND2_X1 U8331 ( .A1(n8028), .A2(n8027), .ZN(n13340) );
  OR2_X1 U8332 ( .A1(n10329), .A2(n8199), .ZN(n8028) );
  NAND2_X1 U8333 ( .A1(n7966), .A2(n7965), .ZN(n11946) );
  AOI21_X1 U8334 ( .B1(n12761), .B2(n15240), .A(n6921), .ZN(n6920) );
  NOR2_X1 U8335 ( .A1(n12802), .A2(n6922), .ZN(n6921) );
  XNOR2_X1 U8336 ( .A(n12801), .B(n12800), .ZN(n6922) );
  NAND2_X1 U8337 ( .A1(n12805), .A2(n12804), .ZN(n6919) );
  INV_X1 U8338 ( .A(n13273), .ZN(n13249) );
  INV_X1 U8339 ( .A(n10918), .ZN(n13058) );
  NAND2_X1 U8340 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7698) );
  NAND2_X1 U8341 ( .A1(n6977), .A2(n6978), .ZN(n6975) );
  INV_X1 U8342 ( .A(n10422), .ZN(n6978) );
  INV_X1 U8343 ( .A(n10421), .ZN(n6977) );
  XNOR2_X1 U8344 ( .A(n11560), .B(n11568), .ZN(n11454) );
  NOR2_X1 U8345 ( .A1(n11454), .A2(n11196), .ZN(n11561) );
  XNOR2_X1 U8346 ( .A(n12057), .B(n13072), .ZN(n13063) );
  NOR2_X1 U8347 ( .A1(n13063), .A2(n7929), .ZN(n13062) );
  XNOR2_X1 U8348 ( .A(n12061), .B(n12060), .ZN(n13098) );
  AOI21_X1 U8349 ( .B1(n13157), .B2(n13156), .A(n13155), .ZN(n13160) );
  XNOR2_X1 U8350 ( .A(n13162), .B(n13161), .ZN(n7064) );
  NAND2_X1 U8351 ( .A1(n13166), .A2(n13167), .ZN(n7063) );
  NAND2_X1 U8352 ( .A1(n6989), .A2(n6988), .ZN(n6987) );
  INV_X1 U8353 ( .A(n13152), .ZN(n6989) );
  OR2_X1 U8354 ( .A1(n12109), .A2(n6860), .ZN(n6985) );
  NAND2_X1 U8355 ( .A1(n8128), .A2(n8127), .ZN(n13372) );
  NAND2_X1 U8356 ( .A1(n8116), .A2(n8115), .ZN(n13375) );
  OR2_X1 U8358 ( .A1(n8199), .A2(n7739), .ZN(n7743) );
  INV_X1 U8359 ( .A(n13341), .ZN(n13322) );
  INV_X1 U8360 ( .A(n7572), .ZN(n7570) );
  NAND2_X1 U8361 ( .A1(n13358), .A2(n13359), .ZN(n7023) );
  NAND2_X1 U8362 ( .A1(n15699), .A2(n15302), .ZN(n13409) );
  NOR2_X1 U8363 ( .A1(n7657), .A2(n9740), .ZN(n9741) );
  OAI21_X1 U8364 ( .B1(n12585), .B2(n8199), .A(n8200), .ZN(n13353) );
  NAND2_X1 U8365 ( .A1(n8231), .A2(n15309), .ZN(n7301) );
  NAND2_X1 U8366 ( .A1(n13357), .A2(n13356), .ZN(n13418) );
  NAND2_X1 U8367 ( .A1(n15309), .A2(n15302), .ZN(n13456) );
  XNOR2_X1 U8368 ( .A(n7692), .B(n7691), .ZN(n12806) );
  NAND2_X1 U8369 ( .A1(n6752), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7692) );
  INV_X1 U8370 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U8371 ( .A1(n9232), .A2(n9231), .ZN(n11505) );
  NAND2_X1 U8372 ( .A1(n9317), .A2(n9316), .ZN(n13896) );
  NOR2_X1 U8373 ( .A1(n7445), .A2(n14999), .ZN(n7443) );
  AND2_X1 U8374 ( .A1(n7448), .A2(n7446), .ZN(n7445) );
  INV_X1 U8375 ( .A(n7449), .ZN(n7446) );
  NAND2_X1 U8376 ( .A1(n7448), .A2(n7451), .ZN(n7447) );
  NAND2_X1 U8377 ( .A1(n7452), .A2(n6751), .ZN(n7451) );
  INV_X1 U8378 ( .A(n13469), .ZN(n7452) );
  OR2_X1 U8379 ( .A1(n11134), .A2(n9370), .ZN(n9348) );
  INV_X1 U8380 ( .A(n15136), .ZN(n9661) );
  NOR2_X1 U8381 ( .A1(n12013), .A2(n12010), .ZN(n7457) );
  NAND2_X1 U8382 ( .A1(n9413), .A2(n9412), .ZN(n13582) );
  AND2_X1 U8383 ( .A1(n9895), .A2(n13957), .ZN(n15085) );
  AND2_X1 U8384 ( .A1(n7072), .A2(n7071), .ZN(n13844) );
  AOI21_X1 U8385 ( .B1(n13657), .B2(n13656), .A(n7472), .ZN(n9703) );
  AND2_X1 U8386 ( .A1(n9701), .A2(n13579), .ZN(n7472) );
  AND3_X1 U8387 ( .A1(n13659), .A2(n15134), .A3(n13658), .ZN(n13850) );
  AND2_X1 U8388 ( .A1(n15155), .A2(n10975), .ZN(n13835) );
  INV_X1 U8389 ( .A(n9511), .ZN(n10975) );
  INV_X1 U8390 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10681) );
  NAND2_X1 U8391 ( .A1(n9858), .A2(n6643), .ZN(n6906) );
  INV_X1 U8392 ( .A(n11700), .ZN(n11703) );
  NAND2_X1 U8393 ( .A1(n8665), .A2(n8664), .ZN(n14039) );
  INV_X1 U8394 ( .A(n14514), .ZN(n14587) );
  XNOR2_X1 U8395 ( .A(n11700), .B(n11701), .ZN(n11765) );
  NAND2_X1 U8396 ( .A1(n14007), .A2(n7644), .ZN(n14073) );
  NOR2_X1 U8397 ( .A1(n12555), .A2(n12554), .ZN(n7177) );
  INV_X1 U8398 ( .A(n13969), .ZN(n14133) );
  INV_X1 U8399 ( .A(n12344), .ZN(n14153) );
  NOR2_X1 U8400 ( .A1(n10084), .A2(n6784), .ZN(n14225) );
  NAND2_X1 U8401 ( .A1(n14225), .A2(n14226), .ZN(n14224) );
  NOR2_X1 U8402 ( .A1(n10275), .A2(n6964), .ZN(n14251) );
  AND2_X1 U8403 ( .A1(n10282), .A2(n10097), .ZN(n6964) );
  NAND2_X1 U8404 ( .A1(n14251), .A2(n14250), .ZN(n14249) );
  NOR2_X1 U8405 ( .A1(n10277), .A2(n10278), .ZN(n10565) );
  OR2_X1 U8406 ( .A1(n10683), .A2(n8741), .ZN(n8697) );
  NAND2_X1 U8407 ( .A1(n10342), .A2(n10341), .ZN(n14507) );
  INV_X1 U8408 ( .A(n12498), .ZN(n12509) );
  NAND2_X1 U8409 ( .A1(n7231), .A2(n9761), .ZN(n9765) );
  AND2_X1 U8410 ( .A1(n7126), .A2(n7124), .ZN(n9761) );
  INV_X1 U8411 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10682) );
  NAND2_X1 U8412 ( .A1(n14711), .A2(n14712), .ZN(n7107) );
  NAND2_X1 U8413 ( .A1(n14719), .A2(n14720), .ZN(n7103) );
  XNOR2_X1 U8414 ( .A(n14732), .B(n14733), .ZN(n14851) );
  OR2_X1 U8415 ( .A1(n14851), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7099) );
  NAND2_X1 U8416 ( .A1(n7094), .A2(n6839), .ZN(n7095) );
  NAND2_X1 U8417 ( .A1(n6762), .A2(n7093), .ZN(n7094) );
  NAND2_X1 U8418 ( .A1(n6762), .A2(n7092), .ZN(n7249) );
  NAND2_X1 U8419 ( .A1(n6962), .A2(n7088), .ZN(n7082) );
  INV_X1 U8420 ( .A(n14780), .ZN(n6962) );
  AOI21_X1 U8421 ( .B1(n14780), .B2(n6848), .A(n7085), .ZN(n7084) );
  OAI21_X1 U8422 ( .B1(n7086), .B2(n7090), .A(n7089), .ZN(n7085) );
  NAND2_X1 U8423 ( .A1(n6836), .A2(n14756), .ZN(n7089) );
  NAND2_X1 U8424 ( .A1(n7082), .A2(n15112), .ZN(n6961) );
  INV_X1 U8425 ( .A(n7084), .ZN(n6963) );
  NAND2_X1 U8426 ( .A1(n7083), .A2(n7088), .ZN(n7087) );
  NAND2_X1 U8427 ( .A1(n14780), .A2(n7090), .ZN(n7083) );
  INV_X1 U8428 ( .A(n9026), .ZN(n7641) );
  NAND2_X1 U8429 ( .A1(n7109), .A2(n12502), .ZN(n12301) );
  OR2_X1 U8430 ( .A1(n9087), .A2(n7630), .ZN(n7629) );
  INV_X1 U8431 ( .A(n9086), .ZN(n7630) );
  OAI21_X1 U8432 ( .B1(n12318), .B2(n12315), .A(n12314), .ZN(n12321) );
  NAND2_X1 U8433 ( .A1(n9123), .A2(n9125), .ZN(n7625) );
  MUX2_X1 U8434 ( .A(n12341), .B(n12340), .S(n12506), .Z(n12352) );
  NAND2_X1 U8435 ( .A1(n9181), .A2(n7627), .ZN(n7626) );
  NAND2_X1 U8436 ( .A1(n7190), .A2(n7189), .ZN(n7188) );
  AND2_X1 U8437 ( .A1(n12402), .A2(n12389), .ZN(n12390) );
  NOR2_X1 U8438 ( .A1(n12386), .A2(n12383), .ZN(n7174) );
  AND2_X1 U8439 ( .A1(n7173), .A2(n12388), .ZN(n7172) );
  AOI21_X1 U8440 ( .B1(n12415), .B2(n6778), .A(n7181), .ZN(n7180) );
  NAND2_X1 U8441 ( .A1(n7431), .A2(n7429), .ZN(n12434) );
  NAND2_X1 U8442 ( .A1(n7433), .A2(n12491), .ZN(n7431) );
  NAND2_X1 U8443 ( .A1(n12431), .A2(n7430), .ZN(n7429) );
  AOI21_X1 U8444 ( .B1(n7185), .B2(n7187), .A(n6650), .ZN(n7184) );
  NAND2_X1 U8445 ( .A1(n12446), .A2(n7434), .ZN(n7435) );
  INV_X1 U8446 ( .A(n12444), .ZN(n7434) );
  NAND2_X1 U8447 ( .A1(n12447), .A2(n12444), .ZN(n7436) );
  INV_X1 U8448 ( .A(n12453), .ZN(n7427) );
  NOR2_X1 U8449 ( .A1(n12453), .A2(n12455), .ZN(n7428) );
  INV_X1 U8450 ( .A(n12071), .ZN(n7058) );
  INV_X1 U8451 ( .A(n13082), .ZN(n7317) );
  INV_X1 U8452 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7665) );
  INV_X1 U8453 ( .A(n8113), .ZN(n7392) );
  INV_X1 U8454 ( .A(n8100), .ZN(n7389) );
  AND2_X1 U8455 ( .A1(n9522), .A2(n9521), .ZN(n7149) );
  NAND2_X1 U8456 ( .A1(n13739), .A2(n13725), .ZN(n7080) );
  NOR2_X1 U8457 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n7025) );
  NOR2_X1 U8458 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7026) );
  AOI21_X1 U8459 ( .B1(n13982), .B2(n7504), .A(n7503), .ZN(n7502) );
  INV_X1 U8460 ( .A(n13983), .ZN(n7504) );
  INV_X1 U8461 ( .A(n14058), .ZN(n7503) );
  OAI21_X1 U8462 ( .B1(n8918), .B2(n12297), .A(n12296), .ZN(n12488) );
  NAND2_X1 U8463 ( .A1(n14158), .A2(n14964), .ZN(n12306) );
  AND2_X1 U8464 ( .A1(n8838), .A2(n10360), .ZN(n7267) );
  INV_X1 U8465 ( .A(n8775), .ZN(n8386) );
  INV_X1 U8466 ( .A(n8382), .ZN(n7162) );
  AND2_X1 U8467 ( .A1(n8363), .A2(n8362), .ZN(n6881) );
  INV_X1 U8468 ( .A(n8706), .ZN(n8363) );
  NOR2_X1 U8469 ( .A1(n8361), .A2(SI_18_), .ZN(n8364) );
  AOI21_X1 U8470 ( .B1(n7410), .B2(n8352), .A(n7407), .ZN(n7406) );
  INV_X1 U8471 ( .A(n8661), .ZN(n7407) );
  INV_X1 U8472 ( .A(n8352), .ZN(n7408) );
  NAND2_X1 U8473 ( .A1(n8353), .A2(n10083), .ZN(n8356) );
  NAND2_X1 U8474 ( .A1(n8543), .A2(n8336), .ZN(n7153) );
  NAND2_X1 U8475 ( .A1(n8333), .A2(SI_9_), .ZN(n8336) );
  NAND2_X1 U8476 ( .A1(n14879), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n6950) );
  INV_X1 U8477 ( .A(n6950), .ZN(n6945) );
  NOR2_X1 U8478 ( .A1(n6949), .A2(n6868), .ZN(n6947) );
  INV_X1 U8479 ( .A(n6946), .ZN(n6942) );
  OR2_X1 U8480 ( .A1(n6944), .A2(n6748), .ZN(n6939) );
  INV_X1 U8481 ( .A(n12997), .ZN(n7356) );
  NAND2_X1 U8482 ( .A1(n13195), .A2(n13217), .ZN(n12794) );
  AOI21_X1 U8483 ( .B1(n12756), .B2(n8227), .A(n12759), .ZN(n7377) );
  NAND2_X1 U8484 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10404), .ZN(n10131) );
  OR2_X1 U8485 ( .A1(n10131), .A2(P3_IR_REG_1__SCAN_IN), .ZN(n7648) );
  NAND2_X1 U8486 ( .A1(n7212), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7211) );
  INV_X1 U8487 ( .A(n7216), .ZN(n7215) );
  NAND2_X1 U8488 ( .A1(n7218), .A2(n10224), .ZN(n7217) );
  NAND2_X1 U8489 ( .A1(n7217), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7216) );
  AOI21_X1 U8490 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10477), .A(n10476), .ZN(
        n10479) );
  INV_X1 U8491 ( .A(n10458), .ZN(n7053) );
  INV_X1 U8492 ( .A(n11229), .ZN(n7001) );
  INV_X1 U8493 ( .A(n11459), .ZN(n6992) );
  AND2_X1 U8494 ( .A1(n7310), .A2(n7050), .ZN(n12084) );
  NAND2_X1 U8495 ( .A1(n12083), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U8496 ( .A1(n8148), .A2(n8147), .ZN(n8163) );
  INV_X1 U8497 ( .A(n8149), .ZN(n8148) );
  OR2_X1 U8498 ( .A1(n8129), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U8499 ( .A1(n8106), .A2(n8105), .ZN(n8117) );
  INV_X1 U8500 ( .A(n8107), .ZN(n8106) );
  OAI21_X1 U8501 ( .B1(n8243), .B2(n7008), .A(n12722), .ZN(n7007) );
  AND2_X1 U8502 ( .A1(n12725), .A2(n12726), .ZN(n12764) );
  OR2_X1 U8503 ( .A1(n8088), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8107) );
  INV_X1 U8504 ( .A(n7288), .ZN(n7287) );
  OAI21_X1 U8505 ( .B1(n8239), .B2(n7289), .A(n12689), .ZN(n7288) );
  AND2_X1 U8506 ( .A1(n7938), .A2(n7919), .ZN(n7547) );
  INV_X1 U8507 ( .A(n12672), .ZN(n7283) );
  INV_X1 U8508 ( .A(n7282), .ZN(n7281) );
  OAI21_X1 U8509 ( .B1(n8237), .B2(n7283), .A(n12781), .ZN(n7282) );
  NOR2_X1 U8510 ( .A1(n7015), .A2(n7843), .ZN(n7013) );
  INV_X1 U8511 ( .A(n7273), .ZN(n7015) );
  NAND2_X1 U8512 ( .A1(n7769), .A2(n10212), .ZN(n7789) );
  NAND2_X1 U8513 ( .A1(n6909), .A2(n6908), .ZN(n12750) );
  INV_X1 U8514 ( .A(n13353), .ZN(n6909) );
  NAND2_X1 U8515 ( .A1(n15245), .A2(n7747), .ZN(n10808) );
  AND2_X1 U8516 ( .A1(n12767), .A2(n10807), .ZN(n7747) );
  NAND2_X1 U8517 ( .A1(n11950), .A2(n15590), .ZN(n7368) );
  AND2_X1 U8518 ( .A1(n7565), .A2(n7303), .ZN(n7302) );
  INV_X1 U8519 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7303) );
  AND2_X1 U8520 ( .A1(n7677), .A2(n7566), .ZN(n7565) );
  INV_X1 U8521 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7566) );
  INV_X1 U8522 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7677) );
  AND2_X1 U8523 ( .A1(n8218), .A2(n7363), .ZN(n7362) );
  NOR2_X1 U8524 ( .A1(n7959), .A2(n10081), .ZN(n7379) );
  XNOR2_X1 U8525 ( .A(n12033), .B(n10654), .ZN(n10523) );
  AND2_X1 U8526 ( .A1(n9145), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9167) );
  INV_X1 U8527 ( .A(n12032), .ZN(n7450) );
  AND2_X1 U8528 ( .A1(n9167), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9183) );
  OAI21_X1 U8529 ( .B1(n11991), .B2(n11990), .A(n13510), .ZN(n11994) );
  OR2_X1 U8530 ( .A1(n13861), .A2(n13526), .ZN(n9627) );
  NAND2_X1 U8531 ( .A1(n9393), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9407) );
  INV_X1 U8532 ( .A(n9394), .ZN(n9393) );
  OAI21_X1 U8533 ( .B1(n7585), .B2(n7583), .A(n9620), .ZN(n7582) );
  AOI21_X1 U8534 ( .B1(n10894), .B2(n7578), .A(n6794), .ZN(n7577) );
  INV_X1 U8535 ( .A(n9601), .ZN(n7578) );
  NOR2_X1 U8536 ( .A1(n9127), .A2(n12118), .ZN(n9145) );
  INV_X1 U8537 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9089) );
  OR2_X1 U8538 ( .A1(n9090), .A2(n9089), .ZN(n9112) );
  NOR2_X1 U8539 ( .A1(n7591), .A2(n9671), .ZN(n7590) );
  INV_X1 U8540 ( .A(n9597), .ZN(n7591) );
  INV_X1 U8541 ( .A(n9598), .ZN(n7593) );
  NOR2_X1 U8542 ( .A1(n10858), .A2(n7035), .ZN(n7032) );
  NOR2_X1 U8543 ( .A1(n9050), .A2(n9049), .ZN(n9074) );
  NAND2_X1 U8544 ( .A1(n11591), .A2(n7077), .ZN(n13831) );
  NAND2_X1 U8545 ( .A1(n8955), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U8546 ( .A1(n9565), .A2(n9566), .ZN(n9570) );
  INV_X1 U8547 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U8548 ( .A1(n7502), .A2(n7505), .ZN(n7500) );
  AND2_X1 U8549 ( .A1(n7502), .A2(n6897), .ZN(n6896) );
  NAND2_X1 U8550 ( .A1(n14083), .A2(n6898), .ZN(n6897) );
  NAND2_X1 U8551 ( .A1(n6896), .A2(n6899), .ZN(n6894) );
  AND2_X1 U8552 ( .A1(n12508), .A2(n12507), .ZN(n12550) );
  NAND2_X1 U8553 ( .A1(n12537), .A2(n8797), .ZN(n7227) );
  OR2_X1 U8554 ( .A1(n14570), .A2(n7199), .ZN(n7198) );
  NAND2_X1 U8555 ( .A1(n12411), .A2(n7262), .ZN(n7261) );
  INV_X1 U8556 ( .A(n12531), .ZN(n7262) );
  AND2_X1 U8557 ( .A1(n12530), .A2(n11602), .ZN(n8599) );
  AND2_X1 U8558 ( .A1(n12527), .A2(n7115), .ZN(n7112) );
  INV_X1 U8559 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8520) );
  INV_X1 U8560 ( .A(n8466), .ZN(n7235) );
  NAND2_X1 U8561 ( .A1(n12306), .A2(n7267), .ZN(n8839) );
  NAND2_X1 U8562 ( .A1(n8380), .A2(n6850), .ZN(n7163) );
  AND2_X1 U8563 ( .A1(n8380), .A2(n6843), .ZN(n7159) );
  NAND2_X1 U8564 ( .A1(n8360), .A2(n8359), .ZN(n8689) );
  NAND2_X1 U8565 ( .A1(n8349), .A2(SI_15_), .ZN(n8644) );
  NAND2_X1 U8566 ( .A1(n8341), .A2(n9881), .ZN(n8604) );
  NAND2_X1 U8567 ( .A1(n8345), .A2(SI_13_), .ZN(n8606) );
  INV_X1 U8568 ( .A(n8340), .ZN(n7416) );
  INV_X1 U8569 ( .A(n7423), .ZN(n7417) );
  INV_X1 U8570 ( .A(n7419), .ZN(n7418) );
  OR2_X1 U8571 ( .A1(n8577), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U8572 ( .A1(n8561), .A2(SI_10_), .ZN(n7422) );
  NAND2_X1 U8573 ( .A1(n7425), .A2(n7424), .ZN(n7423) );
  INV_X1 U8574 ( .A(n8561), .ZN(n7425) );
  NAND2_X1 U8575 ( .A1(n8528), .A2(n7397), .ZN(n7396) );
  INV_X1 U8576 ( .A(n8326), .ZN(n7171) );
  OAI21_X1 U8577 ( .B1(n9829), .B2(n6884), .A(n6883), .ZN(n8323) );
  NAND2_X1 U8578 ( .A1(n9829), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U8579 ( .A1(n8474), .A2(n8316), .ZN(n8481) );
  INV_X1 U8580 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7266) );
  OAI21_X1 U8581 ( .B1(n8317), .B2(n9824), .A(n8306), .ZN(n8308) );
  NAND2_X1 U8582 ( .A1(n14662), .A2(n14661), .ZN(n14663) );
  NAND2_X1 U8583 ( .A1(n14683), .A2(n14684), .ZN(n14662) );
  XNOR2_X1 U8584 ( .A(n14665), .B(n6960), .ZN(n14682) );
  INV_X1 U8585 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n6960) );
  NOR2_X1 U8586 ( .A1(n14674), .A2(n6956), .ZN(n6955) );
  AND2_X1 U8587 ( .A1(n14675), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n6956) );
  OAI21_X1 U8588 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n10030), .A(n14673), .ZN(
        n14714) );
  NAND2_X1 U8589 ( .A1(n14681), .A2(n14680), .ZN(n14673) );
  OAI22_X1 U8590 ( .A1(n14726), .A2(n14676), .B1(P1_ADDR_REG_11__SCAN_IN), 
        .B2(n14725), .ZN(n14731) );
  AND2_X1 U8591 ( .A1(n14740), .A2(n6950), .ZN(n6946) );
  NAND2_X1 U8592 ( .A1(n6938), .A2(n6937), .ZN(n14751) );
  OR2_X1 U8593 ( .A1(n6941), .A2(n6748), .ZN(n6937) );
  OR2_X1 U8594 ( .A1(n14741), .A2(n6939), .ZN(n6938) );
  AOI21_X1 U8595 ( .B1(n6942), .B2(n6943), .A(n6867), .ZN(n6941) );
  INV_X1 U8596 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10501) );
  NOR2_X1 U8597 ( .A1(n12914), .A2(n7359), .ZN(n7358) );
  INV_X1 U8598 ( .A(n12843), .ZN(n7359) );
  CLKBUF_X1 U8599 ( .A(n12920), .Z(n12921) );
  INV_X1 U8600 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11455) );
  INV_X1 U8601 ( .A(n10304), .ZN(n10306) );
  NAND2_X1 U8602 ( .A1(n10126), .A2(n6741), .ZN(n7018) );
  OR2_X1 U8603 ( .A1(n7910), .A2(n7722), .ZN(n7016) );
  OR2_X1 U8604 ( .A1(n10126), .A2(n7728), .ZN(n7017) );
  INV_X1 U8605 ( .A(n7950), .ZN(n7949) );
  OR2_X1 U8606 ( .A1(n7967), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7992) );
  AND2_X1 U8607 ( .A1(n12595), .A2(n12594), .ZN(n13173) );
  OR2_X1 U8608 ( .A1(n7754), .A2(n7730), .ZN(n7731) );
  NOR2_X1 U8609 ( .A1(n6776), .A2(n6738), .ZN(n7293) );
  NAND2_X1 U8610 ( .A1(n7750), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7704) );
  OR2_X1 U8611 ( .A1(n7754), .A2(n7702), .ZN(n7705) );
  OR2_X1 U8612 ( .A1(n10190), .A2(n7684), .ZN(n10192) );
  NAND2_X1 U8613 ( .A1(n7221), .A2(n10143), .ZN(n10144) );
  NAND2_X1 U8614 ( .A1(n10412), .A2(n10411), .ZN(n10410) );
  NAND2_X1 U8615 ( .A1(n7212), .A2(n10175), .ZN(n10149) );
  NAND2_X1 U8616 ( .A1(n7330), .A2(n10166), .ZN(n10136) );
  NAND2_X1 U8617 ( .A1(n10148), .A2(n10147), .ZN(n10175) );
  NAND2_X1 U8618 ( .A1(n7210), .A2(n10175), .ZN(n10177) );
  INV_X1 U8619 ( .A(n7211), .ZN(n7210) );
  OR2_X1 U8620 ( .A1(n7329), .A2(n7328), .ZN(n10168) );
  INV_X1 U8621 ( .A(n10166), .ZN(n7328) );
  NOR2_X1 U8622 ( .A1(n7332), .A2(n10441), .ZN(n10442) );
  NAND2_X1 U8623 ( .A1(n10457), .A2(n10456), .ZN(n7306) );
  NAND2_X1 U8624 ( .A1(n10477), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10456) );
  NAND2_X1 U8625 ( .A1(n7312), .A2(n6771), .ZN(n7061) );
  OR2_X1 U8626 ( .A1(n7985), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7911) );
  XNOR2_X1 U8627 ( .A(n11566), .B(n11572), .ZN(n11466) );
  INV_X1 U8628 ( .A(n11566), .ZN(n11567) );
  XNOR2_X1 U8629 ( .A(n7315), .B(n12092), .ZN(n13074) );
  INV_X1 U8630 ( .A(n7315), .ZN(n12075) );
  NOR2_X1 U8631 ( .A1(n13074), .A2(n15669), .ZN(n13073) );
  NOR2_X1 U8632 ( .A1(n13067), .A2(n6982), .ZN(n13087) );
  NAND2_X1 U8633 ( .A1(n6984), .A2(n6983), .ZN(n6982) );
  INV_X1 U8634 ( .A(n13066), .ZN(n6983) );
  INV_X1 U8635 ( .A(n13065), .ZN(n6984) );
  INV_X1 U8636 ( .A(n12098), .ZN(n12099) );
  NAND2_X1 U8637 ( .A1(n7304), .A2(n7049), .ZN(n13139) );
  NAND2_X1 U8638 ( .A1(n12084), .A2(n13148), .ZN(n7049) );
  INV_X1 U8639 ( .A(n12894), .ZN(n7327) );
  NOR2_X1 U8640 ( .A1(n7321), .A2(n7325), .ZN(n7319) );
  OR2_X1 U8641 ( .A1(n7321), .A2(n6872), .ZN(n7320) );
  INV_X1 U8642 ( .A(n7296), .ZN(n7295) );
  AOI21_X1 U8643 ( .B1(n7297), .B2(n13212), .A(n8249), .ZN(n7296) );
  AOI21_X1 U8644 ( .B1(n7290), .B2(n7004), .A(n7003), .ZN(n7002) );
  INV_X1 U8645 ( .A(n13263), .ZN(n7004) );
  INV_X1 U8646 ( .A(n12733), .ZN(n7003) );
  INV_X1 U8647 ( .A(n12764), .ZN(n13270) );
  AND2_X1 U8648 ( .A1(n12714), .A2(n12702), .ZN(n7294) );
  NAND2_X1 U8649 ( .A1(n7009), .A2(n8243), .ZN(n13304) );
  INV_X1 U8650 ( .A(n13302), .ZN(n7009) );
  NAND2_X1 U8651 ( .A1(n8030), .A2(n8029), .ZN(n8055) );
  INV_X1 U8652 ( .A(n8031), .ZN(n8030) );
  INV_X1 U8653 ( .A(n7543), .ZN(n7542) );
  NAND2_X1 U8654 ( .A1(n7286), .A2(n7284), .ZN(n11849) );
  AOI21_X1 U8655 ( .B1(n7287), .B2(n7289), .A(n7285), .ZN(n7284) );
  NAND2_X1 U8656 ( .A1(n11647), .A2(n7287), .ZN(n7286) );
  INV_X1 U8657 ( .A(n12696), .ZN(n7285) );
  NAND2_X1 U8658 ( .A1(n11316), .A2(n8238), .ZN(n7920) );
  AOI21_X1 U8659 ( .B1(n7281), .B2(n7283), .A(n7278), .ZN(n7277) );
  INV_X1 U8660 ( .A(n12679), .ZN(n7278) );
  AND2_X1 U8661 ( .A1(n12681), .A2(n12680), .ZN(n12783) );
  AND4_X1 U8662 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n11749)
         );
  NAND2_X1 U8663 ( .A1(n7846), .A2(n15587), .ZN(n7865) );
  NAND2_X1 U8664 ( .A1(n7808), .A2(n10501), .ZN(n7826) );
  INV_X1 U8665 ( .A(n7809), .ZN(n7808) );
  OR2_X1 U8666 ( .A1(n7826), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7847) );
  CLKBUF_X1 U8667 ( .A(n10737), .Z(n10916) );
  AND2_X1 U8668 ( .A1(n12642), .A2(n12646), .ZN(n12775) );
  INV_X1 U8669 ( .A(n10846), .ZN(n12771) );
  XNOR2_X1 U8670 ( .A(n12956), .B(n15270), .ZN(n10846) );
  INV_X1 U8671 ( .A(n15246), .ZN(n15236) );
  AND4_X1 U8672 ( .A1(n7293), .A2(n7705), .A3(n7704), .A4(n10248), .ZN(n12619)
         );
  CLKBUF_X1 U8673 ( .A(n10312), .Z(n12772) );
  AND2_X1 U8674 ( .A1(n12750), .A2(n12751), .ZN(n12904) );
  NAND2_X1 U8675 ( .A1(n12588), .A2(n12587), .ZN(n12609) );
  AND3_X1 U8676 ( .A1(n7823), .A2(n7822), .A3(n7821), .ZN(n15283) );
  NAND2_X1 U8677 ( .A1(n7368), .A2(n8275), .ZN(n10299) );
  NAND2_X1 U8678 ( .A1(n9723), .A2(n9722), .ZN(n11954) );
  INV_X1 U8679 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U8680 ( .A1(n8176), .A2(n8175), .ZN(n8191) );
  NAND2_X1 U8681 ( .A1(n8140), .A2(n6936), .ZN(n8143) );
  NAND2_X1 U8682 ( .A1(n8081), .A2(n8080), .ZN(n8084) );
  NAND2_X1 U8683 ( .A1(n8064), .A2(n8063), .ZN(n8067) );
  INV_X1 U8684 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7668) );
  AOI21_X1 U8685 ( .B1(n7385), .B2(n7387), .A(n7384), .ZN(n7383) );
  INV_X1 U8686 ( .A(n8020), .ZN(n7384) );
  NAND2_X1 U8687 ( .A1(n8023), .A2(n8022), .ZN(n8040) );
  NAND2_X1 U8688 ( .A1(n7983), .A2(n7673), .ZN(n8003) );
  NAND2_X1 U8689 ( .A1(n7378), .A2(n7380), .ZN(n7977) );
  INV_X1 U8690 ( .A(n7381), .ZN(n7380) );
  NAND2_X1 U8691 ( .A1(n7923), .A2(n7379), .ZN(n7378) );
  OAI21_X1 U8692 ( .B1(n7940), .B2(n7959), .A(n7961), .ZN(n7381) );
  OR2_X1 U8693 ( .A1(n7911), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n7912) );
  NOR2_X1 U8694 ( .A1(n7912), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n7944) );
  OAI21_X1 U8695 ( .B1(n7834), .B2(n6913), .A(n6802), .ZN(n7886) );
  NAND2_X1 U8696 ( .A1(n6917), .A2(n7832), .ZN(n6913) );
  INV_X1 U8697 ( .A(n6915), .ZN(n6914) );
  AND2_X1 U8698 ( .A1(n7818), .A2(n7800), .ZN(n7815) );
  AND2_X1 U8699 ( .A1(n7803), .A2(n7819), .ZN(n10445) );
  NAND2_X1 U8700 ( .A1(n7779), .A2(n7778), .ZN(n7797) );
  NAND2_X1 U8701 ( .A1(n6926), .A2(n7760), .ZN(n6925) );
  XNOR2_X1 U8702 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7796) );
  NOR2_X1 U8703 ( .A1(n7781), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7802) );
  XNOR2_X1 U8704 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7717) );
  NAND2_X1 U8705 ( .A1(n8948), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7716) );
  NOR2_X1 U8706 ( .A1(n6751), .A2(n7450), .ZN(n7449) );
  OR2_X1 U8707 ( .A1(n13494), .A2(n11983), .ZN(n7463) );
  NAND2_X1 U8708 ( .A1(n9183), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9206) );
  OR2_X1 U8709 ( .A1(n9206), .A2(n14995), .ZN(n9221) );
  INV_X1 U8710 ( .A(n9340), .ZN(n9337) );
  XNOR2_X1 U8711 ( .A(n15175), .B(n10516), .ZN(n12048) );
  NAND2_X1 U8712 ( .A1(n7455), .A2(n7458), .ZN(n7454) );
  NAND2_X1 U8713 ( .A1(n13479), .A2(n7132), .ZN(n7453) );
  NOR2_X1 U8714 ( .A1(n6833), .A2(n7133), .ZN(n7132) );
  INV_X1 U8715 ( .A(n11996), .ZN(n7133) );
  AND2_X1 U8716 ( .A1(n9704), .A2(n9510), .ZN(n9891) );
  OR2_X1 U8717 ( .A1(n11509), .A2(n11508), .ZN(n11510) );
  XNOR2_X1 U8718 ( .A(n13648), .B(n13646), .ZN(n9540) );
  INV_X1 U8719 ( .A(n9531), .ZN(n7621) );
  AND2_X1 U8720 ( .A1(n9478), .A2(n9477), .ZN(n13473) );
  AND2_X1 U8721 ( .A1(n9434), .A2(n9433), .ZN(n12036) );
  NAND4_X1 U8722 ( .A1(n8978), .A2(n8977), .A3(n8976), .A4(n8975), .ZN(n9543)
         );
  NAND2_X1 U8723 ( .A1(n9505), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8976) );
  OR2_X1 U8724 ( .A1(n9213), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9229) );
  INV_X1 U8725 ( .A(n7071), .ZN(n13652) );
  INV_X1 U8726 ( .A(n9702), .ZN(n9632) );
  NAND2_X1 U8727 ( .A1(n13675), .A2(n13851), .ZN(n13659) );
  NAND2_X1 U8728 ( .A1(n13694), .A2(n13526), .ZN(n9700) );
  AND2_X1 U8729 ( .A1(n9471), .A2(n9417), .ZN(n13692) );
  NOR2_X1 U8730 ( .A1(n13754), .A2(n7079), .ZN(n13707) );
  NOR3_X1 U8731 ( .A1(n13754), .A2(n13861), .A3(n7079), .ZN(n13691) );
  AOI21_X1 U8732 ( .B1(n7478), .B2(n7480), .A(n9696), .ZN(n13720) );
  AND2_X1 U8733 ( .A1(n7479), .A2(n9697), .ZN(n7478) );
  OAI21_X1 U8734 ( .B1(n13805), .B2(n7586), .A(n6797), .ZN(n13790) );
  AND2_X1 U8735 ( .A1(n13814), .A2(n13589), .ZN(n7586) );
  OR2_X1 U8736 ( .A1(n9293), .A2(n9292), .ZN(n9310) );
  AND2_X1 U8737 ( .A1(n6763), .A2(n13814), .ZN(n7075) );
  OR2_X1 U8738 ( .A1(n9260), .A2(n9259), .ZN(n9277) );
  NAND2_X1 U8739 ( .A1(n7029), .A2(n9686), .ZN(n11803) );
  NAND2_X1 U8740 ( .A1(n7475), .A2(n7473), .ZN(n7029) );
  NOR2_X1 U8741 ( .A1(n7474), .A2(n6799), .ZN(n7473) );
  NAND2_X1 U8742 ( .A1(n11591), .A2(n9708), .ZN(n11812) );
  NOR2_X1 U8743 ( .A1(n11597), .A2(n7613), .ZN(n7612) );
  NOR2_X1 U8744 ( .A1(n9680), .A2(n7487), .ZN(n7486) );
  NAND2_X1 U8745 ( .A1(n10988), .A2(n9707), .ZN(n11179) );
  OAI21_X1 U8746 ( .B1(n9602), .B2(n9676), .A(n7577), .ZN(n10980) );
  OR2_X1 U8747 ( .A1(n9112), .A2(n9111), .ZN(n9127) );
  INV_X1 U8748 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n12118) );
  NAND2_X1 U8749 ( .A1(n7074), .A2(n7073), .ZN(n10987) );
  INV_X1 U8750 ( .A(n11095), .ZN(n7074) );
  NAND2_X1 U8751 ( .A1(n7068), .A2(n10636), .ZN(n10824) );
  INV_X1 U8752 ( .A(n10634), .ZN(n7068) );
  NAND2_X1 U8753 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9050) );
  NAND2_X1 U8754 ( .A1(n7070), .A2(n7069), .ZN(n10634) );
  INV_X1 U8755 ( .A(n10865), .ZN(n7070) );
  NAND2_X1 U8756 ( .A1(n10866), .A2(n15191), .ZN(n10865) );
  AND2_X1 U8757 ( .A1(n10594), .A2(n10596), .ZN(n10866) );
  INV_X1 U8758 ( .A(n13567), .ZN(n15127) );
  CLKBUF_X1 U8759 ( .A(n9512), .Z(n9659) );
  NAND2_X1 U8760 ( .A1(n9415), .A2(n9414), .ZN(n13866) );
  NAND2_X1 U8761 ( .A1(n9402), .A2(n9401), .ZN(n13871) );
  INV_X1 U8762 ( .A(n15200), .ZN(n15218) );
  AND2_X1 U8763 ( .A1(n9786), .A2(n9890), .ZN(n9790) );
  AND2_X1 U8764 ( .A1(n6816), .A2(n8933), .ZN(n7642) );
  INV_X1 U8765 ( .A(n8956), .ZN(n8934) );
  OR2_X1 U8766 ( .A1(n9580), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n9582) );
  XNOR2_X1 U8767 ( .A(n8967), .B(n8968), .ZN(n8972) );
  INV_X1 U8768 ( .A(n9248), .ZN(n8959) );
  OR2_X1 U8769 ( .A1(n9096), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9098) );
  OR2_X1 U8770 ( .A1(n9056), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9058) );
  CLKBUF_X1 U8771 ( .A(n8981), .Z(n8982) );
  INV_X1 U8772 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8948) );
  INV_X1 U8773 ( .A(n11537), .ZN(n6905) );
  NAND2_X1 U8774 ( .A1(n8566), .A2(n8415), .ZN(n8581) );
  NAND2_X1 U8775 ( .A1(n8698), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8715) );
  NOR2_X1 U8776 ( .A1(n8521), .A2(n8520), .ZN(n8536) );
  NAND2_X1 U8777 ( .A1(n11291), .A2(n7531), .ZN(n7529) );
  OR2_X1 U8778 ( .A1(n8581), .A2(n11887), .ZN(n8592) );
  INV_X1 U8779 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10574) );
  AND2_X1 U8780 ( .A1(n12254), .A2(n12252), .ZN(n14019) );
  INV_X1 U8781 ( .A(n8768), .ZN(n8780) );
  NAND2_X1 U8782 ( .A1(n7509), .A2(n6764), .ZN(n7508) );
  INV_X1 U8783 ( .A(n6749), .ZN(n12265) );
  AOI21_X1 U8784 ( .B1(n7526), .B2(n7525), .A(n7524), .ZN(n7523) );
  INV_X1 U8785 ( .A(n11697), .ZN(n7524) );
  INV_X1 U8786 ( .A(n7531), .ZN(n7525) );
  OAI21_X1 U8787 ( .B1(n8838), .B2(n10622), .A(n10351), .ZN(n10352) );
  INV_X1 U8788 ( .A(n10350), .ZN(n10351) );
  AOI21_X1 U8789 ( .B1(n8837), .B2(n11281), .A(n10347), .ZN(n10619) );
  NAND2_X1 U8790 ( .A1(n10346), .A2(n10345), .ZN(n10347) );
  NAND2_X1 U8791 ( .A1(n10344), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U8792 ( .A1(n10360), .A2(n12262), .ZN(n10346) );
  INV_X1 U8793 ( .A(n14083), .ZN(n6899) );
  NOR2_X1 U8794 ( .A1(n13999), .A2(n7515), .ZN(n7514) );
  INV_X1 U8795 ( .A(n12210), .ZN(n7515) );
  AOI22_X1 U8796 ( .A1(n11281), .A2(n14158), .B1(n10710), .B2(n12262), .ZN(
        n10623) );
  AND3_X1 U8797 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U8798 ( .A1(n6902), .A2(n6900), .ZN(n14027) );
  AOI21_X1 U8799 ( .B1(n7517), .B2(n14005), .A(n6901), .ZN(n6900) );
  NOR2_X1 U8800 ( .A1(n7521), .A2(n7518), .ZN(n7517) );
  INV_X1 U8801 ( .A(n10622), .ZN(n12268) );
  NAND2_X1 U8802 ( .A1(n7440), .A2(n7441), .ZN(n7438) );
  NOR2_X1 U8803 ( .A1(n7441), .A2(n7440), .ZN(n7439) );
  AND4_X1 U8804 ( .A1(n8809), .A2(n8808), .A3(n8807), .A4(n8806), .ZN(n13969)
         );
  AND4_X1 U8805 ( .A1(n8636), .A2(n8635), .A3(n8634), .A4(n8633), .ZN(n12157)
         );
  AND4_X1 U8806 ( .A1(n8509), .A2(n8508), .A3(n8507), .A4(n8506), .ZN(n12344)
         );
  NAND2_X1 U8807 ( .A1(n6639), .A2(n8400), .ZN(n8532) );
  OR2_X1 U8808 ( .A1(n11056), .A2(n11057), .ZN(n6968) );
  AND2_X1 U8809 ( .A1(n6968), .A2(n6967), .ZN(n11776) );
  NAND2_X1 U8810 ( .A1(n11782), .A2(n11775), .ZN(n6967) );
  NOR2_X1 U8811 ( .A1(n14285), .A2(n14284), .ZN(n14287) );
  NOR2_X1 U8812 ( .A1(n14313), .A2(n12475), .ZN(n7193) );
  NAND2_X1 U8813 ( .A1(n8823), .A2(n8821), .ZN(n8824) );
  NOR2_X1 U8814 ( .A1(n12542), .A2(n7245), .ZN(n7244) );
  INV_X1 U8815 ( .A(n8824), .ZN(n7245) );
  NAND2_X1 U8816 ( .A1(n7265), .A2(n8862), .ZN(n14386) );
  INV_X1 U8817 ( .A(n8754), .ZN(n8769) );
  NOR2_X1 U8818 ( .A1(n14511), .A2(n7198), .ZN(n14462) );
  OR2_X1 U8819 ( .A1(n8715), .A2(n15441), .ZN(n8728) );
  NOR2_X1 U8820 ( .A1(n8728), .A2(n8727), .ZN(n8744) );
  OR2_X1 U8821 ( .A1(n14583), .A2(n14047), .ZN(n14479) );
  INV_X1 U8822 ( .A(n14095), .ZN(n14110) );
  AND2_X1 U8823 ( .A1(n14479), .A2(n12430), .ZN(n14490) );
  AND2_X1 U8824 ( .A1(n8682), .A2(n8681), .ZN(n14514) );
  OR2_X1 U8825 ( .A1(n11661), .A2(n12402), .ZN(n11831) );
  NAND2_X1 U8826 ( .A1(n11358), .A2(n8849), .ZN(n11482) );
  NAND2_X1 U8827 ( .A1(n6652), .A2(n7192), .ZN(n11475) );
  OAI21_X1 U8828 ( .B1(n6739), .B2(n6785), .A(n7255), .ZN(n7254) );
  NOR2_X1 U8829 ( .A1(n10339), .A2(n8915), .ZN(n11305) );
  NAND2_X1 U8830 ( .A1(n8846), .A2(n8845), .ZN(n10882) );
  NAND2_X1 U8831 ( .A1(n11306), .A2(n8834), .ZN(n14974) );
  AND2_X1 U8832 ( .A1(n10348), .A2(n8913), .ZN(n10342) );
  NAND2_X1 U8833 ( .A1(n8405), .A2(n8410), .ZN(n7535) );
  XNOR2_X1 U8834 ( .A(n9463), .B(n9462), .ZN(n13944) );
  AND2_X1 U8835 ( .A1(n9500), .A2(n9499), .ZN(n12484) );
  NAND2_X1 U8836 ( .A1(n9456), .A2(n9455), .ZN(n7145) );
  XNOR2_X1 U8837 ( .A(n9492), .B(n9491), .ZN(n13949) );
  OAI21_X1 U8838 ( .B1(n8811), .B2(SI_27_), .A(n7652), .ZN(n8394) );
  INV_X1 U8839 ( .A(n8874), .ZN(n8876) );
  INV_X1 U8840 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8882) );
  OR2_X1 U8841 ( .A1(n8377), .A2(SI_22_), .ZN(n8378) );
  NAND2_X1 U8842 ( .A1(n8724), .A2(n8372), .ZN(n8738) );
  AND2_X1 U8843 ( .A1(n8376), .A2(n8375), .ZN(n8737) );
  NAND2_X1 U8844 ( .A1(n8372), .A2(n8371), .ZN(n8722) );
  AND2_X1 U8845 ( .A1(n8489), .A2(n8517), .ZN(n10042) );
  AND2_X1 U8846 ( .A1(n8316), .A2(n8315), .ZN(n8471) );
  NAND2_X1 U8847 ( .A1(n8472), .A2(n8471), .ZN(n8474) );
  XNOR2_X1 U8848 ( .A(n14663), .B(P3_ADDR_REG_3__SCAN_IN), .ZN(n14693) );
  NAND2_X1 U8849 ( .A1(n14669), .A2(n14668), .ZN(n14703) );
  NAND2_X1 U8850 ( .A1(n14698), .A2(n14699), .ZN(n14668) );
  XNOR2_X1 U8851 ( .A(n14671), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14710) );
  NAND2_X1 U8852 ( .A1(n6954), .A2(n6953), .ZN(n14721) );
  INV_X1 U8853 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6953) );
  INV_X1 U8854 ( .A(n6955), .ZN(n6954) );
  NAND2_X1 U8855 ( .A1(n6955), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n14722) );
  NAND2_X1 U8856 ( .A1(n7106), .A2(n7105), .ZN(n14718) );
  NAND2_X1 U8857 ( .A1(n14713), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7105) );
  OR2_X1 U8858 ( .A1(n14713), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7104) );
  AND2_X1 U8859 ( .A1(n14721), .A2(n6952), .ZN(n14726) );
  NAND2_X1 U8860 ( .A1(n14722), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U8861 ( .A1(n7098), .A2(n7097), .ZN(n14738) );
  NAND2_X1 U8862 ( .A1(n14853), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U8863 ( .A1(n7099), .A2(n6787), .ZN(n7098) );
  AND2_X1 U8864 ( .A1(n7096), .A2(n7095), .ZN(n14747) );
  NAND2_X1 U8865 ( .A1(n6940), .A2(n6943), .ZN(n14749) );
  NAND2_X1 U8866 ( .A1(n14741), .A2(n6946), .ZN(n6940) );
  INV_X1 U8867 ( .A(n7088), .ZN(n7086) );
  NOR2_X2 U8868 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14761) );
  NAND2_X1 U8869 ( .A1(n7091), .A2(n14782), .ZN(n7090) );
  INV_X1 U8870 ( .A(n14781), .ZN(n7091) );
  AOI21_X1 U8871 ( .B1(n7345), .B2(n7352), .A(n7343), .ZN(n7342) );
  NAND2_X1 U8872 ( .A1(n12848), .A2(n7339), .ZN(n7337) );
  NAND2_X1 U8873 ( .A1(n13004), .A2(n7336), .ZN(n7335) );
  AND2_X1 U8874 ( .A1(n12982), .A2(n11742), .ZN(n12871) );
  NAND2_X1 U8875 ( .A1(n10689), .A2(n7364), .ZN(n12882) );
  AND2_X1 U8876 ( .A1(n10690), .A2(n10688), .ZN(n7364) );
  NAND2_X1 U8877 ( .A1(n10689), .A2(n10688), .ZN(n12881) );
  NAND2_X1 U8878 ( .A1(n12893), .A2(n12892), .ZN(n12891) );
  NAND2_X1 U8879 ( .A1(n12996), .A2(n12843), .ZN(n12913) );
  NAND2_X1 U8880 ( .A1(n8087), .A2(n8086), .ZN(n13286) );
  OR2_X1 U8881 ( .A1(n10731), .A2(n8199), .ZN(n8087) );
  NAND2_X1 U8882 ( .A1(n7353), .A2(n12853), .ZN(n12933) );
  NAND2_X1 U8883 ( .A1(n7989), .A2(n7988), .ZN(n12949) );
  OR2_X1 U8884 ( .A1(n10082), .A2(n8199), .ZN(n7989) );
  INV_X1 U8885 ( .A(n7348), .ZN(n12972) );
  NAND2_X1 U8886 ( .A1(n11739), .A2(n11738), .ZN(n12984) );
  AND4_X1 U8887 ( .A1(n8060), .A2(n8059), .A3(n8058), .A4(n8057), .ZN(n13027)
         );
  NAND2_X1 U8888 ( .A1(n12998), .A2(n12997), .ZN(n12996) );
  INV_X1 U8889 ( .A(n13046), .ZN(n12995) );
  NAND2_X1 U8890 ( .A1(n8104), .A2(n8103), .ZN(n13275) );
  OR2_X1 U8891 ( .A1(n10763), .A2(n8199), .ZN(n8104) );
  INV_X1 U8892 ( .A(n13028), .ZN(n13037) );
  INV_X1 U8893 ( .A(n7729), .ZN(n7746) );
  NAND2_X1 U8894 ( .A1(n7341), .A2(n7349), .ZN(n13035) );
  NAND2_X1 U8895 ( .A1(n7353), .A2(n7351), .ZN(n7341) );
  AND2_X1 U8896 ( .A1(n10247), .A2(n10246), .ZN(n13044) );
  AND2_X1 U8897 ( .A1(n12595), .A2(n9732), .ZN(n12608) );
  AND2_X1 U8898 ( .A1(n12595), .A2(n8225), .ZN(n12909) );
  NAND2_X1 U8899 ( .A1(n8187), .A2(n8186), .ZN(n13216) );
  NAND2_X1 U8900 ( .A1(n8169), .A2(n8168), .ZN(n13233) );
  INV_X1 U8901 ( .A(n13256), .ZN(n13232) );
  INV_X1 U8902 ( .A(n13027), .ZN(n13334) );
  INV_X1 U8903 ( .A(n12944), .ZN(n13333) );
  INV_X1 U8904 ( .A(n11744), .ZN(n13016) );
  INV_X1 U8905 ( .A(n11740), .ZN(n12874) );
  INV_X1 U8906 ( .A(n11072), .ZN(n13057) );
  INV_X1 U8907 ( .A(n7745), .ZN(n10809) );
  OR2_X1 U8908 ( .A1(n10236), .A2(n11949), .ZN(n13060) );
  NAND2_X1 U8909 ( .A1(n6973), .A2(n6972), .ZN(n10201) );
  OAI21_X1 U8910 ( .B1(n10422), .B2(n6971), .A(n6970), .ZN(n6973) );
  NAND2_X1 U8911 ( .A1(n10421), .A2(n6974), .ZN(n6972) );
  NAND2_X1 U8912 ( .A1(n7331), .A2(n7333), .ZN(n10211) );
  NAND2_X1 U8913 ( .A1(n10443), .A2(n10444), .ZN(n10457) );
  NAND2_X1 U8914 ( .A1(n7332), .A2(n7331), .ZN(n10443) );
  XNOR2_X1 U8915 ( .A(n7306), .B(n7305), .ZN(n10492) );
  INV_X1 U8916 ( .A(n7220), .ZN(n10962) );
  INV_X1 U8917 ( .A(n10460), .ZN(n7054) );
  INV_X1 U8918 ( .A(n7055), .ZN(n10461) );
  XNOR2_X1 U8919 ( .A(n11208), .B(n7313), .ZN(n10950) );
  INV_X1 U8920 ( .A(n7312), .ZN(n11209) );
  INV_X1 U8921 ( .A(n7059), .ZN(n11465) );
  INV_X1 U8922 ( .A(n7061), .ZN(n11212) );
  AND2_X1 U8923 ( .A1(n6995), .A2(n6993), .ZN(n11460) );
  NOR2_X1 U8924 ( .A1(n11561), .A2(n11562), .ZN(n11565) );
  NOR2_X1 U8925 ( .A1(n13062), .A2(n12058), .ZN(n13081) );
  NOR2_X1 U8926 ( .A1(n13098), .A2(n13099), .ZN(n13097) );
  INV_X1 U8927 ( .A(n7307), .ZN(n13108) );
  NAND2_X1 U8928 ( .A1(n7224), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7223) );
  NAND2_X1 U8929 ( .A1(n12062), .A2(n7224), .ZN(n7222) );
  INV_X1 U8930 ( .A(n13116), .ZN(n7224) );
  INV_X1 U8931 ( .A(n7310), .ZN(n13126) );
  INV_X1 U8932 ( .A(n13157), .ZN(n13135) );
  NAND2_X1 U8933 ( .A1(n13215), .A2(n8248), .ZN(n13202) );
  NAND2_X1 U8934 ( .A1(n8162), .A2(n8161), .ZN(n13361) );
  NAND2_X1 U8935 ( .A1(n8146), .A2(n8145), .ZN(n13368) );
  OR2_X1 U8936 ( .A1(n11422), .A2(n8199), .ZN(n8146) );
  NAND2_X1 U8937 ( .A1(n7553), .A2(n7557), .ZN(n13248) );
  NAND2_X1 U8938 ( .A1(n13266), .A2(n12730), .ZN(n13241) );
  NAND2_X1 U8939 ( .A1(n7563), .A2(n7561), .ZN(n13258) );
  NAND2_X1 U8940 ( .A1(n8070), .A2(n8069), .ZN(n13308) );
  OR2_X1 U8941 ( .A1(n10563), .A2(n8199), .ZN(n8070) );
  NAND2_X1 U8942 ( .A1(n13331), .A2(n8038), .ZN(n13311) );
  NAND2_X1 U8943 ( .A1(n8054), .A2(n8053), .ZN(n13323) );
  OR2_X1 U8944 ( .A1(n10402), .A2(n8199), .ZN(n8054) );
  NAND2_X1 U8945 ( .A1(n8240), .A2(n12701), .ZN(n13338) );
  NAND2_X1 U8946 ( .A1(n7545), .A2(n7974), .ZN(n11845) );
  NAND2_X1 U8947 ( .A1(n11823), .A2(n7973), .ZN(n7545) );
  NAND2_X1 U8948 ( .A1(n11646), .A2(n12686), .ZN(n11822) );
  NAND2_X1 U8949 ( .A1(n7928), .A2(n7927), .ZN(n14789) );
  NAND2_X1 U8950 ( .A1(n7280), .A2(n12672), .ZN(n11320) );
  NAND2_X1 U8951 ( .A1(n11192), .A2(n8237), .ZN(n7280) );
  NAND2_X1 U8952 ( .A1(n11252), .A2(n7845), .ZN(n11071) );
  NAND2_X1 U8953 ( .A1(n10734), .A2(n7273), .ZN(n7014) );
  INV_X1 U8954 ( .A(n11241), .ZN(n15289) );
  NAND2_X1 U8955 ( .A1(n10736), .A2(n12651), .ZN(n10776) );
  OR2_X1 U8956 ( .A1(n10745), .A2(n10744), .ZN(n13341) );
  INV_X1 U8957 ( .A(n15238), .ZN(n13288) );
  NAND2_X1 U8958 ( .A1(n12604), .A2(n12603), .ZN(n13411) );
  INV_X1 U8959 ( .A(n12609), .ZN(n13417) );
  INV_X1 U8960 ( .A(n12949), .ZN(n13457) );
  AND2_X1 U8961 ( .A1(n8273), .A2(n8272), .ZN(n13458) );
  AND2_X1 U8962 ( .A1(n10232), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13459) );
  INV_X1 U8963 ( .A(n7686), .ZN(n11960) );
  NOR2_X1 U8964 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  NOR2_X1 U8965 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8260) );
  NAND2_X1 U8966 ( .A1(n8140), .A2(n8126), .ZN(n8139) );
  NAND2_X1 U8967 ( .A1(n8114), .A2(n8113), .ZN(n8123) );
  INV_X1 U8968 ( .A(n9775), .ZN(n10561) );
  NAND2_X1 U8969 ( .A1(n8001), .A2(n8000), .ZN(n8019) );
  INV_X1 U8970 ( .A(SI_16_), .ZN(n10083) );
  NAND2_X1 U8971 ( .A1(n7941), .A2(n7940), .ZN(n7960) );
  NAND2_X1 U8972 ( .A1(n6932), .A2(n6835), .ZN(n7922) );
  NAND2_X1 U8973 ( .A1(n6932), .A2(n7905), .ZN(n7908) );
  INV_X1 U8974 ( .A(SI_11_), .ZN(n9870) );
  OAI21_X1 U8975 ( .B1(n7854), .B2(n7853), .A(n7855), .ZN(n7871) );
  NAND2_X1 U8976 ( .A1(n7839), .A2(n7838), .ZN(n10963) );
  INV_X1 U8977 ( .A(n10445), .ZN(n10477) );
  NAND2_X1 U8978 ( .A1(n6924), .A2(n7760), .ZN(n7777) );
  NAND2_X1 U8979 ( .A1(n6928), .A2(n6927), .ZN(n6924) );
  INV_X1 U8980 ( .A(n6926), .ZN(n6927) );
  OR2_X1 U8981 ( .A1(n7761), .A2(n13462), .ZN(n7762) );
  NAND2_X1 U8982 ( .A1(n6928), .A2(n7737), .ZN(n7759) );
  NAND2_X1 U8983 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7725) );
  INV_X1 U8984 ( .A(n7221), .ZN(n7699) );
  NAND2_X1 U8985 ( .A1(n12126), .A2(n11010), .ZN(n11085) );
  NAND2_X1 U8986 ( .A1(n12054), .A2(n9803), .ZN(n9815) );
  NAND2_X1 U8987 ( .A1(n10548), .A2(n10549), .ZN(n10551) );
  OAI21_X1 U8988 ( .B1(n10539), .B2(n10540), .A(n10544), .ZN(n10545) );
  AND2_X1 U8989 ( .A1(n7137), .A2(n7136), .ZN(n13512) );
  NAND2_X1 U8990 ( .A1(n11495), .A2(n12576), .ZN(n12582) );
  NAND2_X1 U8991 ( .A1(n9197), .A2(n9196), .ZN(n14815) );
  NAND2_X1 U8992 ( .A1(n11688), .A2(n11687), .ZN(n11689) );
  NAND2_X1 U8993 ( .A1(n13533), .A2(n13532), .ZN(n13521) );
  NAND2_X1 U8994 ( .A1(n13482), .A2(n12000), .ZN(n13533) );
  NAND2_X1 U8995 ( .A1(n7141), .A2(n6767), .ZN(n7138) );
  NAND2_X1 U8996 ( .A1(n12582), .A2(n11499), .ZN(n15000) );
  NAND2_X1 U8997 ( .A1(n9216), .A2(n9215), .ZN(n15005) );
  INV_X1 U8998 ( .A(n9795), .ZN(n9796) );
  AND2_X1 U8999 ( .A1(n9820), .A2(n15132), .ZN(n13539) );
  INV_X1 U9000 ( .A(n13539), .ZN(n15004) );
  INV_X1 U9001 ( .A(n13473), .ZN(n13579) );
  INV_X1 U9002 ( .A(n13526), .ZN(n13581) );
  OR2_X1 U9003 ( .A1(n9506), .A2(n9974), .ZN(n8946) );
  NAND2_X1 U9004 ( .A1(n13645), .A2(n15134), .ZN(n13840) );
  XNOR2_X1 U9005 ( .A(n13651), .B(n13644), .ZN(n13645) );
  INV_X1 U9006 ( .A(n13643), .ZN(n13843) );
  XNOR2_X1 U9007 ( .A(n7048), .B(n9630), .ZN(n13860) );
  OAI21_X1 U9008 ( .B1(n13695), .B2(n7468), .A(n6737), .ZN(n7048) );
  INV_X1 U9009 ( .A(n9700), .ZN(n7468) );
  NAND2_X1 U9010 ( .A1(n7599), .A2(n7600), .ZN(n13715) );
  NOR2_X1 U9011 ( .A1(n7477), .A2(n7476), .ZN(n13734) );
  INV_X1 U9012 ( .A(n7479), .ZN(n7476) );
  INV_X1 U9013 ( .A(n7480), .ZN(n7477) );
  AOI21_X1 U9014 ( .B1(n13743), .B2(n13748), .A(n7605), .ZN(n13729) );
  NAND2_X1 U9015 ( .A1(n7483), .A2(n7484), .ZN(n13747) );
  AND2_X1 U9016 ( .A1(n7483), .A2(n7481), .ZN(n13746) );
  OR2_X1 U9017 ( .A1(n11389), .A2(n9370), .ZN(n9372) );
  NAND2_X1 U9018 ( .A1(n7042), .A2(n7046), .ZN(n13779) );
  NAND2_X1 U9019 ( .A1(n13808), .A2(n7043), .ZN(n7042) );
  NAND2_X1 U9020 ( .A1(n9333), .A2(n9332), .ZN(n13891) );
  OR2_X1 U9021 ( .A1(n10905), .A2(n9370), .ZN(n9333) );
  NAND2_X1 U9022 ( .A1(n13808), .A2(n9691), .ZN(n13801) );
  AND2_X1 U9023 ( .A1(n7490), .A2(n7491), .ZN(n13810) );
  AND2_X1 U9024 ( .A1(n7493), .A2(n9690), .ZN(n13824) );
  NAND2_X1 U9025 ( .A1(n9274), .A2(n9273), .ZN(n13907) );
  NAND2_X1 U9026 ( .A1(n7580), .A2(n7584), .ZN(n13821) );
  NAND2_X1 U9027 ( .A1(n11796), .A2(n7585), .ZN(n7580) );
  NAND2_X1 U9028 ( .A1(n9258), .A2(n9257), .ZN(n13911) );
  AOI21_X1 U9029 ( .B1(n11177), .B2(n7614), .A(n9612), .ZN(n11587) );
  NAND2_X1 U9030 ( .A1(n7488), .A2(n9679), .ZN(n11169) );
  NAND2_X1 U9031 ( .A1(n9158), .A2(n9157), .ZN(n15213) );
  OAI21_X1 U9032 ( .B1(n10856), .B2(n7034), .A(n7033), .ZN(n10632) );
  AOI21_X1 U9033 ( .B1(n7036), .B2(n10858), .A(n7035), .ZN(n7033) );
  NAND2_X1 U9034 ( .A1(n7594), .A2(n9598), .ZN(n10638) );
  NAND2_X1 U9035 ( .A1(n10608), .A2(n9597), .ZN(n7594) );
  NAND2_X1 U9036 ( .A1(n7038), .A2(n9669), .ZN(n10606) );
  NAND2_X1 U9037 ( .A1(n10856), .A2(n9667), .ZN(n7038) );
  NAND2_X1 U9038 ( .A1(n15155), .A2(n9818), .ZN(n13813) );
  NAND2_X1 U9039 ( .A1(n15166), .A2(n10073), .ZN(n15132) );
  CLKBUF_X1 U9040 ( .A(n15151), .Z(n6875) );
  AND3_X2 U9041 ( .A1(n10076), .A2(n11970), .A3(n10661), .ZN(n15233) );
  NOR2_X1 U9042 ( .A1(n13844), .A2(n6774), .ZN(n13846) );
  AND2_X1 U9043 ( .A1(n13852), .A2(n7654), .ZN(n13855) );
  OR2_X1 U9044 ( .A1(n13853), .A2(n15187), .ZN(n13854) );
  AND2_X1 U9045 ( .A1(n9790), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15166) );
  INV_X1 U9046 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13945) );
  NOR2_X1 U9047 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7028) );
  INV_X1 U9048 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10401) );
  INV_X1 U9049 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10369) );
  INV_X1 U9050 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10056) );
  INV_X1 U9051 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9917) );
  INV_X1 U9052 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9865) );
  INV_X1 U9053 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9861) );
  INV_X1 U9054 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9848) );
  INV_X1 U9055 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9035) );
  INV_X1 U9056 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9826) );
  INV_X1 U9057 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9872) );
  CLKBUF_X1 U9058 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n13962) );
  XNOR2_X1 U9059 ( .A(n11536), .B(n6905), .ZN(n11538) );
  AOI21_X1 U9060 ( .B1(n11291), .B2(n11290), .A(n7533), .ZN(n11539) );
  OAI21_X1 U9061 ( .B1(n14106), .B2(n12260), .A(n7497), .ZN(n13964) );
  NAND2_X1 U9062 ( .A1(n14105), .A2(n12261), .ZN(n13965) );
  NAND2_X1 U9063 ( .A1(n7501), .A2(n13982), .ZN(n13980) );
  NAND2_X1 U9064 ( .A1(n13981), .A2(n13983), .ZN(n7501) );
  NAND2_X1 U9065 ( .A1(n7513), .A2(n7510), .ZN(n10722) );
  INV_X1 U9066 ( .A(n7512), .ZN(n7510) );
  AOI21_X1 U9067 ( .B1(n7497), .B2(n12260), .A(n12273), .ZN(n7496) );
  NAND2_X1 U9068 ( .A1(n7529), .A2(n7530), .ZN(n11548) );
  NOR2_X1 U9069 ( .A1(n10621), .A2(n10620), .ZN(n10707) );
  AND2_X1 U9070 ( .A1(n10619), .A2(n12212), .ZN(n10620) );
  OR2_X1 U9071 ( .A1(n14006), .A2(n14005), .ZN(n14007) );
  NAND2_X1 U9072 ( .A1(n7522), .A2(n12188), .ZN(n14093) );
  NAND2_X1 U9073 ( .A1(n6645), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8445) );
  NOR2_X1 U9074 ( .A1(n10085), .A2(n10086), .ZN(n10084) );
  NAND2_X1 U9075 ( .A1(n14224), .A2(n6782), .ZN(n14239) );
  NAND2_X1 U9076 ( .A1(n14249), .A2(n6852), .ZN(n10277) );
  INV_X1 U9077 ( .A(n6968), .ZN(n11774) );
  XNOR2_X1 U9078 ( .A(n11776), .B(n6966), .ZN(n14867) );
  NAND2_X1 U9079 ( .A1(n14867), .A2(n14866), .ZN(n14865) );
  AND2_X1 U9080 ( .A1(n7194), .A2(n14901), .ZN(n14519) );
  XNOR2_X1 U9081 ( .A(n7195), .B(n12505), .ZN(n7194) );
  NAND2_X1 U9082 ( .A1(n14131), .A2(n14111), .ZN(n7127) );
  OR3_X1 U9083 ( .A1(n8835), .A2(n9754), .A3(n14909), .ZN(n14334) );
  AOI21_X1 U9084 ( .B1(n7272), .B2(n14899), .A(n7271), .ZN(n14338) );
  INV_X1 U9085 ( .A(n12281), .ZN(n7271) );
  OR3_X1 U9086 ( .A1(n14347), .A2(n14346), .A3(n14909), .ZN(n14526) );
  NAND2_X1 U9087 ( .A1(n14367), .A2(n8797), .ZN(n14355) );
  NAND2_X1 U9088 ( .A1(n14388), .A2(n8864), .ZN(n14377) );
  NAND2_X1 U9089 ( .A1(n14411), .A2(n8774), .ZN(n14392) );
  NAND2_X1 U9090 ( .A1(n14459), .A2(n8858), .ZN(n14441) );
  NAND2_X1 U9091 ( .A1(n7230), .A2(n8703), .ZN(n14469) );
  NAND2_X1 U9092 ( .A1(n7122), .A2(n7259), .ZN(n14503) );
  NAND2_X1 U9093 ( .A1(n11833), .A2(n12411), .ZN(n11913) );
  OAI21_X1 U9094 ( .B1(n11480), .B2(n7115), .A(n7114), .ZN(n11606) );
  NAND2_X1 U9095 ( .A1(n11300), .A2(n8851), .ZN(n11607) );
  AND2_X1 U9096 ( .A1(n11480), .A2(n8850), .ZN(n11301) );
  AOI21_X1 U9097 ( .B1(n8846), .B2(n7257), .A(n6739), .ZN(n11047) );
  NAND2_X1 U9098 ( .A1(n7236), .A2(n8466), .ZN(n10580) );
  NAND2_X1 U9099 ( .A1(n11344), .A2(n8465), .ZN(n7236) );
  NAND2_X1 U9100 ( .A1(n8580), .A2(n8579), .ZN(n12377) );
  NAND2_X1 U9101 ( .A1(n8565), .A2(n8564), .ZN(n12372) );
  INV_X1 U9102 ( .A(n14596), .ZN(n14602) );
  INV_X1 U9103 ( .A(n14994), .ZN(n14991) );
  AND2_X1 U9104 ( .A1(n8802), .A2(n8801), .ZN(n14616) );
  NAND2_X1 U9105 ( .A1(n8791), .A2(n8790), .ZN(n14619) );
  NAND2_X1 U9106 ( .A1(n8743), .A2(n8742), .ZN(n14632) );
  NAND2_X1 U9107 ( .A1(n10973), .A2(n6643), .ZN(n8714) );
  NAND2_X1 U9108 ( .A1(n8650), .A2(n8649), .ZN(n14647) );
  NAND2_X1 U9109 ( .A1(n8554), .A2(n8553), .ZN(n12368) );
  INV_X1 U9110 ( .A(n14643), .ZN(n14648) );
  INV_X1 U9111 ( .A(n12342), .ZN(n12340) );
  INV_X1 U9112 ( .A(n12327), .ZN(n11331) );
  INV_X1 U9113 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8411) );
  INV_X1 U9114 ( .A(n8419), .ZN(n12561) );
  NOR2_X1 U9115 ( .A1(n8404), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7537) );
  NAND2_X1 U9116 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n8403), .ZN(n8891) );
  NAND2_X1 U9117 ( .A1(n9369), .A2(n8380), .ZN(n8765) );
  NAND2_X1 U9118 ( .A1(n8832), .A2(n8831), .ZN(n12498) );
  NAND2_X1 U9119 ( .A1(n8705), .A2(n8693), .ZN(n10683) );
  INV_X1 U9120 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10399) );
  INV_X1 U9121 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10371) );
  INV_X1 U9122 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10079) );
  INV_X1 U9123 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9915) );
  INV_X1 U9124 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9876) );
  INV_X1 U9125 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U9126 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  NAND2_X1 U9127 ( .A1(n7401), .A2(n7400), .ZN(n8529) );
  OR2_X1 U9128 ( .A1(n8500), .A2(n8499), .ZN(n8501) );
  INV_X1 U9129 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9841) );
  INV_X1 U9130 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9857) );
  INV_X1 U9131 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9862) );
  NAND2_X1 U9132 ( .A1(n7130), .A2(n8305), .ZN(n8449) );
  XNOR2_X1 U9133 ( .A(n6969), .B(n8448), .ZN(n14180) );
  NAND2_X1 U9134 ( .A1(n6808), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6969) );
  INV_X1 U9135 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14687) );
  INV_X1 U9136 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7100) );
  XNOR2_X1 U9137 ( .A(n14705), .B(n14702), .ZN(n14775) );
  XNOR2_X1 U9138 ( .A(n14709), .B(n14708), .ZN(n15707) );
  NAND2_X1 U9139 ( .A1(n7102), .A2(n7101), .ZN(n14848) );
  NAND2_X1 U9140 ( .A1(n14724), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7101) );
  AND2_X1 U9141 ( .A1(n14738), .A2(n14737), .ZN(n14856) );
  AND2_X1 U9142 ( .A1(n14747), .A2(n14746), .ZN(n14862) );
  NAND2_X1 U9143 ( .A1(n11120), .A2(n11119), .ZN(n11123) );
  AND3_X1 U9144 ( .A1(n6810), .A2(n6920), .A3(n6919), .ZN(n12813) );
  NAND2_X1 U9145 ( .A1(n13166), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10406) );
  NAND2_X1 U9146 ( .A1(n6975), .A2(n6757), .ZN(n10162) );
  AOI21_X1 U9147 ( .B1(n7064), .B2(n13093), .A(n7062), .ZN(n13168) );
  AOI21_X1 U9148 ( .B1(n6986), .B2(n13132), .A(n6985), .ZN(n12110) );
  XNOR2_X1 U9149 ( .A(n6987), .B(n12108), .ZN(n6986) );
  INV_X1 U9150 ( .A(n9782), .ZN(n9783) );
  OAI22_X1 U9151 ( .A1(n13181), .A2(n13409), .B1(n15699), .B2(n9781), .ZN(
        n9782) );
  OR2_X1 U9152 ( .A1(n7572), .A2(n15699), .ZN(n7569) );
  AOI21_X1 U9153 ( .B1(n13418), .B2(n15699), .A(n7021), .ZN(n13360) );
  NAND2_X1 U9154 ( .A1(n7023), .A2(n7022), .ZN(n7021) );
  NOR2_X1 U9155 ( .A1(n9743), .A2(n9745), .ZN(n9746) );
  NAND2_X1 U9156 ( .A1(n8299), .A2(n8298), .ZN(P3_U3455) );
  NAND2_X1 U9157 ( .A1(n13353), .A2(n13410), .ZN(n8298) );
  NAND2_X1 U9158 ( .A1(n7300), .A2(n7299), .ZN(n8299) );
  NAND2_X1 U9159 ( .A1(n7447), .A2(n13552), .ZN(n7444) );
  INV_X1 U9160 ( .A(n9717), .ZN(n9718) );
  NAND2_X1 U9161 ( .A1(n7158), .A2(n7156), .ZN(P2_U3528) );
  OR2_X1 U9162 ( .A1(n15233), .A2(n7157), .ZN(n7156) );
  NAND2_X1 U9163 ( .A1(n13928), .A2(n15233), .ZN(n7158) );
  INV_X1 U9164 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7157) );
  NAND2_X1 U9165 ( .A1(n14071), .A2(n12162), .ZN(n14825) );
  NAND2_X1 U9166 ( .A1(n6865), .A2(n7176), .ZN(n7175) );
  INV_X1 U9167 ( .A(n12559), .ZN(n7176) );
  OAI21_X1 U9168 ( .B1(n14321), .B2(n14596), .A(n9767), .ZN(n9768) );
  XNOR2_X1 U9169 ( .A(n7107), .B(n14713), .ZN(n14776) );
  XNOR2_X1 U9170 ( .A(n7103), .B(n14724), .ZN(n14778) );
  NOR2_X1 U9171 ( .A1(n14854), .A2(n14853), .ZN(n14852) );
  AND2_X1 U9172 ( .A1(n7099), .A2(n6765), .ZN(n14854) );
  INV_X1 U9173 ( .A(n7249), .ZN(n14859) );
  NAND2_X1 U9174 ( .A1(n14780), .A2(n14781), .ZN(n14779) );
  NAND2_X1 U9175 ( .A1(n7084), .A2(n7082), .ZN(n14767) );
  XNOR2_X1 U9176 ( .A(n7247), .B(n6844), .ZN(SUB_1596_U4) );
  OAI21_X1 U9177 ( .B1(n6963), .B2(n6961), .A(n7087), .ZN(n7247) );
  INV_X1 U9178 ( .A(n14339), .ZN(n7242) );
  INV_X1 U9179 ( .A(n12402), .ZN(n8637) );
  AND2_X1 U9180 ( .A1(n12397), .A2(n12391), .ZN(n12402) );
  NAND2_X1 U9181 ( .A1(n13861), .A2(n13581), .ZN(n6737) );
  NOR2_X1 U9182 ( .A1(n7749), .A2(n15623), .ZN(n6738) );
  AND2_X1 U9183 ( .A1(n12348), .A2(n14153), .ZN(n6739) );
  OAI21_X1 U9184 ( .B1(n13264), .B2(n7291), .A(n7002), .ZN(n13228) );
  AND2_X1 U9185 ( .A1(n8810), .A2(n7227), .ZN(n6740) );
  INV_X1 U9186 ( .A(n12777), .ZN(n12650) );
  NAND2_X1 U9187 ( .A1(n9348), .A2(n9347), .ZN(n13886) );
  INV_X1 U9188 ( .A(n13886), .ZN(n7485) );
  AND2_X1 U9189 ( .A1(n9828), .A2(n6873), .ZN(n6741) );
  AND4_X1 U9190 ( .A1(n7026), .A2(n7025), .A3(n7024), .A4(n8926), .ZN(n6742)
         );
  AND2_X1 U9191 ( .A1(n7277), .A2(n12681), .ZN(n6743) );
  AND2_X1 U9192 ( .A1(n13891), .A2(n13587), .ZN(n6744) );
  AND2_X1 U9193 ( .A1(n12658), .A2(n12659), .ZN(n12770) );
  INV_X1 U9194 ( .A(n12770), .ZN(n7843) );
  AND2_X1 U9195 ( .A1(n13851), .A2(n9714), .ZN(n6745) );
  INV_X1 U9196 ( .A(n6895), .ZN(n13981) );
  OR2_X1 U9197 ( .A1(n7041), .A2(n7653), .ZN(n6746) );
  OR2_X1 U9198 ( .A1(n14853), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6747) );
  AND2_X1 U9199 ( .A1(n9303), .A2(n9302), .ZN(n13814) );
  INV_X1 U9200 ( .A(n13814), .ZN(n13902) );
  AND4_X1 U9201 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n13968)
         );
  NAND2_X1 U9202 ( .A1(n8630), .A2(n8629), .ZN(n14832) );
  INV_X1 U9203 ( .A(n14832), .ZN(n7202) );
  OR2_X1 U9204 ( .A1(n13165), .A2(n7322), .ZN(n7321) );
  INV_X1 U9205 ( .A(n14921), .ZN(n14899) );
  AND2_X1 U9206 ( .A1(n14750), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n6748) );
  AND2_X1 U9207 ( .A1(n8833), .A2(n12502), .ZN(n6749) );
  INV_X2 U9208 ( .A(n11281), .ZN(n12274) );
  AND2_X1 U9209 ( .A1(n8996), .A2(n8995), .ZN(n6750) );
  NAND2_X1 U9210 ( .A1(n7736), .A2(n7735), .ZN(n6928) );
  INV_X1 U9211 ( .A(n7567), .ZN(n8259) );
  XOR2_X1 U9212 ( .A(n13851), .B(n12035), .Z(n6751) );
  INV_X1 U9213 ( .A(n14148), .ZN(n6885) );
  NAND2_X1 U9214 ( .A1(n7567), .A2(n7302), .ZN(n6752) );
  NAND2_X1 U9215 ( .A1(n10217), .A2(n10216), .ZN(n6753) );
  AND2_X1 U9216 ( .A1(n7292), .A2(n7539), .ZN(n7761) );
  NOR2_X1 U9217 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7724) );
  XNOR2_X1 U9218 ( .A(n7741), .B(n7740), .ZN(n10147) );
  INV_X1 U9219 ( .A(n10147), .ZN(n7213) );
  AND2_X1 U9220 ( .A1(n7453), .A2(n7454), .ZN(n6754) );
  OR2_X1 U9221 ( .A1(n12367), .A2(n12366), .ZN(n6755) );
  NAND2_X1 U9222 ( .A1(n9465), .A2(n9464), .ZN(n13648) );
  INV_X1 U9223 ( .A(n9690), .ZN(n13825) );
  AND4_X1 U9224 ( .A1(n15674), .A2(n7663), .A3(n7780), .A4(n7662), .ZN(n6756)
         );
  OR2_X1 U9225 ( .A1(n10123), .A2(n7728), .ZN(n6757) );
  NAND2_X1 U9226 ( .A1(n13275), .A2(n13049), .ZN(n6758) );
  AND2_X1 U9227 ( .A1(n11687), .A2(n7459), .ZN(n6759) );
  INV_X1 U9228 ( .A(n9607), .ZN(n11174) );
  INV_X1 U9229 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13462) );
  NOR2_X1 U9230 ( .A1(n9029), .A2(n9973), .ZN(n6760) );
  INV_X1 U9231 ( .A(n10364), .ZN(n10244) );
  NAND2_X1 U9232 ( .A1(n14073), .A2(n14072), .ZN(n14071) );
  XNOR2_X1 U9233 ( .A(n13358), .B(n13216), .ZN(n13195) );
  OR2_X1 U9234 ( .A1(n13754), .A2(n13876), .ZN(n6761) );
  OR2_X1 U9235 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n14856), .ZN(n6762) );
  AOI21_X1 U9236 ( .B1(n9690), .B2(n9689), .A(n7492), .ZN(n7491) );
  AND2_X1 U9237 ( .A1(n7077), .A2(n7076), .ZN(n6763) );
  NAND2_X1 U9238 ( .A1(n10941), .A2(n10940), .ZN(n6764) );
  XNOR2_X1 U9239 ( .A(n14351), .B(n8821), .ZN(n14339) );
  OR2_X1 U9240 ( .A1(n14732), .A2(n14733), .ZN(n6765) );
  AND2_X1 U9241 ( .A1(n8332), .A2(n8331), .ZN(n8528) );
  AND2_X1 U9242 ( .A1(n13809), .A2(n7491), .ZN(n6766) );
  AND2_X1 U9243 ( .A1(n13562), .A2(n11984), .ZN(n6767) );
  AND2_X1 U9244 ( .A1(n14657), .A2(n9884), .ZN(n14628) );
  INV_X1 U9245 ( .A(n13532), .ZN(n7456) );
  AND2_X1 U9246 ( .A1(n13911), .A2(n12286), .ZN(n6768) );
  INV_X1 U9247 ( .A(n12493), .ZN(n7441) );
  OR2_X1 U9248 ( .A1(n14321), .A2(n14643), .ZN(n6769) );
  NAND2_X1 U9249 ( .A1(n13479), .A2(n11996), .ZN(n13482) );
  NAND2_X1 U9250 ( .A1(n7516), .A2(n12210), .ZN(n13997) );
  INV_X1 U9251 ( .A(n9182), .ZN(n7627) );
  INV_X1 U9252 ( .A(n12376), .ZN(n7189) );
  AND3_X1 U9253 ( .A1(n7150), .A2(n7146), .A3(n7621), .ZN(n6770) );
  OR2_X1 U9254 ( .A1(n7313), .A2(n11208), .ZN(n6771) );
  OR2_X1 U9255 ( .A1(n12288), .A2(n11978), .ZN(n6772) );
  AND2_X1 U9256 ( .A1(n10654), .A2(n10537), .ZN(n6773) );
  NAND2_X1 U9257 ( .A1(n9252), .A2(n9251), .ZN(n13918) );
  AND2_X1 U9258 ( .A1(n13845), .A2(n15196), .ZN(n6774) );
  NOR2_X1 U9259 ( .A1(n15197), .A2(n13603), .ZN(n6775) );
  NAND2_X1 U9260 ( .A1(n8215), .A2(n8218), .ZN(n8257) );
  NOR2_X1 U9261 ( .A1(n6732), .A2(n7703), .ZN(n6776) );
  NOR2_X1 U9262 ( .A1(n13097), .A2(n12062), .ZN(n6777) );
  AND2_X1 U9263 ( .A1(n12398), .A2(n12491), .ZN(n6778) );
  INV_X1 U9264 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n15475) );
  AND2_X1 U9265 ( .A1(n7126), .A2(n7127), .ZN(n6779) );
  AND2_X1 U9266 ( .A1(n14058), .A2(n12233), .ZN(n13982) );
  INV_X1 U9267 ( .A(n13982), .ZN(n7505) );
  INV_X1 U9268 ( .A(n9670), .ZN(n7035) );
  INV_X1 U9269 ( .A(n10224), .ZN(n10216) );
  AND2_X1 U9270 ( .A1(n7784), .A2(n7783), .ZN(n10224) );
  AND2_X1 U9271 ( .A1(n7045), .A2(n7043), .ZN(n6780) );
  AND2_X1 U9272 ( .A1(n12996), .A2(n7358), .ZN(n6781) );
  OR2_X1 U9273 ( .A1(n10022), .A2(n10021), .ZN(n6782) );
  AND2_X1 U9274 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n6783) );
  AND2_X1 U9275 ( .A1(n10087), .A2(n10020), .ZN(n6784) );
  INV_X1 U9276 ( .A(n9374), .ZN(n7636) );
  NOR2_X1 U9277 ( .A1(n12342), .A2(n12341), .ZN(n6785) );
  INV_X1 U9278 ( .A(n9532), .ZN(n7622) );
  INV_X1 U9279 ( .A(n9714), .ZN(n13845) );
  AND2_X1 U9280 ( .A1(n9494), .A2(n9493), .ZN(n9714) );
  AND2_X1 U9281 ( .A1(n7259), .A2(n8855), .ZN(n6786) );
  INV_X1 U9282 ( .A(n12475), .ZN(n14321) );
  NAND2_X1 U9283 ( .A1(n9749), .A2(n9748), .ZN(n12475) );
  INV_X1 U9284 ( .A(n7607), .ZN(n7605) );
  INV_X1 U9285 ( .A(n7584), .ZN(n7583) );
  NAND2_X1 U9286 ( .A1(n7587), .A2(n6768), .ZN(n7584) );
  AND2_X1 U9287 ( .A1(n6765), .A2(n6747), .ZN(n6787) );
  AND2_X1 U9288 ( .A1(n13266), .A2(n7290), .ZN(n6788) );
  AND2_X1 U9289 ( .A1(n12165), .A2(n12164), .ZN(n6789) );
  OR2_X1 U9290 ( .A1(n14724), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6790) );
  INV_X1 U9291 ( .A(n7047), .ZN(n7046) );
  NOR2_X1 U9292 ( .A1(n13799), .A2(n13569), .ZN(n7047) );
  NOR2_X1 U9293 ( .A1(n12377), .A2(n6885), .ZN(n6791) );
  NOR2_X1 U9294 ( .A1(n14647), .A2(n14144), .ZN(n6792) );
  NOR2_X1 U9295 ( .A1(n14616), .A2(n13969), .ZN(n6793) );
  NOR2_X1 U9296 ( .A1(n11033), .A2(n9603), .ZN(n6794) );
  INV_X1 U9297 ( .A(n13325), .ZN(n8061) );
  AND2_X1 U9298 ( .A1(n12714), .A2(n12713), .ZN(n13325) );
  AND2_X1 U9299 ( .A1(n13375), .A2(n13249), .ZN(n6795) );
  INV_X1 U9300 ( .A(n7258), .ZN(n7257) );
  NAND2_X1 U9301 ( .A1(n7658), .A2(n8845), .ZN(n7258) );
  OR2_X1 U9302 ( .A1(n13678), .A2(n12036), .ZN(n6796) );
  AND2_X1 U9303 ( .A1(n12662), .A2(n12663), .ZN(n12774) );
  NAND2_X1 U9304 ( .A1(n13902), .A2(n13488), .ZN(n6797) );
  INV_X1 U9305 ( .A(n9630), .ZN(n13680) );
  INV_X1 U9306 ( .A(n7653), .ZN(n7045) );
  NAND2_X1 U9307 ( .A1(n13215), .A2(n7297), .ZN(n6798) );
  AND2_X1 U9308 ( .A1(n11505), .A2(n13593), .ZN(n6799) );
  AND2_X1 U9309 ( .A1(n12450), .A2(n7436), .ZN(n6800) );
  NAND2_X1 U9310 ( .A1(n12438), .A2(n12436), .ZN(n6801) );
  INV_X1 U9311 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9824) );
  INV_X1 U9312 ( .A(n7291), .ZN(n7290) );
  NAND2_X1 U9313 ( .A1(n8246), .A2(n12730), .ZN(n7291) );
  INV_X1 U9314 ( .A(n7527), .ZN(n7526) );
  NAND2_X1 U9315 ( .A1(n7530), .A2(n7528), .ZN(n7527) );
  AND2_X1 U9316 ( .A1(n6914), .A2(n6911), .ZN(n6802) );
  AND2_X1 U9317 ( .A1(n6751), .A2(n7450), .ZN(n6803) );
  OR2_X1 U9318 ( .A1(n13754), .A2(n7080), .ZN(n6804) );
  AND2_X1 U9319 ( .A1(n7433), .A2(n12431), .ZN(n14468) );
  INV_X1 U9320 ( .A(n14468), .ZN(n7432) );
  INV_X1 U9321 ( .A(n7410), .ZN(n7409) );
  NAND2_X1 U9322 ( .A1(n8348), .A2(n8644), .ZN(n7410) );
  AND2_X1 U9323 ( .A1(n9425), .A2(n9424), .ZN(n13694) );
  INV_X1 U9324 ( .A(n13694), .ZN(n13861) );
  INV_X1 U9325 ( .A(n7598), .ZN(n7597) );
  NAND2_X1 U9326 ( .A1(n9626), .A2(n7600), .ZN(n7598) );
  NOR2_X1 U9327 ( .A1(n13725), .A2(n13583), .ZN(n6805) );
  AND2_X1 U9328 ( .A1(n14332), .A2(n14131), .ZN(n6806) );
  NAND2_X1 U9329 ( .A1(n9826), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6807) );
  INV_X1 U9330 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8405) );
  OR2_X1 U9331 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6808) );
  AND3_X1 U9332 ( .A1(n7651), .A2(n15475), .A3(n7191), .ZN(n6809) );
  OR2_X1 U9333 ( .A1(n9776), .A2(n12761), .ZN(n6810) );
  OR2_X1 U9334 ( .A1(n14701), .A2(n14700), .ZN(n6811) );
  AND2_X1 U9335 ( .A1(n7651), .A2(n15475), .ZN(n6812) );
  AND2_X1 U9336 ( .A1(n7213), .A2(n10134), .ZN(n6813) );
  AND2_X1 U9337 ( .A1(n10160), .A2(n7213), .ZN(n6814) );
  AND2_X1 U9338 ( .A1(n7735), .A2(n7760), .ZN(n6815) );
  INV_X1 U9339 ( .A(n12537), .ZN(n14376) );
  AND2_X1 U9340 ( .A1(n8935), .A2(n8951), .ZN(n6816) );
  AND2_X1 U9341 ( .A1(n13201), .A2(n8171), .ZN(n6817) );
  AND2_X1 U9342 ( .A1(n11121), .A2(n11119), .ZN(n6818) );
  AND2_X1 U9343 ( .A1(n12190), .A2(n12188), .ZN(n6819) );
  OR2_X1 U9344 ( .A1(n9219), .A2(n9217), .ZN(n6820) );
  OR2_X1 U9345 ( .A1(n7636), .A2(n9373), .ZN(n6821) );
  OR2_X1 U9346 ( .A1(n9405), .A2(n9403), .ZN(n6822) );
  OR2_X1 U9347 ( .A1(n7627), .A2(n9181), .ZN(n6823) );
  OR2_X1 U9348 ( .A1(n12460), .A2(n12459), .ZN(n6824) );
  OR2_X1 U9349 ( .A1(n9088), .A2(n9086), .ZN(n6825) );
  AND2_X1 U9350 ( .A1(n7576), .A2(n10978), .ZN(n6826) );
  OR2_X1 U9351 ( .A1(n9125), .A2(n9123), .ZN(n6827) );
  OR2_X1 U9352 ( .A1(n7190), .A2(n7189), .ZN(n6828) );
  AND2_X1 U9353 ( .A1(n7302), .A2(n7691), .ZN(n6829) );
  AND2_X1 U9354 ( .A1(n6894), .A2(n7499), .ZN(n6830) );
  INV_X1 U9355 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10404) );
  INV_X1 U9356 ( .A(n7534), .ZN(n7533) );
  NAND2_X1 U9357 ( .A1(n11288), .A2(n11289), .ZN(n7534) );
  INV_X1 U9358 ( .A(n8513), .ZN(n8327) );
  NAND2_X1 U9359 ( .A1(n7171), .A2(n9838), .ZN(n8513) );
  NAND2_X1 U9360 ( .A1(n11988), .A2(n11987), .ZN(n6831) );
  OR2_X1 U9361 ( .A1(n14583), .A2(n14141), .ZN(n6832) );
  NAND2_X1 U9362 ( .A1(n13532), .A2(n7458), .ZN(n6833) );
  OR2_X1 U9363 ( .A1(n12550), .A2(n12548), .ZN(n6834) );
  INV_X1 U9364 ( .A(n15134), .ZN(n13753) );
  INV_X1 U9365 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7363) );
  AND2_X1 U9366 ( .A1(n6933), .A2(n7905), .ZN(n6835) );
  XNOR2_X1 U9367 ( .A(n7820), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10478) );
  INV_X1 U9368 ( .A(n10478), .ZN(n7305) );
  AND2_X1 U9369 ( .A1(n14781), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6836) );
  AOI21_X1 U9370 ( .B1(n13185), .B2(n8209), .A(n8208), .ZN(n13198) );
  NAND2_X1 U9371 ( .A1(n10963), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6837) );
  OR2_X1 U9372 ( .A1(n13571), .A2(n7463), .ZN(n6838) );
  XNOR2_X1 U9373 ( .A(n14744), .B(n14742), .ZN(n6839) );
  AND2_X1 U9374 ( .A1(n9878), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n6840) );
  AND2_X1 U9375 ( .A1(n7001), .A2(n10957), .ZN(n6841) );
  NAND2_X1 U9376 ( .A1(n12855), .A2(n13042), .ZN(n6842) );
  INV_X1 U9377 ( .A(n10964), .ZN(n7313) );
  INV_X1 U9378 ( .A(n13049), .ZN(n13285) );
  AOI21_X1 U9379 ( .B1(n14027), .B2(n12181), .A(n12180), .ZN(n14042) );
  OAI21_X1 U9380 ( .B1(n11765), .B2(n11764), .A(n11704), .ZN(n11882) );
  AOI21_X1 U9381 ( .B1(n13790), .B2(n9622), .A(n9621), .ZN(n13775) );
  NAND2_X1 U9382 ( .A1(n13304), .A2(n12718), .ZN(n13281) );
  NAND2_X1 U9383 ( .A1(n11177), .A2(n9609), .ZN(n11263) );
  NAND2_X1 U9384 ( .A1(n11796), .A2(n9616), .ZN(n11808) );
  NAND2_X1 U9385 ( .A1(n7475), .A2(n9685), .ZN(n11596) );
  NAND2_X1 U9386 ( .A1(n13336), .A2(n12702), .ZN(n13324) );
  OR2_X1 U9387 ( .A1(n8381), .A2(n10998), .ZN(n6843) );
  INV_X1 U9388 ( .A(n6877), .ZN(n14445) );
  NAND2_X1 U9389 ( .A1(n8778), .A2(n8777), .ZN(n14623) );
  INV_X1 U9390 ( .A(n14623), .ZN(n7200) );
  INV_X1 U9391 ( .A(n14082), .ZN(n6898) );
  XOR2_X1 U9392 ( .A(n14766), .B(n14765), .Z(n6844) );
  NAND2_X1 U9393 ( .A1(n8614), .A2(n8613), .ZN(n12387) );
  OR2_X1 U9394 ( .A1(n14511), .A2(n14583), .ZN(n6845) );
  NAND2_X1 U9395 ( .A1(n7490), .A2(n6766), .ZN(n13808) );
  NAND2_X1 U9396 ( .A1(n7920), .A2(n7919), .ZN(n11676) );
  OR2_X1 U9397 ( .A1(n14511), .A2(n7199), .ZN(n6846) );
  INV_X1 U9398 ( .A(n9335), .ZN(n7633) );
  NOR2_X1 U9399 ( .A1(n11592), .A2(n11505), .ZN(n11591) );
  INV_X1 U9400 ( .A(n7561), .ZN(n7559) );
  NOR2_X1 U9401 ( .A1(n13263), .A2(n7562), .ZN(n7561) );
  AND2_X1 U9402 ( .A1(n12844), .A2(n13274), .ZN(n6847) );
  XNOR2_X1 U9403 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n7832) );
  AND2_X1 U9404 ( .A1(n7090), .A2(n14756), .ZN(n6848) );
  INV_X1 U9405 ( .A(n12854), .ZN(n7347) );
  AND2_X1 U9406 ( .A1(n7307), .A2(n7309), .ZN(n6849) );
  NAND2_X1 U9407 ( .A1(n11591), .A2(n6763), .ZN(n7078) );
  AND2_X1 U9408 ( .A1(n6843), .A2(n9366), .ZN(n6850) );
  INV_X1 U9409 ( .A(n7352), .ZN(n7351) );
  NAND2_X1 U9410 ( .A1(n6842), .A2(n12853), .ZN(n7352) );
  NAND2_X1 U9411 ( .A1(n11464), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6851) );
  INV_X1 U9412 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6884) );
  OR2_X1 U9413 ( .A1(n14252), .A2(n10276), .ZN(n6852) );
  NAND2_X1 U9414 ( .A1(n13411), .A2(n13173), .ZN(n6853) );
  AND2_X1 U9415 ( .A1(n6841), .A2(n6992), .ZN(n6854) );
  INV_X1 U9416 ( .A(n7201), .ZN(n14413) );
  AND2_X1 U9417 ( .A1(n7137), .A2(n7138), .ZN(n6855) );
  INV_X1 U9418 ( .A(n6994), .ZN(n6993) );
  NAND2_X1 U9419 ( .A1(n6996), .A2(n11457), .ZN(n6994) );
  NOR2_X1 U9420 ( .A1(n13073), .A2(n12076), .ZN(n6856) );
  INV_X1 U9421 ( .A(n12718), .ZN(n7008) );
  OR2_X1 U9422 ( .A1(n7633), .A2(n9334), .ZN(n6857) );
  AND2_X1 U9423 ( .A1(n7540), .A2(n7998), .ZN(n6858) );
  INV_X1 U9424 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9873) );
  INV_X1 U9425 ( .A(n14999), .ZN(n13552) );
  AND2_X1 U9426 ( .A1(n15234), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U9427 ( .A1(n9602), .A2(n9601), .ZN(n10893) );
  NAND2_X1 U9428 ( .A1(n7014), .A2(n7274), .ZN(n11249) );
  NAND2_X1 U9429 ( .A1(n7279), .A2(n7277), .ZN(n11675) );
  AND2_X1 U9430 ( .A1(n13166), .A2(n12613), .ZN(n6860) );
  NAND2_X1 U9431 ( .A1(n11358), .A2(n7269), .ZN(n11480) );
  NAND2_X1 U9432 ( .A1(n8215), .A2(n7362), .ZN(n8289) );
  NAND2_X1 U9433 ( .A1(n11480), .A2(n7268), .ZN(n11300) );
  NOR2_X1 U9434 ( .A1(n8045), .A2(n8003), .ZN(n8050) );
  INV_X1 U9435 ( .A(n7205), .ZN(n11604) );
  AND2_X1 U9436 ( .A1(n7529), .A2(n7526), .ZN(n6861) );
  INV_X1 U9437 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10081) );
  AND2_X1 U9438 ( .A1(n8124), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6862) );
  AND2_X1 U9439 ( .A1(n7513), .A2(n7511), .ZN(n6863) );
  NOR2_X1 U9440 ( .A1(n6859), .A2(n7327), .ZN(n6864) );
  INV_X1 U9441 ( .A(n12382), .ZN(n7204) );
  INV_X1 U9442 ( .A(n15197), .ZN(n7069) );
  NAND2_X1 U9443 ( .A1(n8535), .A2(n8534), .ZN(n12363) );
  INV_X1 U9444 ( .A(n12363), .ZN(n7192) );
  BUF_X1 U9445 ( .A(n9543), .Z(n13606) );
  NAND2_X1 U9446 ( .A1(n9136), .A2(n9135), .ZN(n11033) );
  INV_X1 U9447 ( .A(n11033), .ZN(n7073) );
  OR3_X1 U9448 ( .A1(n12558), .A2(n14065), .A3(n12557), .ZN(n6865) );
  INV_X1 U9449 ( .A(n14909), .ZN(n14901) );
  NAND2_X1 U9450 ( .A1(n9179), .A2(n9178), .ZN(n11200) );
  AND2_X1 U9451 ( .A1(n7144), .A2(n9455), .ZN(n6866) );
  INV_X1 U9452 ( .A(n7108), .ZN(n12515) );
  NAND2_X1 U9453 ( .A1(n12300), .A2(n7109), .ZN(n7108) );
  NOR2_X1 U9454 ( .A1(n7326), .A2(n12088), .ZN(n7325) );
  NOR2_X1 U9455 ( .A1(n14750), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n6867) );
  AND2_X1 U9456 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14743), .ZN(n6868) );
  AND2_X1 U9457 ( .A1(n7055), .A2(n7054), .ZN(n6869) );
  AND2_X1 U9458 ( .A1(n7215), .A2(n6753), .ZN(n6870) );
  AND2_X1 U9459 ( .A1(n10426), .A2(n10308), .ZN(n6871) );
  INV_X1 U9460 ( .A(n6944), .ZN(n6943) );
  NOR2_X1 U9461 ( .A1(n6947), .A2(n6945), .ZN(n6944) );
  INV_X1 U9462 ( .A(n6951), .ZN(n6949) );
  NAND2_X1 U9463 ( .A1(n14739), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n6951) );
  NOR2_X1 U9464 ( .A1(n13161), .A2(n12106), .ZN(n6872) );
  INV_X1 U9465 ( .A(n11785), .ZN(n6966) );
  AND2_X1 U9466 ( .A1(n10210), .A2(n10216), .ZN(n10441) );
  NAND2_X1 U9467 ( .A1(n10135), .A2(n10147), .ZN(n10166) );
  INV_X1 U9468 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n12886) );
  XOR2_X1 U9469 ( .A(n7736), .B(n7721), .Z(n6873) );
  INV_X1 U9470 ( .A(SI_10_), .ZN(n7424) );
  NAND2_X1 U9471 ( .A1(n15696), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U9472 ( .A1(n15696), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U9473 ( .A1(n15307), .A2(n15532), .ZN(n7299) );
  INV_X1 U9474 ( .A(n8839), .ZN(n12303) );
  OAI22_X1 U9475 ( .A1(n7426), .A2(n7428), .B1(n12454), .B2(n7427), .ZN(n12457) );
  NAND2_X1 U9476 ( .A1(n11617), .A2(n8623), .ZN(n11661) );
  NAND2_X1 U9477 ( .A1(n7233), .A2(n7232), .ZN(n10752) );
  NAND3_X1 U9478 ( .A1(n6874), .A2(n7639), .A3(n9013), .ZN(n6880) );
  NAND2_X1 U9479 ( .A1(n9008), .A2(n9007), .ZN(n6874) );
  NAND2_X1 U9480 ( .A1(n7234), .A2(n11344), .ZN(n7233) );
  AOI21_X1 U9481 ( .B1(n14336), .B2(n14918), .A(n8836), .ZN(n8873) );
  NAND2_X1 U9482 ( .A1(n7825), .A2(n7824), .ZN(n11251) );
  NAND2_X1 U9483 ( .A1(n13246), .A2(n8138), .ZN(n13231) );
  NAND2_X1 U9484 ( .A1(n7788), .A2(n7787), .ZN(n10737) );
  OAI21_X2 U9485 ( .B1(n9737), .B2(n13310), .A(n9736), .ZN(n13183) );
  AND2_X2 U9486 ( .A1(n7675), .A2(n7676), .ZN(n7567) );
  NAND2_X1 U9487 ( .A1(n6876), .A2(n6891), .ZN(n8461) );
  NAND2_X1 U9488 ( .A1(n6889), .A2(n8450), .ZN(n6876) );
  OAI22_X1 U9489 ( .A1(n13761), .A2(n9623), .B1(n13886), .B2(n13558), .ZN(
        n13743) );
  INV_X1 U9490 ( .A(n7267), .ZN(n7109) );
  INV_X1 U9491 ( .A(n7538), .ZN(n8708) );
  NAND2_X1 U9492 ( .A1(n12297), .A2(n8918), .ZN(n12296) );
  NAND2_X2 U9493 ( .A1(n7340), .A2(n7354), .ZN(n7348) );
  OAI21_X1 U9494 ( .B1(n12943), .B2(n12828), .A(n12830), .ZN(n12963) );
  INV_X1 U9495 ( .A(n12880), .ZN(n10690) );
  NAND2_X1 U9496 ( .A1(n11238), .A2(n11237), .ZN(n12816) );
  NAND3_X1 U9497 ( .A1(n7368), .A2(n8275), .A3(n10300), .ZN(n10303) );
  NAND2_X1 U9498 ( .A1(n14371), .A2(n14616), .ZN(n14356) );
  NAND3_X1 U9499 ( .A1(n12301), .A2(n12300), .A3(n12491), .ZN(n12302) );
  NAND2_X1 U9500 ( .A1(n12400), .A2(n12390), .ZN(n12395) );
  INV_X2 U9501 ( .A(n7750), .ZN(n8112) );
  NAND2_X1 U9502 ( .A1(n11120), .A2(n6818), .ZN(n11238) );
  NAND2_X1 U9503 ( .A1(n12827), .A2(n12826), .ZN(n12943) );
  NAND2_X1 U9504 ( .A1(n13004), .A2(n13285), .ZN(n7340) );
  NAND2_X1 U9505 ( .A1(n12963), .A2(n12962), .ZN(n12834) );
  NAND2_X1 U9506 ( .A1(n6878), .A2(n7626), .ZN(n9200) );
  NAND3_X1 U9507 ( .A1(n9166), .A2(n9165), .A3(n6823), .ZN(n6878) );
  NAND2_X1 U9508 ( .A1(n6879), .A2(n7623), .ZN(n9235) );
  NAND3_X1 U9509 ( .A1(n9205), .A2(n9204), .A3(n6820), .ZN(n6879) );
  OAI21_X2 U9510 ( .B1(n9291), .B2(n9290), .A(n9289), .ZN(n9306) );
  NAND2_X1 U9511 ( .A1(n6880), .A2(n7640), .ZN(n9042) );
  OAI211_X1 U9512 ( .C1(n13848), .C2(n15187), .A(n13847), .B(n13846), .ZN(
        n13928) );
  INV_X1 U9513 ( .A(n9367), .ZN(n7166) );
  NAND2_X1 U9514 ( .A1(n8232), .A2(n12635), .ZN(n12767) );
  NAND2_X1 U9515 ( .A1(n13317), .A2(n8062), .ZN(n13294) );
  NAND2_X1 U9516 ( .A1(n8096), .A2(n8095), .ZN(n13271) );
  NAND2_X1 U9517 ( .A1(n15243), .A2(n15266), .ZN(n12635) );
  NAND2_X1 U9518 ( .A1(n11641), .A2(n7957), .ZN(n11640) );
  AOI21_X1 U9519 ( .B1(n12542), .B2(n8825), .A(n9747), .ZN(n14336) );
  NAND2_X1 U9520 ( .A1(n8601), .A2(n8602), .ZN(n7246) );
  NAND2_X1 U9521 ( .A1(n7538), .A2(n7537), .ZN(n6886) );
  NAND2_X1 U9522 ( .A1(n11522), .A2(n8603), .ZN(n11618) );
  NAND2_X1 U9523 ( .A1(n7240), .A2(n7239), .ZN(n11916) );
  NAND2_X1 U9524 ( .A1(n14345), .A2(n8824), .ZN(n8825) );
  NAND2_X1 U9525 ( .A1(n14761), .A2(n7695), .ZN(n6888) );
  NAND2_X1 U9526 ( .A1(n6890), .A2(n8305), .ZN(n6889) );
  NAND3_X1 U9527 ( .A1(n8303), .A2(SI_0_), .A3(n8304), .ZN(n6890) );
  AND2_X1 U9528 ( .A1(n6892), .A2(n6891), .ZN(n8450) );
  NAND2_X1 U9529 ( .A1(n8307), .A2(n7722), .ZN(n6892) );
  NAND2_X1 U9530 ( .A1(n13998), .A2(n6896), .ZN(n6893) );
  NAND2_X1 U9531 ( .A1(n6893), .A2(n6830), .ZN(n14018) );
  AOI21_X1 U9532 ( .B1(n13998), .B2(n14082), .A(n6899), .ZN(n6895) );
  NAND2_X1 U9533 ( .A1(n14006), .A2(n7517), .ZN(n6902) );
  NAND2_X1 U9534 ( .A1(n7981), .A2(n7385), .ZN(n7382) );
  NAND2_X1 U9535 ( .A1(n7977), .A2(n7976), .ZN(n6907) );
  INV_X1 U9536 ( .A(n13198), .ZN(n6908) );
  NAND2_X1 U9537 ( .A1(n8198), .A2(n9723), .ZN(n12585) );
  NAND2_X1 U9538 ( .A1(n7736), .A2(n6815), .ZN(n6923) );
  NAND3_X1 U9539 ( .A1(n6925), .A2(n6923), .A3(n7776), .ZN(n7779) );
  NAND2_X1 U9540 ( .A1(n7904), .A2(n6835), .ZN(n6931) );
  NAND3_X1 U9541 ( .A1(n12755), .A2(n12746), .A3(n12763), .ZN(n6935) );
  NAND2_X1 U9542 ( .A1(n8126), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U9543 ( .A1(n8143), .A2(n8142), .ZN(n8159) );
  AOI22_X1 U9544 ( .A1(n10184), .A2(n10403), .B1(n7221), .B2(n10122), .ZN(
        n10421) );
  AOI21_X1 U9545 ( .B1(n6976), .B2(n10161), .A(n6814), .ZN(n6970) );
  INV_X1 U9546 ( .A(n10161), .ZN(n6971) );
  NAND2_X1 U9547 ( .A1(n12104), .A2(n13167), .ZN(n6988) );
  NAND2_X1 U9548 ( .A1(n6995), .A2(n6996), .ZN(n11458) );
  NAND2_X1 U9549 ( .A1(n6998), .A2(n10957), .ZN(n11231) );
  OR2_X1 U9550 ( .A1(n10959), .A2(n10958), .ZN(n6998) );
  NAND2_X1 U9551 ( .A1(n13302), .A2(n12718), .ZN(n7005) );
  NAND2_X1 U9552 ( .A1(n7005), .A2(n7006), .ZN(n8244) );
  NAND2_X1 U9553 ( .A1(n7010), .A2(n7011), .ZN(n11077) );
  NAND2_X1 U9554 ( .A1(n7013), .A2(n10734), .ZN(n7010) );
  NAND3_X1 U9555 ( .A1(n7017), .A2(n7018), .A3(n7016), .ZN(n7729) );
  NAND2_X1 U9556 ( .A1(n10809), .A2(n7746), .ZN(n12633) );
  NAND2_X1 U9557 ( .A1(n8240), .A2(n7020), .ZN(n13336) );
  NAND2_X1 U9558 ( .A1(n13336), .A2(n7294), .ZN(n8242) );
  XNOR2_X1 U9559 ( .A(n13605), .B(n15183), .ZN(n10598) );
  OAI21_X1 U9560 ( .B1(n10491), .B2(n7052), .A(n7051), .ZN(n11208) );
  NAND2_X1 U9561 ( .A1(n11570), .A2(n7058), .ZN(n7057) );
  NOR2_X1 U9562 ( .A1(n11570), .A2(n11569), .ZN(n12072) );
  NAND2_X1 U9563 ( .A1(n10413), .A2(n10134), .ZN(n10135) );
  NAND2_X1 U9564 ( .A1(n10413), .A2(n6813), .ZN(n7330) );
  NAND3_X1 U9565 ( .A1(n13163), .A2(n13164), .A3(n7063), .ZN(n7062) );
  AOI21_X1 U9566 ( .B1(n13659), .B2(n13845), .A(n12009), .ZN(n7072) );
  NAND2_X1 U9567 ( .A1(n11591), .A2(n7075), .ZN(n13811) );
  INV_X1 U9568 ( .A(n7078), .ZN(n13834) );
  NAND2_X1 U9569 ( .A1(n8932), .A2(n8957), .ZN(n8956) );
  NAND3_X1 U9570 ( .A1(n8932), .A2(n8957), .A3(n8933), .ZN(n8955) );
  OAI21_X1 U9571 ( .B1(n15705), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6811), .ZN(
        n7081) );
  XNOR2_X1 U9572 ( .A(n14701), .B(n14700), .ZN(n15705) );
  NOR2_X1 U9573 ( .A1(n14857), .A2(n6839), .ZN(n7092) );
  INV_X1 U9574 ( .A(n14857), .ZN(n7093) );
  NAND2_X1 U9575 ( .A1(n7249), .A2(n7248), .ZN(n7096) );
  INV_X1 U9576 ( .A(n7095), .ZN(n14860) );
  NAND2_X1 U9577 ( .A1(n15712), .A2(n15713), .ZN(n14689) );
  XNOR2_X1 U9578 ( .A(n14688), .B(n7100), .ZN(n15712) );
  XNOR2_X1 U9579 ( .A(n14685), .B(n14686), .ZN(n14688) );
  NAND2_X1 U9580 ( .A1(n7103), .A2(n6790), .ZN(n7102) );
  NAND2_X1 U9581 ( .A1(n7107), .A2(n7104), .ZN(n7106) );
  NAND2_X1 U9582 ( .A1(n11480), .A2(n7114), .ZN(n7110) );
  NAND2_X1 U9583 ( .A1(n7110), .A2(n7111), .ZN(n11526) );
  NAND2_X1 U9584 ( .A1(n14388), .A2(n7116), .ZN(n14379) );
  NAND2_X1 U9585 ( .A1(n14457), .A2(n8858), .ZN(n7119) );
  NAND2_X2 U9586 ( .A1(n11968), .A2(n14169), .ZN(n9884) );
  XNOR2_X2 U9587 ( .A(n7123), .B(n8410), .ZN(n11968) );
  XNOR2_X1 U9588 ( .A(n9753), .B(n12540), .ZN(n7128) );
  NAND2_X1 U9589 ( .A1(n7128), .A2(n14899), .ZN(n7126) );
  NOR2_X2 U9590 ( .A1(n9760), .A2(n7125), .ZN(n7124) );
  NAND2_X1 U9591 ( .A1(n7461), .A2(n6772), .ZN(n7460) );
  XNOR2_X1 U9592 ( .A(n11686), .B(n11684), .ZN(n11512) );
  NAND4_X1 U9593 ( .A1(n8303), .A2(n8304), .A3(n8305), .A4(SI_0_), .ZN(n7130)
         );
  NAND2_X1 U9594 ( .A1(n8304), .A2(SI_0_), .ZN(n8430) );
  NAND2_X1 U9595 ( .A1(n8303), .A2(n8305), .ZN(n8429) );
  NAND2_X1 U9596 ( .A1(n12582), .A2(n7134), .ZN(n12130) );
  NAND2_X1 U9597 ( .A1(n7137), .A2(n7135), .ZN(n13510) );
  NAND3_X1 U9598 ( .A1(n7143), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7142) );
  NAND2_X1 U9599 ( .A1(n7145), .A2(n9498), .ZN(n9499) );
  NAND3_X1 U9600 ( .A1(n9523), .A2(n7149), .A3(n9540), .ZN(n7148) );
  NAND3_X1 U9601 ( .A1(n7396), .A2(n7398), .A3(n8332), .ZN(n8544) );
  AOI21_X2 U9602 ( .B1(n9640), .B2(n15131), .A(n9639), .ZN(n13847) );
  NAND2_X1 U9603 ( .A1(n9367), .A2(n7159), .ZN(n7164) );
  NAND3_X1 U9604 ( .A1(n7164), .A2(n7163), .A3(n8382), .ZN(n8776) );
  INV_X1 U9605 ( .A(n8800), .ZN(n7168) );
  MUX2_X1 U9606 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8407), .Z(n8326) );
  OAI21_X1 U9607 ( .B1(n12384), .B2(n7174), .A(n7172), .ZN(n12400) );
  OAI21_X1 U9608 ( .B1(n12399), .B2(n6651), .A(n7180), .ZN(n7179) );
  INV_X1 U9609 ( .A(n12461), .ZN(n12464) );
  NAND2_X1 U9610 ( .A1(n12437), .A2(n7185), .ZN(n7183) );
  NAND2_X1 U9611 ( .A1(n7183), .A2(n7184), .ZN(n12441) );
  INV_X1 U9612 ( .A(n12375), .ZN(n7190) );
  NAND2_X1 U9613 ( .A1(n8647), .A2(n6812), .ZN(n8874) );
  AND2_X1 U9614 ( .A1(n8647), .A2(n6809), .ZN(n8828) );
  INV_X2 U9615 ( .A(n12495), .ZN(n8712) );
  NAND2_X1 U9616 ( .A1(n9754), .A2(n14321), .ZN(n14314) );
  NAND2_X1 U9617 ( .A1(n9754), .A2(n7193), .ZN(n7195) );
  INV_X1 U9618 ( .A(n7195), .ZN(n14312) );
  NOR2_X2 U9619 ( .A1(n14396), .A2(n14619), .ZN(n14371) );
  NAND2_X1 U9620 ( .A1(n7211), .A2(n10175), .ZN(n10173) );
  INV_X1 U9621 ( .A(n10148), .ZN(n7214) );
  INV_X1 U9622 ( .A(n10217), .ZN(n7218) );
  NAND2_X1 U9623 ( .A1(n7221), .A2(n10131), .ZN(n10132) );
  XNOR2_X1 U9624 ( .A(n10121), .B(n7221), .ZN(n10184) );
  NAND2_X1 U9625 ( .A1(n13166), .A2(n7221), .ZN(n10196) );
  OAI21_X1 U9626 ( .B1(n13098), .B2(n7223), .A(n7222), .ZN(n13115) );
  NAND2_X1 U9627 ( .A1(n14368), .A2(n6740), .ZN(n7225) );
  NAND2_X1 U9628 ( .A1(n14327), .A2(n14918), .ZN(n7231) );
  OAI21_X1 U9629 ( .B1(n7235), .B2(n8479), .A(n8478), .ZN(n7232) );
  AND2_X1 U9630 ( .A1(n8465), .A2(n8478), .ZN(n7234) );
  NAND2_X1 U9631 ( .A1(n11661), .A2(n8659), .ZN(n7240) );
  INV_X1 U9632 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7248) );
  XNOR2_X1 U9633 ( .A(n14718), .B(n14717), .ZN(n14777) );
  NAND2_X1 U9634 ( .A1(n8647), .A2(n7251), .ZN(n8893) );
  NAND2_X1 U9635 ( .A1(n8846), .A2(n7256), .ZN(n7253) );
  NAND2_X1 U9636 ( .A1(n7253), .A2(n7254), .ZN(n11354) );
  NAND2_X1 U9637 ( .A1(n14405), .A2(n14410), .ZN(n7265) );
  NAND3_X1 U9638 ( .A1(n8448), .A2(n7266), .A3(n8432), .ZN(n8458) );
  XNOR2_X1 U9639 ( .A(n9752), .B(n12542), .ZN(n7272) );
  NAND2_X1 U9640 ( .A1(n11192), .A2(n7281), .ZN(n7279) );
  INV_X1 U9641 ( .A(n12686), .ZN(n7289) );
  NAND2_X1 U9642 ( .A1(n11647), .A2(n8239), .ZN(n11646) );
  NAND3_X1 U9643 ( .A1(n7293), .A2(n7705), .A3(n7704), .ZN(n13061) );
  NAND2_X1 U9644 ( .A1(n13061), .A2(n10248), .ZN(n10674) );
  AOI21_X1 U9645 ( .B1(n13213), .B2(n7297), .A(n7295), .ZN(n9739) );
  OR2_X1 U9646 ( .A1(n13213), .A2(n13212), .ZN(n13215) );
  NAND2_X1 U9647 ( .A1(n7567), .A2(n6829), .ZN(n7680) );
  INV_X1 U9648 ( .A(n7304), .ZN(n12085) );
  OR2_X1 U9649 ( .A1(n12084), .A2(n13148), .ZN(n7304) );
  MUX2_X1 U9650 ( .A(n13468), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  MUX2_X1 U9651 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13468), .S(n7723), .Z(n10248)
         );
  OR2_X1 U9652 ( .A1(n13109), .A2(n13110), .ZN(n7307) );
  OAI211_X1 U9653 ( .C1(n12081), .C2(P3_REG1_REG_15__SCAN_IN), .A(n7308), .B(
        n7311), .ZN(n7310) );
  NAND2_X1 U9654 ( .A1(n7309), .A2(n13109), .ZN(n7308) );
  INV_X1 U9655 ( .A(n12081), .ZN(n7309) );
  INV_X1 U9656 ( .A(n13127), .ZN(n7311) );
  XNOR2_X1 U9657 ( .A(n12080), .B(n13107), .ZN(n13109) );
  OAI21_X1 U9658 ( .B1(n13074), .B2(n7316), .A(n7314), .ZN(n12079) );
  OAI211_X1 U9659 ( .C1(n13162), .C2(n7320), .A(n7318), .B(n6864), .ZN(n12109)
         );
  NAND2_X1 U9660 ( .A1(n13162), .A2(n7319), .ZN(n7318) );
  INV_X1 U9661 ( .A(n12106), .ZN(n7326) );
  NAND2_X1 U9662 ( .A1(n7329), .A2(n10166), .ZN(n10164) );
  INV_X1 U9663 ( .A(n10441), .ZN(n7331) );
  OAI211_X1 U9664 ( .C1(n6871), .C2(n10674), .A(n10427), .B(n10314), .ZN(
        n10315) );
  NAND3_X1 U9665 ( .A1(n7337), .A2(n7342), .A3(n7335), .ZN(n12902) );
  NAND2_X1 U9666 ( .A1(n8215), .A2(n7361), .ZN(n7360) );
  NAND2_X1 U9667 ( .A1(n7360), .A2(n8258), .ZN(n8263) );
  NAND2_X1 U9668 ( .A1(n12982), .A2(n7365), .ZN(n12869) );
  NAND2_X1 U9669 ( .A1(n12745), .A2(n12794), .ZN(n7369) );
  NAND2_X1 U9670 ( .A1(n7370), .A2(n7369), .ZN(n7373) );
  NAND2_X1 U9671 ( .A1(n7371), .A2(n7374), .ZN(n7370) );
  INV_X1 U9672 ( .A(n12794), .ZN(n7371) );
  NAND3_X1 U9673 ( .A1(n12752), .A2(n12753), .A3(n7372), .ZN(n12755) );
  NAND3_X1 U9674 ( .A1(n7373), .A2(n12904), .A3(n12748), .ZN(n7372) );
  OAI21_X1 U9675 ( .B1(n12739), .B2(n12740), .A(n12738), .ZN(n7374) );
  NAND2_X1 U9676 ( .A1(n7382), .A2(n7383), .ZN(n8023) );
  NAND3_X1 U9677 ( .A1(n7393), .A2(n7395), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n7394) );
  INV_X1 U9678 ( .A(n7400), .ZN(n7397) );
  NAND3_X1 U9679 ( .A1(n8528), .A2(n8500), .A3(n7399), .ZN(n7398) );
  NAND2_X1 U9680 ( .A1(n8640), .A2(n7406), .ZN(n7404) );
  NAND2_X1 U9681 ( .A1(n12452), .A2(n12451), .ZN(n7426) );
  INV_X2 U9682 ( .A(n12491), .ZN(n7430) );
  INV_X1 U9683 ( .A(n12492), .ZN(n7440) );
  NAND2_X1 U9684 ( .A1(n13470), .A2(n7443), .ZN(n7442) );
  OAI211_X1 U9685 ( .C1(n13470), .C2(n7444), .A(n12042), .B(n7442), .ZN(
        P2_U3192) );
  INV_X1 U9686 ( .A(n13522), .ZN(n7458) );
  INV_X1 U9687 ( .A(n7461), .ZN(n12291) );
  NAND2_X1 U9688 ( .A1(n7460), .A2(n12289), .ZN(n12295) );
  NAND2_X1 U9689 ( .A1(n9796), .A2(n13504), .ZN(n13502) );
  NAND3_X1 U9690 ( .A1(n12054), .A2(n9803), .A3(n9808), .ZN(n10549) );
  NAND3_X1 U9691 ( .A1(n12126), .A2(n11010), .A3(n11015), .ZN(n11017) );
  NAND3_X1 U9692 ( .A1(n11017), .A2(n11016), .A3(n11026), .ZN(n11493) );
  AND3_X2 U9693 ( .A1(n8958), .A2(n6742), .A3(n7465), .ZN(n8932) );
  NAND3_X1 U9694 ( .A1(n8979), .A2(n9829), .A3(n7467), .ZN(n7466) );
  INV_X1 U9695 ( .A(n9874), .ZN(n7467) );
  NAND2_X2 U9696 ( .A1(n8979), .A2(n9829), .ZN(n9370) );
  NOR2_X1 U9697 ( .A1(n13748), .A2(n7482), .ZN(n7481) );
  NAND2_X1 U9698 ( .A1(n7488), .A2(n7486), .ZN(n9682) );
  NAND3_X1 U9699 ( .A1(n8979), .A2(n9828), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n8986) );
  OAI22_X1 U9700 ( .A1(n8979), .A2(n9935), .B1(n9872), .B2(n7489), .ZN(n9004)
         );
  OAI22_X1 U9701 ( .A1(n8979), .A2(n10011), .B1(n9826), .B2(n7489), .ZN(n9019)
         );
  OAI22_X1 U9702 ( .A1(n8979), .A2(n9941), .B1(n9843), .B2(n7489), .ZN(n9062)
         );
  OAI22_X1 U9703 ( .A1(n8979), .A2(n15010), .B1(n9827), .B2(n7489), .ZN(n9037)
         );
  OAI22_X1 U9704 ( .A1(n8979), .A2(n9972), .B1(n9848), .B2(n7489), .ZN(n9084)
         );
  OAI22_X1 U9705 ( .A1(n15037), .A2(n8979), .B1(n9861), .B2(n7489), .ZN(n9100)
         );
  OAI22_X1 U9706 ( .A1(n8979), .A2(n10260), .B1(n9878), .B2(n7489), .ZN(n9134)
         );
  OAI22_X1 U9707 ( .A1(n8979), .A2(n10375), .B1(n9889), .B2(n7489), .ZN(n9156)
         );
  OAI22_X1 U9708 ( .A1(n8979), .A2(n10834), .B1(n9917), .B2(n7489), .ZN(n9177)
         );
  OAI22_X1 U9709 ( .A1(n8979), .A2(n11442), .B1(n10395), .B2(n7489), .ZN(n9250) );
  OAI22_X1 U9710 ( .A1(n8979), .A2(n13627), .B1(n10326), .B2(n7489), .ZN(n9256) );
  NAND2_X1 U9711 ( .A1(n11819), .A2(n9690), .ZN(n7490) );
  INV_X1 U9712 ( .A(n7493), .ZN(n13826) );
  AND3_X2 U9713 ( .A1(n6639), .A2(n8400), .A3(n6640), .ZN(n8647) );
  NAND2_X1 U9714 ( .A1(n7495), .A2(n7496), .ZN(n12280) );
  NAND2_X1 U9715 ( .A1(n14106), .A2(n7497), .ZN(n7495) );
  NAND2_X1 U9716 ( .A1(n14106), .A2(n14107), .ZN(n14105) );
  INV_X1 U9717 ( .A(n10720), .ZN(n7509) );
  NAND2_X1 U9718 ( .A1(n7507), .A2(n6764), .ZN(n7506) );
  XNOR2_X1 U9719 ( .A(n11140), .B(n11138), .ZN(n10945) );
  NAND2_X1 U9720 ( .A1(n7516), .A2(n7514), .ZN(n13998) );
  NAND2_X1 U9721 ( .A1(n7522), .A2(n6819), .ZN(n13988) );
  OAI21_X1 U9722 ( .B1(n11823), .B2(n7542), .A(n6858), .ZN(n7546) );
  INV_X1 U9723 ( .A(n7546), .ZN(n11924) );
  NAND2_X1 U9724 ( .A1(n7920), .A2(n7547), .ZN(n11641) );
  NAND2_X1 U9725 ( .A1(n7550), .A2(n6817), .ZN(n13193) );
  OAI21_X2 U9726 ( .B1(n13271), .B2(n7556), .A(n7554), .ZN(n13246) );
  NAND2_X1 U9727 ( .A1(n8231), .A2(n7570), .ZN(n7568) );
  OAI21_X1 U9728 ( .B1(n7571), .B2(n7568), .A(n7569), .ZN(n13354) );
  AND2_X1 U9729 ( .A1(n8231), .A2(n8230), .ZN(n13192) );
  NAND2_X1 U9730 ( .A1(n9602), .A2(n7577), .ZN(n7575) );
  INV_X1 U9731 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8927) );
  NAND3_X1 U9732 ( .A1(n7589), .A2(n7588), .A3(n8927), .ZN(n8962) );
  NOR2_X2 U9733 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7588) );
  NAND2_X1 U9734 ( .A1(n9624), .A2(n13585), .ZN(n7607) );
  INV_X2 U9735 ( .A(n8944), .ZN(n13951) );
  NAND2_X2 U9736 ( .A1(n8944), .A2(n8943), .ZN(n9506) );
  AND2_X4 U9737 ( .A1(n7608), .A2(n13946), .ZN(n8944) );
  NAND2_X1 U9738 ( .A1(n15138), .A2(n15126), .ZN(n15125) );
  NAND3_X1 U9739 ( .A1(n7610), .A2(n9593), .A3(n7609), .ZN(n10599) );
  NAND2_X1 U9740 ( .A1(n10065), .A2(n7611), .ZN(n7609) );
  INV_X1 U9741 ( .A(n9591), .ZN(n7611) );
  NAND2_X1 U9742 ( .A1(n10063), .A2(n10065), .ZN(n10064) );
  NAND2_X1 U9743 ( .A1(n15125), .A2(n9591), .ZN(n10063) );
  OAI21_X1 U9744 ( .B1(n11177), .B2(n9612), .A(n7612), .ZN(n9614) );
  NAND2_X4 U9745 ( .A1(n7615), .A2(n8944), .ZN(n9482) );
  INV_X1 U9746 ( .A(n9442), .ZN(n7618) );
  INV_X1 U9747 ( .A(n9443), .ZN(n7620) );
  AND2_X2 U9748 ( .A1(n7616), .A2(n6770), .ZN(n9564) );
  NAND3_X1 U9749 ( .A1(n7620), .A2(n7618), .A3(n7619), .ZN(n7616) );
  NAND2_X1 U9750 ( .A1(n7624), .A2(n7625), .ZN(n9139) );
  NAND3_X1 U9751 ( .A1(n9110), .A2(n6827), .A3(n9109), .ZN(n7624) );
  NAND2_X1 U9752 ( .A1(n7628), .A2(n7629), .ZN(n9105) );
  NAND3_X1 U9753 ( .A1(n9072), .A2(n6825), .A3(n9071), .ZN(n7628) );
  NAND2_X1 U9754 ( .A1(n7631), .A2(n7632), .ZN(n9351) );
  NAND3_X1 U9755 ( .A1(n9325), .A2(n6857), .A3(n9324), .ZN(n7631) );
  NAND2_X1 U9756 ( .A1(n7634), .A2(n7635), .ZN(n9387) );
  NAND3_X1 U9757 ( .A1(n9356), .A2(n6821), .A3(n9355), .ZN(n7634) );
  NAND2_X1 U9758 ( .A1(n7637), .A2(n7638), .ZN(n9428) );
  NAND3_X1 U9759 ( .A1(n9392), .A2(n6822), .A3(n9391), .ZN(n7637) );
  OR2_X1 U9760 ( .A1(n9026), .A2(n9028), .ZN(n7639) );
  OR2_X1 U9761 ( .A1(n7641), .A2(n9027), .ZN(n7640) );
  NAND2_X1 U9762 ( .A1(n8934), .A2(n7642), .ZN(n8941) );
  XNOR2_X1 U9763 ( .A(n8576), .B(n8575), .ZN(n9914) );
  XNOR2_X1 U9764 ( .A(n12614), .B(n12800), .ZN(n12805) );
  INV_X2 U9765 ( .A(n12849), .ZN(n12856) );
  NAND2_X1 U9766 ( .A1(n12856), .A2(n12624), .ZN(n10305) );
  INV_X1 U9767 ( .A(n11997), .ZN(n11999) );
  INV_X1 U9768 ( .A(n13195), .ZN(n13201) );
  CLKBUF_X1 U9769 ( .A(n11641), .Z(n11677) );
  NAND2_X1 U9770 ( .A1(n10848), .A2(n12885), .ZN(n8232) );
  INV_X1 U9771 ( .A(n13790), .ZN(n13791) );
  NAND2_X1 U9772 ( .A1(n12625), .A2(n12624), .ZN(n10312) );
  NAND2_X1 U9773 ( .A1(n8412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8413) );
  OAI21_X1 U9774 ( .B1(n13848), .B2(n15139), .A(n9716), .ZN(n9717) );
  OR2_X1 U9775 ( .A1(n8112), .A2(n10120), .ZN(n7734) );
  AND3_X2 U9776 ( .A1(n7733), .A2(n7732), .A3(n7731), .ZN(n7655) );
  NOR2_X1 U9777 ( .A1(n12612), .A2(n12611), .ZN(n12614) );
  OR2_X1 U9778 ( .A1(n8953), .A2(n13945), .ZN(n8938) );
  OR2_X1 U9779 ( .A1(n13661), .A2(n9482), .ZN(n9478) );
  OR2_X1 U9780 ( .A1(n13534), .A2(n9482), .ZN(n9400) );
  INV_X1 U9781 ( .A(n9482), .ZN(n9429) );
  OR2_X1 U9782 ( .A1(n9482), .A2(n15133), .ZN(n8978) );
  OR2_X1 U9783 ( .A1(n9482), .A2(n9978), .ZN(n8945) );
  AND2_X2 U9784 ( .A1(n10669), .A2(n9780), .ZN(n15699) );
  INV_X2 U9785 ( .A(n15307), .ZN(n15309) );
  XOR2_X1 U9786 ( .A(n14917), .B(n14916), .Z(n7643) );
  NAND3_X1 U9787 ( .A1(n11970), .A2(n10661), .A3(n10660), .ZN(n15222) );
  OR2_X1 U9788 ( .A1(n12151), .A2(n12150), .ZN(n7644) );
  AND2_X1 U9789 ( .A1(n6769), .A2(n9763), .ZN(n7645) );
  AND2_X2 U9790 ( .A1(n9764), .A2(n8922), .ZN(n14987) );
  INV_X1 U9791 ( .A(n14301), .ZN(n8918) );
  AND2_X1 U9792 ( .A1(n14977), .A2(n14976), .ZN(n7646) );
  NOR3_X1 U9793 ( .A1(n13691), .A2(n13690), .A3(n9794), .ZN(n7647) );
  NAND2_X1 U9794 ( .A1(n8959), .A2(n8927), .ZN(n9253) );
  XOR2_X1 U9795 ( .A(n14894), .B(n14893), .Z(n7649) );
  AND2_X1 U9796 ( .A1(n10626), .A2(n10625), .ZN(n7650) );
  AND4_X1 U9797 ( .A1(n8402), .A2(n8678), .A3(n8662), .A4(n8401), .ZN(n7651)
         );
  OR2_X1 U9798 ( .A1(n9446), .A2(n9447), .ZN(n7652) );
  INV_X1 U9799 ( .A(n15298), .ZN(n9740) );
  INV_X1 U9800 ( .A(n13339), .ZN(n8241) );
  AND2_X1 U9801 ( .A1(n9693), .A2(n13513), .ZN(n7653) );
  INV_X1 U9802 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9111) );
  INV_X1 U9803 ( .A(n10549), .ZN(n9809) );
  NAND2_X1 U9804 ( .A1(n8876), .A2(n8875), .ZN(n8884) );
  INV_X1 U9805 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14708) );
  OR2_X1 U9806 ( .A1(n13851), .A2(n15215), .ZN(n7654) );
  INV_X1 U9807 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8300) );
  NOR2_X1 U9808 ( .A1(n13181), .A2(n13456), .ZN(n9743) );
  INV_X1 U9809 ( .A(n13301), .ZN(n8243) );
  INV_X1 U9810 ( .A(n12785), .ZN(n8239) );
  INV_X1 U9811 ( .A(n13107), .ZN(n12060) );
  AND2_X1 U9812 ( .A1(n9269), .A2(n9688), .ZN(n7656) );
  XNOR2_X1 U9813 ( .A(n12607), .B(n12749), .ZN(n7657) );
  OR2_X1 U9814 ( .A1(n12348), .A2(n14153), .ZN(n7658) );
  INV_X1 U9815 ( .A(n13918), .ZN(n9708) );
  INV_X1 U9816 ( .A(n12518), .ZN(n8497) );
  NOR3_X1 U9817 ( .A1(n13675), .A2(n13674), .A3(n9794), .ZN(n7659) );
  OR2_X1 U9818 ( .A1(n11140), .A2(n11139), .ZN(n7660) );
  AND2_X1 U9819 ( .A1(n14971), .A2(n14970), .ZN(n7661) );
  INV_X1 U9820 ( .A(n12524), .ZN(n11481) );
  INV_X1 U9821 ( .A(n9027), .ZN(n9028) );
  NAND2_X1 U9822 ( .A1(n12491), .A2(n12306), .ZN(n12307) );
  NAND2_X1 U9823 ( .A1(n12312), .A2(n12311), .ZN(n12317) );
  INV_X1 U9824 ( .A(n12317), .ZN(n12315) );
  INV_X1 U9825 ( .A(n12391), .ZN(n12392) );
  AND2_X1 U9826 ( .A1(n12414), .A2(n12413), .ZN(n12415) );
  AND3_X1 U9827 ( .A1(n9266), .A2(n9688), .A3(n9265), .ZN(n9291) );
  INV_X1 U9828 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8397) );
  INV_X1 U9829 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7664) );
  INV_X1 U9830 ( .A(n8691), .ZN(n8361) );
  INV_X1 U9831 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8951) );
  INV_X1 U9832 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8401) );
  INV_X1 U9833 ( .A(n12783), .ZN(n7938) );
  INV_X1 U9834 ( .A(n12775), .ZN(n7787) );
  AND2_X1 U9835 ( .A1(n8049), .A2(n7674), .ZN(n7675) );
  OAI22_X1 U9836 ( .A1(n12274), .A2(n14908), .B1(n10349), .B2(n10348), .ZN(
        n10350) );
  NAND2_X1 U9837 ( .A1(n8800), .A2(n11557), .ZN(n8393) );
  INV_X1 U9838 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15543) );
  INV_X1 U9839 ( .A(n11963), .ZN(n7685) );
  INV_X1 U9840 ( .A(n12742), .ZN(n8249) );
  INV_X1 U9841 ( .A(n12789), .ZN(n8016) );
  INV_X1 U9842 ( .A(n7847), .ZN(n7846) );
  INV_X1 U9843 ( .A(n9277), .ZN(n9275) );
  INV_X1 U9844 ( .A(n9814), .ZN(n9808) );
  INV_X1 U9845 ( .A(n9407), .ZN(n9406) );
  INV_X1 U9846 ( .A(n9243), .ZN(n9241) );
  OR2_X1 U9847 ( .A1(n9416), .A2(n12018), .ZN(n9471) );
  NOR2_X1 U9848 ( .A1(n13711), .A2(n12011), .ZN(n9698) );
  AND2_X1 U9849 ( .A1(n14021), .A2(n12242), .ZN(n14056) );
  INV_X1 U9850 ( .A(n14351), .ZN(n8823) );
  INV_X1 U9851 ( .A(n14385), .ZN(n8863) );
  INV_X1 U9852 ( .A(n14146), .ZN(n12389) );
  INV_X1 U9853 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8403) );
  AND2_X1 U9854 ( .A1(n8351), .A2(n8643), .ZN(n8352) );
  NAND2_X1 U9855 ( .A1(n8317), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U9856 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n14177), .ZN(n14661) );
  NAND2_X1 U9857 ( .A1(n7949), .A2(n15543), .ZN(n7967) );
  OR2_X1 U9858 ( .A1(n8010), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8031) );
  INV_X1 U9859 ( .A(n8073), .ZN(n8072) );
  INV_X1 U9860 ( .A(n11124), .ZN(n11121) );
  NAND2_X2 U9861 ( .A1(n11960), .A2(n11963), .ZN(n7754) );
  OAI22_X1 U9862 ( .A1(n7724), .A2(n7725), .B1(P3_IR_REG_2__SCAN_IN), .B2(
        P3_IR_REG_31__SCAN_IN), .ZN(n7727) );
  NOR2_X1 U9863 ( .A1(n11216), .A2(n11215), .ZN(n11219) );
  AND2_X1 U9864 ( .A1(n12083), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12064) );
  INV_X1 U9865 ( .A(n13247), .ZN(n8246) );
  OR2_X1 U9866 ( .A1(n8055), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8073) );
  NOR2_X1 U9867 ( .A1(n13198), .A2(n13314), .ZN(n9735) );
  NAND2_X1 U9868 ( .A1(n8174), .A2(n8173), .ZN(n8176) );
  XNOR2_X1 U9869 ( .A(n11099), .B(n12033), .ZN(n12112) );
  NAND2_X1 U9870 ( .A1(n9275), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9293) );
  XNOR2_X1 U9871 ( .A(n11033), .B(n12033), .ZN(n11007) );
  INV_X1 U9872 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9049) );
  INV_X1 U9873 ( .A(n8972), .ZN(n9510) );
  NAND2_X1 U9874 ( .A1(n9406), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U9875 ( .A1(n9241), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9260) );
  AND2_X1 U9876 ( .A1(n9505), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8942) );
  INV_X1 U9877 ( .A(n10639), .ZN(n9671) );
  INV_X1 U9878 ( .A(n11972), .ZN(n8971) );
  AND2_X1 U9879 ( .A1(n14826), .A2(n14824), .ZN(n12162) );
  NAND2_X1 U9880 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  OR2_X1 U9881 ( .A1(n8653), .A2(n8652), .ZN(n8669) );
  INV_X1 U9882 ( .A(n8779), .ZN(n8803) );
  NOR2_X1 U9883 ( .A1(n8669), .A2(n8668), .ZN(n8683) );
  NAND2_X1 U9884 ( .A1(n6654), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8440) );
  INV_X1 U9885 ( .A(n14632), .ZN(n14446) );
  OR2_X1 U9886 ( .A1(n8592), .A2(n10574), .ZN(n8616) );
  AND2_X1 U9887 ( .A1(n8536), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8566) );
  INV_X1 U9888 ( .A(n14502), .ZN(n8855) );
  NOR2_X1 U9889 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n8885) );
  NAND2_X1 U9890 ( .A1(n8337), .A2(n9870), .ZN(n8340) );
  INV_X1 U9891 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U9892 ( .A1(n8072), .A2(n8071), .ZN(n8088) );
  OAI21_X1 U9893 ( .B1(n12903), .B2(n10306), .A(n10305), .ZN(n10426) );
  AND2_X1 U9894 ( .A1(n8156), .A2(n8155), .ZN(n13042) );
  AND4_X2 U9895 ( .A1(n7715), .A2(n7714), .A3(n7713), .A4(n7712), .ZN(n7745)
         );
  OAI21_X1 U9896 ( .B1(n9739), .B2(n9738), .A(n12751), .ZN(n12607) );
  INV_X1 U9897 ( .A(n13295), .ZN(n13274) );
  INV_X1 U9898 ( .A(n13052), .ZN(n12940) );
  OR2_X1 U9899 ( .A1(n13173), .A2(n13172), .ZN(n13412) );
  AND2_X1 U9900 ( .A1(n8293), .A2(n12615), .ZN(n13310) );
  INV_X1 U9901 ( .A(n12885), .ZN(n15266) );
  INV_X1 U9902 ( .A(n10319), .ZN(n10243) );
  NAND2_X1 U9903 ( .A1(n11956), .A2(n11955), .ZN(n12598) );
  INV_X1 U9904 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U9905 ( .A1(n8040), .A2(n8039), .ZN(n8043) );
  OR2_X1 U9906 ( .A1(n9375), .A2(n13484), .ZN(n9394) );
  NAND2_X1 U9907 ( .A1(n9337), .A2(n9336), .ZN(n9359) );
  OR2_X1 U9908 ( .A1(n11686), .A2(n11685), .ZN(n11687) );
  NAND2_X1 U9909 ( .A1(n11999), .A2(n11998), .ZN(n12000) );
  AND2_X1 U9910 ( .A1(n10931), .A2(n10929), .ZN(n10999) );
  INV_X1 U9911 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n14995) );
  AND2_X1 U9912 ( .A1(n13592), .A2(n12009), .ZN(n11511) );
  AND2_X1 U9913 ( .A1(n9416), .A2(n9408), .ZN(n13708) );
  OR2_X1 U9914 ( .A1(n9310), .A2(n9309), .ZN(n9340) );
  OR2_X1 U9915 ( .A1(n9221), .A2(n9220), .ZN(n9243) );
  OR2_X1 U9916 ( .A1(n9952), .A2(n9951), .ZN(n10267) );
  INV_X1 U9917 ( .A(n13648), .ZN(n13644) );
  NAND2_X1 U9918 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  INV_X1 U9919 ( .A(n9688), .ZN(n11816) );
  INV_X1 U9920 ( .A(n10988), .ZN(n11165) );
  INV_X1 U9921 ( .A(n9626), .ZN(n13719) );
  AND2_X1 U9922 ( .A1(n9635), .A2(n9634), .ZN(n11793) );
  OR2_X1 U9923 ( .A1(n9659), .A2(n9704), .ZN(n15200) );
  OR2_X1 U9924 ( .A1(n9175), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n9192) );
  NOR2_X1 U9925 ( .A1(n8616), .A2(n8615), .ZN(n8631) );
  AND2_X1 U9926 ( .A1(n13983), .A2(n12223), .ZN(n14083) );
  AND2_X1 U9927 ( .A1(n8744), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8753) );
  AND2_X1 U9928 ( .A1(n8683), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8698) );
  INV_X1 U9929 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11887) );
  INV_X1 U9930 ( .A(n12533), .ZN(n11834) );
  INV_X1 U9931 ( .A(n14065), .ZN(n14111) );
  NAND2_X1 U9932 ( .A1(n14923), .A2(n14301), .ZN(n14477) );
  OR2_X1 U9933 ( .A1(n14987), .A2(n9762), .ZN(n9763) );
  OR3_X1 U9934 ( .A1(n14600), .A2(n14599), .A3(n14598), .ZN(n14645) );
  INV_X1 U9935 ( .A(n12526), .ZN(n11310) );
  AND2_X1 U9936 ( .A1(n12296), .A2(n12482), .ZN(n14921) );
  NAND2_X1 U9937 ( .A1(n9500), .A2(n9460), .ZN(n9463) );
  NOR2_X1 U9938 ( .A1(n8879), .A2(n8885), .ZN(n8886) );
  AND2_X1 U9939 ( .A1(n8604), .A2(n8343), .ZN(n8587) );
  AND2_X1 U9940 ( .A1(n8511), .A2(n8325), .ZN(n8499) );
  NAND2_X1 U9941 ( .A1(n10241), .A2(n10240), .ZN(n13038) );
  INV_X1 U9942 ( .A(n13042), .ZN(n13250) );
  AND4_X1 U9943 ( .A1(n8078), .A2(n8077), .A3(n8076), .A4(n8075), .ZN(n13313)
         );
  INV_X1 U9944 ( .A(n11749), .ZN(n13015) );
  INV_X1 U9945 ( .A(n13314), .ZN(n15244) );
  INV_X1 U9946 ( .A(n13310), .ZN(n15248) );
  INV_X1 U9947 ( .A(n13305), .ZN(n13347) );
  NAND2_X1 U9948 ( .A1(n10671), .A2(n10670), .ZN(n15238) );
  AND2_X1 U9949 ( .A1(n9773), .A2(n9772), .ZN(n10669) );
  AND2_X1 U9950 ( .A1(n13389), .A2(n13388), .ZN(n13438) );
  OR2_X1 U9951 ( .A1(n13204), .A2(n15303), .ZN(n15298) );
  AND2_X1 U9952 ( .A1(n15240), .A2(n12617), .ZN(n15303) );
  INV_X1 U9953 ( .A(n12617), .ZN(n12809) );
  INV_X1 U9954 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8218) );
  INV_X1 U9955 ( .A(n13504), .ZN(n13500) );
  NOR2_X1 U9956 ( .A1(n12116), .A2(n11003), .ZN(n11004) );
  NAND2_X1 U9957 ( .A1(n9074), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9090) );
  AND2_X1 U9958 ( .A1(n9811), .A2(n15166), .ZN(n9819) );
  AND2_X1 U9959 ( .A1(n9299), .A2(n9298), .ZN(n13488) );
  OR2_X1 U9960 ( .A1(n10269), .A2(n10268), .ZN(n10373) );
  INV_X1 U9961 ( .A(n15105), .ZN(n15091) );
  AND2_X1 U9962 ( .A1(n15201), .A2(n15200), .ZN(n15187) );
  INV_X1 U9963 ( .A(n10075), .ZN(n10661) );
  AND2_X1 U9964 ( .A1(n9653), .A2(n9652), .ZN(n15158) );
  NOR2_X1 U9965 ( .A1(n10705), .A2(n7650), .ZN(n10721) );
  INV_X1 U9966 ( .A(n14103), .ZN(n14828) );
  INV_X1 U9967 ( .A(n9755), .ZN(n12481) );
  AND3_X1 U9968 ( .A1(n8702), .A2(n8701), .A3(n8700), .ZN(n14047) );
  INV_X1 U9969 ( .A(n6653), .ZN(n14923) );
  AND2_X1 U9970 ( .A1(n14929), .A2(n11312), .ZN(n14843) );
  INV_X1 U9971 ( .A(n14925), .ZN(n14900) );
  INV_X1 U9972 ( .A(n14477), .ZN(n14911) );
  AND2_X1 U9973 ( .A1(n11305), .A2(n8919), .ZN(n9764) );
  AND2_X1 U9974 ( .A1(n8895), .A2(n8920), .ZN(n10252) );
  NAND2_X1 U9975 ( .A1(n14697), .A2(n14696), .ZN(n14701) );
  INV_X1 U9976 ( .A(n14716), .ZN(n14717) );
  AND2_X1 U9977 ( .A1(n10153), .A2(n10152), .ZN(n15234) );
  INV_X1 U9978 ( .A(n13038), .ZN(n13031) );
  NAND2_X1 U9979 ( .A1(n10230), .A2(n10671), .ZN(n13046) );
  INV_X1 U9980 ( .A(n13313), .ZN(n13050) );
  INV_X1 U9981 ( .A(n13012), .ZN(n13056) );
  OR2_X1 U9982 ( .A1(n10140), .A2(n12807), .ZN(n13165) );
  OR2_X1 U9983 ( .A1(n10140), .A2(n10139), .ZN(n13150) );
  INV_X1 U9984 ( .A(n13344), .ZN(n13328) );
  INV_X1 U9985 ( .A(n13344), .ZN(n15258) );
  INV_X1 U9986 ( .A(n15699), .ZN(n15696) );
  AND2_X1 U9987 ( .A1(n8297), .A2(n8296), .ZN(n15307) );
  OR2_X1 U9988 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  INV_X1 U9989 ( .A(SI_12_), .ZN(n9881) );
  INV_X1 U9990 ( .A(n11568), .ZN(n11572) );
  OR2_X1 U9991 ( .A1(n14999), .A2(n15134), .ZN(n13561) );
  NAND2_X1 U9992 ( .A1(n9792), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15007) );
  INV_X1 U9993 ( .A(n12038), .ZN(n13578) );
  NAND2_X1 U9994 ( .A1(n9400), .A2(n9399), .ZN(n13583) );
  OR2_X1 U9995 ( .A1(n9212), .A2(n9211), .ZN(n13594) );
  INV_X1 U9996 ( .A(n15085), .ZN(n15103) );
  INV_X1 U9997 ( .A(n15089), .ZN(n15107) );
  OR2_X1 U9998 ( .A1(n9894), .A2(P2_U3088), .ZN(n15111) );
  NAND2_X1 U9999 ( .A1(n15155), .A2(n9706), .ZN(n15139) );
  INV_X1 U10000 ( .A(n15233), .ZN(n15231) );
  INV_X1 U10001 ( .A(n15159), .ZN(n15160) );
  INV_X1 U10002 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10326) );
  INV_X1 U10003 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U10004 ( .A1(n10355), .A2(n10354), .ZN(n14103) );
  NAND2_X1 U10005 ( .A1(n10715), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14836) );
  INV_X1 U10006 ( .A(n13968), .ZN(n14131) );
  NAND2_X1 U10007 ( .A1(n14923), .A2(n11307), .ZN(n14925) );
  INV_X1 U10008 ( .A(n14843), .ZN(n14518) );
  NAND2_X1 U10009 ( .A1(n14320), .A2(n14507), .ZN(n14929) );
  NAND2_X1 U10010 ( .A1(n14994), .A2(n14974), .ZN(n14596) );
  AND2_X2 U10011 ( .A1(n9764), .A2(n11303), .ZN(n14994) );
  NAND2_X1 U10012 ( .A1(n14987), .A2(n14974), .ZN(n14643) );
  INV_X1 U10013 ( .A(n14987), .ZN(n14985) );
  CLKBUF_X1 U10014 ( .A(n14943), .Z(n14959) );
  INV_X1 U10015 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10328) );
  INV_X1 U10016 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10054) );
  OAI21_X1 U10017 ( .B1(n9784), .B2(n15307), .A(n9746), .ZN(P3_U3456) );
  INV_X1 U10018 ( .A(n14159), .ZN(P1_U4016) );
  NOR2_X1 U10019 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n7666) );
  NAND4_X1 U10020 ( .A1(n7666), .A2(n7665), .A3(n8290), .A4(n7664), .ZN(n7667)
         );
  NOR2_X1 U10021 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), 
        .ZN(n7672) );
  NOR2_X1 U10022 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), 
        .ZN(n7671) );
  NOR2_X1 U10023 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), 
        .ZN(n7670) );
  INV_X1 U10024 ( .A(n8003), .ZN(n7674) );
  INV_X1 U10025 ( .A(n7680), .ZN(n7678) );
  NAND2_X1 U10026 ( .A1(n7678), .A2(n7681), .ZN(n13463) );
  XNOR2_X2 U10027 ( .A(n7679), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U10028 ( .A1(n7680), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7682) );
  INV_X1 U10029 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7683) );
  OR2_X1 U10030 ( .A1(n7754), .A2(n7683), .ZN(n7690) );
  NAND2_X1 U10031 ( .A1(n7750), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7689) );
  INV_X1 U10032 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n7684) );
  OR2_X1 U10033 ( .A1(n7749), .A2(n7684), .ZN(n7688) );
  INV_X1 U10034 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10673) );
  AND4_X2 U10035 ( .A1(n7690), .A2(n7689), .A3(n7688), .A4(n7687), .ZN(n10364)
         );
  NAND2_X1 U10036 ( .A1(n8268), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7693) );
  NAND2_X2 U10037 ( .A1(n12806), .A2(n6647), .ZN(n7723) );
  XNOR2_X1 U10038 ( .A(n7717), .B(n7716), .ZN(n9830) );
  INV_X1 U10039 ( .A(SI_1_), .ZN(n7697) );
  OR2_X1 U10040 ( .A1(n7723), .A2(n7699), .ZN(n7700) );
  INV_X1 U10041 ( .A(n10307), .ZN(n7709) );
  NAND2_X1 U10042 ( .A1(n10364), .A2(n10307), .ZN(n12624) );
  INV_X1 U10043 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n7702) );
  INV_X1 U10044 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10908) );
  INV_X1 U10045 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n15623) );
  INV_X1 U10046 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n7703) );
  INV_X1 U10047 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n7706) );
  NAND2_X1 U10048 ( .A1(n7706), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U10049 ( .A1(n7716), .A2(n7707), .ZN(n7708) );
  MUX2_X1 U10050 ( .A(n7708), .B(SI_0_), .S(n9829), .Z(n13468) );
  NAND2_X1 U10051 ( .A1(n10312), .A2(n10674), .ZN(n7710) );
  NAND2_X1 U10052 ( .A1(n10364), .A2(n7709), .ZN(n10304) );
  NAND2_X1 U10053 ( .A1(n7710), .A2(n10304), .ZN(n15247) );
  INV_X1 U10054 ( .A(n8112), .ZN(n8131) );
  NAND2_X1 U10055 ( .A1(n7750), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7715) );
  INV_X1 U10056 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n7711) );
  OR2_X1 U10057 ( .A1(n7754), .A2(n7711), .ZN(n7714) );
  INV_X1 U10058 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15239) );
  OR2_X1 U10059 ( .A1(n6732), .A2(n15239), .ZN(n7713) );
  INV_X1 U10060 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10133) );
  OR2_X1 U10061 ( .A1(n7749), .A2(n10133), .ZN(n7712) );
  INV_X1 U10062 ( .A(n7716), .ZN(n7718) );
  NAND2_X1 U10063 ( .A1(n7718), .A2(n7717), .ZN(n7720) );
  NAND2_X1 U10064 ( .A1(n9873), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7719) );
  XNOR2_X1 U10065 ( .A(n9872), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n7721) );
  INV_X1 U10066 ( .A(SI_2_), .ZN(n7722) );
  NOR2_X2 U10067 ( .A1(n7727), .A2(n7726), .ZN(n10130) );
  INV_X1 U10068 ( .A(n10130), .ZN(n7728) );
  NAND2_X1 U10069 ( .A1(n7745), .A2(n7729), .ZN(n12629) );
  NAND2_X1 U10070 ( .A1(n15247), .A2(n15246), .ZN(n15245) );
  INV_X1 U10071 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10120) );
  OR2_X1 U10072 ( .A1(n6732), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n7733) );
  INV_X1 U10073 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10119) );
  OR2_X1 U10074 ( .A1(n7749), .A2(n10119), .ZN(n7732) );
  INV_X1 U10075 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n7730) );
  INV_X1 U10076 ( .A(n15243), .ZN(n10848) );
  INV_X1 U10077 ( .A(SI_3_), .ZN(n9833) );
  NAND2_X1 U10078 ( .A1(n7836), .A2(n9833), .ZN(n7744) );
  NAND2_X1 U10079 ( .A1(n9824), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U10080 ( .A1(n9872), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7737) );
  XNOR2_X1 U10081 ( .A(n9826), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n7738) );
  XNOR2_X1 U10082 ( .A(n7759), .B(n7738), .ZN(n9834) );
  INV_X1 U10083 ( .A(n9834), .ZN(n7739) );
  OR2_X1 U10084 ( .A1(n7726), .A2(n13462), .ZN(n7741) );
  NAND2_X1 U10085 ( .A1(n7745), .A2(n7746), .ZN(n10807) );
  NAND2_X1 U10086 ( .A1(n15243), .A2(n12885), .ZN(n7748) );
  NAND2_X1 U10087 ( .A1(n10808), .A2(n7748), .ZN(n10847) );
  NAND2_X1 U10088 ( .A1(n8205), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7758) );
  INV_X1 U10089 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10172) );
  OR2_X1 U10090 ( .A1(n8112), .A2(n10172), .ZN(n7757) );
  INV_X1 U10091 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n7751) );
  NAND2_X1 U10092 ( .A1(n12886), .A2(n7751), .ZN(n7770) );
  NAND2_X1 U10093 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7752) );
  AND2_X1 U10094 ( .A1(n7770), .A2(n7752), .ZN(n10845) );
  OR2_X1 U10095 ( .A1(n6732), .A2(n10845), .ZN(n7756) );
  INV_X1 U10096 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n7753) );
  OR2_X1 U10097 ( .A1(n7754), .A2(n7753), .ZN(n7755) );
  NAND2_X1 U10098 ( .A1(n9862), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7760) );
  XNOR2_X1 U10099 ( .A(n7777), .B(n7776), .ZN(n9844) );
  NAND2_X1 U10100 ( .A1(n12601), .A2(n9844), .ZN(n7764) );
  NAND2_X1 U10101 ( .A1(n8052), .A2(n10213), .ZN(n7763) );
  OAI211_X1 U10102 ( .C1(n7910), .C2(SI_4_), .A(n7764), .B(n7763), .ZN(n15270)
         );
  NAND2_X1 U10103 ( .A1(n10847), .A2(n10846), .ZN(n7766) );
  INV_X1 U10104 ( .A(n15270), .ZN(n10697) );
  NAND2_X1 U10105 ( .A1(n12956), .A2(n10697), .ZN(n7765) );
  NAND2_X1 U10106 ( .A1(n7766), .A2(n7765), .ZN(n10914) );
  INV_X1 U10107 ( .A(n10914), .ZN(n7788) );
  NAND2_X1 U10108 ( .A1(n9727), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7775) );
  INV_X1 U10109 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10923) );
  OR2_X1 U10110 ( .A1(n8112), .A2(n10923), .ZN(n7774) );
  INV_X1 U10111 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15697) );
  OR2_X1 U10112 ( .A1(n7767), .A2(n15697), .ZN(n7773) );
  INV_X1 U10113 ( .A(n7770), .ZN(n7769) );
  NAND2_X1 U10114 ( .A1(n7770), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n7771) );
  AND2_X1 U10115 ( .A1(n7789), .A2(n7771), .ZN(n10924) );
  OR2_X1 U10116 ( .A1(n6732), .A2(n10924), .ZN(n7772) );
  NAND2_X1 U10117 ( .A1(n9857), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7778) );
  XNOR2_X1 U10118 ( .A(n7797), .B(n7796), .ZN(n9855) );
  NAND2_X1 U10119 ( .A1(n7836), .A2(SI_5_), .ZN(n7786) );
  NAND2_X1 U10120 ( .A1(n7761), .A2(n7780), .ZN(n7781) );
  INV_X1 U10121 ( .A(n7802), .ZN(n7784) );
  NAND2_X1 U10122 ( .A1(n7781), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7782) );
  MUX2_X1 U10123 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7782), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n7783) );
  NAND2_X1 U10124 ( .A1(n8052), .A2(n10224), .ZN(n7785) );
  OAI211_X1 U10125 ( .C1(n8199), .C2(n9855), .A(n7786), .B(n7785), .ZN(n15274)
         );
  NAND2_X1 U10126 ( .A1(n11117), .A2(n15274), .ZN(n12642) );
  INV_X1 U10127 ( .A(n11117), .ZN(n13059) );
  INV_X1 U10128 ( .A(n15274), .ZN(n11115) );
  NAND2_X1 U10129 ( .A1(n13059), .A2(n11115), .ZN(n12646) );
  NAND2_X1 U10130 ( .A1(n8131), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7795) );
  INV_X1 U10131 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10433) );
  OR2_X1 U10132 ( .A1(n7767), .A2(n10433), .ZN(n7794) );
  NAND2_X1 U10133 ( .A1(n7789), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7790) );
  AND2_X1 U10134 ( .A1(n7809), .A2(n7790), .ZN(n10746) );
  OR2_X1 U10135 ( .A1(n6732), .A2(n10746), .ZN(n7793) );
  INV_X1 U10136 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n7791) );
  OR2_X1 U10137 ( .A1(n7754), .A2(n7791), .ZN(n7792) );
  NAND2_X1 U10138 ( .A1(n9841), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U10139 ( .A1(n6884), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7800) );
  XNOR2_X1 U10140 ( .A(n7817), .B(n7815), .ZN(n9836) );
  NAND2_X1 U10141 ( .A1(n7836), .A2(SI_6_), .ZN(n7805) );
  OR2_X1 U10142 ( .A1(n7802), .A2(n13462), .ZN(n7801) );
  MUX2_X1 U10143 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7801), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n7803) );
  NAND2_X1 U10144 ( .A1(n7802), .A2(n15674), .ZN(n7819) );
  NAND2_X1 U10145 ( .A1(n8052), .A2(n10445), .ZN(n7804) );
  OAI211_X1 U10146 ( .C1(n8199), .C2(n9836), .A(n7805), .B(n7804), .ZN(n11126)
         );
  NAND2_X1 U10147 ( .A1(n10918), .A2(n11126), .ZN(n12651) );
  INV_X1 U10148 ( .A(n11126), .ZN(n15279) );
  NAND2_X1 U10149 ( .A1(n13058), .A2(n15279), .ZN(n12648) );
  NAND2_X1 U10150 ( .A1(n12651), .A2(n12648), .ZN(n12766) );
  NAND2_X1 U10151 ( .A1(n11117), .A2(n11115), .ZN(n10738) );
  AND2_X1 U10152 ( .A1(n12766), .A2(n10738), .ZN(n7806) );
  NAND2_X1 U10153 ( .A1(n10737), .A2(n7806), .ZN(n10739) );
  NAND2_X1 U10154 ( .A1(n13058), .A2(n11126), .ZN(n7807) );
  NAND2_X1 U10155 ( .A1(n10739), .A2(n7807), .ZN(n10777) );
  NAND2_X1 U10156 ( .A1(n9727), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7814) );
  INV_X1 U10157 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10464) );
  OR2_X1 U10158 ( .A1(n8112), .A2(n10464), .ZN(n7813) );
  INV_X1 U10159 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10463) );
  OR2_X1 U10160 ( .A1(n7767), .A2(n10463), .ZN(n7812) );
  NAND2_X1 U10161 ( .A1(n7809), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7810) );
  AND2_X1 U10162 ( .A1(n7826), .A2(n7810), .ZN(n10782) );
  OR2_X1 U10163 ( .A1(n6732), .A2(n10782), .ZN(n7811) );
  NAND4_X1 U10164 ( .A1(n7814), .A2(n7813), .A3(n7812), .A4(n7811), .ZN(n12652) );
  NAND2_X1 U10165 ( .A1(n7836), .A2(SI_7_), .ZN(n7823) );
  XNOR2_X1 U10166 ( .A(n7834), .B(n7832), .ZN(n9837) );
  NAND2_X1 U10167 ( .A1(n12601), .A2(n9837), .ZN(n7822) );
  NAND2_X1 U10168 ( .A1(n7819), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7820) );
  NAND2_X1 U10169 ( .A1(n8052), .A2(n10478), .ZN(n7821) );
  XNOR2_X1 U10170 ( .A(n12652), .B(n15283), .ZN(n12777) );
  NAND2_X1 U10171 ( .A1(n10777), .A2(n12777), .ZN(n7825) );
  INV_X1 U10172 ( .A(n15283), .ZN(n12818) );
  NAND2_X1 U10173 ( .A1(n12652), .A2(n12818), .ZN(n7824) );
  INV_X1 U10174 ( .A(n11251), .ZN(n7844) );
  NAND2_X1 U10175 ( .A1(n9727), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7831) );
  INV_X1 U10176 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15639) );
  OR2_X1 U10177 ( .A1(n7767), .A2(n15639), .ZN(n7830) );
  NAND2_X1 U10178 ( .A1(n7826), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7827) );
  AND2_X1 U10179 ( .A1(n7847), .A2(n7827), .ZN(n11250) );
  OR2_X1 U10180 ( .A1(n6732), .A2(n11250), .ZN(n7829) );
  INV_X1 U10181 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10468) );
  OR2_X1 U10182 ( .A1(n8112), .A2(n10468), .ZN(n7828) );
  INV_X1 U10183 ( .A(n7832), .ZN(n7833) );
  XNOR2_X1 U10184 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7835) );
  XNOR2_X1 U10185 ( .A(n7854), .B(n7835), .ZN(n9846) );
  NAND2_X1 U10186 ( .A1(n12601), .A2(n9846), .ZN(n7842) );
  INV_X1 U10187 ( .A(SI_8_), .ZN(n9847) );
  NAND2_X1 U10188 ( .A1(n7836), .A2(n9847), .ZN(n7841) );
  NOR2_X1 U10189 ( .A1(n8045), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7859) );
  INV_X1 U10190 ( .A(n7859), .ZN(n7839) );
  NAND2_X1 U10191 ( .A1(n8045), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7837) );
  MUX2_X1 U10192 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7837), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n7838) );
  NAND2_X1 U10193 ( .A1(n8052), .A2(n10963), .ZN(n7840) );
  NAND2_X1 U10194 ( .A1(n11072), .A2(n11241), .ZN(n12658) );
  NAND2_X1 U10195 ( .A1(n13057), .A2(n15289), .ZN(n12659) );
  NAND2_X1 U10196 ( .A1(n11072), .A2(n15289), .ZN(n7845) );
  NAND2_X1 U10197 ( .A1(n9727), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7852) );
  INV_X1 U10198 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10953) );
  OR2_X1 U10199 ( .A1(n8112), .A2(n10953), .ZN(n7851) );
  INV_X1 U10200 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10952) );
  OR2_X1 U10201 ( .A1(n7767), .A2(n10952), .ZN(n7850) );
  NAND2_X1 U10202 ( .A1(n7847), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n7848) );
  AND2_X1 U10203 ( .A1(n7865), .A2(n7848), .ZN(n12989) );
  OR2_X1 U10204 ( .A1(n6732), .A2(n12989), .ZN(n7849) );
  NAND2_X1 U10205 ( .A1(n9865), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7855) );
  XNOR2_X1 U10206 ( .A(n9876), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n7856) );
  XNOR2_X1 U10207 ( .A(n7871), .B(n7856), .ZN(n9832) );
  NAND2_X1 U10208 ( .A1(n12601), .A2(n9832), .ZN(n7863) );
  INV_X1 U10209 ( .A(SI_9_), .ZN(n9831) );
  NAND2_X1 U10210 ( .A1(n12602), .A2(n9831), .ZN(n7862) );
  OR2_X1 U10211 ( .A1(n7859), .A2(n13462), .ZN(n7857) );
  MUX2_X1 U10212 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7857), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n7860) );
  INV_X1 U10213 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10214 ( .A1(n7859), .A2(n7858), .ZN(n7985) );
  NAND2_X1 U10215 ( .A1(n7860), .A2(n7985), .ZN(n10964) );
  NAND2_X1 U10216 ( .A1(n8052), .A2(n10964), .ZN(n7861) );
  NAND2_X1 U10217 ( .A1(n11740), .A2(n12988), .ZN(n12662) );
  INV_X1 U10218 ( .A(n12988), .ZN(n15296) );
  NAND2_X1 U10219 ( .A1(n12874), .A2(n15296), .ZN(n12663) );
  NAND2_X1 U10220 ( .A1(n12874), .A2(n12988), .ZN(n7864) );
  NAND2_X1 U10221 ( .A1(n9727), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7870) );
  INV_X1 U10222 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11223) );
  OR2_X1 U10223 ( .A1(n7767), .A2(n11223), .ZN(n7869) );
  INV_X1 U10224 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11224) );
  OR2_X1 U10225 ( .A1(n8112), .A2(n11224), .ZN(n7868) );
  OR2_X2 U10226 ( .A1(n7865), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10227 ( .A1(n7865), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7866) );
  AND2_X1 U10228 ( .A1(n7897), .A2(n7866), .ZN(n11158) );
  OR2_X1 U10229 ( .A1(n6732), .A2(n11158), .ZN(n7867) );
  NAND2_X1 U10230 ( .A1(n9876), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7872) );
  XNOR2_X1 U10231 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7885) );
  XNOR2_X1 U10232 ( .A(n7886), .B(n7885), .ZN(n9853) );
  NAND2_X1 U10233 ( .A1(n12602), .A2(SI_10_), .ZN(n7876) );
  NAND2_X1 U10234 ( .A1(n7985), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7874) );
  INV_X1 U10235 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7873) );
  XNOR2_X1 U10236 ( .A(n7874), .B(n7873), .ZN(n11464) );
  INV_X1 U10237 ( .A(n11464), .ZN(n11225) );
  NAND2_X1 U10238 ( .A1(n8052), .A2(n11225), .ZN(n7875) );
  OAI211_X1 U10239 ( .C1(n8199), .C2(n9853), .A(n7876), .B(n7875), .ZN(n15301)
         );
  NAND2_X1 U10240 ( .A1(n11744), .A2(n15301), .ZN(n12668) );
  INV_X1 U10241 ( .A(n15301), .ZN(n11743) );
  NAND2_X1 U10242 ( .A1(n13016), .A2(n11743), .ZN(n12667) );
  NAND2_X1 U10243 ( .A1(n12668), .A2(n12667), .ZN(n12776) );
  NAND2_X1 U10244 ( .A1(n11153), .A2(n12776), .ZN(n7878) );
  NAND2_X1 U10245 ( .A1(n13016), .A2(n15301), .ZN(n7877) );
  NAND2_X1 U10246 ( .A1(n7878), .A2(n7877), .ZN(n11188) );
  NAND2_X1 U10247 ( .A1(n9727), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7883) );
  INV_X1 U10248 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11196) );
  OR2_X1 U10249 ( .A1(n8112), .A2(n11196), .ZN(n7882) );
  INV_X1 U10250 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n7879) );
  OR2_X1 U10251 ( .A1(n7767), .A2(n7879), .ZN(n7881) );
  XNOR2_X1 U10252 ( .A(n7897), .B(n11455), .ZN(n11194) );
  OR2_X1 U10253 ( .A1(n6732), .A2(n11194), .ZN(n7880) );
  NAND2_X1 U10254 ( .A1(n7911), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7884) );
  XNOR2_X1 U10255 ( .A(n7884), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11568) );
  INV_X1 U10256 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U10257 ( .A1(n9887), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7887) );
  XNOR2_X1 U10258 ( .A(n9917), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n7889) );
  XNOR2_X1 U10259 ( .A(n7904), .B(n7889), .ZN(n9868) );
  NAND2_X1 U10260 ( .A1(n9868), .A2(n12601), .ZN(n7891) );
  NAND2_X1 U10261 ( .A1(n12602), .A2(SI_11_), .ZN(n7890) );
  OAI211_X1 U10262 ( .C1(n10126), .C2(n11572), .A(n7891), .B(n7890), .ZN(
        n14799) );
  NAND2_X1 U10263 ( .A1(n13012), .A2(n14799), .ZN(n12672) );
  INV_X1 U10264 ( .A(n14799), .ZN(n7892) );
  NAND2_X1 U10265 ( .A1(n13056), .A2(n7892), .ZN(n12675) );
  NAND2_X1 U10266 ( .A1(n12672), .A2(n12675), .ZN(n12669) );
  NAND2_X1 U10267 ( .A1(n11188), .A2(n12669), .ZN(n7894) );
  NAND2_X1 U10268 ( .A1(n13056), .A2(n14799), .ZN(n7893) );
  NAND2_X1 U10269 ( .A1(n7894), .A2(n7893), .ZN(n11316) );
  NAND2_X1 U10270 ( .A1(n9727), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7902) );
  INV_X1 U10271 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n7895) );
  OR2_X1 U10272 ( .A1(n7767), .A2(n7895), .ZN(n7901) );
  INV_X1 U10273 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11579) );
  NAND2_X1 U10274 ( .A1(n11455), .A2(n11579), .ZN(n7896) );
  OAI21_X1 U10275 ( .B1(n7897), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n7898) );
  AND2_X1 U10276 ( .A1(n7932), .A2(n7898), .ZN(n11321) );
  OR2_X1 U10277 ( .A1(n6732), .A2(n11321), .ZN(n7900) );
  INV_X1 U10278 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11323) );
  OR2_X1 U10279 ( .A1(n8112), .A2(n11323), .ZN(n7899) );
  AND2_X1 U10280 ( .A1(n9915), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U10281 ( .A1(n9917), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U10282 ( .A1(n10054), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10283 ( .A1(n10056), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U10284 ( .A1(n7921), .A2(n7906), .ZN(n7907) );
  NAND2_X1 U10285 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  AND2_X1 U10286 ( .A1(n7922), .A2(n7909), .ZN(n9879) );
  NAND2_X1 U10287 ( .A1(n9879), .A2(n12601), .ZN(n7917) );
  INV_X1 U10288 ( .A(n7944), .ZN(n7915) );
  NAND2_X1 U10289 ( .A1(n7912), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7913) );
  MUX2_X1 U10290 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7913), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7914) );
  NAND2_X1 U10291 ( .A1(n7915), .A2(n7914), .ZN(n12073) );
  INV_X1 U10292 ( .A(n12073), .ZN(n12090) );
  AOI22_X1 U10293 ( .A1(n12602), .A2(SI_12_), .B1(n8052), .B2(n12090), .ZN(
        n7916) );
  NAND2_X1 U10294 ( .A1(n7917), .A2(n7916), .ZN(n14794) );
  NAND2_X1 U10295 ( .A1(n11749), .A2(n14794), .ZN(n12679) );
  INV_X1 U10296 ( .A(n14794), .ZN(n7918) );
  NAND2_X1 U10297 ( .A1(n7918), .A2(n13015), .ZN(n12677) );
  NAND2_X1 U10298 ( .A1(n12679), .A2(n12677), .ZN(n8238) );
  NAND2_X1 U10299 ( .A1(n14794), .A2(n13015), .ZN(n7919) );
  INV_X1 U10300 ( .A(n7923), .ZN(n7924) );
  NAND2_X1 U10301 ( .A1(n7924), .A2(n10081), .ZN(n7925) );
  NAND2_X1 U10302 ( .A1(n7941), .A2(n7925), .ZN(n9912) );
  NAND2_X1 U10303 ( .A1(n9912), .A2(n12601), .ZN(n7928) );
  INV_X1 U10304 ( .A(SI_13_), .ZN(n9913) );
  OR2_X1 U10305 ( .A1(n7944), .A2(n13462), .ZN(n7926) );
  XNOR2_X1 U10306 ( .A(n7926), .B(P3_IR_REG_13__SCAN_IN), .ZN(n13072) );
  INV_X1 U10307 ( .A(n13072), .ZN(n12092) );
  AOI22_X1 U10308 ( .A1(n12602), .A2(n9913), .B1(n8052), .B2(n12092), .ZN(
        n7927) );
  NAND2_X1 U10309 ( .A1(n9727), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7937) );
  INV_X1 U10310 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n7929) );
  OR2_X1 U10311 ( .A1(n8112), .A2(n7929), .ZN(n7936) );
  OR2_X1 U10312 ( .A1(n7767), .A2(n15669), .ZN(n7935) );
  INV_X1 U10313 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10314 ( .A1(n7932), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7933) );
  AND2_X1 U10315 ( .A1(n7950), .A2(n7933), .ZN(n11757) );
  OR2_X1 U10316 ( .A1(n6732), .A2(n11757), .ZN(n7934) );
  NAND4_X1 U10317 ( .A1(n7937), .A2(n7936), .A3(n7935), .A4(n7934), .ZN(n13055) );
  NAND2_X1 U10318 ( .A1(n14789), .A2(n13055), .ZN(n12680) );
  NAND2_X1 U10319 ( .A1(n10371), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U10320 ( .A1(n10369), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U10321 ( .A1(n7961), .A2(n7942), .ZN(n7959) );
  XNOR2_X1 U10322 ( .A(n7960), .B(n7959), .ZN(n10012) );
  NAND2_X1 U10323 ( .A1(n10012), .A2(n12601), .ZN(n7948) );
  INV_X1 U10324 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U10325 ( .A1(n7944), .A2(n7943), .ZN(n7963) );
  NAND2_X1 U10326 ( .A1(n7963), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7946) );
  INV_X1 U10327 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7945) );
  XNOR2_X1 U10328 ( .A(n7946), .B(n7945), .ZN(n12077) );
  INV_X1 U10329 ( .A(n12077), .ZN(n13083) );
  AOI22_X1 U10330 ( .A1(n12602), .A2(SI_14_), .B1(n8052), .B2(n13083), .ZN(
        n7947) );
  NAND2_X1 U10331 ( .A1(n7948), .A2(n7947), .ZN(n11858) );
  NAND2_X1 U10332 ( .A1(n8131), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7956) );
  INV_X1 U10333 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14788) );
  OR2_X1 U10334 ( .A1(n7767), .A2(n14788), .ZN(n7955) );
  NAND2_X1 U10335 ( .A1(n7950), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7951) );
  AND2_X1 U10336 ( .A1(n7967), .A2(n7951), .ZN(n11861) );
  OR2_X1 U10337 ( .A1(n6732), .A2(n11861), .ZN(n7954) );
  INV_X1 U10338 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n7952) );
  OR2_X1 U10339 ( .A1(n7754), .A2(n7952), .ZN(n7953) );
  OR2_X1 U10340 ( .A1(n11858), .A2(n11941), .ZN(n12687) );
  NAND2_X1 U10341 ( .A1(n11858), .A2(n11941), .ZN(n12686) );
  NAND2_X1 U10342 ( .A1(n12687), .A2(n12686), .ZN(n12785) );
  INV_X1 U10343 ( .A(n13055), .ZN(n11734) );
  NAND2_X1 U10344 ( .A1(n14789), .A2(n11734), .ZN(n11642) );
  AND2_X1 U10345 ( .A1(n12785), .A2(n11642), .ZN(n7957) );
  INV_X1 U10346 ( .A(n11941), .ZN(n13054) );
  NAND2_X1 U10347 ( .A1(n11858), .A2(n13054), .ZN(n7958) );
  NAND2_X2 U10348 ( .A1(n11640), .A2(n7958), .ZN(n11823) );
  INV_X1 U10349 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U10350 ( .A1(n10397), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7978) );
  INV_X1 U10351 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U10352 ( .A1(n10395), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7962) );
  NAND2_X1 U10353 ( .A1(n7978), .A2(n7962), .ZN(n7975) );
  XNOR2_X1 U10354 ( .A(n7977), .B(n7975), .ZN(n10057) );
  NAND2_X1 U10355 ( .A1(n10057), .A2(n12601), .ZN(n7966) );
  OAI21_X1 U10356 ( .B1(n7963), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7964) );
  XNOR2_X1 U10357 ( .A(n7964), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U10358 ( .A1(n12602), .A2(SI_15_), .B1(n8052), .B2(n13107), .ZN(
        n7965) );
  NAND2_X1 U10359 ( .A1(n9727), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7972) );
  INV_X1 U10360 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13110) );
  OR2_X1 U10361 ( .A1(n7767), .A2(n13110), .ZN(n7971) );
  INV_X1 U10362 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13099) );
  OR2_X1 U10363 ( .A1(n8112), .A2(n13099), .ZN(n7970) );
  NAND2_X1 U10364 ( .A1(n7967), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7968) );
  AND2_X1 U10365 ( .A1(n7992), .A2(n7968), .ZN(n11944) );
  OR2_X1 U10366 ( .A1(n6732), .A2(n11944), .ZN(n7969) );
  NAND4_X1 U10367 ( .A1(n7972), .A2(n7971), .A3(n7970), .A4(n7969), .ZN(n13053) );
  OR2_X1 U10368 ( .A1(n11946), .A2(n13053), .ZN(n7973) );
  NAND2_X1 U10369 ( .A1(n11946), .A2(n13053), .ZN(n7974) );
  INV_X1 U10370 ( .A(n7975), .ZN(n7976) );
  NAND2_X1 U10371 ( .A1(n10328), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10372 ( .A1(n10326), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7979) );
  AND2_X1 U10373 ( .A1(n8000), .A2(n7979), .ZN(n7980) );
  OR2_X1 U10374 ( .A1(n7981), .A2(n7980), .ZN(n7982) );
  NAND2_X1 U10375 ( .A1(n8001), .A2(n7982), .ZN(n10082) );
  INV_X1 U10376 ( .A(n7983), .ZN(n7984) );
  OAI21_X1 U10377 ( .B1(n7985), .B2(n7984), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7987) );
  INV_X1 U10378 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7986) );
  XNOR2_X1 U10379 ( .A(n7987), .B(n7986), .ZN(n12083) );
  INV_X1 U10380 ( .A(n12083), .ZN(n13122) );
  AOI22_X1 U10381 ( .A1(n12602), .A2(SI_16_), .B1(n8052), .B2(n13122), .ZN(
        n7988) );
  NAND2_X1 U10382 ( .A1(n9727), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7997) );
  INV_X1 U10383 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12100) );
  OR2_X1 U10384 ( .A1(n8112), .A2(n12100), .ZN(n7996) );
  INV_X1 U10385 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n15443) );
  OR2_X1 U10386 ( .A1(n7767), .A2(n15443), .ZN(n7995) );
  INV_X1 U10387 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U10388 ( .A1(n7992), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7993) );
  AND2_X1 U10389 ( .A1(n8010), .A2(n7993), .ZN(n12947) );
  OR2_X1 U10390 ( .A1(n6732), .A2(n12947), .ZN(n7994) );
  NAND4_X1 U10391 ( .A1(n7997), .A2(n7996), .A3(n7995), .A4(n7994), .ZN(n13052) );
  AND2_X1 U10392 ( .A1(n12949), .A2(n13052), .ZN(n7999) );
  NAND2_X1 U10393 ( .A1(n13457), .A2(n12940), .ZN(n7998) );
  NAND2_X1 U10394 ( .A1(n10399), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U10395 ( .A1(n10401), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U10396 ( .A1(n8020), .A2(n8002), .ZN(n8017) );
  XNOR2_X1 U10397 ( .A(n8019), .B(n8017), .ZN(n10293) );
  NAND2_X1 U10398 ( .A1(n10293), .A2(n12601), .ZN(n8009) );
  OR2_X1 U10399 ( .A1(n8045), .A2(n8003), .ZN(n8005) );
  NAND2_X1 U10400 ( .A1(n8005), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8004) );
  MUX2_X1 U10401 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8004), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8007) );
  NAND2_X1 U10402 ( .A1(n6642), .A2(n8006), .ZN(n8025) );
  NAND2_X1 U10403 ( .A1(n8007), .A2(n8025), .ZN(n12102) );
  INV_X1 U10404 ( .A(n12102), .ZN(n13148) );
  AOI22_X1 U10405 ( .A1(n12602), .A2(SI_17_), .B1(n8052), .B2(n13148), .ZN(
        n8008) );
  NAND2_X1 U10406 ( .A1(n9727), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8015) );
  INV_X1 U10407 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13137) );
  OR2_X1 U10408 ( .A1(n8112), .A2(n13137), .ZN(n8014) );
  INV_X1 U10409 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13404) );
  OR2_X1 U10410 ( .A1(n7767), .A2(n13404), .ZN(n8013) );
  NAND2_X1 U10411 ( .A1(n8010), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8011) );
  AND2_X1 U10412 ( .A1(n8031), .A2(n8011), .ZN(n12966) );
  OR2_X1 U10413 ( .A1(n6732), .A2(n12966), .ZN(n8012) );
  OR2_X1 U10414 ( .A1(n12968), .A2(n12944), .ZN(n12704) );
  NAND2_X1 U10415 ( .A1(n12968), .A2(n12944), .ZN(n12701) );
  NAND2_X1 U10416 ( .A1(n11924), .A2(n8016), .ZN(n13330) );
  INV_X1 U10417 ( .A(n8017), .ZN(n8018) );
  NAND2_X1 U10418 ( .A1(n10682), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U10419 ( .A1(n10681), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8021) );
  AND2_X1 U10420 ( .A1(n8039), .A2(n8021), .ZN(n8022) );
  OR2_X1 U10421 ( .A1(n8023), .A2(n8022), .ZN(n8024) );
  NAND2_X1 U10422 ( .A1(n8040), .A2(n8024), .ZN(n10329) );
  NAND2_X1 U10423 ( .A1(n8025), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8026) );
  XNOR2_X1 U10424 ( .A(n8026), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13167) );
  AOI22_X1 U10425 ( .A1(n12602), .A2(SI_18_), .B1(n8052), .B2(n13167), .ZN(
        n8027) );
  NAND2_X1 U10426 ( .A1(n8205), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8036) );
  INV_X1 U10427 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13343) );
  OR2_X1 U10428 ( .A1(n8112), .A2(n13343), .ZN(n8035) );
  INV_X1 U10429 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10430 ( .A1(n8031), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8032) );
  AND2_X1 U10431 ( .A1(n8055), .A2(n8032), .ZN(n13342) );
  OR2_X1 U10432 ( .A1(n6732), .A2(n13342), .ZN(n8034) );
  INV_X1 U10433 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13446) );
  OR2_X1 U10434 ( .A1(n7754), .A2(n13446), .ZN(n8033) );
  NAND2_X1 U10435 ( .A1(n13340), .A2(n13315), .ZN(n12708) );
  NAND2_X1 U10436 ( .A1(n12702), .A2(n12708), .ZN(n13339) );
  NAND2_X1 U10437 ( .A1(n12968), .A2(n13333), .ZN(n13329) );
  AND2_X1 U10438 ( .A1(n13339), .A2(n13329), .ZN(n8037) );
  INV_X1 U10439 ( .A(n13315), .ZN(n13051) );
  OR2_X1 U10440 ( .A1(n13340), .A2(n13051), .ZN(n8038) );
  INV_X1 U10441 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U10442 ( .A1(n10974), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8063) );
  INV_X1 U10443 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10977) );
  NAND2_X1 U10444 ( .A1(n10977), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8041) );
  AND2_X1 U10445 ( .A1(n8063), .A2(n8041), .ZN(n8042) );
  OR2_X1 U10446 ( .A1(n8043), .A2(n8042), .ZN(n8044) );
  NAND2_X1 U10447 ( .A1(n8064), .A2(n8044), .ZN(n10402) );
  NAND2_X1 U10448 ( .A1(n6642), .A2(n8046), .ZN(n8047) );
  NAND2_X1 U10449 ( .A1(n8047), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8048) );
  MUX2_X1 U10450 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8048), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8051) );
  NAND2_X1 U10451 ( .A1(n6642), .A2(n8049), .ZN(n8211) );
  NAND2_X1 U10452 ( .A1(n8051), .A2(n8211), .ZN(n12800) );
  AOI22_X1 U10453 ( .A1(n12602), .A2(SI_19_), .B1(n8052), .B2(n12613), .ZN(
        n8053) );
  NAND2_X1 U10454 ( .A1(n9727), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8060) );
  INV_X1 U10455 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13320) );
  OR2_X1 U10456 ( .A1(n8112), .A2(n13320), .ZN(n8059) );
  INV_X1 U10457 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13395) );
  OR2_X1 U10458 ( .A1(n7767), .A2(n13395), .ZN(n8058) );
  NAND2_X1 U10459 ( .A1(n8055), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8056) );
  AND2_X1 U10460 ( .A1(n8073), .A2(n8056), .ZN(n13319) );
  OR2_X1 U10461 ( .A1(n6732), .A2(n13319), .ZN(n8057) );
  NAND2_X1 U10462 ( .A1(n13323), .A2(n13027), .ZN(n12713) );
  NAND2_X1 U10463 ( .A1(n13323), .A2(n13334), .ZN(n8062) );
  INV_X1 U10464 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10904) );
  NAND2_X1 U10465 ( .A1(n10904), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8080) );
  INV_X1 U10466 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U10467 ( .A1(n10907), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8065) );
  AND2_X1 U10468 ( .A1(n8080), .A2(n8065), .ZN(n8066) );
  OR2_X1 U10469 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U10470 ( .A1(n8081), .A2(n8068), .ZN(n10563) );
  NAND2_X1 U10471 ( .A1(n12602), .A2(SI_20_), .ZN(n8069) );
  INV_X1 U10472 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10473 ( .A1(n8073), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10474 ( .A1(n8088), .A2(n8074), .ZN(n13298) );
  NAND2_X1 U10475 ( .A1(n8209), .A2(n13298), .ZN(n8078) );
  INV_X1 U10476 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13390) );
  OR2_X1 U10477 ( .A1(n7767), .A2(n13390), .ZN(n8077) );
  INV_X1 U10478 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13300) );
  OR2_X1 U10479 ( .A1(n8112), .A2(n13300), .ZN(n8076) );
  INV_X1 U10480 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13437) );
  OR2_X1 U10481 ( .A1(n7754), .A2(n13437), .ZN(n8075) );
  XNOR2_X1 U10482 ( .A(n13308), .B(n13313), .ZN(n13301) );
  NAND2_X1 U10483 ( .A1(n13294), .A2(n13301), .ZN(n13293) );
  NAND2_X1 U10484 ( .A1(n13308), .A2(n13050), .ZN(n8079) );
  NAND2_X1 U10485 ( .A1(n13293), .A2(n8079), .ZN(n13283) );
  INV_X1 U10486 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11040) );
  NAND2_X1 U10487 ( .A1(n11040), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8097) );
  INV_X1 U10488 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U10489 ( .A1(n11136), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8082) );
  AND2_X1 U10490 ( .A1(n8097), .A2(n8082), .ZN(n8083) );
  OR2_X1 U10491 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  NAND2_X1 U10492 ( .A1(n8098), .A2(n8085), .ZN(n10731) );
  NAND2_X1 U10493 ( .A1(n12602), .A2(SI_21_), .ZN(n8086) );
  NAND2_X1 U10494 ( .A1(n8088), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10495 ( .A1(n8107), .A2(n8089), .ZN(n13287) );
  NAND2_X1 U10496 ( .A1(n13287), .A2(n8209), .ZN(n8093) );
  NAND2_X1 U10497 ( .A1(n8131), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8092) );
  INV_X1 U10498 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13385) );
  OR2_X1 U10499 ( .A1(n7767), .A2(n13385), .ZN(n8091) );
  NAND2_X1 U10500 ( .A1(n9727), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8090) );
  NAND4_X1 U10501 ( .A1(n8093), .A2(n8092), .A3(n8091), .A4(n8090), .ZN(n13295) );
  OR2_X1 U10502 ( .A1(n13286), .A2(n13295), .ZN(n8094) );
  NAND2_X1 U10503 ( .A1(n13283), .A2(n8094), .ZN(n8096) );
  NAND2_X1 U10504 ( .A1(n13286), .A2(n13295), .ZN(n8095) );
  INV_X1 U10505 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U10506 ( .A1(n8379), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8113) );
  INV_X1 U10507 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11391) );
  NAND2_X1 U10508 ( .A1(n11391), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8099) );
  AND2_X1 U10509 ( .A1(n8113), .A2(n8099), .ZN(n8100) );
  OR2_X1 U10510 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  NAND2_X1 U10511 ( .A1(n8114), .A2(n8102), .ZN(n10763) );
  NAND2_X1 U10512 ( .A1(n12602), .A2(SI_22_), .ZN(n8103) );
  INV_X1 U10513 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8111) );
  INV_X1 U10514 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U10515 ( .A1(n8107), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U10516 ( .A1(n8117), .A2(n8108), .ZN(n13276) );
  NAND2_X1 U10517 ( .A1(n13276), .A2(n8209), .ZN(n8110) );
  AOI22_X1 U10518 ( .A1(n8205), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n9727), .B2(
        P3_REG0_REG_22__SCAN_IN), .ZN(n8109) );
  OAI211_X1 U10519 ( .C1(n8112), .C2(n8111), .A(n8110), .B(n8109), .ZN(n13049)
         );
  INV_X1 U10520 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8124) );
  XNOR2_X1 U10521 ( .A(n8124), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n8122) );
  XNOR2_X1 U10522 ( .A(n8123), .B(n8122), .ZN(n10996) );
  NAND2_X1 U10523 ( .A1(n10996), .A2(n12601), .ZN(n8116) );
  NAND2_X1 U10524 ( .A1(n12602), .A2(SI_23_), .ZN(n8115) );
  NAND2_X1 U10525 ( .A1(n8117), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U10526 ( .A1(n8129), .A2(n8118), .ZN(n13260) );
  NAND2_X1 U10527 ( .A1(n13260), .A2(n8209), .ZN(n8121) );
  AOI22_X1 U10528 ( .A1(n8205), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n8131), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U10529 ( .A1(n9727), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10530 ( .A1(n13375), .A2(n13273), .ZN(n12729) );
  NAND2_X1 U10531 ( .A1(n8125), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8126) );
  XNOR2_X1 U10532 ( .A(n8139), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11260) );
  NAND2_X1 U10533 ( .A1(n11260), .A2(n12601), .ZN(n8128) );
  NAND2_X1 U10534 ( .A1(n12602), .A2(SI_24_), .ZN(n8127) );
  NAND2_X1 U10535 ( .A1(n8129), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8130) );
  NAND2_X1 U10536 ( .A1(n8149), .A2(n8130), .ZN(n13242) );
  NAND2_X1 U10537 ( .A1(n13242), .A2(n8209), .ZN(n8137) );
  INV_X1 U10538 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U10539 ( .A1(n8131), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10540 ( .A1(n9727), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8132) );
  OAI211_X1 U10541 ( .C1(n7767), .C2(n8134), .A(n8133), .B(n8132), .ZN(n8135)
         );
  INV_X1 U10542 ( .A(n8135), .ZN(n8136) );
  XNOR2_X1 U10543 ( .A(n13372), .B(n13256), .ZN(n13247) );
  NAND2_X1 U10544 ( .A1(n13372), .A2(n13232), .ZN(n8138) );
  INV_X1 U10545 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11631) );
  INV_X1 U10546 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11721) );
  NAND2_X1 U10547 ( .A1(n11721), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8158) );
  INV_X1 U10548 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11724) );
  NAND2_X1 U10549 ( .A1(n11724), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8141) );
  AND2_X1 U10550 ( .A1(n8158), .A2(n8141), .ZN(n8142) );
  OR2_X1 U10551 ( .A1(n8143), .A2(n8142), .ZN(n8144) );
  NAND2_X1 U10552 ( .A1(n8159), .A2(n8144), .ZN(n11422) );
  NAND2_X1 U10553 ( .A1(n12602), .A2(SI_25_), .ZN(n8145) );
  INV_X1 U10554 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U10555 ( .A1(n8149), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U10556 ( .A1(n8163), .A2(n8150), .ZN(n13236) );
  NAND2_X1 U10557 ( .A1(n13236), .A2(n8209), .ZN(n8156) );
  INV_X1 U10558 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U10559 ( .A1(n9727), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U10560 ( .A1(n8131), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8151) );
  OAI211_X1 U10561 ( .C1(n7767), .C2(n8153), .A(n8152), .B(n8151), .ZN(n8154)
         );
  INV_X1 U10562 ( .A(n8154), .ZN(n8155) );
  OR2_X1 U10563 ( .A1(n13368), .A2(n13042), .ZN(n12736) );
  NAND2_X1 U10564 ( .A1(n13368), .A2(n13042), .ZN(n12737) );
  NAND2_X1 U10565 ( .A1(n12736), .A2(n12737), .ZN(n13230) );
  NAND2_X1 U10566 ( .A1(n13231), .A2(n13230), .ZN(n13229) );
  NAND2_X1 U10567 ( .A1(n13368), .A2(n13250), .ZN(n8157) );
  NAND2_X1 U10568 ( .A1(n13229), .A2(n8157), .ZN(n13218) );
  INV_X1 U10569 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15601) );
  NAND2_X1 U10570 ( .A1(n15601), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8175) );
  INV_X1 U10571 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11876) );
  NAND2_X1 U10572 ( .A1(n11876), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U10573 ( .A1(n8175), .A2(n8160), .ZN(n8172) );
  XNOR2_X1 U10574 ( .A(n8174), .B(n8172), .ZN(n11556) );
  NAND2_X1 U10575 ( .A1(n11556), .A2(n12601), .ZN(n8162) );
  NAND2_X1 U10576 ( .A1(n12602), .A2(SI_26_), .ZN(n8161) );
  NAND2_X1 U10577 ( .A1(n8163), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10578 ( .A1(n8180), .A2(n8164), .ZN(n13222) );
  NAND2_X1 U10579 ( .A1(n13222), .A2(n8209), .ZN(n8169) );
  INV_X1 U10580 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13365) );
  NAND2_X1 U10581 ( .A1(n8131), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10582 ( .A1(n9727), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8165) );
  OAI211_X1 U10583 ( .C1(n7767), .C2(n13365), .A(n8166), .B(n8165), .ZN(n8167)
         );
  INV_X1 U10584 ( .A(n8167), .ZN(n8168) );
  OR2_X1 U10585 ( .A1(n13361), .A2(n13233), .ZN(n8170) );
  XNOR2_X1 U10586 ( .A(n13361), .B(n13233), .ZN(n13217) );
  NAND2_X1 U10587 ( .A1(n13217), .A2(n13361), .ZN(n8171) );
  INV_X1 U10588 ( .A(n8172), .ZN(n8173) );
  INV_X1 U10589 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11966) );
  NAND2_X1 U10590 ( .A1(n11966), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8192) );
  INV_X1 U10591 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13959) );
  NAND2_X1 U10592 ( .A1(n13959), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8177) );
  NAND2_X1 U10593 ( .A1(n8192), .A2(n8177), .ZN(n8189) );
  XNOR2_X1 U10594 ( .A(n8191), .B(n8189), .ZN(n11637) );
  NAND2_X1 U10595 ( .A1(n11637), .A2(n12601), .ZN(n8179) );
  NAND2_X1 U10596 ( .A1(n12602), .A2(SI_27_), .ZN(n8178) );
  NAND2_X1 U10597 ( .A1(n8180), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10598 ( .A1(n8203), .A2(n8181), .ZN(n13207) );
  NAND2_X1 U10599 ( .A1(n13207), .A2(n8209), .ZN(n8187) );
  INV_X1 U10600 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n15474) );
  NAND2_X1 U10601 ( .A1(n8205), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8184) );
  INV_X1 U10602 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8182) );
  OR2_X1 U10603 ( .A1(n8112), .A2(n8182), .ZN(n8183) );
  OAI211_X1 U10604 ( .C1(n15474), .C2(n7754), .A(n8184), .B(n8183), .ZN(n8185)
         );
  INV_X1 U10605 ( .A(n8185), .ZN(n8186) );
  OR2_X1 U10606 ( .A1(n13358), .A2(n13216), .ZN(n8188) );
  NAND2_X1 U10607 ( .A1(n13193), .A2(n8188), .ZN(n8210) );
  INV_X1 U10608 ( .A(n8189), .ZN(n8190) );
  NAND2_X1 U10609 ( .A1(n8191), .A2(n8190), .ZN(n8193) );
  NAND2_X1 U10610 ( .A1(n8193), .A2(n8192), .ZN(n8197) );
  INV_X1 U10611 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11969) );
  NAND2_X1 U10612 ( .A1(n11969), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9722) );
  INV_X1 U10613 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U10614 ( .A1(n8194), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8195) );
  AND2_X1 U10615 ( .A1(n9722), .A2(n8195), .ZN(n8196) );
  NAND2_X1 U10616 ( .A1(n8197), .A2(n8196), .ZN(n9723) );
  OR2_X1 U10617 ( .A1(n8197), .A2(n8196), .ZN(n8198) );
  NAND2_X1 U10618 ( .A1(n12602), .A2(SI_28_), .ZN(n8200) );
  INV_X1 U10619 ( .A(n8203), .ZN(n8202) );
  INV_X1 U10620 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8201) );
  NAND2_X1 U10621 ( .A1(n8202), .A2(n8201), .ZN(n13174) );
  NAND2_X1 U10622 ( .A1(n8203), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8204) );
  NAND2_X1 U10623 ( .A1(n13174), .A2(n8204), .ZN(n13185) );
  INV_X1 U10624 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n15532) );
  NAND2_X1 U10625 ( .A1(n8205), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U10626 ( .A1(n8131), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8206) );
  OAI211_X1 U10627 ( .C1(n15532), .C2(n7754), .A(n8207), .B(n8206), .ZN(n8208)
         );
  NAND2_X1 U10628 ( .A1(n13353), .A2(n13198), .ZN(n12751) );
  NOR2_X2 U10629 ( .A1(n8210), .A2(n12904), .ZN(n9719) );
  NAND2_X1 U10630 ( .A1(n8210), .A2(n12904), .ZN(n8220) );
  NAND2_X1 U10631 ( .A1(n8257), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U10632 ( .A1(n12809), .A2(n12613), .ZN(n8293) );
  NAND2_X1 U10633 ( .A1(n8211), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8213) );
  MUX2_X1 U10634 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8213), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8214) );
  INV_X1 U10635 ( .A(n8214), .ZN(n8216) );
  NOR2_X1 U10636 ( .A1(n8216), .A2(n8215), .ZN(n9775) );
  INV_X1 U10637 ( .A(n8215), .ZN(n8217) );
  XNOR2_X2 U10638 ( .A(n8219), .B(n8218), .ZN(n12618) );
  INV_X1 U10639 ( .A(n12618), .ZN(n8226) );
  NAND2_X1 U10640 ( .A1(n9775), .A2(n8226), .ZN(n12615) );
  NAND2_X1 U10641 ( .A1(n8220), .A2(n15248), .ZN(n8221) );
  OR2_X1 U10642 ( .A1(n9719), .A2(n8221), .ZN(n8231) );
  OR2_X1 U10643 ( .A1(n13174), .A2(n6732), .ZN(n12595) );
  INV_X1 U10644 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U10645 ( .A1(n8131), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U10646 ( .A1(n9727), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8222) );
  OAI211_X1 U10647 ( .C1(n7767), .C2(n9781), .A(n8223), .B(n8222), .ZN(n8224)
         );
  INV_X1 U10648 ( .A(n8224), .ZN(n8225) );
  INV_X1 U10649 ( .A(n12806), .ZN(n10128) );
  INV_X1 U10650 ( .A(n12105), .ZN(n12807) );
  NAND2_X1 U10651 ( .A1(n10128), .A2(n12807), .ZN(n10139) );
  NAND2_X1 U10652 ( .A1(n10126), .A2(n10139), .ZN(n8228) );
  AND2_X2 U10653 ( .A1(n12809), .A2(n8226), .ZN(n8227) );
  INV_X1 U10654 ( .A(n13216), .ZN(n12900) );
  INV_X1 U10655 ( .A(n8228), .ZN(n10316) );
  NAND2_X1 U10656 ( .A1(n10316), .A2(n8227), .ZN(n13314) );
  OAI22_X1 U10657 ( .A1(n12909), .A2(n13312), .B1(n12900), .B2(n13314), .ZN(
        n8229) );
  INV_X1 U10658 ( .A(n8229), .ZN(n8230) );
  INV_X1 U10659 ( .A(n10248), .ZN(n10912) );
  NAND2_X1 U10660 ( .A1(n12625), .A2(n12619), .ZN(n10310) );
  NAND2_X1 U10661 ( .A1(n10310), .A2(n12624), .ZN(n15237) );
  NAND2_X1 U10662 ( .A1(n15236), .A2(n15237), .ZN(n15235) );
  NAND2_X1 U10663 ( .A1(n15235), .A2(n12629), .ZN(n10804) );
  INV_X1 U10664 ( .A(n12767), .ZN(n10803) );
  NAND2_X1 U10665 ( .A1(n10804), .A2(n10803), .ZN(n10806) );
  NAND2_X1 U10666 ( .A1(n10806), .A2(n8232), .ZN(n10842) );
  NAND2_X1 U10667 ( .A1(n10842), .A2(n12771), .ZN(n10844) );
  INV_X1 U10668 ( .A(n12956), .ZN(n11111) );
  NAND2_X1 U10669 ( .A1(n11111), .A2(n10697), .ZN(n12637) );
  NAND2_X1 U10670 ( .A1(n10844), .A2(n12637), .ZN(n10913) );
  NAND2_X1 U10671 ( .A1(n10913), .A2(n12646), .ZN(n8233) );
  NAND2_X1 U10672 ( .A1(n8233), .A2(n12642), .ZN(n10734) );
  INV_X1 U10673 ( .A(n12766), .ZN(n10733) );
  INV_X1 U10674 ( .A(n12652), .ZN(n11244) );
  NAND2_X1 U10675 ( .A1(n11244), .A2(n12818), .ZN(n12653) );
  INV_X1 U10676 ( .A(n12662), .ZN(n11150) );
  INV_X1 U10677 ( .A(n12668), .ZN(n8236) );
  OR2_X1 U10678 ( .A1(n11150), .A2(n8236), .ZN(n8234) );
  INV_X1 U10679 ( .A(n12669), .ZN(n12782) );
  AND2_X1 U10680 ( .A1(n12667), .A2(n12663), .ZN(n8235) );
  OR2_X1 U10681 ( .A1(n8236), .A2(n8235), .ZN(n11191) );
  AND2_X1 U10682 ( .A1(n12782), .A2(n11191), .ZN(n8237) );
  OR2_X1 U10683 ( .A1(n11946), .A2(n12824), .ZN(n12691) );
  NAND2_X1 U10684 ( .A1(n11946), .A2(n12824), .ZN(n12696) );
  NAND2_X1 U10685 ( .A1(n13457), .A2(n13052), .ZN(n12698) );
  NAND2_X1 U10686 ( .A1(n12949), .A2(n12940), .ZN(n12697) );
  NAND2_X1 U10687 ( .A1(n11849), .A2(n11848), .ZN(n11847) );
  NAND2_X1 U10688 ( .A1(n11847), .A2(n12697), .ZN(n11923) );
  NAND2_X1 U10689 ( .A1(n11923), .A2(n12789), .ZN(n8240) );
  NAND2_X1 U10690 ( .A1(n8242), .A2(n12713), .ZN(n13302) );
  OR2_X1 U10691 ( .A1(n13308), .A2(n13313), .ZN(n12718) );
  NAND2_X1 U10692 ( .A1(n13286), .A2(n13274), .ZN(n12722) );
  OR2_X1 U10693 ( .A1(n13286), .A2(n13274), .ZN(n12721) );
  NAND2_X1 U10694 ( .A1(n8244), .A2(n12721), .ZN(n13269) );
  NAND2_X1 U10695 ( .A1(n13275), .A2(n13285), .ZN(n12726) );
  NAND2_X1 U10696 ( .A1(n13269), .A2(n12726), .ZN(n8245) );
  NAND2_X1 U10697 ( .A1(n8245), .A2(n12725), .ZN(n13264) );
  NAND2_X1 U10698 ( .A1(n13372), .A2(n13256), .ZN(n12733) );
  INV_X1 U10699 ( .A(n13230), .ZN(n12792) );
  NAND2_X1 U10700 ( .A1(n8247), .A2(n12737), .ZN(n13213) );
  INV_X1 U10701 ( .A(n13217), .ZN(n13212) );
  OR2_X1 U10702 ( .A1(n13361), .A2(n13197), .ZN(n8248) );
  NAND2_X1 U10703 ( .A1(n13358), .A2(n12900), .ZN(n12742) );
  INV_X1 U10704 ( .A(n12904), .ZN(n12795) );
  XNOR2_X1 U10705 ( .A(n9739), .B(n12795), .ZN(n13189) );
  NAND2_X1 U10706 ( .A1(n12618), .A2(n10561), .ZN(n8250) );
  XNOR2_X1 U10707 ( .A(n12809), .B(n8250), .ZN(n8252) );
  NAND2_X1 U10708 ( .A1(n12618), .A2(n12800), .ZN(n8251) );
  NAND2_X1 U10709 ( .A1(n8252), .A2(n8251), .ZN(n10231) );
  NAND2_X1 U10710 ( .A1(n10561), .A2(n12800), .ZN(n9776) );
  INV_X1 U10711 ( .A(n9776), .ZN(n12616) );
  AND2_X1 U10712 ( .A1(n15295), .A2(n12616), .ZN(n8253) );
  NAND2_X1 U10713 ( .A1(n10231), .A2(n8253), .ZN(n8255) );
  NOR2_X1 U10714 ( .A1(n10561), .A2(n12613), .ZN(n8254) );
  NAND2_X1 U10715 ( .A1(n12809), .A2(n8254), .ZN(n9774) );
  NAND2_X1 U10716 ( .A1(n8255), .A2(n9774), .ZN(n13204) );
  NAND2_X1 U10717 ( .A1(n10561), .A2(n12613), .ZN(n12803) );
  INV_X1 U10718 ( .A(n12803), .ZN(n15240) );
  NAND2_X1 U10719 ( .A1(n13189), .A2(n15298), .ZN(n8256) );
  NAND2_X1 U10720 ( .A1(n8263), .A2(n8262), .ZN(n8274) );
  XNOR2_X1 U10721 ( .A(n8274), .B(P3_B_REG_SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10722 ( .A1(n8259), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8264) );
  MUX2_X1 U10723 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8264), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8266) );
  NAND2_X1 U10724 ( .A1(n8266), .A2(n8265), .ZN(n11423) );
  NAND2_X1 U10725 ( .A1(n8265), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8267) );
  MUX2_X1 U10726 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8267), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8269) );
  NAND2_X1 U10727 ( .A1(n8269), .A2(n8268), .ZN(n11559) );
  INV_X1 U10728 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U10729 ( .A1(n11950), .A2(n8271), .ZN(n8273) );
  NAND2_X1 U10730 ( .A1(n11559), .A2(n11423), .ZN(n8272) );
  INV_X1 U10731 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n15590) );
  NAND2_X1 U10732 ( .A1(n8274), .A2(n11559), .ZN(n8275) );
  NOR2_X1 U10733 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .ZN(
        n8279) );
  NOR4_X1 U10734 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8278) );
  NOR4_X1 U10735 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n8277) );
  NOR4_X1 U10736 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n8276) );
  NAND4_X1 U10737 ( .A1(n8279), .A2(n8278), .A3(n8277), .A4(n8276), .ZN(n8285)
         );
  NOR4_X1 U10738 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8283) );
  NOR4_X1 U10739 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n8282) );
  NOR4_X1 U10740 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8281) );
  NOR4_X1 U10741 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8280) );
  NAND4_X1 U10742 ( .A1(n8283), .A2(n8282), .A3(n8281), .A4(n8280), .ZN(n8284)
         );
  OAI21_X1 U10743 ( .B1(n8285), .B2(n8284), .A(n11950), .ZN(n9771) );
  NAND2_X1 U10744 ( .A1(n10299), .A2(n9771), .ZN(n8286) );
  INV_X1 U10745 ( .A(n8274), .ZN(n8288) );
  NOR2_X1 U10746 ( .A1(n11559), .A2(n11423), .ZN(n8287) );
  NAND2_X1 U10747 ( .A1(n8288), .A2(n8287), .ZN(n10236) );
  NAND2_X1 U10748 ( .A1(n8289), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8291) );
  XNOR2_X1 U10749 ( .A(n8291), .B(n8290), .ZN(n10232) );
  AND2_X1 U10750 ( .A1(n10671), .A2(n10231), .ZN(n8292) );
  NAND2_X1 U10751 ( .A1(n10243), .A2(n8292), .ZN(n8297) );
  INV_X1 U10752 ( .A(n10299), .ZN(n13460) );
  NAND3_X1 U10753 ( .A1(n13460), .A2(n13458), .A3(n9771), .ZN(n10245) );
  AND2_X1 U10754 ( .A1(n8227), .A2(n12616), .ZN(n10363) );
  NAND2_X1 U10755 ( .A1(n10671), .A2(n10363), .ZN(n12808) );
  NAND2_X1 U10756 ( .A1(n9775), .A2(n12618), .ZN(n12802) );
  NOR2_X1 U10757 ( .A1(n8293), .A2(n12802), .ZN(n10234) );
  NAND2_X1 U10758 ( .A1(n10671), .A2(n10234), .ZN(n8294) );
  AND2_X1 U10759 ( .A1(n12808), .A2(n8294), .ZN(n8295) );
  OR2_X1 U10760 ( .A1(n10245), .A2(n8295), .ZN(n8296) );
  INV_X1 U10761 ( .A(n13456), .ZN(n13410) );
  MUX2_X1 U10762 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n8317), .Z(n8304) );
  INV_X1 U10763 ( .A(n8308), .ZN(n8307) );
  MUX2_X1 U10764 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8317), .Z(n8309) );
  NAND2_X1 U10765 ( .A1(n8309), .A2(SI_3_), .ZN(n8312) );
  INV_X1 U10766 ( .A(n8309), .ZN(n8310) );
  NAND2_X1 U10767 ( .A1(n8310), .A2(n9833), .ZN(n8311) );
  AND2_X1 U10768 ( .A1(n8312), .A2(n8311), .ZN(n8460) );
  NAND2_X1 U10769 ( .A1(n8461), .A2(n8460), .ZN(n8463) );
  NAND2_X1 U10770 ( .A1(n8463), .A2(n8312), .ZN(n8472) );
  MUX2_X1 U10771 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8317), .Z(n8313) );
  NAND2_X1 U10772 ( .A1(n8313), .A2(SI_4_), .ZN(n8316) );
  INV_X1 U10773 ( .A(n8313), .ZN(n8314) );
  INV_X1 U10774 ( .A(SI_4_), .ZN(n9845) );
  NAND2_X1 U10775 ( .A1(n8314), .A2(n9845), .ZN(n8315) );
  MUX2_X1 U10776 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8317), .Z(n8318) );
  NAND2_X1 U10777 ( .A1(n8318), .A2(SI_5_), .ZN(n8322) );
  INV_X1 U10778 ( .A(n8318), .ZN(n8319) );
  INV_X1 U10779 ( .A(SI_5_), .ZN(n15673) );
  NAND2_X1 U10780 ( .A1(n8319), .A2(n15673), .ZN(n8320) );
  NAND2_X1 U10781 ( .A1(n8322), .A2(n8320), .ZN(n8480) );
  INV_X1 U10782 ( .A(n8480), .ZN(n8321) );
  NAND2_X1 U10783 ( .A1(n8323), .A2(SI_6_), .ZN(n8511) );
  INV_X1 U10784 ( .A(n8323), .ZN(n8324) );
  INV_X1 U10785 ( .A(SI_6_), .ZN(n9835) );
  NAND2_X1 U10786 ( .A1(n8324), .A2(n9835), .ZN(n8325) );
  NAND2_X1 U10787 ( .A1(n8326), .A2(SI_7_), .ZN(n8514) );
  INV_X1 U10788 ( .A(SI_7_), .ZN(n9838) );
  MUX2_X1 U10789 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9829), .Z(n8329) );
  NAND2_X1 U10790 ( .A1(n8329), .A2(SI_8_), .ZN(n8332) );
  INV_X1 U10791 ( .A(n8329), .ZN(n8330) );
  NAND2_X1 U10792 ( .A1(n8330), .A2(n9847), .ZN(n8331) );
  MUX2_X1 U10793 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9829), .Z(n8333) );
  INV_X1 U10794 ( .A(n8333), .ZN(n8334) );
  NAND2_X1 U10795 ( .A1(n8334), .A2(n9831), .ZN(n8335) );
  NAND2_X1 U10796 ( .A1(n8336), .A2(n8335), .ZN(n8543) );
  MUX2_X1 U10797 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9829), .Z(n8561) );
  MUX2_X1 U10798 ( .A(n9915), .B(n9917), .S(n9829), .Z(n8337) );
  INV_X1 U10799 ( .A(n8337), .ZN(n8338) );
  NAND2_X1 U10800 ( .A1(n8338), .A2(SI_11_), .ZN(n8339) );
  MUX2_X1 U10801 ( .A(n10054), .B(n10056), .S(n9829), .Z(n8341) );
  INV_X1 U10802 ( .A(n8341), .ZN(n8342) );
  NAND2_X1 U10803 ( .A1(n8342), .A2(SI_12_), .ZN(n8343) );
  MUX2_X1 U10804 ( .A(n10079), .B(n10081), .S(n9829), .Z(n8344) );
  NAND2_X1 U10805 ( .A1(n8344), .A2(n9913), .ZN(n8607) );
  INV_X1 U10806 ( .A(n8344), .ZN(n8345) );
  MUX2_X1 U10807 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n9829), .Z(n8349) );
  MUX2_X1 U10808 ( .A(n10371), .B(n10369), .S(n9829), .Z(n8624) );
  INV_X1 U10809 ( .A(n8624), .ZN(n8638) );
  NAND2_X1 U10810 ( .A1(n8638), .A2(SI_14_), .ZN(n8348) );
  INV_X1 U10811 ( .A(SI_14_), .ZN(n10013) );
  NAND3_X1 U10812 ( .A1(n8644), .A2(n10013), .A3(n8624), .ZN(n8351) );
  INV_X1 U10813 ( .A(n8349), .ZN(n8350) );
  INV_X1 U10814 ( .A(SI_15_), .ZN(n10058) );
  NAND2_X1 U10815 ( .A1(n8350), .A2(n10058), .ZN(n8643) );
  MUX2_X1 U10816 ( .A(n10328), .B(n10326), .S(n9829), .Z(n8353) );
  INV_X1 U10817 ( .A(n8353), .ZN(n8354) );
  NAND2_X1 U10818 ( .A1(n8354), .A2(SI_16_), .ZN(n8355) );
  MUX2_X1 U10819 ( .A(n10399), .B(n10401), .S(n9829), .Z(n8676) );
  INV_X1 U10820 ( .A(n8676), .ZN(n8357) );
  NAND2_X1 U10821 ( .A1(n8357), .A2(SI_17_), .ZN(n8358) );
  NAND2_X1 U10822 ( .A1(n8675), .A2(n8358), .ZN(n8360) );
  INV_X1 U10823 ( .A(SI_17_), .ZN(n10294) );
  NAND2_X1 U10824 ( .A1(n8676), .A2(n10294), .ZN(n8359) );
  MUX2_X1 U10825 ( .A(n10682), .B(n10681), .S(n9829), .Z(n8691) );
  MUX2_X1 U10826 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9829), .Z(n8365) );
  NAND2_X1 U10827 ( .A1(n8361), .A2(SI_18_), .ZN(n8362) );
  INV_X1 U10828 ( .A(n8365), .ZN(n8366) );
  INV_X1 U10829 ( .A(SI_19_), .ZN(n15620) );
  NAND2_X1 U10830 ( .A1(n8366), .A2(n15620), .ZN(n8367) );
  INV_X1 U10831 ( .A(SI_20_), .ZN(n10562) );
  NAND2_X1 U10832 ( .A1(n8369), .A2(n10562), .ZN(n8371) );
  INV_X1 U10833 ( .A(n8369), .ZN(n8370) );
  MUX2_X1 U10834 ( .A(n10904), .B(n10907), .S(n9829), .Z(n8721) );
  MUX2_X1 U10835 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9829), .Z(n8373) );
  NAND2_X1 U10836 ( .A1(n8373), .A2(SI_21_), .ZN(n8376) );
  INV_X1 U10837 ( .A(n8373), .ZN(n8374) );
  INV_X1 U10838 ( .A(SI_21_), .ZN(n10732) );
  NAND2_X1 U10839 ( .A1(n8374), .A2(n10732), .ZN(n8375) );
  MUX2_X1 U10840 ( .A(n8379), .B(n11391), .S(n9829), .Z(n9366) );
  MUX2_X1 U10841 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9829), .Z(n8763) );
  INV_X1 U10842 ( .A(SI_23_), .ZN(n10998) );
  NAND2_X1 U10843 ( .A1(n8381), .A2(n10998), .ZN(n8382) );
  MUX2_X1 U10844 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9829), .Z(n8383) );
  NAND2_X1 U10845 ( .A1(n8383), .A2(SI_24_), .ZN(n8387) );
  INV_X1 U10846 ( .A(n8383), .ZN(n8384) );
  INV_X1 U10847 ( .A(SI_24_), .ZN(n11261) );
  NAND2_X1 U10848 ( .A1(n8384), .A2(n11261), .ZN(n8385) );
  MUX2_X1 U10849 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9829), .Z(n8389) );
  XNOR2_X1 U10850 ( .A(n8389), .B(SI_25_), .ZN(n8788) );
  INV_X1 U10851 ( .A(n8389), .ZN(n8390) );
  INV_X1 U10852 ( .A(SI_25_), .ZN(n15454) );
  NAND2_X1 U10853 ( .A1(n8390), .A2(n15454), .ZN(n8391) );
  INV_X1 U10854 ( .A(SI_26_), .ZN(n11557) );
  MUX2_X1 U10855 ( .A(n15601), .B(n11876), .S(n9829), .Z(n8798) );
  INV_X1 U10856 ( .A(n8798), .ZN(n8392) );
  MUX2_X1 U10857 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9829), .Z(n9447) );
  INV_X1 U10858 ( .A(n8394), .ZN(n8396) );
  MUX2_X1 U10859 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n9829), .Z(n9448) );
  XNOR2_X1 U10860 ( .A(n9448), .B(SI_28_), .ZN(n8395) );
  INV_X1 U10861 ( .A(n8458), .ZN(n8400) );
  NAND2_X1 U10862 ( .A1(n11967), .A2(n6643), .ZN(n8409) );
  OR2_X1 U10863 ( .A1(n12495), .A2(n11969), .ZN(n8408) );
  NAND2_X1 U10864 ( .A1(n9755), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8423) );
  OR2_X1 U10865 ( .A1(n8453), .A2(n6681), .ZN(n8422) );
  NAND2_X1 U10866 ( .A1(n8505), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8521) );
  AND2_X1 U10867 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n8415) );
  INV_X1 U10868 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U10869 ( .A1(n8631), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8653) );
  INV_X1 U10870 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8652) );
  INV_X1 U10871 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8668) );
  INV_X1 U10872 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n15441) );
  INV_X1 U10873 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U10874 ( .A1(n8753), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U10875 ( .A1(n8769), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U10876 ( .A1(n8780), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8779) );
  NAND3_X1 U10877 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG3_REG_26__SCAN_IN), 
        .A3(n8803), .ZN(n8814) );
  INV_X1 U10878 ( .A(n8814), .ZN(n8416) );
  NAND2_X1 U10879 ( .A1(n8416), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8816) );
  INV_X1 U10880 ( .A(n8816), .ZN(n8417) );
  NAND2_X1 U10881 ( .A1(n8417), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14318) );
  INV_X1 U10882 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n15462) );
  NAND2_X1 U10883 ( .A1(n8816), .A2(n15462), .ZN(n8418) );
  NAND2_X1 U10884 ( .A1(n14318), .A2(n8418), .ZN(n14329) );
  OR2_X1 U10885 ( .A1(n8868), .A2(n14329), .ZN(n8421) );
  INV_X1 U10886 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14330) );
  OR2_X1 U10887 ( .A1(n8781), .A2(n14330), .ZN(n8420) );
  NAND2_X1 U10888 ( .A1(n9755), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10889 ( .A1(n6654), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U10890 ( .A1(n8437), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10891 ( .A1(n8443), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8424) );
  XNOR2_X1 U10892 ( .A(n8429), .B(n8430), .ZN(n9874) );
  OR2_X1 U10893 ( .A1(n8741), .A2(n9874), .ZN(n8435) );
  OR2_X1 U10894 ( .A1(n12495), .A2(n8300), .ZN(n8434) );
  INV_X1 U10895 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U10896 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8431) );
  XNOR2_X1 U10897 ( .A(n8432), .B(n8431), .ZN(n10035) );
  OR2_X1 U10898 ( .A1(n9884), .A2(n10035), .ZN(n8433) );
  NAND2_X1 U10899 ( .A1(n8437), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10900 ( .A1(n8443), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8438) );
  INV_X1 U10901 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10349) );
  INV_X1 U10902 ( .A(SI_0_), .ZN(n8441) );
  NOR2_X1 U10903 ( .A1(n9829), .A2(n8441), .ZN(n8442) );
  XNOR2_X1 U10904 ( .A(n8442), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14658) );
  MUX2_X1 U10905 ( .A(n10349), .B(n14658), .S(n9884), .Z(n14908) );
  INV_X1 U10906 ( .A(n14908), .ZN(n10360) );
  AND2_X1 U10907 ( .A1(n8837), .A2(n10360), .ZN(n14915) );
  NAND2_X1 U10908 ( .A1(n8437), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8446) );
  NAND2_X1 U10909 ( .A1(n9755), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8444) );
  XNOR2_X1 U10910 ( .A(n8449), .B(n8450), .ZN(n9871) );
  NAND2_X1 U10911 ( .A1(n14157), .A2(n14969), .ZN(n8451) );
  INV_X1 U10912 ( .A(n14890), .ZN(n14894) );
  NAND2_X1 U10913 ( .A1(n14893), .A2(n14894), .ZN(n8452) );
  NAND2_X1 U10914 ( .A1(n8452), .A2(n12311), .ZN(n11344) );
  NAND2_X1 U10915 ( .A1(n8443), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10916 ( .A1(n6733), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10917 ( .A1(n9755), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8455) );
  OR2_X1 U10918 ( .A1(n8868), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8454) );
  INV_X2 U10919 ( .A(n9884), .ZN(n8711) );
  NAND2_X1 U10920 ( .A1(n8458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8459) );
  XNOR2_X1 U10921 ( .A(n8459), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14195) );
  OR2_X1 U10922 ( .A1(n8461), .A2(n8460), .ZN(n8462) );
  AND2_X1 U10923 ( .A1(n8463), .A2(n8462), .ZN(n9825) );
  NAND2_X1 U10924 ( .A1(n9825), .A2(n12497), .ZN(n8464) );
  XNOR2_X2 U10925 ( .A(n14975), .B(n14156), .ZN(n12514) );
  INV_X1 U10926 ( .A(n12514), .ZN(n8465) );
  INV_X1 U10927 ( .A(n14156), .ZN(n12322) );
  NAND2_X1 U10928 ( .A1(n12322), .A2(n11340), .ZN(n8466) );
  NAND2_X1 U10929 ( .A1(n9755), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10930 ( .A1(n12478), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8469) );
  XNOR2_X1 U10931 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11330) );
  OR2_X1 U10932 ( .A1(n8868), .A2(n11330), .ZN(n8468) );
  NAND2_X1 U10933 ( .A1(n6645), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8467) );
  NAND4_X1 U10934 ( .A1(n8470), .A2(n8469), .A3(n8468), .A4(n8467), .ZN(n14155) );
  OR2_X1 U10935 ( .A1(n8472), .A2(n8471), .ZN(n8473) );
  NAND2_X1 U10936 ( .A1(n8474), .A2(n8473), .ZN(n9856) );
  OR2_X1 U10937 ( .A1(n9856), .A2(n8741), .ZN(n8477) );
  OR2_X1 U10938 ( .A1(n8458), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U10939 ( .A1(n8482), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8475) );
  XNOR2_X1 U10940 ( .A(n8475), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14210) );
  AOI22_X1 U10941 ( .A1(n8712), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8711), .B2(
        n14210), .ZN(n8476) );
  NAND2_X1 U10942 ( .A1(n8477), .A2(n8476), .ZN(n12327) );
  NOR2_X1 U10943 ( .A1(n14155), .A2(n12327), .ZN(n8479) );
  NAND2_X1 U10944 ( .A1(n14155), .A2(n12327), .ZN(n8478) );
  XNOR2_X1 U10945 ( .A(n8481), .B(n8480), .ZN(n9840) );
  NAND2_X1 U10946 ( .A1(n9840), .A2(n6643), .ZN(n8491) );
  INV_X1 U10947 ( .A(n8482), .ZN(n8484) );
  INV_X1 U10948 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U10949 ( .A1(n8484), .A2(n8483), .ZN(n8486) );
  NAND2_X1 U10950 ( .A1(n8486), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8485) );
  MUX2_X1 U10951 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8485), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n8489) );
  INV_X1 U10952 ( .A(n8486), .ZN(n8488) );
  NAND2_X1 U10953 ( .A1(n8488), .A2(n8487), .ZN(n8517) );
  AOI22_X1 U10954 ( .A1(n8712), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8711), .B2(
        n10042), .ZN(n8490) );
  NAND2_X1 U10955 ( .A1(n8491), .A2(n8490), .ZN(n12331) );
  NAND2_X1 U10956 ( .A1(n12478), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10957 ( .A1(n6645), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8495) );
  AOI21_X1 U10958 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8492) );
  NOR2_X1 U10959 ( .A1(n8492), .A2(n8505), .ZN(n11137) );
  NAND2_X1 U10960 ( .A1(n8437), .A2(n11137), .ZN(n8494) );
  NAND2_X1 U10961 ( .A1(n9755), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8493) );
  NAND4_X1 U10962 ( .A1(n8496), .A2(n8495), .A3(n8494), .A4(n8493), .ZN(n14154) );
  XNOR2_X1 U10963 ( .A(n12331), .B(n14154), .ZN(n12518) );
  OR2_X1 U10964 ( .A1(n12331), .A2(n14154), .ZN(n8498) );
  OR2_X1 U10965 ( .A1(n9849), .A2(n8741), .ZN(n8504) );
  NAND2_X1 U10966 ( .A1(n8517), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8502) );
  XNOR2_X1 U10967 ( .A(n8502), .B(P1_IR_REG_6__SCAN_IN), .ZN(n14223) );
  AOI22_X1 U10968 ( .A1(n8712), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8711), .B2(
        n14223), .ZN(n8503) );
  AND2_X2 U10969 ( .A1(n8504), .A2(n8503), .ZN(n12348) );
  INV_X1 U10970 ( .A(n12348), .ZN(n12343) );
  NAND2_X1 U10971 ( .A1(n9755), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8509) );
  INV_X1 U10972 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10021) );
  OR2_X1 U10973 ( .A1(n8453), .A2(n10021), .ZN(n8508) );
  OAI21_X1 U10974 ( .B1(n8505), .B2(P1_REG3_REG_6__SCAN_IN), .A(n8521), .ZN(
        n11371) );
  OR2_X1 U10975 ( .A1(n8868), .A2(n11371), .ZN(n8507) );
  INV_X1 U10976 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11370) );
  OR2_X1 U10977 ( .A1(n8781), .A2(n11370), .ZN(n8506) );
  XNOR2_X1 U10978 ( .A(n12343), .B(n14153), .ZN(n12520) );
  INV_X1 U10979 ( .A(n12520), .ZN(n10881) );
  NAND2_X1 U10980 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  OAI21_X1 U10981 ( .B1(n8517), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8518) );
  XNOR2_X1 U10982 ( .A(n8518), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10043) );
  AOI22_X1 U10983 ( .A1(n8712), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8711), .B2(
        n10043), .ZN(n8519) );
  NAND2_X1 U10984 ( .A1(n9755), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U10985 ( .A1(n12478), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8525) );
  AND2_X1 U10986 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  OR2_X1 U10987 ( .A1(n8522), .A2(n8536), .ZN(n11394) );
  OR2_X1 U10988 ( .A1(n8868), .A2(n11394), .ZN(n8524) );
  NAND2_X1 U10989 ( .A1(n6645), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8523) );
  NAND4_X1 U10990 ( .A1(n8526), .A2(n8525), .A3(n8524), .A4(n8523), .ZN(n14152) );
  XNOR2_X1 U10991 ( .A(n12342), .B(n12341), .ZN(n12522) );
  NOR2_X1 U10992 ( .A1(n12342), .A2(n14152), .ZN(n12349) );
  INV_X1 U10993 ( .A(n12349), .ZN(n8527) );
  NAND2_X1 U10994 ( .A1(n11043), .A2(n8527), .ZN(n11353) );
  OR2_X1 U10995 ( .A1(n8529), .A2(n8528), .ZN(n8531) );
  NAND2_X1 U10996 ( .A1(n8531), .A2(n8530), .ZN(n9866) );
  OR2_X1 U10997 ( .A1(n9866), .A2(n8741), .ZN(n8535) );
  NAND2_X1 U10998 ( .A1(n8532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8533) );
  XNOR2_X1 U10999 ( .A(n8533), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11000 ( .A1(n8712), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8711), .B2(
        n10103), .ZN(n8534) );
  NAND2_X1 U11001 ( .A1(n9755), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U11002 ( .A1(n12478), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U11003 ( .A1(n6645), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8539) );
  NOR2_X1 U11004 ( .A1(n8536), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8537) );
  OR2_X1 U11005 ( .A1(n8566), .A2(n8537), .ZN(n11552) );
  OR2_X1 U11006 ( .A1(n8868), .A2(n11552), .ZN(n8538) );
  NAND4_X1 U11007 ( .A1(n8541), .A2(n8540), .A3(n8539), .A4(n8538), .ZN(n14151) );
  INV_X1 U11008 ( .A(n14151), .ZN(n11543) );
  OR2_X1 U11009 ( .A1(n12363), .A2(n11543), .ZN(n8849) );
  NAND2_X1 U11010 ( .A1(n12363), .A2(n11543), .ZN(n8542) );
  NAND2_X1 U11011 ( .A1(n8849), .A2(n8542), .ZN(n12523) );
  NAND2_X1 U11012 ( .A1(n11353), .A2(n12523), .ZN(n11352) );
  OR2_X1 U11013 ( .A1(n12363), .A2(n14151), .ZN(n12355) );
  NAND2_X1 U11014 ( .A1(n11352), .A2(n12355), .ZN(n11477) );
  XNOR2_X1 U11015 ( .A(n8544), .B(n8543), .ZN(n9875) );
  NAND2_X1 U11016 ( .A1(n9875), .A2(n6643), .ZN(n8554) );
  INV_X1 U11017 ( .A(n8532), .ZN(n8546) );
  INV_X1 U11018 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U11019 ( .A1(n8546), .A2(n8545), .ZN(n8548) );
  NAND2_X1 U11020 ( .A1(n8548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8547) );
  MUX2_X1 U11021 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8547), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n8551) );
  INV_X1 U11022 ( .A(n8548), .ZN(n8550) );
  INV_X1 U11023 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U11024 ( .A1(n8550), .A2(n8549), .ZN(n8577) );
  NAND2_X1 U11025 ( .A1(n8551), .A2(n8577), .ZN(n10282) );
  INV_X1 U11026 ( .A(n10282), .ZN(n8552) );
  AOI22_X1 U11027 ( .A1(n8712), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8711), .B2(
        n8552), .ZN(n8553) );
  NAND2_X1 U11028 ( .A1(n12478), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U11029 ( .A1(n6645), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8557) );
  XNOR2_X1 U11030 ( .A(n8566), .B(P1_REG3_REG_9__SCAN_IN), .ZN(n14881) );
  OR2_X1 U11031 ( .A1(n8868), .A2(n14881), .ZN(n8556) );
  NAND2_X1 U11032 ( .A1(n9755), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8555) );
  NAND4_X1 U11033 ( .A1(n8558), .A2(n8557), .A3(n8556), .A4(n8555), .ZN(n14150) );
  XNOR2_X1 U11034 ( .A(n12368), .B(n14150), .ZN(n12524) );
  OR2_X1 U11035 ( .A1(n12368), .A2(n14150), .ZN(n8559) );
  XNOR2_X1 U11036 ( .A(n8561), .B(SI_10_), .ZN(n8562) );
  XNOR2_X1 U11037 ( .A(n8560), .B(n8562), .ZN(n9886) );
  NAND2_X1 U11038 ( .A1(n9886), .A2(n6643), .ZN(n8565) );
  NAND2_X1 U11039 ( .A1(n8577), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8563) );
  XNOR2_X1 U11040 ( .A(n8563), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14256) );
  AOI22_X1 U11041 ( .A1(n8712), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8711), 
        .B2(n14256), .ZN(n8564) );
  NAND2_X1 U11042 ( .A1(n9755), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11043 ( .A1(n12478), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U11044 ( .A1(n8566), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8568) );
  INV_X1 U11045 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U11046 ( .A1(n8568), .A2(n8567), .ZN(n8569) );
  NAND2_X1 U11047 ( .A1(n8569), .A2(n8581), .ZN(n11715) );
  OR2_X1 U11048 ( .A1(n8868), .A2(n11715), .ZN(n8571) );
  NAND2_X1 U11049 ( .A1(n6645), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8570) );
  NAND4_X1 U11050 ( .A1(n8573), .A2(n8572), .A3(n8571), .A4(n8570), .ZN(n14149) );
  INV_X1 U11051 ( .A(n14149), .ZN(n12374) );
  OR2_X1 U11052 ( .A1(n12372), .A2(n12374), .ZN(n8851) );
  NAND2_X1 U11053 ( .A1(n12372), .A2(n12374), .ZN(n8574) );
  NAND2_X1 U11054 ( .A1(n9914), .A2(n6643), .ZN(n8580) );
  NAND2_X1 U11055 ( .A1(n8589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8578) );
  XNOR2_X1 U11056 ( .A(n8578), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U11057 ( .A1(n8712), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8711), 
        .B2(n10571), .ZN(n8579) );
  NAND2_X1 U11058 ( .A1(n9755), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U11059 ( .A1(n12478), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U11060 ( .A1(n6645), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U11061 ( .A1(n8581), .A2(n11887), .ZN(n8582) );
  NAND2_X1 U11062 ( .A1(n8592), .A2(n8582), .ZN(n11886) );
  OR2_X1 U11063 ( .A1(n8868), .A2(n11886), .ZN(n8583) );
  NAND4_X1 U11064 ( .A1(n8586), .A2(n8585), .A3(n8584), .A4(n8583), .ZN(n14148) );
  XNOR2_X1 U11065 ( .A(n8588), .B(n8587), .ZN(n10053) );
  NAND2_X1 U11066 ( .A1(n10053), .A2(n6643), .ZN(n8591) );
  OAI21_X1 U11067 ( .B1(n8589), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8611) );
  XNOR2_X1 U11068 ( .A(n8611), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U11069 ( .A1(n8712), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8711), 
        .B2(n10793), .ZN(n8590) );
  NAND2_X1 U11070 ( .A1(n9755), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11071 ( .A1(n12478), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U11072 ( .A1(n6645), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U11073 ( .A1(n8592), .A2(n10574), .ZN(n8593) );
  NAND2_X1 U11074 ( .A1(n8616), .A2(n8593), .ZN(n14009) );
  OR2_X1 U11075 ( .A1(n8868), .A2(n14009), .ZN(n8594) );
  NAND4_X1 U11076 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n14147) );
  INV_X1 U11077 ( .A(n14147), .ZN(n12144) );
  XNOR2_X1 U11078 ( .A(n12382), .B(n12144), .ZN(n12530) );
  AND2_X1 U11079 ( .A1(n11310), .A2(n8599), .ZN(n8598) );
  INV_X1 U11080 ( .A(n8599), .ZN(n8600) );
  OR2_X1 U11081 ( .A1(n12372), .A2(n14149), .ZN(n11519) );
  OR2_X1 U11082 ( .A1(n8600), .A2(n11519), .ZN(n8601) );
  INV_X1 U11083 ( .A(n12530), .ZN(n11525) );
  OR2_X1 U11084 ( .A1(n12377), .A2(n14148), .ZN(n11521) );
  OR2_X1 U11085 ( .A1(n11525), .A2(n11521), .ZN(n8602) );
  OR2_X1 U11086 ( .A1(n12382), .A2(n14147), .ZN(n8603) );
  NAND2_X1 U11087 ( .A1(n8605), .A2(n8604), .ZN(n8609) );
  AND2_X1 U11088 ( .A1(n8607), .A2(n8606), .ZN(n8608) );
  XNOR2_X1 U11089 ( .A(n8609), .B(n8608), .ZN(n10078) );
  NAND2_X1 U11090 ( .A1(n10078), .A2(n6643), .ZN(n8614) );
  NAND2_X1 U11091 ( .A1(n8611), .A2(n8610), .ZN(n8612) );
  NAND2_X1 U11092 ( .A1(n8612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8626) );
  XNOR2_X1 U11093 ( .A(n8626), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U11094 ( .A1(n8712), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10794), 
        .B2(n8711), .ZN(n8613) );
  NAND2_X1 U11095 ( .A1(n12478), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8621) );
  AND2_X1 U11096 ( .A1(n8616), .A2(n8615), .ZN(n8617) );
  OR2_X1 U11097 ( .A1(n8617), .A2(n8631), .ZN(n14074) );
  OR2_X1 U11098 ( .A1(n8868), .A2(n14074), .ZN(n8620) );
  NAND2_X1 U11099 ( .A1(n6645), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U11100 ( .A1(n9755), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8618) );
  NAND4_X1 U11101 ( .A1(n8621), .A2(n8620), .A3(n8619), .A4(n8618), .ZN(n14146) );
  OR2_X1 U11102 ( .A1(n12387), .A2(n12389), .ZN(n8853) );
  NAND2_X1 U11103 ( .A1(n12387), .A2(n12389), .ZN(n8622) );
  NAND2_X1 U11104 ( .A1(n8853), .A2(n8622), .ZN(n12529) );
  NAND2_X1 U11105 ( .A1(n11618), .A2(n12529), .ZN(n11617) );
  OR2_X1 U11106 ( .A1(n12387), .A2(n14146), .ZN(n8623) );
  XNOR2_X1 U11107 ( .A(n8640), .B(SI_14_), .ZN(n8639) );
  XNOR2_X1 U11108 ( .A(n8639), .B(n8624), .ZN(n10368) );
  NAND2_X1 U11109 ( .A1(n10368), .A2(n6643), .ZN(n8630) );
  INV_X1 U11110 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U11111 ( .A1(n8626), .A2(n8625), .ZN(n8627) );
  NAND2_X1 U11112 ( .A1(n8627), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8628) );
  XNOR2_X1 U11113 ( .A(n8628), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U11114 ( .A1(n11063), .A2(n8711), .B1(n8712), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11115 ( .A1(n9755), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8636) );
  OR2_X1 U11116 ( .A1(n8631), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U11117 ( .A1(n8653), .A2(n8632), .ZN(n14835) );
  OR2_X1 U11118 ( .A1(n8868), .A2(n14835), .ZN(n8635) );
  INV_X1 U11119 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11783) );
  OR2_X1 U11120 ( .A1(n8781), .A2(n11783), .ZN(n8634) );
  INV_X1 U11121 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11775) );
  OR2_X1 U11122 ( .A1(n8453), .A2(n11775), .ZN(n8633) );
  NAND2_X1 U11123 ( .A1(n14832), .A2(n12157), .ZN(n12391) );
  NAND2_X1 U11124 ( .A1(n8639), .A2(n8638), .ZN(n8642) );
  OR2_X1 U11125 ( .A1(n8640), .A2(n10013), .ZN(n8641) );
  NAND2_X1 U11126 ( .A1(n8642), .A2(n8641), .ZN(n8646) );
  NAND2_X1 U11127 ( .A1(n8644), .A2(n8643), .ZN(n8645) );
  NAND2_X1 U11128 ( .A1(n10394), .A2(n6643), .ZN(n8650) );
  OR2_X1 U11129 ( .A1(n8647), .A2(n8411), .ZN(n8648) );
  XNOR2_X1 U11130 ( .A(n8648), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U11131 ( .A1(n8712), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8711), 
        .B2(n11785), .ZN(n8649) );
  NAND2_X1 U11132 ( .A1(n9755), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8658) );
  INV_X1 U11133 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14866) );
  OR2_X1 U11134 ( .A1(n8453), .A2(n14866), .ZN(n8657) );
  INV_X1 U11135 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8651) );
  OR2_X1 U11136 ( .A1(n8781), .A2(n8651), .ZN(n8656) );
  NAND2_X1 U11137 ( .A1(n8653), .A2(n8652), .ZN(n8654) );
  NAND2_X1 U11138 ( .A1(n8669), .A2(n8654), .ZN(n11839) );
  OR2_X1 U11139 ( .A1(n8868), .A2(n11839), .ZN(n8655) );
  NAND2_X1 U11140 ( .A1(n14647), .A2(n11666), .ZN(n12412) );
  NAND2_X1 U11141 ( .A1(n12411), .A2(n12412), .ZN(n12533) );
  INV_X1 U11142 ( .A(n12157), .ZN(n14145) );
  NAND2_X1 U11143 ( .A1(n14832), .A2(n14145), .ZN(n11830) );
  AND2_X1 U11144 ( .A1(n12533), .A2(n11830), .ZN(n8659) );
  INV_X1 U11145 ( .A(n11666), .ZN(n14144) );
  XNOR2_X1 U11146 ( .A(n8660), .B(n8661), .ZN(n10325) );
  NAND2_X1 U11147 ( .A1(n10325), .A2(n6643), .ZN(n8665) );
  AND2_X1 U11148 ( .A1(n8647), .A2(n8662), .ZN(n8679) );
  OR2_X1 U11149 ( .A1(n8679), .A2(n8411), .ZN(n8663) );
  XNOR2_X1 U11150 ( .A(n8663), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U11151 ( .A1(n8712), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8711), 
        .B2(n11906), .ZN(n8664) );
  INV_X1 U11152 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8673) );
  NAND2_X1 U11153 ( .A1(n12478), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8667) );
  INV_X1 U11154 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15640) );
  OR2_X1 U11155 ( .A1(n12481), .A2(n15640), .ZN(n8666) );
  AND2_X1 U11156 ( .A1(n8667), .A2(n8666), .ZN(n8672) );
  AND2_X1 U11157 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  NOR2_X1 U11158 ( .A1(n8683), .A2(n8670), .ZN(n14034) );
  NAND2_X1 U11159 ( .A1(n14034), .A2(n8437), .ZN(n8671) );
  OAI211_X1 U11160 ( .C1(n8781), .C2(n8673), .A(n8672), .B(n8671), .ZN(n14143)
         );
  INV_X1 U11161 ( .A(n14143), .ZN(n14046) );
  XNOR2_X1 U11162 ( .A(n14039), .B(n14046), .ZN(n12531) );
  NAND2_X1 U11163 ( .A1(n11916), .A2(n12531), .ZN(n11915) );
  OR2_X1 U11164 ( .A1(n14039), .A2(n14143), .ZN(n8674) );
  XNOR2_X1 U11165 ( .A(n8676), .B(SI_17_), .ZN(n8677) );
  XNOR2_X1 U11166 ( .A(n8675), .B(n8677), .ZN(n10398) );
  NAND2_X1 U11167 ( .A1(n10398), .A2(n6643), .ZN(n8682) );
  NAND2_X1 U11168 ( .A1(n8679), .A2(n8678), .ZN(n8694) );
  NAND2_X1 U11169 ( .A1(n8694), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8680) );
  XNOR2_X1 U11170 ( .A(n8680), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14270) );
  AOI22_X1 U11171 ( .A1(n8712), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8711), 
        .B2(n14270), .ZN(n8681) );
  NOR2_X1 U11172 ( .A1(n8683), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8684) );
  OR2_X1 U11173 ( .A1(n8698), .A2(n8684), .ZN(n14508) );
  AOI22_X1 U11174 ( .A1(n9755), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n12478), 
        .B2(P1_REG1_REG_17__SCAN_IN), .ZN(n8686) );
  NAND2_X1 U11175 ( .A1(n6645), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8685) );
  OAI211_X1 U11176 ( .C1(n14508), .C2(n8868), .A(n8686), .B(n8685), .ZN(n14142) );
  INV_X1 U11177 ( .A(n14142), .ZN(n12406) );
  AND2_X1 U11178 ( .A1(n14514), .A2(n12406), .ZN(n8688) );
  OR2_X1 U11179 ( .A1(n14514), .A2(n12406), .ZN(n8687) );
  INV_X1 U11180 ( .A(SI_18_), .ZN(n10330) );
  OR2_X1 U11181 ( .A1(n8689), .A2(n10330), .ZN(n8704) );
  NAND2_X1 U11182 ( .A1(n8689), .A2(n10330), .ZN(n8690) );
  NAND2_X1 U11183 ( .A1(n8704), .A2(n8690), .ZN(n8692) );
  NAND2_X1 U11184 ( .A1(n8692), .A2(n8691), .ZN(n8693) );
  OAI21_X1 U11185 ( .B1(n8694), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8695) );
  XNOR2_X1 U11186 ( .A(n8695), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14289) );
  AOI22_X1 U11187 ( .A1(n8712), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8711), 
        .B2(n14289), .ZN(n8696) );
  NAND2_X2 U11188 ( .A1(n8697), .A2(n8696), .ZN(n14583) );
  OR2_X1 U11189 ( .A1(n8698), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8699) );
  AND2_X1 U11190 ( .A1(n8715), .A2(n8699), .ZN(n14494) );
  NAND2_X1 U11191 ( .A1(n14494), .A2(n8437), .ZN(n8702) );
  AOI22_X1 U11192 ( .A1(n9755), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n12478), 
        .B2(P1_REG1_REG_18__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U11193 ( .A1(n6645), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8700) );
  INV_X1 U11194 ( .A(n14047), .ZN(n14141) );
  NAND2_X1 U11195 ( .A1(n14583), .A2(n14141), .ZN(n8703) );
  NAND2_X1 U11196 ( .A1(n8705), .A2(n8704), .ZN(n8707) );
  XNOR2_X1 U11197 ( .A(n8707), .B(n8706), .ZN(n10973) );
  NAND2_X1 U11198 ( .A1(n8708), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8709) );
  MUX2_X1 U11199 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8709), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n8710) );
  AOI22_X1 U11200 ( .A1(n8712), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8918), 
        .B2(n8711), .ZN(n8713) );
  NAND2_X1 U11201 ( .A1(n8715), .A2(n15441), .ZN(n8716) );
  AND2_X1 U11202 ( .A1(n8728), .A2(n8716), .ZN(n14474) );
  INV_X1 U11203 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14286) );
  NAND2_X1 U11204 ( .A1(n9755), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11205 ( .A1(n6645), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8717) );
  OAI211_X1 U11206 ( .C1(n8453), .C2(n14286), .A(n8718), .B(n8717), .ZN(n8719)
         );
  AOI21_X1 U11207 ( .B1(n14474), .B2(n8437), .A(n8719), .ZN(n14096) );
  INV_X1 U11208 ( .A(n14096), .ZN(n14140) );
  OR2_X1 U11209 ( .A1(n14637), .A2(n14140), .ZN(n8720) );
  NAND2_X1 U11210 ( .A1(n14471), .A2(n8720), .ZN(n14455) );
  NAND2_X1 U11211 ( .A1(n8722), .A2(n8721), .ZN(n8723) );
  NAND2_X1 U11212 ( .A1(n8724), .A2(n8723), .ZN(n10905) );
  OR2_X1 U11213 ( .A1(n10905), .A2(n8741), .ZN(n8726) );
  OR2_X1 U11214 ( .A1(n12495), .A2(n10904), .ZN(n8725) );
  AND2_X1 U11215 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  OR2_X1 U11216 ( .A1(n8729), .A2(n8744), .ZN(n14461) );
  INV_X1 U11217 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11218 ( .A1(n12478), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11219 ( .A1(n6645), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8730) );
  OAI211_X1 U11220 ( .C1(n12481), .C2(n8732), .A(n8731), .B(n8730), .ZN(n8733)
         );
  INV_X1 U11221 ( .A(n8733), .ZN(n8734) );
  OAI21_X1 U11222 ( .B1(n14461), .B2(n8868), .A(n8734), .ZN(n14139) );
  INV_X1 U11223 ( .A(n14139), .ZN(n12203) );
  OR2_X1 U11224 ( .A1(n14570), .A2(n12203), .ZN(n8858) );
  NAND2_X1 U11225 ( .A1(n14570), .A2(n12203), .ZN(n8735) );
  NAND2_X1 U11226 ( .A1(n8858), .A2(n8735), .ZN(n14456) );
  INV_X1 U11227 ( .A(n14456), .ZN(n14454) );
  NAND2_X1 U11228 ( .A1(n14570), .A2(n14139), .ZN(n8736) );
  OR2_X1 U11229 ( .A1(n8738), .A2(n8737), .ZN(n8739) );
  NAND2_X1 U11230 ( .A1(n8740), .A2(n8739), .ZN(n11134) );
  OR2_X1 U11231 ( .A1(n11134), .A2(n8741), .ZN(n8743) );
  OR2_X1 U11232 ( .A1(n12495), .A2(n11040), .ZN(n8742) );
  NOR2_X1 U11233 ( .A1(n8744), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8745) );
  OR2_X1 U11234 ( .A1(n8753), .A2(n8745), .ZN(n14447) );
  INV_X1 U11235 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11236 ( .A1(n6645), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U11237 ( .A1(n12478), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8746) );
  OAI211_X1 U11238 ( .C1(n12481), .C2(n8748), .A(n8747), .B(n8746), .ZN(n8749)
         );
  INV_X1 U11239 ( .A(n8749), .ZN(n8750) );
  OAI21_X1 U11240 ( .B1(n14447), .B2(n8868), .A(n8750), .ZN(n14138) );
  INV_X1 U11241 ( .A(n14138), .ZN(n14066) );
  NAND2_X1 U11242 ( .A1(n14632), .A2(n14066), .ZN(n8751) );
  NAND2_X1 U11243 ( .A1(n14421), .A2(n8751), .ZN(n14440) );
  INV_X1 U11244 ( .A(n14440), .ZN(n14442) );
  OR2_X1 U11245 ( .A1(n9367), .A2(n9829), .ZN(n8752) );
  XNOR2_X1 U11246 ( .A(n8752), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14657) );
  INV_X1 U11247 ( .A(n14628), .ZN(n14091) );
  OR2_X1 U11248 ( .A1(n8753), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8755) );
  AND2_X1 U11249 ( .A1(n8755), .A2(n8754), .ZN(n14429) );
  NAND2_X1 U11250 ( .A1(n14429), .A2(n8437), .ZN(n8761) );
  INV_X1 U11251 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11252 ( .A1(n6645), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U11253 ( .A1(n12478), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8756) );
  OAI211_X1 U11254 ( .C1(n12481), .C2(n8758), .A(n8757), .B(n8756), .ZN(n8759)
         );
  INV_X1 U11255 ( .A(n8759), .ZN(n8760) );
  NAND2_X1 U11256 ( .A1(n8761), .A2(n8760), .ZN(n14137) );
  XNOR2_X1 U11257 ( .A(n14091), .B(n14137), .ZN(n14430) );
  NAND2_X1 U11258 ( .A1(n14431), .A2(n14430), .ZN(n14433) );
  OR2_X1 U11259 ( .A1(n14628), .A2(n14137), .ZN(n8762) );
  XNOR2_X1 U11260 ( .A(n8763), .B(SI_23_), .ZN(n8764) );
  XNOR2_X1 U11261 ( .A(n8765), .B(n8764), .ZN(n11472) );
  NAND2_X1 U11262 ( .A1(n11472), .A2(n6643), .ZN(n8767) );
  INV_X1 U11263 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n15499) );
  OR2_X1 U11264 ( .A1(n12495), .A2(n15499), .ZN(n8766) );
  NAND2_X1 U11265 ( .A1(n9755), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U11266 ( .A1(n12478), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8772) );
  OAI21_X1 U11267 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8769), .A(n8768), .ZN(
        n14408) );
  OR2_X1 U11268 ( .A1(n8868), .A2(n14408), .ZN(n8771) );
  NAND2_X1 U11269 ( .A1(n6645), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8770) );
  NAND4_X1 U11270 ( .A1(n8773), .A2(n8772), .A3(n8771), .A4(n8770), .ZN(n14136) );
  XNOR2_X1 U11271 ( .A(n14553), .B(n14136), .ZN(n14410) );
  NAND2_X1 U11272 ( .A1(n14553), .A2(n14136), .ZN(n8774) );
  XNOR2_X1 U11273 ( .A(n8776), .B(n8775), .ZN(n11630) );
  NAND2_X1 U11274 ( .A1(n11630), .A2(n6643), .ZN(n8778) );
  INV_X1 U11275 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11634) );
  OR2_X1 U11276 ( .A1(n12495), .A2(n11634), .ZN(n8777) );
  NAND2_X1 U11277 ( .A1(n12478), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8785) );
  INV_X1 U11278 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15437) );
  OR2_X1 U11279 ( .A1(n12481), .A2(n15437), .ZN(n8784) );
  OAI21_X1 U11280 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8780), .A(n8779), .ZN(
        n14398) );
  OR2_X1 U11281 ( .A1(n8868), .A2(n14398), .ZN(n8783) );
  INV_X1 U11282 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14399) );
  OR2_X1 U11283 ( .A1(n8781), .A2(n14399), .ZN(n8782) );
  NAND4_X1 U11284 ( .A1(n8785), .A2(n8784), .A3(n8783), .A4(n8782), .ZN(n14135) );
  INV_X1 U11285 ( .A(n14135), .ZN(n13977) );
  OR2_X1 U11286 ( .A1(n14623), .A2(n13977), .ZN(n8864) );
  NAND2_X1 U11287 ( .A1(n14623), .A2(n13977), .ZN(n8786) );
  NAND2_X1 U11288 ( .A1(n8864), .A2(n8786), .ZN(n14385) );
  OR2_X1 U11289 ( .A1(n14623), .A2(n14135), .ZN(n8787) );
  NAND2_X1 U11290 ( .A1(n11719), .A2(n6643), .ZN(n8791) );
  OR2_X1 U11291 ( .A1(n12495), .A2(n11721), .ZN(n8790) );
  NAND2_X1 U11292 ( .A1(n9755), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11293 ( .A1(n12478), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8794) );
  XNOR2_X1 U11294 ( .A(P1_REG3_REG_25__SCAN_IN), .B(n8803), .ZN(n14372) );
  OR2_X1 U11295 ( .A1(n8868), .A2(n14372), .ZN(n8793) );
  NAND2_X1 U11296 ( .A1(n6645), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8792) );
  NAND4_X1 U11297 ( .A1(n8795), .A2(n8794), .A3(n8793), .A4(n8792), .ZN(n14134) );
  NAND2_X1 U11298 ( .A1(n14619), .A2(n14134), .ZN(n8797) );
  OR2_X1 U11299 ( .A1(n14619), .A2(n14134), .ZN(n8796) );
  NAND2_X1 U11300 ( .A1(n8797), .A2(n8796), .ZN(n12537) );
  XNOR2_X1 U11301 ( .A(n8798), .B(SI_26_), .ZN(n8799) );
  XNOR2_X1 U11302 ( .A(n8800), .B(n8799), .ZN(n11874) );
  NAND2_X1 U11303 ( .A1(n11874), .A2(n6643), .ZN(n8802) );
  OR2_X1 U11304 ( .A1(n12495), .A2(n15601), .ZN(n8801) );
  NAND2_X1 U11305 ( .A1(n6645), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8809) );
  INV_X1 U11306 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n15558) );
  OR2_X1 U11307 ( .A1(n12481), .A2(n15558), .ZN(n8808) );
  INV_X1 U11308 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n14536) );
  OR2_X1 U11309 ( .A1(n8453), .A2(n14536), .ZN(n8807) );
  INV_X1 U11310 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n15531) );
  NAND2_X1 U11311 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8803), .ZN(n8804) );
  NAND2_X1 U11312 ( .A1(n15531), .A2(n8804), .ZN(n8805) );
  NAND2_X1 U11313 ( .A1(n8814), .A2(n8805), .ZN(n14109) );
  OR2_X1 U11314 ( .A1(n8868), .A2(n14109), .ZN(n8806) );
  INV_X1 U11315 ( .A(n14361), .ZN(n8810) );
  NAND2_X1 U11316 ( .A1(n11965), .A2(n6643), .ZN(n8813) );
  OR2_X1 U11317 ( .A1(n12495), .A2(n11966), .ZN(n8812) );
  INV_X1 U11318 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15449) );
  OR2_X1 U11319 ( .A1(n12481), .A2(n15449), .ZN(n8820) );
  NAND2_X1 U11320 ( .A1(n8443), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8819) );
  INV_X1 U11321 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n15574) );
  NAND2_X1 U11322 ( .A1(n8814), .A2(n15574), .ZN(n8815) );
  NAND2_X1 U11323 ( .A1(n8816), .A2(n8815), .ZN(n14348) );
  OR2_X1 U11324 ( .A1(n8868), .A2(n14348), .ZN(n8818) );
  NAND2_X1 U11325 ( .A1(n6645), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8817) );
  NAND4_X1 U11326 ( .A1(n8820), .A2(n8819), .A3(n8818), .A4(n8817), .ZN(n14132) );
  INV_X1 U11327 ( .A(n14132), .ZN(n8821) );
  NAND2_X1 U11328 ( .A1(n8831), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8829) );
  NAND2_X1 U11329 ( .A1(n12297), .A2(n12489), .ZN(n12501) );
  NAND2_X1 U11330 ( .A1(n12297), .A2(n14301), .ZN(n8833) );
  NAND2_X1 U11331 ( .A1(n8874), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8830) );
  MUX2_X1 U11332 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8830), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8832) );
  NAND2_X1 U11333 ( .A1(n12501), .A2(n12212), .ZN(n14895) );
  OR2_X1 U11334 ( .A1(n11414), .A2(n12498), .ZN(n11306) );
  OR2_X1 U11335 ( .A1(n11414), .A2(n14301), .ZN(n8834) );
  INV_X1 U11336 ( .A(n14974), .ZN(n14982) );
  INV_X1 U11337 ( .A(n12372), .ZN(n12373) );
  NAND2_X1 U11338 ( .A1(n14510), .A2(n14514), .ZN(n14511) );
  INV_X1 U11339 ( .A(n14570), .ZN(n12204) );
  NOR2_X2 U11340 ( .A1(n14351), .A2(n14356), .ZN(n14347) );
  NOR2_X1 U11341 ( .A1(n12467), .A2(n14347), .ZN(n8835) );
  AND2_X2 U11342 ( .A1(n12467), .A2(n14347), .ZN(n9754) );
  OAI21_X1 U11343 ( .B1(n12467), .B2(n14982), .A(n14334), .ZN(n8836) );
  NAND2_X1 U11344 ( .A1(n8839), .A2(n12305), .ZN(n14891) );
  NAND2_X1 U11345 ( .A1(n14891), .A2(n14890), .ZN(n14889) );
  INV_X1 U11346 ( .A(n14969), .ZN(n12316) );
  OR2_X1 U11347 ( .A1(n14157), .A2(n12316), .ZN(n8840) );
  NAND2_X1 U11348 ( .A1(n14889), .A2(n8840), .ZN(n11343) );
  NAND2_X1 U11349 ( .A1(n11343), .A2(n12514), .ZN(n11342) );
  NAND2_X1 U11350 ( .A1(n12322), .A2(n14975), .ZN(n8841) );
  NAND2_X1 U11351 ( .A1(n11342), .A2(n8841), .ZN(n10581) );
  NAND2_X1 U11352 ( .A1(n11331), .A2(n14155), .ZN(n8842) );
  NAND2_X1 U11353 ( .A1(n10581), .A2(n8842), .ZN(n8844) );
  INV_X1 U11354 ( .A(n14155), .ZN(n10942) );
  NAND2_X1 U11355 ( .A1(n10942), .A2(n12327), .ZN(n8843) );
  NAND2_X1 U11356 ( .A1(n8844), .A2(n8843), .ZN(n10754) );
  NAND2_X1 U11357 ( .A1(n10754), .A2(n12518), .ZN(n8846) );
  INV_X1 U11358 ( .A(n14154), .ZN(n11143) );
  NAND2_X1 U11359 ( .A1(n12331), .A2(n11143), .ZN(n8845) );
  AND2_X1 U11360 ( .A1(n12342), .A2(n12341), .ZN(n8847) );
  INV_X1 U11361 ( .A(n12523), .ZN(n8848) );
  NAND2_X1 U11362 ( .A1(n11354), .A2(n8848), .ZN(n11358) );
  INV_X1 U11363 ( .A(n14150), .ZN(n12369) );
  NAND2_X1 U11364 ( .A1(n12368), .A2(n12369), .ZN(n8850) );
  NAND2_X1 U11365 ( .A1(n11526), .A2(n11525), .ZN(n11524) );
  OR2_X1 U11366 ( .A1(n12382), .A2(n12144), .ZN(n8852) );
  NAND2_X1 U11367 ( .A1(n11524), .A2(n8852), .ZN(n11621) );
  INV_X1 U11368 ( .A(n12529), .ZN(n11620) );
  NAND2_X1 U11369 ( .A1(n11621), .A2(n11620), .ZN(n11619) );
  NAND2_X1 U11370 ( .A1(n11619), .A2(n8853), .ZN(n11664) );
  NAND2_X1 U11371 ( .A1(n11664), .A2(n12402), .ZN(n11663) );
  NAND2_X1 U11372 ( .A1(n14039), .A2(n14046), .ZN(n8854) );
  XNOR2_X1 U11373 ( .A(n14587), .B(n12406), .ZN(n14502) );
  NAND2_X1 U11374 ( .A1(n14514), .A2(n14142), .ZN(n8856) );
  NAND2_X1 U11375 ( .A1(n14505), .A2(n8856), .ZN(n14489) );
  NAND2_X1 U11376 ( .A1(n14583), .A2(n14047), .ZN(n12430) );
  NAND2_X1 U11377 ( .A1(n14489), .A2(n14490), .ZN(n14478) );
  AND2_X1 U11378 ( .A1(n14468), .A2(n14479), .ZN(n8857) );
  NAND2_X1 U11379 ( .A1(n14478), .A2(n8857), .ZN(n14481) );
  NAND2_X1 U11380 ( .A1(n14481), .A2(n12431), .ZN(n14457) );
  INV_X1 U11381 ( .A(n14421), .ZN(n8859) );
  NOR2_X1 U11382 ( .A1(n14430), .A2(n8859), .ZN(n8860) );
  NAND2_X1 U11383 ( .A1(n14420), .A2(n8860), .ZN(n14423) );
  INV_X1 U11384 ( .A(n14137), .ZN(n13978) );
  NAND2_X1 U11385 ( .A1(n14628), .A2(n13978), .ZN(n8861) );
  NAND2_X1 U11386 ( .A1(n14423), .A2(n8861), .ZN(n14405) );
  INV_X1 U11387 ( .A(n14136), .ZN(n12227) );
  NAND2_X1 U11388 ( .A1(n14553), .A2(n12227), .ZN(n8862) );
  INV_X1 U11389 ( .A(n14134), .ZN(n12246) );
  NAND2_X1 U11390 ( .A1(n14619), .A2(n12246), .ZN(n8865) );
  NOR2_X1 U11391 ( .A1(n14616), .A2(n14133), .ZN(n8866) );
  NAND2_X1 U11392 ( .A1(n12489), .A2(n12509), .ZN(n12482) );
  OR2_X1 U11393 ( .A1(n12501), .A2(n11968), .ZN(n14065) );
  NAND2_X1 U11394 ( .A1(n9755), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U11395 ( .A1(n12478), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8871) );
  OR2_X1 U11396 ( .A1(n8868), .A2(n14318), .ZN(n8870) );
  NAND2_X1 U11397 ( .A1(n6645), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8869) );
  NAND4_X1 U11398 ( .A1(n8872), .A2(n8871), .A3(n8870), .A4(n8869), .ZN(n14130) );
  INV_X1 U11399 ( .A(n11968), .ZN(n14172) );
  OR2_X1 U11400 ( .A1(n12501), .A2(n14172), .ZN(n14095) );
  AOI22_X1 U11401 ( .A1(n14111), .A2(n14132), .B1(n14130), .B2(n14110), .ZN(
        n12281) );
  NAND2_X1 U11402 ( .A1(n8884), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8877) );
  MUX2_X1 U11403 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8877), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8880) );
  INV_X1 U11404 ( .A(n8884), .ZN(n8879) );
  NAND2_X1 U11405 ( .A1(n8879), .A2(n8878), .ZN(n8889) );
  NAND2_X1 U11406 ( .A1(n8880), .A2(n8889), .ZN(n11720) );
  NAND2_X1 U11407 ( .A1(n11720), .A2(P1_B_REG_SCAN_IN), .ZN(n8888) );
  INV_X1 U11408 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U11409 ( .A1(n8908), .A2(n8881), .ZN(n8911) );
  NAND2_X1 U11410 ( .A1(n8911), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8883) );
  MUX2_X1 U11411 ( .A(n8888), .B(P1_B_REG_SCAN_IN), .S(n11633), .Z(n8895) );
  NAND2_X1 U11412 ( .A1(n8889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11413 ( .A1(n8890), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11414 ( .A1(n8892), .A2(n8891), .ZN(n8894) );
  NAND2_X1 U11415 ( .A1(n8894), .A2(n8893), .ZN(n11875) );
  INV_X1 U11416 ( .A(n11875), .ZN(n8920) );
  NOR2_X1 U11417 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .ZN(
        n8899) );
  NOR4_X1 U11418 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n8898) );
  NOR4_X1 U11419 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8897) );
  NOR4_X1 U11420 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n8896) );
  AND4_X1 U11421 ( .A1(n8899), .A2(n8898), .A3(n8897), .A4(n8896), .ZN(n8905)
         );
  NOR4_X1 U11422 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n8903) );
  NOR4_X1 U11423 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n8902) );
  NOR4_X1 U11424 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8901) );
  NOR4_X1 U11425 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n8900) );
  AND4_X1 U11426 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), .ZN(n8904)
         );
  NAND2_X1 U11427 ( .A1(n8905), .A2(n8904), .ZN(n8906) );
  NAND2_X1 U11428 ( .A1(n10252), .A2(n8906), .ZN(n10332) );
  INV_X1 U11429 ( .A(n8908), .ZN(n8909) );
  NAND2_X1 U11430 ( .A1(n8909), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8910) );
  MUX2_X1 U11431 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8910), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8912) );
  NAND2_X1 U11432 ( .A1(n8912), .A2(n8911), .ZN(n10335) );
  NAND2_X1 U11433 ( .A1(n10335), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10257) );
  INV_X1 U11434 ( .A(n10257), .ZN(n8913) );
  NAND2_X1 U11435 ( .A1(n10332), .A2(n10342), .ZN(n10339) );
  AND2_X1 U11436 ( .A1(n12498), .A2(n14301), .ZN(n8914) );
  OR2_X1 U11437 ( .A1(n12501), .A2(n8914), .ZN(n10334) );
  INV_X1 U11438 ( .A(n10334), .ZN(n8915) );
  INV_X1 U11439 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U11440 ( .A1(n10252), .A2(n8916), .ZN(n8917) );
  NAND2_X1 U11441 ( .A1(n11875), .A2(n11720), .ZN(n10256) );
  NAND2_X1 U11442 ( .A1(n8917), .A2(n10256), .ZN(n11302) );
  NAND2_X1 U11443 ( .A1(n14901), .A2(n8918), .ZN(n10340) );
  AND2_X1 U11444 ( .A1(n11302), .A2(n10340), .ZN(n8919) );
  INV_X1 U11445 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8921) );
  NOR2_X1 U11446 ( .A1(n11633), .A2(n8920), .ZN(n10253) );
  INV_X1 U11447 ( .A(n11303), .ZN(n8922) );
  INV_X1 U11448 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8923) );
  OR2_X1 U11449 ( .A1(n14987), .A2(n8923), .ZN(n8924) );
  NAND2_X1 U11450 ( .A1(n8925), .A2(n8924), .ZN(P1_U3524) );
  INV_X1 U11451 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8926) );
  INV_X1 U11452 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8933) );
  INV_X1 U11453 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8935) );
  INV_X1 U11454 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8936) );
  XNOR2_X2 U11455 ( .A(n8937), .B(n8936), .ZN(n8943) );
  NAND2_X1 U11456 ( .A1(n8938), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8940) );
  AND2_X4 U11457 ( .A1(n8943), .A2(n13951), .ZN(n9505) );
  INV_X1 U11458 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9973) );
  NOR2_X1 U11459 ( .A1(n8942), .A2(n6760), .ZN(n8947) );
  INV_X1 U11460 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9974) );
  INV_X1 U11461 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9978) );
  NAND3_X2 U11462 ( .A1(n8947), .A2(n8946), .A3(n8945), .ZN(n11972) );
  INV_X1 U11463 ( .A(n13962), .ZN(n9907) );
  NAND2_X1 U11464 ( .A1(n9829), .A2(SI_0_), .ZN(n8949) );
  XNOR2_X1 U11465 ( .A(n8949), .B(n8948), .ZN(n13961) );
  INV_X1 U11466 ( .A(n8953), .ZN(n8954) );
  MUX2_X1 U11467 ( .A(n9907), .B(n13961), .S(n8979), .Z(n15136) );
  NAND2_X1 U11468 ( .A1(n11972), .A2(n15136), .ZN(n11976) );
  NOR2_X2 U11469 ( .A1(n9253), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n9271) );
  NAND2_X1 U11470 ( .A1(n9271), .A2(n8960), .ZN(n9300) );
  XNOR2_X1 U11471 ( .A(n8961), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9511) );
  NOR2_X2 U11472 ( .A1(n9248), .A2(n8962), .ZN(n8966) );
  INV_X1 U11473 ( .A(n8966), .ZN(n8963) );
  NAND2_X1 U11474 ( .A1(n8963), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8965) );
  INV_X1 U11475 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8964) );
  XNOR2_X1 U11476 ( .A(n8965), .B(n8964), .ZN(n10906) );
  NAND2_X1 U11477 ( .A1(n9511), .A2(n10906), .ZN(n9512) );
  OR2_X1 U11478 ( .A1(n9512), .A2(n11135), .ZN(n15151) );
  OR2_X2 U11479 ( .A1(n9565), .A2(n13945), .ZN(n8970) );
  XNOR2_X2 U11480 ( .A(n8970), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9704) );
  INV_X2 U11481 ( .A(n9006), .ZN(n9515) );
  XNOR2_X1 U11482 ( .A(n11976), .B(n6646), .ZN(n8974) );
  AND2_X2 U11483 ( .A1(n8971), .A2(n9661), .ZN(n15126) );
  INV_X1 U11484 ( .A(n15126), .ZN(n9541) );
  NAND2_X1 U11485 ( .A1(n9541), .A2(n9793), .ZN(n8973) );
  NAND2_X1 U11486 ( .A1(n8974), .A2(n8973), .ZN(n8989) );
  INV_X1 U11487 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n15133) );
  NAND2_X1 U11488 ( .A1(n9262), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8977) );
  INV_X1 U11489 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9903) );
  OR2_X1 U11490 ( .A1(n9029), .A2(n9903), .ZN(n8975) );
  NAND2_X1 U11491 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n13962), .ZN(n8980) );
  MUX2_X1 U11492 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8980), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8984) );
  INV_X1 U11493 ( .A(n8982), .ZN(n8983) );
  NAND2_X1 U11494 ( .A1(n8984), .A2(n8983), .ZN(n9911) );
  INV_X1 U11495 ( .A(n9911), .ZN(n9931) );
  NAND2_X1 U11496 ( .A1(n9120), .A2(n9931), .ZN(n8985) );
  MUX2_X1 U11497 ( .A(n13606), .B(n15143), .S(n9006), .Z(n8990) );
  NAND2_X1 U11498 ( .A1(n8989), .A2(n8990), .ZN(n8988) );
  MUX2_X1 U11499 ( .A(n13606), .B(n15143), .S(n6735), .Z(n8987) );
  NAND2_X1 U11500 ( .A1(n8988), .A2(n8987), .ZN(n8994) );
  INV_X1 U11501 ( .A(n8989), .ZN(n8992) );
  INV_X1 U11502 ( .A(n8990), .ZN(n8991) );
  NAND2_X1 U11503 ( .A1(n8992), .A2(n8991), .ZN(n8993) );
  NAND2_X1 U11504 ( .A1(n8994), .A2(n8993), .ZN(n9009) );
  NAND2_X1 U11505 ( .A1(n9262), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8998) );
  INV_X1 U11506 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12043) );
  OR2_X1 U11507 ( .A1(n9482), .A2(n12043), .ZN(n8997) );
  INV_X1 U11508 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9934) );
  OR2_X1 U11509 ( .A1(n9029), .A2(n9934), .ZN(n8995) );
  OR2_X1 U11510 ( .A1(n9871), .A2(n9370), .ZN(n9005) );
  NOR2_X1 U11511 ( .A1(n8982), .A2(n13945), .ZN(n8999) );
  MUX2_X1 U11512 ( .A(n13945), .B(n8999), .S(P2_IR_REG_2__SCAN_IN), .Z(n9000)
         );
  INV_X1 U11513 ( .A(n9000), .ZN(n9003) );
  INV_X1 U11514 ( .A(n9017), .ZN(n9002) );
  NAND2_X1 U11515 ( .A1(n9003), .A2(n9002), .ZN(n9935) );
  MUX2_X1 U11516 ( .A(n15129), .B(n12047), .S(n6735), .Z(n9010) );
  NAND2_X1 U11517 ( .A1(n9009), .A2(n9010), .ZN(n9008) );
  MUX2_X1 U11518 ( .A(n12047), .B(n15129), .S(n9515), .Z(n9007) );
  INV_X1 U11519 ( .A(n9009), .ZN(n9012) );
  INV_X1 U11520 ( .A(n9010), .ZN(n9011) );
  NAND2_X1 U11521 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  NOR2_X1 U11522 ( .A1(n9017), .A2(n13945), .ZN(n9014) );
  MUX2_X1 U11523 ( .A(n13945), .B(n9014), .S(P2_IR_REG_3__SCAN_IN), .Z(n9015)
         );
  INV_X1 U11524 ( .A(n9015), .ZN(n9018) );
  NAND2_X1 U11525 ( .A1(n9017), .A2(n9016), .ZN(n9056) );
  NAND2_X1 U11526 ( .A1(n9018), .A2(n9056), .ZN(n10011) );
  INV_X1 U11527 ( .A(n9019), .ZN(n9020) );
  NAND2_X1 U11528 ( .A1(n9505), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9025) );
  INV_X1 U11529 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10603) );
  OR2_X1 U11530 ( .A1(n9029), .A2(n10603), .ZN(n9024) );
  INV_X1 U11531 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9021) );
  OR2_X1 U11532 ( .A1(n9506), .A2(n9021), .ZN(n9023) );
  OR2_X1 U11533 ( .A1(n9482), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9022) );
  MUX2_X1 U11534 ( .A(n15183), .B(n13605), .S(n9515), .Z(n9027) );
  MUX2_X1 U11535 ( .A(n13605), .B(n15183), .S(n9515), .Z(n9026) );
  NAND2_X1 U11536 ( .A1(n9505), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9034) );
  INV_X1 U11537 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9939) );
  OR2_X1 U11538 ( .A1(n9029), .A2(n9939), .ZN(n9033) );
  OAI21_X1 U11539 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9050), .ZN(n13544) );
  OR2_X1 U11540 ( .A1(n9482), .A2(n13544), .ZN(n9032) );
  INV_X1 U11541 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9030) );
  OR2_X1 U11542 ( .A1(n9506), .A2(n9030), .ZN(n9031) );
  NAND4_X1 U11543 ( .A1(n9034), .A2(n9033), .A3(n9032), .A4(n9031), .ZN(n13604) );
  OR2_X1 U11544 ( .A1(n9856), .A2(n9370), .ZN(n9039) );
  INV_X1 U11545 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U11546 ( .A1(n9056), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9036) );
  XNOR2_X1 U11547 ( .A(n9036), .B(n9035), .ZN(n15010) );
  INV_X1 U11548 ( .A(n9037), .ZN(n9038) );
  NAND2_X1 U11549 ( .A1(n9039), .A2(n9038), .ZN(n13543) );
  MUX2_X1 U11550 ( .A(n13604), .B(n13543), .S(n6735), .Z(n9043) );
  NAND2_X1 U11551 ( .A1(n9042), .A2(n9043), .ZN(n9041) );
  MUX2_X1 U11552 ( .A(n13543), .B(n13604), .S(n9515), .Z(n9040) );
  NAND2_X1 U11553 ( .A1(n9041), .A2(n9040), .ZN(n9047) );
  INV_X1 U11554 ( .A(n9042), .ZN(n9045) );
  INV_X1 U11555 ( .A(n9043), .ZN(n9044) );
  NAND2_X1 U11556 ( .A1(n9045), .A2(n9044), .ZN(n9046) );
  NAND2_X1 U11557 ( .A1(n9047), .A2(n9046), .ZN(n9067) );
  NAND2_X1 U11558 ( .A1(n9483), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9055) );
  INV_X1 U11559 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9048) );
  OR2_X1 U11560 ( .A1(n9487), .A2(n9048), .ZN(n9054) );
  INV_X1 U11561 ( .A(n9074), .ZN(n9076) );
  NAND2_X1 U11562 ( .A1(n9050), .A2(n9049), .ZN(n9051) );
  NAND2_X1 U11563 ( .A1(n9076), .A2(n9051), .ZN(n10764) );
  OR2_X1 U11564 ( .A1(n9482), .A2(n10764), .ZN(n9053) );
  INV_X1 U11565 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9922) );
  OR2_X1 U11566 ( .A1(n9506), .A2(n9922), .ZN(n9052) );
  NAND4_X1 U11567 ( .A1(n9055), .A2(n9054), .A3(n9053), .A4(n9052), .ZN(n13603) );
  NAND2_X1 U11568 ( .A1(n9840), .A2(n9501), .ZN(n9064) );
  INV_X1 U11569 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U11570 ( .A1(n9058), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9057) );
  MUX2_X1 U11571 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9057), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9061) );
  INV_X1 U11572 ( .A(n9058), .ZN(n9060) );
  INV_X1 U11573 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U11574 ( .A1(n9060), .A2(n9059), .ZN(n9096) );
  NAND2_X1 U11575 ( .A1(n9061), .A2(n9096), .ZN(n9941) );
  INV_X1 U11576 ( .A(n9062), .ZN(n9063) );
  NAND2_X1 U11577 ( .A1(n9064), .A2(n9063), .ZN(n15197) );
  INV_X1 U11578 ( .A(n9515), .ZN(n9180) );
  MUX2_X1 U11579 ( .A(n13603), .B(n15197), .S(n9180), .Z(n9068) );
  NAND2_X1 U11580 ( .A1(n9067), .A2(n9068), .ZN(n9066) );
  MUX2_X1 U11581 ( .A(n13603), .B(n15197), .S(n9515), .Z(n9065) );
  NAND2_X1 U11582 ( .A1(n9066), .A2(n9065), .ZN(n9072) );
  INV_X1 U11583 ( .A(n9067), .ZN(n9070) );
  INV_X1 U11584 ( .A(n9068), .ZN(n9069) );
  NAND2_X1 U11585 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  NAND2_X1 U11586 ( .A1(n9483), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9081) );
  INV_X1 U11587 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9073) );
  OR2_X1 U11588 ( .A1(n9487), .A2(n9073), .ZN(n9080) );
  INV_X1 U11589 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U11590 ( .A1(n9076), .A2(n9075), .ZN(n9077) );
  NAND2_X1 U11591 ( .A1(n9090), .A2(n9077), .ZN(n10635) );
  OR2_X1 U11592 ( .A1(n9482), .A2(n10635), .ZN(n9079) );
  INV_X1 U11593 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9923) );
  OR2_X1 U11594 ( .A1(n9506), .A2(n9923), .ZN(n9078) );
  NAND4_X1 U11595 ( .A1(n9081), .A2(n9080), .A3(n9079), .A4(n9078), .ZN(n13602) );
  NAND2_X1 U11596 ( .A1(n9096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9083) );
  INV_X1 U11597 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9082) );
  XNOR2_X1 U11598 ( .A(n9083), .B(n9082), .ZN(n9972) );
  INV_X1 U11599 ( .A(n9084), .ZN(n9085) );
  MUX2_X1 U11600 ( .A(n13602), .B(n10654), .S(n6735), .Z(n9087) );
  MUX2_X1 U11601 ( .A(n10654), .B(n13602), .S(n9515), .Z(n9086) );
  INV_X1 U11602 ( .A(n9087), .ZN(n9088) );
  NAND2_X1 U11603 ( .A1(n9505), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9095) );
  INV_X1 U11604 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n15115) );
  OR2_X1 U11605 ( .A1(n9029), .A2(n15115), .ZN(n9094) );
  NAND2_X1 U11606 ( .A1(n9090), .A2(n9089), .ZN(n9091) );
  NAND2_X1 U11607 ( .A1(n9112), .A2(n9091), .ZN(n15114) );
  OR2_X1 U11608 ( .A1(n9482), .A2(n15114), .ZN(n9093) );
  INV_X1 U11609 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9924) );
  OR2_X1 U11610 ( .A1(n9506), .A2(n9924), .ZN(n9092) );
  NAND4_X1 U11611 ( .A1(n9095), .A2(n9094), .A3(n9093), .A4(n9092), .ZN(n13601) );
  NAND2_X1 U11612 ( .A1(n9858), .A2(n9501), .ZN(n9102) );
  NAND2_X1 U11613 ( .A1(n9098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9097) );
  MUX2_X1 U11614 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9097), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n9099) );
  NAND2_X1 U11615 ( .A1(n9099), .A2(n9118), .ZN(n15037) );
  INV_X1 U11616 ( .A(n9100), .ZN(n9101) );
  INV_X1 U11617 ( .A(n9515), .ZN(n9528) );
  MUX2_X1 U11618 ( .A(n13601), .B(n15117), .S(n9528), .Z(n9106) );
  NAND2_X1 U11619 ( .A1(n9105), .A2(n9106), .ZN(n9104) );
  MUX2_X1 U11620 ( .A(n13601), .B(n15117), .S(n9515), .Z(n9103) );
  NAND2_X1 U11621 ( .A1(n9104), .A2(n9103), .ZN(n9110) );
  INV_X1 U11622 ( .A(n9105), .ZN(n9108) );
  INV_X1 U11623 ( .A(n9106), .ZN(n9107) );
  NAND2_X1 U11624 ( .A1(n9108), .A2(n9107), .ZN(n9109) );
  NAND2_X1 U11625 ( .A1(n9505), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9117) );
  INV_X1 U11626 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9946) );
  OR2_X1 U11627 ( .A1(n9029), .A2(n9946), .ZN(n9116) );
  NAND2_X1 U11628 ( .A1(n9112), .A2(n9111), .ZN(n9113) );
  NAND2_X1 U11629 ( .A1(n9127), .A2(n9113), .ZN(n11097) );
  OR2_X1 U11630 ( .A1(n9482), .A2(n11097), .ZN(n9115) );
  INV_X1 U11631 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9925) );
  OR2_X1 U11632 ( .A1(n9506), .A2(n9925), .ZN(n9114) );
  NAND4_X1 U11633 ( .A1(n9117), .A2(n9116), .A3(n9115), .A4(n9114), .ZN(n13600) );
  NAND2_X1 U11634 ( .A1(n9118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9119) );
  XNOR2_X1 U11635 ( .A(n9119), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U11636 ( .A1(n9502), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9947), .B2(
        n9120), .ZN(n9121) );
  MUX2_X1 U11637 ( .A(n13600), .B(n11099), .S(n9515), .Z(n9124) );
  MUX2_X1 U11638 ( .A(n13600), .B(n11099), .S(n9528), .Z(n9123) );
  INV_X1 U11639 ( .A(n9124), .ZN(n9125) );
  NAND2_X1 U11640 ( .A1(n9483), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9132) );
  INV_X1 U11641 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9126) );
  OR2_X1 U11642 ( .A1(n9487), .A2(n9126), .ZN(n9131) );
  INV_X1 U11643 ( .A(n9145), .ZN(n9147) );
  NAND2_X1 U11644 ( .A1(n9127), .A2(n12118), .ZN(n9128) );
  NAND2_X1 U11645 ( .A1(n9147), .A2(n9128), .ZN(n12119) );
  OR2_X1 U11646 ( .A1(n9482), .A2(n12119), .ZN(n9130) );
  INV_X1 U11647 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9926) );
  OR2_X1 U11648 ( .A1(n9506), .A2(n9926), .ZN(n9129) );
  NAND4_X1 U11649 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n13598) );
  NAND2_X1 U11650 ( .A1(n9875), .A2(n9501), .ZN(n9136) );
  OR2_X1 U11651 ( .A1(n8957), .A2(n13945), .ZN(n9133) );
  INV_X1 U11652 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9153) );
  XNOR2_X1 U11653 ( .A(n9133), .B(n9153), .ZN(n10260) );
  INV_X1 U11654 ( .A(n9134), .ZN(n9135) );
  MUX2_X1 U11655 ( .A(n13598), .B(n11033), .S(n9528), .Z(n9140) );
  NAND2_X1 U11656 ( .A1(n9139), .A2(n9140), .ZN(n9138) );
  MUX2_X1 U11657 ( .A(n13598), .B(n11033), .S(n6735), .Z(n9137) );
  NAND2_X1 U11658 ( .A1(n9138), .A2(n9137), .ZN(n9144) );
  INV_X1 U11659 ( .A(n9139), .ZN(n9142) );
  INV_X1 U11660 ( .A(n9140), .ZN(n9141) );
  NAND2_X1 U11661 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  NAND2_X1 U11662 ( .A1(n9144), .A2(n9143), .ZN(n9161) );
  NAND2_X1 U11663 ( .A1(n9505), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9152) );
  INV_X1 U11664 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10990) );
  OR2_X1 U11665 ( .A1(n9029), .A2(n10990), .ZN(n9151) );
  INV_X1 U11666 ( .A(n9167), .ZN(n9169) );
  INV_X1 U11667 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U11668 ( .A1(n9147), .A2(n9146), .ZN(n9148) );
  NAND2_X1 U11669 ( .A1(n9169), .A2(n9148), .ZN(n11083) );
  OR2_X1 U11670 ( .A1(n9482), .A2(n11083), .ZN(n9150) );
  INV_X1 U11671 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10261) );
  OR2_X1 U11672 ( .A1(n9506), .A2(n10261), .ZN(n9149) );
  NAND4_X1 U11673 ( .A1(n9152), .A2(n9151), .A3(n9150), .A4(n9149), .ZN(n13597) );
  NAND2_X1 U11674 ( .A1(n9886), .A2(n9501), .ZN(n9158) );
  INV_X1 U11675 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U11676 ( .A1(n8957), .A2(n9153), .ZN(n9175) );
  NAND2_X1 U11677 ( .A1(n9175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9155) );
  INV_X1 U11678 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9154) );
  XNOR2_X1 U11679 ( .A(n9155), .B(n9154), .ZN(n10375) );
  INV_X1 U11680 ( .A(n9156), .ZN(n9157) );
  MUX2_X1 U11681 ( .A(n13597), .B(n15213), .S(n9515), .Z(n9162) );
  NAND2_X1 U11682 ( .A1(n9161), .A2(n9162), .ZN(n9160) );
  MUX2_X1 U11683 ( .A(n13597), .B(n15213), .S(n9528), .Z(n9159) );
  NAND2_X1 U11684 ( .A1(n9160), .A2(n9159), .ZN(n9166) );
  INV_X1 U11685 ( .A(n9161), .ZN(n9164) );
  INV_X1 U11686 ( .A(n9162), .ZN(n9163) );
  NAND2_X1 U11687 ( .A1(n9164), .A2(n9163), .ZN(n9165) );
  NAND2_X1 U11688 ( .A1(n9505), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9174) );
  INV_X1 U11689 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10386) );
  OR2_X1 U11690 ( .A1(n9029), .A2(n10386), .ZN(n9173) );
  INV_X1 U11691 ( .A(n9183), .ZN(n9185) );
  INV_X1 U11692 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U11693 ( .A1(n9169), .A2(n9168), .ZN(n9170) );
  NAND2_X1 U11694 ( .A1(n9185), .A2(n9170), .ZN(n11019) );
  OR2_X1 U11695 ( .A1(n9482), .A2(n11019), .ZN(n9172) );
  INV_X1 U11696 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10379) );
  OR2_X1 U11697 ( .A1(n9506), .A2(n10379), .ZN(n9171) );
  NAND4_X1 U11698 ( .A1(n9174), .A2(n9173), .A3(n9172), .A4(n9171), .ZN(n13596) );
  NAND2_X1 U11699 ( .A1(n9914), .A2(n9501), .ZN(n9179) );
  NAND2_X1 U11700 ( .A1(n9192), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9176) );
  INV_X1 U11701 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9193) );
  XNOR2_X1 U11702 ( .A(n9176), .B(n9193), .ZN(n10834) );
  INV_X1 U11703 ( .A(n9177), .ZN(n9178) );
  MUX2_X1 U11704 ( .A(n13596), .B(n11200), .S(n9528), .Z(n9182) );
  MUX2_X1 U11705 ( .A(n13596), .B(n11200), .S(n9515), .Z(n9181) );
  NAND2_X1 U11706 ( .A1(n9505), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9191) );
  OR2_X1 U11707 ( .A1(n9029), .A2(n15546), .ZN(n9190) );
  INV_X1 U11708 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9184) );
  NAND2_X1 U11709 ( .A1(n9185), .A2(n9184), .ZN(n9186) );
  NAND2_X1 U11710 ( .A1(n9206), .A2(n9186), .ZN(n12574) );
  OR2_X1 U11711 ( .A1(n9482), .A2(n12574), .ZN(n9189) );
  INV_X1 U11712 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9187) );
  OR2_X1 U11713 ( .A1(n9506), .A2(n9187), .ZN(n9188) );
  NAND4_X1 U11714 ( .A1(n9191), .A2(n9190), .A3(n9189), .A4(n9188), .ZN(n13595) );
  NAND2_X1 U11715 ( .A1(n10053), .A2(n9501), .ZN(n9197) );
  INV_X1 U11716 ( .A(n9192), .ZN(n9194) );
  NAND2_X1 U11717 ( .A1(n9194), .A2(n9193), .ZN(n9213) );
  NAND2_X1 U11718 ( .A1(n9213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9195) );
  XNOR2_X1 U11719 ( .A(n9195), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U11720 ( .A1(n9502), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9120), 
        .B2(n11436), .ZN(n9196) );
  MUX2_X1 U11721 ( .A(n13595), .B(n14815), .S(n9515), .Z(n9201) );
  NAND2_X1 U11722 ( .A1(n9200), .A2(n9201), .ZN(n9199) );
  MUX2_X1 U11723 ( .A(n13595), .B(n14815), .S(n9528), .Z(n9198) );
  NAND2_X1 U11724 ( .A1(n9199), .A2(n9198), .ZN(n9205) );
  INV_X1 U11725 ( .A(n9200), .ZN(n9203) );
  INV_X1 U11726 ( .A(n9201), .ZN(n9202) );
  NAND2_X1 U11727 ( .A1(n9203), .A2(n9202), .ZN(n9204) );
  NAND2_X1 U11728 ( .A1(n9206), .A2(n14995), .ZN(n9207) );
  NAND2_X1 U11729 ( .A1(n9221), .A2(n9207), .ZN(n15008) );
  INV_X1 U11730 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11424) );
  OR2_X1 U11731 ( .A1(n9029), .A2(n11424), .ZN(n9208) );
  OAI21_X1 U11732 ( .B1(n9482), .B2(n15008), .A(n9208), .ZN(n9212) );
  INV_X1 U11733 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9210) );
  INV_X1 U11734 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11439) );
  OR2_X1 U11735 ( .A1(n9506), .A2(n11439), .ZN(n9209) );
  OAI21_X1 U11736 ( .B1(n9487), .B2(n9210), .A(n9209), .ZN(n9211) );
  NAND2_X1 U11737 ( .A1(n10078), .A2(n9501), .ZN(n9216) );
  NAND2_X1 U11738 ( .A1(n9229), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9214) );
  XNOR2_X1 U11739 ( .A(n9214), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15050) );
  AOI22_X1 U11740 ( .A1(n9502), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n15050), 
        .B2(n9120), .ZN(n9215) );
  MUX2_X1 U11741 ( .A(n13594), .B(n15005), .S(n9528), .Z(n9218) );
  MUX2_X1 U11742 ( .A(n13594), .B(n15005), .S(n6735), .Z(n9217) );
  INV_X1 U11743 ( .A(n9218), .ZN(n9219) );
  INV_X1 U11744 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11745 ( .A1(n9221), .A2(n9220), .ZN(n9222) );
  NAND2_X1 U11746 ( .A1(n9243), .A2(n9222), .ZN(n12129) );
  INV_X1 U11747 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9223) );
  OR2_X1 U11748 ( .A1(n9487), .A2(n9223), .ZN(n9226) );
  INV_X1 U11749 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9224) );
  OR2_X1 U11750 ( .A1(n9029), .A2(n9224), .ZN(n9225) );
  AND2_X1 U11751 ( .A1(n9226), .A2(n9225), .ZN(n9228) );
  INV_X1 U11752 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n15541) );
  OR2_X1 U11753 ( .A1(n9506), .A2(n15541), .ZN(n9227) );
  OAI211_X1 U11754 ( .C1(n12129), .C2(n9482), .A(n9228), .B(n9227), .ZN(n13593) );
  NAND2_X1 U11755 ( .A1(n10368), .A2(n9501), .ZN(n9232) );
  OAI21_X1 U11756 ( .B1(n9229), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9230) );
  XNOR2_X1 U11757 ( .A(n9230), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U11758 ( .A1(n11428), .A2(n9120), .B1(n9502), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n9231) );
  MUX2_X1 U11759 ( .A(n13593), .B(n11505), .S(n6735), .Z(n9236) );
  NAND2_X1 U11760 ( .A1(n9235), .A2(n9236), .ZN(n9234) );
  MUX2_X1 U11761 ( .A(n13593), .B(n11505), .S(n9528), .Z(n9233) );
  NAND2_X1 U11762 ( .A1(n9234), .A2(n9233), .ZN(n9240) );
  INV_X1 U11763 ( .A(n9235), .ZN(n9238) );
  INV_X1 U11764 ( .A(n9236), .ZN(n9237) );
  NAND2_X1 U11765 ( .A1(n9238), .A2(n9237), .ZN(n9239) );
  NAND2_X1 U11766 ( .A1(n9240), .A2(n9239), .ZN(n9267) );
  INV_X1 U11767 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9247) );
  INV_X1 U11768 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U11769 ( .A1(n9243), .A2(n9242), .ZN(n9244) );
  NAND2_X1 U11770 ( .A1(n9260), .A2(n9244), .ZN(n11800) );
  OR2_X1 U11771 ( .A1(n11800), .A2(n9482), .ZN(n9246) );
  AOI22_X1 U11772 ( .A1(n9505), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n9483), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n9245) );
  OAI211_X1 U11773 ( .C1(n9506), .C2(n9247), .A(n9246), .B(n9245), .ZN(n13592)
         );
  NAND2_X1 U11774 ( .A1(n10394), .A2(n9501), .ZN(n9252) );
  NAND2_X1 U11775 ( .A1(n9248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9249) );
  XNOR2_X1 U11776 ( .A(n9249), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15073) );
  INV_X1 U11777 ( .A(n15073), .ZN(n11442) );
  INV_X1 U11778 ( .A(n9250), .ZN(n9251) );
  MUX2_X1 U11779 ( .A(n13592), .B(n13918), .S(n9180), .Z(n9268) );
  NAND2_X1 U11780 ( .A1(n9267), .A2(n9268), .ZN(n9266) );
  NAND2_X1 U11781 ( .A1(n10325), .A2(n9501), .ZN(n9258) );
  NAND2_X1 U11782 ( .A1(n9253), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9255) );
  INV_X1 U11783 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9254) );
  XNOR2_X1 U11784 ( .A(n9255), .B(n9254), .ZN(n13627) );
  INV_X1 U11785 ( .A(n9256), .ZN(n9257) );
  INV_X1 U11786 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U11787 ( .A1(n9260), .A2(n9259), .ZN(n9261) );
  NAND2_X1 U11788 ( .A1(n9277), .A2(n9261), .ZN(n11811) );
  AOI22_X1 U11789 ( .A1(n9505), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n9483), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U11790 ( .A1(n9262), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9263) );
  OAI211_X1 U11791 ( .C1(n11811), .C2(n9482), .A(n9264), .B(n9263), .ZN(n13591) );
  XNOR2_X1 U11792 ( .A(n13911), .B(n13591), .ZN(n9688) );
  MUX2_X1 U11793 ( .A(n13592), .B(n13918), .S(n9515), .Z(n9265) );
  INV_X1 U11794 ( .A(n9267), .ZN(n9270) );
  INV_X1 U11795 ( .A(n9268), .ZN(n9269) );
  NAND2_X1 U11796 ( .A1(n9270), .A2(n7656), .ZN(n9288) );
  NAND2_X1 U11797 ( .A1(n10398), .A2(n9501), .ZN(n9274) );
  OR2_X1 U11798 ( .A1(n9271), .A2(n13945), .ZN(n9272) );
  XNOR2_X1 U11799 ( .A(n9272), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15088) );
  AOI22_X1 U11800 ( .A1(n9502), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9120), 
        .B2(n15088), .ZN(n9273) );
  INV_X1 U11801 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11802 ( .A1(n9277), .A2(n9276), .ZN(n9278) );
  NAND2_X1 U11803 ( .A1(n9293), .A2(n9278), .ZN(n13828) );
  OR2_X1 U11804 ( .A1(n13828), .A2(n9482), .ZN(n9283) );
  INV_X1 U11805 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13829) );
  NAND2_X1 U11806 ( .A1(n9505), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9280) );
  INV_X1 U11807 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13629) );
  OR2_X1 U11808 ( .A1(n9506), .A2(n13629), .ZN(n9279) );
  OAI211_X1 U11809 ( .C1(n9029), .C2(n13829), .A(n9280), .B(n9279), .ZN(n9281)
         );
  INV_X1 U11810 ( .A(n9281), .ZN(n9282) );
  OR2_X1 U11811 ( .A1(n13907), .A2(n13568), .ZN(n9620) );
  NAND2_X1 U11812 ( .A1(n13907), .A2(n13568), .ZN(n9618) );
  AND2_X1 U11813 ( .A1(n13591), .A2(n9528), .ZN(n9285) );
  OAI21_X1 U11814 ( .B1(n9528), .B2(n13591), .A(n13911), .ZN(n9284) );
  OAI21_X1 U11815 ( .B1(n9285), .B2(n13911), .A(n9284), .ZN(n9286) );
  AND3_X1 U11816 ( .A1(n9620), .A2(n9618), .A3(n9286), .ZN(n9287) );
  NAND2_X1 U11817 ( .A1(n9288), .A2(n9287), .ZN(n9290) );
  MUX2_X1 U11818 ( .A(n9618), .B(n9620), .S(n6646), .Z(n9289) );
  INV_X1 U11819 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U11820 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  NAND2_X1 U11821 ( .A1(n9310), .A2(n9294), .ZN(n13815) );
  OR2_X1 U11822 ( .A1(n13815), .A2(n9482), .ZN(n9299) );
  INV_X1 U11823 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13816) );
  NAND2_X1 U11824 ( .A1(n9505), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U11825 ( .A1(n9262), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9295) );
  OAI211_X1 U11826 ( .C1(n9029), .C2(n13816), .A(n9296), .B(n9295), .ZN(n9297)
         );
  INV_X1 U11827 ( .A(n9297), .ZN(n9298) );
  NAND2_X1 U11828 ( .A1(n9300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9301) );
  XNOR2_X1 U11829 ( .A(n9301), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13631) );
  AOI22_X1 U11830 ( .A1(n9502), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n13631), 
        .B2(n9120), .ZN(n9302) );
  MUX2_X1 U11831 ( .A(n13488), .B(n13814), .S(n9515), .Z(n9305) );
  INV_X1 U11832 ( .A(n13488), .ZN(n13589) );
  MUX2_X1 U11833 ( .A(n13589), .B(n13902), .S(n9180), .Z(n9304) );
  OAI21_X1 U11834 ( .B1(n9306), .B2(n9305), .A(n9304), .ZN(n9308) );
  NAND2_X1 U11835 ( .A1(n9306), .A2(n9305), .ZN(n9307) );
  NAND2_X1 U11836 ( .A1(n9308), .A2(n9307), .ZN(n9320) );
  INV_X1 U11837 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11838 ( .A1(n9310), .A2(n9309), .ZN(n9311) );
  NAND2_X1 U11839 ( .A1(n9340), .A2(n9311), .ZN(n13796) );
  INV_X1 U11840 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n15561) );
  NAND2_X1 U11841 ( .A1(n9262), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U11842 ( .A1(n9483), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9312) );
  OAI211_X1 U11843 ( .C1(n9487), .C2(n15561), .A(n9313), .B(n9312), .ZN(n9314)
         );
  INV_X1 U11844 ( .A(n9314), .ZN(n9315) );
  OAI21_X1 U11845 ( .B1(n13796), .B2(n9482), .A(n9315), .ZN(n13588) );
  NAND2_X1 U11846 ( .A1(n10973), .A2(n9501), .ZN(n9317) );
  AOI22_X1 U11847 ( .A1(n13638), .A2(n9120), .B1(n9502), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n9316) );
  MUX2_X1 U11848 ( .A(n13588), .B(n13896), .S(n9180), .Z(n9321) );
  NAND2_X1 U11849 ( .A1(n9320), .A2(n9321), .ZN(n9319) );
  MUX2_X1 U11850 ( .A(n13588), .B(n13896), .S(n9515), .Z(n9318) );
  NAND2_X1 U11851 ( .A1(n9319), .A2(n9318), .ZN(n9325) );
  INV_X1 U11852 ( .A(n9320), .ZN(n9323) );
  INV_X1 U11853 ( .A(n9321), .ZN(n9322) );
  NAND2_X1 U11854 ( .A1(n9323), .A2(n9322), .ZN(n9324) );
  XNOR2_X1 U11855 ( .A(n9340), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13557) );
  NAND2_X1 U11856 ( .A1(n13557), .A2(n9429), .ZN(n9331) );
  INV_X1 U11857 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U11858 ( .A1(n9262), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U11859 ( .A1(n9483), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9326) );
  OAI211_X1 U11860 ( .C1(n9487), .C2(n9328), .A(n9327), .B(n9326), .ZN(n9329)
         );
  INV_X1 U11861 ( .A(n9329), .ZN(n9330) );
  NAND2_X1 U11862 ( .A1(n9331), .A2(n9330), .ZN(n13587) );
  NAND2_X1 U11863 ( .A1(n9502), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9332) );
  MUX2_X1 U11864 ( .A(n13587), .B(n13891), .S(n6735), .Z(n9335) );
  MUX2_X1 U11865 ( .A(n13587), .B(n13891), .S(n9528), .Z(n9334) );
  AND2_X1 U11866 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n9336) );
  INV_X1 U11867 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9339) );
  INV_X1 U11868 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9338) );
  OAI21_X1 U11869 ( .B1(n9340), .B2(n9339), .A(n9338), .ZN(n9341) );
  AND2_X1 U11870 ( .A1(n9359), .A2(n9341), .ZN(n13766) );
  NAND2_X1 U11871 ( .A1(n13766), .A2(n9429), .ZN(n9346) );
  INV_X1 U11872 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13769) );
  NAND2_X1 U11873 ( .A1(n9505), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U11874 ( .A1(n9262), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9342) );
  OAI211_X1 U11875 ( .C1(n9029), .C2(n13769), .A(n9343), .B(n9342), .ZN(n9344)
         );
  INV_X1 U11876 ( .A(n9344), .ZN(n9345) );
  NAND2_X1 U11877 ( .A1(n9346), .A2(n9345), .ZN(n13586) );
  NAND2_X1 U11878 ( .A1(n9502), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9347) );
  MUX2_X1 U11879 ( .A(n13586), .B(n13886), .S(n9180), .Z(n9352) );
  NAND2_X1 U11880 ( .A1(n9351), .A2(n9352), .ZN(n9350) );
  MUX2_X1 U11881 ( .A(n13586), .B(n13886), .S(n6735), .Z(n9349) );
  NAND2_X1 U11882 ( .A1(n9350), .A2(n9349), .ZN(n9356) );
  INV_X1 U11883 ( .A(n9351), .ZN(n9354) );
  INV_X1 U11884 ( .A(n9352), .ZN(n9353) );
  NAND2_X1 U11885 ( .A1(n9354), .A2(n9353), .ZN(n9355) );
  INV_X1 U11886 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11887 ( .A1(n9359), .A2(n9358), .ZN(n9360) );
  NAND2_X1 U11888 ( .A1(n9375), .A2(n9360), .ZN(n13750) );
  OR2_X1 U11889 ( .A1(n13750), .A2(n9482), .ZN(n9365) );
  INV_X1 U11890 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13751) );
  NAND2_X1 U11891 ( .A1(n9505), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U11892 ( .A1(n9262), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9361) );
  OAI211_X1 U11893 ( .C1(n9029), .C2(n13751), .A(n9362), .B(n9361), .ZN(n9363)
         );
  INV_X1 U11894 ( .A(n9363), .ZN(n9364) );
  NAND2_X1 U11895 ( .A1(n9365), .A2(n9364), .ZN(n13585) );
  NAND2_X1 U11896 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  NAND2_X1 U11897 ( .A1(n9369), .A2(n9368), .ZN(n11389) );
  NAND2_X1 U11898 ( .A1(n9502), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9371) );
  MUX2_X1 U11899 ( .A(n13585), .B(n13881), .S(n6646), .Z(n9374) );
  MUX2_X1 U11900 ( .A(n13585), .B(n13881), .S(n9528), .Z(n9373) );
  INV_X1 U11901 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13484) );
  NAND2_X1 U11902 ( .A1(n9375), .A2(n13484), .ZN(n9376) );
  AND2_X1 U11903 ( .A1(n9394), .A2(n9376), .ZN(n13736) );
  NAND2_X1 U11904 ( .A1(n13736), .A2(n9429), .ZN(n9382) );
  INV_X1 U11905 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9379) );
  NAND2_X1 U11906 ( .A1(n9262), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U11907 ( .A1(n9483), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9377) );
  OAI211_X1 U11908 ( .C1(n9487), .C2(n9379), .A(n9378), .B(n9377), .ZN(n9380)
         );
  INV_X1 U11909 ( .A(n9380), .ZN(n9381) );
  NAND2_X1 U11910 ( .A1(n9382), .A2(n9381), .ZN(n13584) );
  NAND2_X1 U11911 ( .A1(n11472), .A2(n9501), .ZN(n9384) );
  NAND2_X1 U11912 ( .A1(n9502), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9383) );
  MUX2_X1 U11913 ( .A(n13584), .B(n13876), .S(n9180), .Z(n9388) );
  NAND2_X1 U11914 ( .A1(n9387), .A2(n9388), .ZN(n9386) );
  MUX2_X1 U11915 ( .A(n13584), .B(n13876), .S(n6646), .Z(n9385) );
  NAND2_X1 U11916 ( .A1(n9386), .A2(n9385), .ZN(n9392) );
  INV_X1 U11917 ( .A(n9387), .ZN(n9390) );
  INV_X1 U11918 ( .A(n9388), .ZN(n9389) );
  NAND2_X1 U11919 ( .A1(n9390), .A2(n9389), .ZN(n9391) );
  INV_X1 U11920 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13535) );
  NAND2_X1 U11921 ( .A1(n9394), .A2(n13535), .ZN(n9395) );
  NAND2_X1 U11922 ( .A1(n9407), .A2(n9395), .ZN(n13534) );
  INV_X1 U11923 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n15589) );
  NAND2_X1 U11924 ( .A1(n9505), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U11925 ( .A1(n9483), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9396) );
  OAI211_X1 U11926 ( .C1(n15589), .C2(n9506), .A(n9397), .B(n9396), .ZN(n9398)
         );
  INV_X1 U11927 ( .A(n9398), .ZN(n9399) );
  NAND2_X1 U11928 ( .A1(n11630), .A2(n9501), .ZN(n9402) );
  NAND2_X1 U11929 ( .A1(n9502), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9401) );
  MUX2_X1 U11930 ( .A(n13583), .B(n13871), .S(n6735), .Z(n9404) );
  MUX2_X1 U11931 ( .A(n13583), .B(n13871), .S(n9528), .Z(n9403) );
  INV_X1 U11932 ( .A(n9404), .ZN(n9405) );
  INV_X1 U11933 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U11934 ( .A1(n9407), .A2(n13527), .ZN(n9408) );
  NAND2_X1 U11935 ( .A1(n13708), .A2(n9429), .ZN(n9413) );
  INV_X1 U11936 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n15431) );
  NAND2_X1 U11937 ( .A1(n9483), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9410) );
  NAND2_X1 U11938 ( .A1(n9262), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9409) );
  OAI211_X1 U11939 ( .C1(n9487), .C2(n15431), .A(n9410), .B(n9409), .ZN(n9411)
         );
  INV_X1 U11940 ( .A(n9411), .ZN(n9412) );
  NAND2_X1 U11941 ( .A1(n11719), .A2(n9501), .ZN(n9415) );
  NAND2_X1 U11942 ( .A1(n9502), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9414) );
  MUX2_X1 U11943 ( .A(n13582), .B(n13866), .S(n9180), .Z(n9427) );
  INV_X1 U11944 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n12018) );
  NAND2_X1 U11945 ( .A1(n9416), .A2(n12018), .ZN(n9417) );
  NAND2_X1 U11946 ( .A1(n13692), .A2(n9429), .ZN(n9423) );
  INV_X1 U11947 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9420) );
  NAND2_X1 U11948 ( .A1(n9262), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9419) );
  NAND2_X1 U11949 ( .A1(n9483), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9418) );
  OAI211_X1 U11950 ( .C1(n9487), .C2(n9420), .A(n9419), .B(n9418), .ZN(n9421)
         );
  INV_X1 U11951 ( .A(n9421), .ZN(n9422) );
  NAND2_X1 U11952 ( .A1(n11874), .A2(n9501), .ZN(n9425) );
  NAND2_X1 U11953 ( .A1(n9502), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9424) );
  MUX2_X1 U11954 ( .A(n13526), .B(n13694), .S(n9515), .Z(n9438) );
  MUX2_X1 U11955 ( .A(n13581), .B(n13861), .S(n9180), .Z(n9437) );
  OAI22_X1 U11956 ( .A1(n9428), .A2(n9427), .B1(n9438), .B2(n9437), .ZN(n9443)
         );
  INV_X1 U11957 ( .A(n13582), .ZN(n12011) );
  INV_X1 U11958 ( .A(n13866), .ZN(n13711) );
  MUX2_X1 U11959 ( .A(n12011), .B(n13711), .S(n6735), .Z(n9426) );
  AOI21_X1 U11960 ( .B1(n9428), .B2(n9427), .A(n9426), .ZN(n9442) );
  XNOR2_X1 U11961 ( .A(n9471), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13676) );
  NAND2_X1 U11962 ( .A1(n13676), .A2(n9429), .ZN(n9434) );
  INV_X1 U11963 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n15560) );
  NAND2_X1 U11964 ( .A1(n9505), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U11965 ( .A1(n9483), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9430) );
  OAI211_X1 U11966 ( .C1(n9506), .C2(n15560), .A(n9431), .B(n9430), .ZN(n9432)
         );
  INV_X1 U11967 ( .A(n9432), .ZN(n9433) );
  INV_X1 U11968 ( .A(n12036), .ZN(n13580) );
  NAND2_X1 U11969 ( .A1(n11965), .A2(n9501), .ZN(n9436) );
  NAND2_X1 U11970 ( .A1(n9502), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9435) );
  MUX2_X1 U11971 ( .A(n13580), .B(n13857), .S(n6646), .Z(n9480) );
  INV_X1 U11972 ( .A(n9480), .ZN(n9440) );
  MUX2_X1 U11973 ( .A(n12036), .B(n13678), .S(n9528), .Z(n9481) );
  INV_X1 U11974 ( .A(n9481), .ZN(n9439) );
  AOI22_X1 U11975 ( .A1(n9440), .A2(n9439), .B1(n9438), .B2(n9437), .ZN(n9441)
         );
  INV_X1 U11976 ( .A(n9447), .ZN(n9449) );
  INV_X1 U11977 ( .A(SI_27_), .ZN(n11638) );
  NAND2_X1 U11978 ( .A1(n9448), .A2(SI_28_), .ZN(n9444) );
  OAI21_X1 U11979 ( .B1(n9449), .B2(n11638), .A(n9444), .ZN(n9445) );
  OAI21_X1 U11980 ( .B1(n9447), .B2(SI_27_), .A(SI_28_), .ZN(n9452) );
  INV_X1 U11981 ( .A(n9448), .ZN(n9451) );
  NOR2_X1 U11982 ( .A1(SI_27_), .A2(SI_28_), .ZN(n9450) );
  AOI22_X1 U11983 ( .A1(n9452), .A2(n9451), .B1(n9450), .B2(n9449), .ZN(n9453)
         );
  INV_X1 U11984 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14656) );
  INV_X1 U11985 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13950) );
  MUX2_X1 U11986 ( .A(n14656), .B(n13950), .S(n9829), .Z(n9454) );
  XNOR2_X1 U11987 ( .A(n9454), .B(SI_29_), .ZN(n9491) );
  INV_X1 U11988 ( .A(SI_29_), .ZN(n11962) );
  NAND2_X1 U11989 ( .A1(n9454), .A2(n11962), .ZN(n9455) );
  MUX2_X1 U11990 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9829), .Z(n9457) );
  NAND2_X1 U11991 ( .A1(n9457), .A2(SI_30_), .ZN(n9460) );
  INV_X1 U11992 ( .A(n9457), .ZN(n9458) );
  INV_X1 U11993 ( .A(SI_30_), .ZN(n11959) );
  NAND2_X1 U11994 ( .A1(n9458), .A2(n11959), .ZN(n9459) );
  NAND2_X1 U11995 ( .A1(n9460), .A2(n9459), .ZN(n9498) );
  MUX2_X1 U11996 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9829), .Z(n9461) );
  XNOR2_X1 U11997 ( .A(n9461), .B(SI_31_), .ZN(n9462) );
  NAND2_X1 U11998 ( .A1(n13944), .A2(n9501), .ZN(n9465) );
  NAND2_X1 U11999 ( .A1(n9502), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9464) );
  INV_X1 U12000 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U12001 ( .A1(n9483), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U12002 ( .A1(n9262), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9466) );
  OAI211_X1 U12003 ( .C1(n9487), .C2(n9468), .A(n9467), .B(n9466), .ZN(n13646)
         );
  INV_X1 U12004 ( .A(n9471), .ZN(n9470) );
  AND2_X1 U12005 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n9469) );
  NAND2_X1 U12006 ( .A1(n9470), .A2(n9469), .ZN(n9711) );
  INV_X1 U12007 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13474) );
  INV_X1 U12008 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12039) );
  OAI21_X1 U12009 ( .B1(n9471), .B2(n13474), .A(n12039), .ZN(n9472) );
  NAND2_X1 U12010 ( .A1(n9711), .A2(n9472), .ZN(n13661) );
  INV_X1 U12011 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U12012 ( .A1(n9262), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U12013 ( .A1(n9483), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9473) );
  OAI211_X1 U12014 ( .C1(n9487), .C2(n9475), .A(n9474), .B(n9473), .ZN(n9476)
         );
  INV_X1 U12015 ( .A(n9476), .ZN(n9477) );
  NAND2_X1 U12016 ( .A1(n9502), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9479) );
  MUX2_X1 U12017 ( .A(n13473), .B(n13851), .S(n9528), .Z(n9520) );
  MUX2_X1 U12018 ( .A(n13579), .B(n9701), .S(n9515), .Z(n9519) );
  NAND2_X1 U12019 ( .A1(n9520), .A2(n9519), .ZN(n9496) );
  NAND2_X1 U12020 ( .A1(n9481), .A2(n9480), .ZN(n9495) );
  OR2_X1 U12021 ( .A1(n9711), .A2(n9482), .ZN(n9490) );
  INV_X1 U12022 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U12023 ( .A1(n9483), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U12024 ( .A1(n9262), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9484) );
  OAI211_X1 U12025 ( .C1(n9487), .C2(n9486), .A(n9485), .B(n9484), .ZN(n9488)
         );
  INV_X1 U12026 ( .A(n9488), .ZN(n9489) );
  AND2_X1 U12027 ( .A1(n9490), .A2(n9489), .ZN(n12038) );
  NAND2_X1 U12028 ( .A1(n13949), .A2(n9501), .ZN(n9494) );
  NAND2_X1 U12029 ( .A1(n9502), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U12030 ( .A(n12038), .B(n9714), .S(n9180), .Z(n9517) );
  MUX2_X1 U12031 ( .A(n13578), .B(n13845), .S(n9515), .Z(n9516) );
  NAND2_X1 U12032 ( .A1(n9517), .A2(n9516), .ZN(n9521) );
  NAND2_X1 U12033 ( .A1(n12484), .A2(n9501), .ZN(n9504) );
  NAND2_X1 U12034 ( .A1(n9502), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9503) );
  INV_X1 U12035 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9509) );
  NAND2_X1 U12036 ( .A1(n9505), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9508) );
  INV_X1 U12037 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n15603) );
  OR2_X1 U12038 ( .A1(n9506), .A2(n15603), .ZN(n9507) );
  OAI211_X1 U12039 ( .C1(n9029), .C2(n9509), .A(n9508), .B(n9507), .ZN(n13577)
         );
  NAND2_X1 U12040 ( .A1(n9515), .A2(n13646), .ZN(n9513) );
  NAND2_X1 U12041 ( .A1(n10975), .A2(n10906), .ZN(n9816) );
  INV_X1 U12042 ( .A(n9704), .ZN(n11390) );
  OR2_X1 U12043 ( .A1(n9659), .A2(n11390), .ZN(n9533) );
  NAND4_X1 U12044 ( .A1(n9513), .A2(n9510), .A3(n9816), .A4(n9533), .ZN(n9514)
         );
  AOI22_X1 U12045 ( .A1(n13643), .A2(n9528), .B1(n13577), .B2(n9514), .ZN(
        n9526) );
  MUX2_X1 U12046 ( .A(n13577), .B(n13643), .S(n6735), .Z(n9525) );
  OAI22_X1 U12047 ( .A1(n9526), .A2(n9525), .B1(n9517), .B2(n9516), .ZN(n9518)
         );
  NAND2_X1 U12048 ( .A1(n9518), .A2(n9540), .ZN(n9524) );
  INV_X1 U12049 ( .A(n9519), .ZN(n9523) );
  INV_X1 U12050 ( .A(n9520), .ZN(n9522) );
  NAND2_X1 U12051 ( .A1(n9526), .A2(n9525), .ZN(n9532) );
  INV_X1 U12052 ( .A(n13646), .ZN(n9527) );
  AND2_X1 U12053 ( .A1(n13648), .A2(n9527), .ZN(n9530) );
  NOR2_X1 U12054 ( .A1(n13648), .A2(n9527), .ZN(n9529) );
  MUX2_X1 U12055 ( .A(n9530), .B(n9529), .S(n9180), .Z(n9531) );
  INV_X1 U12056 ( .A(n10906), .ZN(n9710) );
  NAND2_X1 U12057 ( .A1(n9510), .A2(n9710), .ZN(n9634) );
  OAI21_X1 U12058 ( .B1(n10975), .B2(n9634), .A(n9533), .ZN(n9534) );
  INV_X1 U12059 ( .A(n9534), .ZN(n9539) );
  INV_X1 U12060 ( .A(n9793), .ZN(n9535) );
  NAND2_X1 U12061 ( .A1(n11390), .A2(n9535), .ZN(n9536) );
  AOI22_X1 U12062 ( .A1(n9536), .A2(n13638), .B1(n9710), .B2(n11135), .ZN(
        n9537) );
  NAND2_X1 U12063 ( .A1(n9564), .A2(n9537), .ZN(n9538) );
  OAI21_X1 U12064 ( .B1(n9564), .B2(n9539), .A(n9538), .ZN(n9569) );
  INV_X1 U12065 ( .A(n9659), .ZN(n15150) );
  INV_X1 U12066 ( .A(n9540), .ZN(n9561) );
  XNOR2_X1 U12067 ( .A(n13643), .B(n13577), .ZN(n9558) );
  NAND2_X1 U12068 ( .A1(n13861), .A2(n13526), .ZN(n9628) );
  NAND2_X1 U12069 ( .A1(n9627), .A2(n9628), .ZN(n13696) );
  XNOR2_X1 U12070 ( .A(n13871), .B(n13583), .ZN(n9626) );
  INV_X1 U12071 ( .A(n13586), .ZN(n13558) );
  XNOR2_X1 U12072 ( .A(n13886), .B(n13558), .ZN(n13770) );
  XNOR2_X1 U12073 ( .A(n13891), .B(n13513), .ZN(n13778) );
  INV_X1 U12074 ( .A(n13588), .ZN(n13569) );
  XNOR2_X1 U12075 ( .A(n13896), .B(n13569), .ZN(n13800) );
  XNOR2_X1 U12076 ( .A(n13902), .B(n13488), .ZN(n13809) );
  XNOR2_X1 U12077 ( .A(n13907), .B(n13568), .ZN(n9690) );
  INV_X1 U12078 ( .A(n13593), .ZN(n11513) );
  XNOR2_X1 U12079 ( .A(n11505), .B(n11513), .ZN(n11597) );
  INV_X1 U12080 ( .A(n13594), .ZN(n12131) );
  OR2_X1 U12081 ( .A1(n15005), .A2(n12131), .ZN(n9610) );
  NAND2_X1 U12082 ( .A1(n15005), .A2(n12131), .ZN(n9611) );
  AND2_X1 U12083 ( .A1(n9610), .A2(n9611), .ZN(n11265) );
  INV_X1 U12084 ( .A(n13596), .ZN(n11176) );
  XNOR2_X1 U12085 ( .A(n11200), .B(n11176), .ZN(n11168) );
  INV_X1 U12086 ( .A(n13597), .ZN(n9604) );
  XNOR2_X1 U12087 ( .A(n15213), .B(n9604), .ZN(n10981) );
  INV_X1 U12088 ( .A(n13598), .ZN(n9603) );
  XNOR2_X1 U12089 ( .A(n11033), .B(n9603), .ZN(n9676) );
  INV_X1 U12090 ( .A(n13601), .ZN(n9599) );
  XNOR2_X1 U12091 ( .A(n15117), .B(n9599), .ZN(n10821) );
  XNOR2_X1 U12092 ( .A(n11099), .B(n13600), .ZN(n11091) );
  INV_X1 U12093 ( .A(n13604), .ZN(n9668) );
  XNOR2_X1 U12094 ( .A(n13543), .B(n9668), .ZN(n9667) );
  NAND2_X1 U12095 ( .A1(n9541), .A2(n11976), .ZN(n15170) );
  NOR2_X1 U12096 ( .A1(n15170), .A2(n10906), .ZN(n9545) );
  INV_X1 U12097 ( .A(n9543), .ZN(n9542) );
  NAND2_X1 U12098 ( .A1(n9542), .A2(n15143), .ZN(n9591) );
  INV_X1 U12099 ( .A(n15143), .ZN(n15175) );
  NAND2_X1 U12100 ( .A1(n9543), .A2(n15175), .ZN(n9544) );
  NAND4_X1 U12101 ( .A1(n9545), .A2(n15138), .A3(n10598), .A4(n10065), .ZN(
        n9546) );
  NOR2_X1 U12102 ( .A1(n9667), .A2(n9546), .ZN(n9547) );
  XNOR2_X1 U12103 ( .A(n15197), .B(n13603), .ZN(n10607) );
  XNOR2_X1 U12104 ( .A(n10654), .B(n13602), .ZN(n10639) );
  NAND4_X1 U12105 ( .A1(n11091), .A2(n9547), .A3(n10607), .A4(n10639), .ZN(
        n9548) );
  OR4_X1 U12106 ( .A1(n10981), .A2(n9676), .A3(n10821), .A4(n9548), .ZN(n9549)
         );
  NOR2_X1 U12107 ( .A1(n11168), .A2(n9549), .ZN(n9550) );
  XNOR2_X1 U12108 ( .A(n14815), .B(n13595), .ZN(n9607) );
  NAND4_X1 U12109 ( .A1(n9688), .A2(n11265), .A3(n9550), .A4(n9607), .ZN(n9552) );
  INV_X1 U12110 ( .A(n13592), .ZN(n11691) );
  NAND2_X1 U12111 ( .A1(n13918), .A2(n11691), .ZN(n9551) );
  NAND2_X1 U12112 ( .A1(n9616), .A2(n9551), .ZN(n11804) );
  OR4_X1 U12113 ( .A1(n9690), .A2(n11597), .A3(n9552), .A4(n11804), .ZN(n9553)
         );
  OR4_X1 U12114 ( .A1(n13778), .A2(n13800), .A3(n13809), .A4(n9553), .ZN(n9554) );
  NOR2_X1 U12115 ( .A1(n13770), .A2(n9554), .ZN(n9555) );
  OR2_X1 U12116 ( .A1(n13876), .A2(n13584), .ZN(n9695) );
  NAND2_X1 U12117 ( .A1(n13876), .A2(n13584), .ZN(n9697) );
  NAND2_X1 U12118 ( .A1(n9695), .A2(n9697), .ZN(n13733) );
  NAND4_X1 U12119 ( .A1(n9626), .A2(n9555), .A3(n13733), .A4(n13748), .ZN(
        n9556) );
  NOR2_X1 U12120 ( .A1(n13696), .A2(n9556), .ZN(n9557) );
  XNOR2_X1 U12121 ( .A(n13866), .B(n13582), .ZN(n13703) );
  NAND4_X1 U12122 ( .A1(n9558), .A2(n9557), .A3(n9702), .A4(n13703), .ZN(n9560) );
  NAND2_X1 U12123 ( .A1(n9701), .A2(n13473), .ZN(n9559) );
  NOR4_X1 U12124 ( .A1(n9561), .A2(n9560), .A3(n13656), .A4(n9630), .ZN(n9562)
         );
  XNOR2_X1 U12125 ( .A(n9562), .B(n13638), .ZN(n9563) );
  INV_X1 U12126 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U12127 ( .A1(n9570), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9576) );
  INV_X1 U12128 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9575) );
  XNOR2_X1 U12129 ( .A(n9576), .B(n9575), .ZN(n9890) );
  OR2_X1 U12130 ( .A1(n9890), .A2(P2_U3088), .ZN(n11450) );
  INV_X1 U12131 ( .A(n11450), .ZN(n9567) );
  OAI21_X1 U12132 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9590) );
  INV_X1 U12133 ( .A(n9570), .ZN(n9572) );
  NOR2_X1 U12134 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n9571) );
  NAND2_X1 U12135 ( .A1(n9572), .A2(n9571), .ZN(n9580) );
  NAND2_X1 U12136 ( .A1(n9582), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9573) );
  MUX2_X1 U12137 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9573), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9574) );
  NAND2_X1 U12138 ( .A1(n9574), .A2(n8956), .ZN(n11878) );
  INV_X1 U12139 ( .A(n11878), .ZN(n9653) );
  NAND2_X1 U12140 ( .A1(n9576), .A2(n9575), .ZN(n9577) );
  NAND2_X1 U12141 ( .A1(n9577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9579) );
  INV_X1 U12142 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9578) );
  XNOR2_X1 U12143 ( .A(n9579), .B(n9578), .ZN(n11632) );
  NAND2_X1 U12144 ( .A1(n9580), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9581) );
  MUX2_X1 U12145 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9581), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9583) );
  NAND2_X1 U12146 ( .A1(n9583), .A2(n9582), .ZN(n11722) );
  NOR2_X1 U12147 ( .A1(n11632), .A2(n11722), .ZN(n9584) );
  NAND2_X1 U12148 ( .A1(n9653), .A2(n9584), .ZN(n9786) );
  INV_X1 U12149 ( .A(n15166), .ZN(n15163) );
  INV_X1 U12150 ( .A(n9585), .ZN(n9586) );
  NAND2_X1 U12151 ( .A1(n9891), .A2(n9586), .ZN(n13567) );
  NOR4_X1 U12152 ( .A1(n15163), .A2(n13957), .A3(n9816), .A4(n13567), .ZN(
        n9588) );
  OAI21_X1 U12153 ( .B1(n11450), .B2(n9704), .A(P2_B_REG_SCAN_IN), .ZN(n9587)
         );
  OR2_X1 U12154 ( .A1(n9588), .A2(n9587), .ZN(n9589) );
  NAND2_X1 U12155 ( .A1(n9590), .A2(n9589), .ZN(P2_U3328) );
  INV_X1 U12156 ( .A(n15129), .ZN(n9592) );
  NAND2_X1 U12157 ( .A1(n9592), .A2(n12047), .ZN(n9593) );
  NAND2_X1 U12158 ( .A1(n10599), .A2(n10598), .ZN(n9595) );
  INV_X1 U12159 ( .A(n13605), .ZN(n10861) );
  NAND2_X1 U12160 ( .A1(n10861), .A2(n15183), .ZN(n9594) );
  NAND2_X1 U12161 ( .A1(n9595), .A2(n9594), .ZN(n10859) );
  INV_X1 U12162 ( .A(n9667), .ZN(n10858) );
  NAND2_X1 U12163 ( .A1(n13543), .A2(n9668), .ZN(n9596) );
  INV_X1 U12164 ( .A(n13603), .ZN(n10860) );
  OR2_X1 U12165 ( .A1(n15197), .A2(n10860), .ZN(n9597) );
  NAND2_X1 U12166 ( .A1(n15197), .A2(n10860), .ZN(n9598) );
  INV_X1 U12167 ( .A(n13602), .ZN(n10537) );
  AND2_X1 U12168 ( .A1(n15117), .A2(n9599), .ZN(n9600) );
  OAI22_X1 U12169 ( .A1(n10820), .A2(n9600), .B1(n9599), .B2(n15117), .ZN(
        n11102) );
  INV_X1 U12170 ( .A(n13600), .ZN(n12114) );
  OR2_X1 U12171 ( .A1(n11099), .A2(n12114), .ZN(n9601) );
  INV_X1 U12172 ( .A(n9676), .ZN(n10894) );
  INV_X1 U12173 ( .A(n10981), .ZN(n10978) );
  OR2_X1 U12174 ( .A1(n15213), .A2(n9604), .ZN(n9605) );
  NAND2_X1 U12175 ( .A1(n11200), .A2(n11176), .ZN(n9606) );
  INV_X1 U12176 ( .A(n13595), .ZN(n11022) );
  OR2_X1 U12177 ( .A1(n14815), .A2(n11022), .ZN(n9609) );
  INV_X1 U12178 ( .A(n9611), .ZN(n9612) );
  NAND2_X1 U12179 ( .A1(n11505), .A2(n11513), .ZN(n9613) );
  INV_X1 U12180 ( .A(n11804), .ZN(n9615) );
  INV_X1 U12181 ( .A(n13591), .ZN(n12286) );
  INV_X1 U12182 ( .A(n13911), .ZN(n9617) );
  INV_X1 U12183 ( .A(n9618), .ZN(n9619) );
  INV_X1 U12184 ( .A(n13896), .ZN(n13799) );
  INV_X1 U12185 ( .A(n13891), .ZN(n9693) );
  OAI22_X1 U12186 ( .A1(n13775), .A2(n13778), .B1(n9693), .B2(n13587), .ZN(
        n13761) );
  NOR2_X1 U12187 ( .A1(n7485), .A2(n13586), .ZN(n9623) );
  INV_X1 U12188 ( .A(n13881), .ZN(n9624) );
  INV_X1 U12189 ( .A(n13876), .ZN(n13739) );
  NAND2_X1 U12190 ( .A1(n13739), .A2(n13584), .ZN(n9625) );
  INV_X1 U12191 ( .A(n13584), .ZN(n13480) );
  INV_X1 U12192 ( .A(n13871), .ZN(n13725) );
  INV_X1 U12193 ( .A(n9627), .ZN(n9629) );
  INV_X1 U12194 ( .A(n13656), .ZN(n13666) );
  NAND2_X1 U12195 ( .A1(n13857), .A2(n12036), .ZN(n13667) );
  XNOR2_X1 U12196 ( .A(n9633), .B(n9632), .ZN(n9640) );
  NAND2_X1 U12197 ( .A1(n13638), .A2(n9704), .ZN(n9635) );
  INV_X2 U12198 ( .A(n11793), .ZN(n15131) );
  NAND2_X1 U12199 ( .A1(n13579), .A2(n15127), .ZN(n9638) );
  NAND2_X1 U12200 ( .A1(n9891), .A2(n9585), .ZN(n15148) );
  INV_X1 U12201 ( .A(P2_B_REG_SCAN_IN), .ZN(n9650) );
  NOR2_X1 U12202 ( .A1(n13957), .A2(n9650), .ZN(n9636) );
  NOR2_X1 U12203 ( .A1(n15148), .A2(n9636), .ZN(n13647) );
  NAND2_X1 U12204 ( .A1(n13647), .A2(n13577), .ZN(n9637) );
  NOR4_X1 U12205 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n9649) );
  OR4_X1 U12206 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9646) );
  NOR4_X1 U12207 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n9644) );
  NOR4_X1 U12208 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n9643) );
  NOR4_X1 U12209 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9642) );
  NOR4_X1 U12210 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9641) );
  NAND4_X1 U12211 ( .A1(n9644), .A2(n9643), .A3(n9642), .A4(n9641), .ZN(n9645)
         );
  NOR4_X1 U12212 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n9646), .A4(n9645), .ZN(n9648) );
  NOR4_X1 U12213 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n9647) );
  NAND3_X1 U12214 ( .A1(n9649), .A2(n9648), .A3(n9647), .ZN(n9654) );
  XOR2_X1 U12215 ( .A(n11632), .B(n9650), .Z(n9651) );
  NAND2_X1 U12216 ( .A1(n11722), .A2(n9651), .ZN(n9652) );
  AND2_X1 U12217 ( .A1(n9654), .A2(n15158), .ZN(n10075) );
  INV_X1 U12218 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15164) );
  NAND2_X1 U12219 ( .A1(n15158), .A2(n15164), .ZN(n9656) );
  NAND2_X1 U12220 ( .A1(n11878), .A2(n11722), .ZN(n9655) );
  NAND2_X1 U12221 ( .A1(n9656), .A2(n9655), .ZN(n15165) );
  NOR2_X1 U12222 ( .A1(n10075), .A2(n15165), .ZN(n9788) );
  NAND2_X1 U12223 ( .A1(n9816), .A2(n9891), .ZN(n9789) );
  INV_X1 U12224 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15161) );
  NAND2_X1 U12225 ( .A1(n15158), .A2(n15161), .ZN(n9658) );
  NAND2_X1 U12226 ( .A1(n11878), .A2(n11632), .ZN(n9657) );
  NAND2_X1 U12227 ( .A1(n9658), .A2(n9657), .ZN(n15162) );
  NAND3_X1 U12228 ( .A1(n9788), .A2(n11970), .A3(n15162), .ZN(n9660) );
  NAND2_X1 U12229 ( .A1(n15218), .A2(n11135), .ZN(n10659) );
  INV_X1 U12230 ( .A(n10659), .ZN(n10073) );
  NAND2_X2 U12231 ( .A1(n9660), .A2(n15132), .ZN(n15155) );
  INV_X2 U12232 ( .A(n15155), .ZN(n15157) );
  INV_X1 U12233 ( .A(n13568), .ZN(n13590) );
  INV_X1 U12234 ( .A(n10065), .ZN(n10060) );
  NAND2_X1 U12235 ( .A1(n11972), .A2(n9661), .ZN(n15137) );
  INV_X1 U12236 ( .A(n15137), .ZN(n13499) );
  OAI22_X1 U12237 ( .A1(n15138), .A2(n13499), .B1(n13606), .B2(n15143), .ZN(
        n10061) );
  NAND2_X1 U12238 ( .A1(n10060), .A2(n10061), .ZN(n9663) );
  OR2_X1 U12239 ( .A1(n12047), .A2(n15129), .ZN(n9662) );
  NAND2_X1 U12240 ( .A1(n9663), .A2(n9662), .ZN(n10593) );
  INV_X1 U12241 ( .A(n10598), .ZN(n9664) );
  NAND2_X1 U12242 ( .A1(n10593), .A2(n9664), .ZN(n9666) );
  OR2_X1 U12243 ( .A1(n15183), .A2(n13605), .ZN(n9665) );
  NAND2_X1 U12244 ( .A1(n9666), .A2(n9665), .ZN(n10856) );
  INV_X1 U12245 ( .A(n13543), .ZN(n15191) );
  NAND2_X1 U12246 ( .A1(n15191), .A2(n9668), .ZN(n9669) );
  NAND2_X1 U12247 ( .A1(n15197), .A2(n13603), .ZN(n9670) );
  NAND2_X1 U12248 ( .A1(n9672), .A2(n9671), .ZN(n10630) );
  OR2_X1 U12249 ( .A1(n10654), .A2(n13602), .ZN(n9673) );
  NAND2_X1 U12250 ( .A1(n10630), .A2(n9673), .ZN(n10819) );
  NAND2_X1 U12251 ( .A1(n10819), .A2(n10821), .ZN(n10818) );
  INV_X1 U12252 ( .A(n11091), .ZN(n11101) );
  OR2_X1 U12253 ( .A1(n15117), .A2(n13601), .ZN(n11090) );
  AND2_X1 U12254 ( .A1(n11101), .A2(n11090), .ZN(n9674) );
  NAND2_X1 U12255 ( .A1(n10818), .A2(n9674), .ZN(n11094) );
  NAND2_X1 U12256 ( .A1(n11099), .A2(n13600), .ZN(n9675) );
  NAND2_X1 U12257 ( .A1(n11094), .A2(n9675), .ZN(n10892) );
  NAND2_X1 U12258 ( .A1(n10892), .A2(n9676), .ZN(n9678) );
  NAND2_X1 U12259 ( .A1(n11033), .A2(n13598), .ZN(n9677) );
  NAND2_X1 U12260 ( .A1(n9678), .A2(n9677), .ZN(n10979) );
  NAND2_X1 U12261 ( .A1(n15213), .A2(n13597), .ZN(n9679) );
  AND2_X1 U12262 ( .A1(n11200), .A2(n13596), .ZN(n9680) );
  OR2_X1 U12263 ( .A1(n11200), .A2(n13596), .ZN(n9681) );
  NAND2_X1 U12264 ( .A1(n9682), .A2(n9681), .ZN(n11173) );
  NOR2_X1 U12265 ( .A1(n14815), .A2(n13595), .ZN(n9683) );
  OR2_X1 U12266 ( .A1(n15005), .A2(n13594), .ZN(n9684) );
  NAND2_X1 U12267 ( .A1(n15005), .A2(n13594), .ZN(n9685) );
  OR2_X1 U12268 ( .A1(n11505), .A2(n13593), .ZN(n9686) );
  NOR2_X1 U12269 ( .A1(n13918), .A2(n13592), .ZN(n9687) );
  NAND2_X1 U12270 ( .A1(n13814), .A2(n13488), .ZN(n9691) );
  NOR2_X1 U12271 ( .A1(n13896), .A2(n13588), .ZN(n9692) );
  INV_X1 U12272 ( .A(n13770), .ZN(n13760) );
  INV_X1 U12273 ( .A(n9695), .ZN(n9696) );
  AOI22_X1 U12274 ( .A1(n13720), .A2(n13719), .B1(n13871), .B2(n13583), .ZN(
        n13704) );
  INV_X1 U12275 ( .A(n13704), .ZN(n9699) );
  XNOR2_X1 U12276 ( .A(n9703), .B(n9702), .ZN(n13848) );
  NAND2_X1 U12277 ( .A1(n15201), .A2(n6875), .ZN(n9706) );
  INV_X1 U12278 ( .A(n15005), .ZN(n14811) );
  INV_X1 U12279 ( .A(n11099), .ZN(n15208) );
  INV_X1 U12280 ( .A(n10654), .ZN(n10636) );
  NOR2_X1 U12281 ( .A1(n9661), .A2(n15143), .ZN(n10062) );
  INV_X1 U12282 ( .A(n12047), .ZN(n10645) );
  AND2_X1 U12283 ( .A1(n10062), .A2(n10645), .ZN(n10594) );
  INV_X1 U12284 ( .A(n15183), .ZN(n10596) );
  NAND2_X1 U12285 ( .A1(n15208), .A2(n11096), .ZN(n11095) );
  INV_X1 U12286 ( .A(n11200), .ZN(n9707) );
  NAND2_X1 U12287 ( .A1(n14811), .A2(n11267), .ZN(n11592) );
  NAND2_X1 U12288 ( .A1(n7485), .A2(n13785), .ZN(n13765) );
  NAND2_X1 U12289 ( .A1(n11390), .A2(n11135), .ZN(n9709) );
  OR2_X2 U12290 ( .A1(n9709), .A2(n9710), .ZN(n9794) );
  INV_X1 U12291 ( .A(n9709), .ZN(n15149) );
  AND2_X1 U12292 ( .A1(n15149), .A2(n9710), .ZN(n9818) );
  INV_X1 U12293 ( .A(n9711), .ZN(n9712) );
  INV_X1 U12294 ( .A(n15132), .ZN(n15154) );
  AOI22_X1 U12295 ( .A1(n9712), .A2(n15154), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n15157), .ZN(n9713) );
  OAI21_X1 U12296 ( .B1(n9714), .B2(n13813), .A(n9713), .ZN(n9715) );
  AOI21_X1 U12297 ( .B1(n13844), .B2(n13835), .A(n9715), .ZN(n9716) );
  OAI21_X1 U12298 ( .B1(n13847), .B2(n15157), .A(n9718), .ZN(P2_U3236) );
  INV_X1 U12299 ( .A(n9719), .ZN(n9721) );
  NAND2_X1 U12300 ( .A1(n13353), .A2(n6908), .ZN(n9720) );
  NAND2_X1 U12301 ( .A1(n9721), .A2(n9720), .ZN(n9726) );
  XNOR2_X1 U12302 ( .A(n14656), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n11952) );
  XNOR2_X1 U12303 ( .A(n11954), .B(n11952), .ZN(n11961) );
  NAND2_X1 U12304 ( .A1(n11961), .A2(n12601), .ZN(n9725) );
  NAND2_X1 U12305 ( .A1(n12602), .A2(SI_29_), .ZN(n9724) );
  NAND2_X1 U12306 ( .A1(n9725), .A2(n9724), .ZN(n9742) );
  NAND2_X1 U12307 ( .A1(n9742), .A2(n12909), .ZN(n12754) );
  NAND2_X1 U12308 ( .A1(n12763), .A2(n12754), .ZN(n12749) );
  XNOR2_X1 U12309 ( .A(n9726), .B(n12749), .ZN(n9737) );
  INV_X1 U12310 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U12311 ( .A1(n8131), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U12312 ( .A1(n9727), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9728) );
  OAI211_X1 U12313 ( .C1(n7767), .C2(n9730), .A(n9729), .B(n9728), .ZN(n9731)
         );
  INV_X1 U12314 ( .A(n9731), .ZN(n9732) );
  NAND2_X1 U12315 ( .A1(n10128), .A2(P3_B_REG_SCAN_IN), .ZN(n9733) );
  NAND2_X1 U12316 ( .A1(n15242), .A2(n9733), .ZN(n13172) );
  NOR2_X1 U12317 ( .A1(n12608), .A2(n13172), .ZN(n9734) );
  INV_X1 U12318 ( .A(n12750), .ZN(n9738) );
  NOR2_X2 U12319 ( .A1(n13183), .A2(n9741), .ZN(n9784) );
  INV_X1 U12320 ( .A(n9742), .ZN(n13181) );
  INV_X1 U12321 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9744) );
  NOR2_X1 U12322 ( .A1(n15309), .A2(n9744), .ZN(n9745) );
  NAND2_X1 U12323 ( .A1(n13949), .A2(n6643), .ZN(n9749) );
  OR2_X1 U12324 ( .A1(n12495), .A2(n14656), .ZN(n9748) );
  XNOR2_X1 U12325 ( .A(n12475), .B(n14130), .ZN(n12472) );
  INV_X1 U12326 ( .A(n12472), .ZN(n12540) );
  NOR2_X1 U12327 ( .A1(n12467), .A2(n14131), .ZN(n9751) );
  OAI22_X1 U12328 ( .A1(n9752), .A2(n9751), .B1(n13968), .B2(n14332), .ZN(
        n9753) );
  OAI211_X1 U12329 ( .C1(n9754), .C2(n14321), .A(n14901), .B(n14314), .ZN(
        n14325) );
  INV_X1 U12330 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n15557) );
  NAND2_X1 U12331 ( .A1(n6645), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U12332 ( .A1(n9755), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9756) );
  OAI211_X1 U12333 ( .C1(n8453), .C2(n15557), .A(n9757), .B(n9756), .ZN(n14129) );
  INV_X1 U12334 ( .A(P1_B_REG_SCAN_IN), .ZN(n9758) );
  NOR2_X1 U12335 ( .A1(n6734), .A2(n9758), .ZN(n9759) );
  NOR2_X1 U12336 ( .A1(n14095), .A2(n9759), .ZN(n14307) );
  NAND2_X1 U12337 ( .A1(n14129), .A2(n14307), .ZN(n14319) );
  NAND2_X1 U12338 ( .A1(n14325), .A2(n14319), .ZN(n9760) );
  INV_X1 U12339 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9762) );
  NAND2_X1 U12340 ( .A1(n9765), .A2(n14994), .ZN(n9770) );
  INV_X1 U12341 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9766) );
  OR2_X1 U12342 ( .A1(n14994), .A2(n9766), .ZN(n9767) );
  INV_X1 U12343 ( .A(n9768), .ZN(n9769) );
  NAND2_X1 U12344 ( .A1(n9770), .A2(n9769), .ZN(P1_U3557) );
  XNOR2_X1 U12345 ( .A(n10299), .B(n13458), .ZN(n9773) );
  AND2_X1 U12346 ( .A1(n9771), .A2(n10671), .ZN(n9772) );
  NAND2_X1 U12347 ( .A1(n8227), .A2(n9776), .ZN(n10233) );
  NAND2_X1 U12348 ( .A1(n12746), .A2(n9774), .ZN(n10664) );
  AND2_X1 U12349 ( .A1(n10233), .A2(n10664), .ZN(n10666) );
  OAI22_X1 U12350 ( .A1(n15295), .A2(n9775), .B1(n12613), .B2(n12617), .ZN(
        n9777) );
  AOI21_X1 U12351 ( .B1(n9777), .B2(n9776), .A(n8227), .ZN(n9779) );
  INV_X1 U12352 ( .A(n13458), .ZN(n9778) );
  MUX2_X1 U12353 ( .A(n10666), .B(n9779), .S(n9778), .Z(n9780) );
  OAI21_X1 U12354 ( .B1(n9784), .B2(n15696), .A(n9783), .ZN(P3_U3488) );
  INV_X1 U12355 ( .A(n9890), .ZN(n9785) );
  NOR2_X1 U12356 ( .A1(n9786), .A2(n9785), .ZN(n9893) );
  AND2_X1 U12357 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9893), .ZN(P2_U3947) );
  OR2_X2 U12358 ( .A1(n10348), .A2(n10257), .ZN(n14159) );
  INV_X1 U12359 ( .A(n13459), .ZN(n11949) );
  INV_X2 U12360 ( .A(n13060), .ZN(P3_U3897) );
  INV_X1 U12361 ( .A(n15162), .ZN(n9787) );
  NAND2_X1 U12362 ( .A1(n9788), .A2(n9787), .ZN(n9810) );
  NAND2_X1 U12363 ( .A1(n9810), .A2(n10659), .ZN(n11971) );
  AND2_X1 U12364 ( .A1(n9790), .A2(n9789), .ZN(n9791) );
  NAND2_X1 U12365 ( .A1(n11971), .A2(n9791), .ZN(n9792) );
  INV_X1 U12366 ( .A(n15007), .ZN(n13546) );
  MUX2_X1 U12367 ( .A(n13546), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n9823) );
  NAND2_X1 U12368 ( .A1(n13606), .A2(n9794), .ZN(n9797) );
  NAND2_X1 U12369 ( .A1(n15201), .A2(n9793), .ZN(n10516) );
  NAND2_X1 U12370 ( .A1(n10928), .A2(n15136), .ZN(n13503) );
  OAI21_X1 U12371 ( .B1(n15137), .B2(n15134), .A(n13503), .ZN(n9795) );
  NAND2_X1 U12372 ( .A1(n12048), .A2(n9797), .ZN(n9798) );
  NAND2_X1 U12373 ( .A1(n13502), .A2(n9798), .ZN(n9799) );
  XNOR2_X1 U12374 ( .A(n12033), .B(n12047), .ZN(n9800) );
  NAND2_X1 U12375 ( .A1(n15129), .A2(n9794), .ZN(n9801) );
  XNOR2_X1 U12376 ( .A(n9800), .B(n9801), .ZN(n12049) );
  NAND2_X1 U12377 ( .A1(n9799), .A2(n12049), .ZN(n12054) );
  INV_X1 U12378 ( .A(n9800), .ZN(n9802) );
  NAND2_X1 U12379 ( .A1(n9802), .A2(n9801), .ZN(n9803) );
  XNOR2_X1 U12380 ( .A(n10928), .B(n15183), .ZN(n13540) );
  NAND2_X1 U12381 ( .A1(n13605), .A2(n12009), .ZN(n9804) );
  NAND2_X1 U12382 ( .A1(n13540), .A2(n9804), .ZN(n9807) );
  INV_X1 U12383 ( .A(n13540), .ZN(n9806) );
  INV_X1 U12384 ( .A(n9804), .ZN(n9805) );
  NAND2_X1 U12385 ( .A1(n9806), .A2(n9805), .ZN(n10513) );
  NAND2_X1 U12386 ( .A1(n9807), .A2(n10513), .ZN(n9814) );
  INV_X1 U12387 ( .A(n9809), .ZN(n13549) );
  INV_X1 U12388 ( .A(n9810), .ZN(n9811) );
  NAND2_X1 U12389 ( .A1(n15149), .A2(n9816), .ZN(n15215) );
  INV_X1 U12390 ( .A(n9891), .ZN(n9812) );
  AND2_X1 U12391 ( .A1(n15215), .A2(n9812), .ZN(n9813) );
  NAND2_X2 U12392 ( .A1(n9819), .A2(n9813), .ZN(n14999) );
  AOI211_X1 U12393 ( .C1(n9815), .C2(n9814), .A(n9809), .B(n14999), .ZN(n9822)
         );
  INV_X1 U12394 ( .A(n15148), .ZN(n15128) );
  AOI22_X1 U12395 ( .A1(n15128), .A2(n13604), .B1(n15129), .B2(n15127), .ZN(
        n10600) );
  INV_X1 U12396 ( .A(n9819), .ZN(n9817) );
  NOR2_X2 U12397 ( .A1(n9817), .A2(n9816), .ZN(n13515) );
  INV_X1 U12398 ( .A(n13515), .ZN(n14997) );
  NAND2_X1 U12399 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  OAI22_X1 U12400 ( .A1(n10600), .A2(n14997), .B1(n13539), .B2(n10596), .ZN(
        n9821) );
  OR3_X1 U12401 ( .A1(n9823), .A2(n9822), .A3(n9821), .ZN(P2_U3190) );
  AND2_X1 U12402 ( .A1(n9829), .A2(P1_U3086), .ZN(n14651) );
  INV_X2 U12403 ( .A(n14651), .ZN(n12562) );
  AND2_X1 U12404 ( .A1(n9828), .A2(P1_U3086), .ZN(n11471) );
  OAI222_X1 U12405 ( .A1(n12562), .A2(n9824), .B1(n6656), .B2(n9871), .C1(
        P1_U3086), .C2(n14180), .ZN(P1_U3353) );
  OAI222_X1 U12406 ( .A1(P1_U3086), .A2(n10035), .B1(n6656), .B2(n9874), .C1(
        n8300), .C2(n12562), .ZN(P1_U3354) );
  INV_X1 U12407 ( .A(n9825), .ZN(n9863) );
  NOR2_X1 U12408 ( .A1(n9829), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13953) );
  INV_X2 U12409 ( .A(n13953), .ZN(n13960) );
  OAI222_X1 U12410 ( .A1(P2_U3088), .A2(n10011), .B1(n13955), .B2(n9863), .C1(
        n9826), .C2(n13960), .ZN(P2_U3324) );
  OAI222_X1 U12411 ( .A1(P2_U3088), .A2(n15010), .B1(n13955), .B2(n9856), .C1(
        n9827), .C2(n13960), .ZN(P2_U3323) );
  AND2_X1 U12412 ( .A1(n9828), .A2(P3_U3151), .ZN(n10995) );
  AND2_X1 U12413 ( .A1(n9829), .A2(P3_U3151), .ZN(n13465) );
  OAI222_X1 U12414 ( .A1(n6655), .A2(n9830), .B1(n12584), .B2(n7697), .C1(
        P3_U3151), .C2(n7699), .ZN(P3_U3294) );
  OAI222_X1 U12415 ( .A1(n10964), .A2(P3_U3151), .B1(n6655), .B2(n9832), .C1(
        n9831), .C2(n12584), .ZN(P3_U3286) );
  OAI222_X1 U12416 ( .A1(P3_U3151), .A2(n10147), .B1(n6655), .B2(n9834), .C1(
        n9833), .C2(n12584), .ZN(P3_U3292) );
  OAI222_X1 U12417 ( .A1(P3_U3151), .A2(n10477), .B1(n6655), .B2(n9836), .C1(
        n9835), .C2(n12584), .ZN(P3_U3289) );
  INV_X1 U12418 ( .A(n9837), .ZN(n9839) );
  OAI222_X1 U12419 ( .A1(P3_U3151), .A2(n7305), .B1(n6655), .B2(n9839), .C1(
        n9838), .C2(n12584), .ZN(P3_U3288) );
  INV_X1 U12420 ( .A(n9840), .ZN(n9842) );
  INV_X1 U12421 ( .A(n10042), .ZN(n10087) );
  OAI222_X1 U12422 ( .A1(n12562), .A2(n9841), .B1(n6656), .B2(n9842), .C1(
        P1_U3086), .C2(n10087), .ZN(P1_U3350) );
  OAI222_X1 U12423 ( .A1(n13960), .A2(n9843), .B1(n13955), .B2(n9842), .C1(
        P2_U3088), .C2(n9941), .ZN(P2_U3322) );
  OAI222_X1 U12424 ( .A1(P3_U3151), .A2(n10213), .B1(n12584), .B2(n9845), .C1(
        n6655), .C2(n9844), .ZN(P3_U3291) );
  OAI222_X1 U12425 ( .A1(P3_U3151), .A2(n10963), .B1(n12584), .B2(n9847), .C1(
        n6655), .C2(n9846), .ZN(P3_U3287) );
  OAI222_X1 U12426 ( .A1(P2_U3088), .A2(n9972), .B1(n13955), .B2(n9849), .C1(
        n9848), .C2(n13960), .ZN(P2_U3321) );
  INV_X1 U12427 ( .A(n14223), .ZN(n10022) );
  OAI222_X1 U12428 ( .A1(n12562), .A2(n6884), .B1(n6656), .B2(n9849), .C1(
        n10022), .C2(P1_U3086), .ZN(P1_U3349) );
  NAND2_X1 U12429 ( .A1(n13465), .A2(n7722), .ZN(n9851) );
  OR2_X1 U12430 ( .A1(n10130), .A2(P3_U3151), .ZN(n9850) );
  OAI211_X1 U12431 ( .C1(n6873), .C2(n6655), .A(n9851), .B(n9850), .ZN(n9852)
         );
  INV_X1 U12432 ( .A(n9852), .ZN(P3_U3293) );
  OAI222_X1 U12433 ( .A1(P3_U3151), .A2(n11464), .B1(n12584), .B2(n7424), .C1(
        n6655), .C2(n9853), .ZN(P3_U3285) );
  OAI22_X1 U12434 ( .A1(n10224), .A2(P3_U3151), .B1(SI_5_), .B2(n12584), .ZN(
        n9854) );
  AOI21_X1 U12435 ( .B1(n10995), .B2(n9855), .A(n9854), .ZN(P3_U3290) );
  INV_X1 U12436 ( .A(n14210), .ZN(n10018) );
  OAI222_X1 U12437 ( .A1(n12562), .A2(n9857), .B1(n6656), .B2(n9856), .C1(
        n10018), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U12438 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9859) );
  INV_X1 U12439 ( .A(n9858), .ZN(n9860) );
  INV_X1 U12440 ( .A(n10043), .ZN(n14235) );
  OAI222_X1 U12441 ( .A1(n12562), .A2(n9859), .B1(n6656), .B2(n9860), .C1(
        P1_U3086), .C2(n14235), .ZN(P1_U3348) );
  OAI222_X1 U12442 ( .A1(n13960), .A2(n9861), .B1(n13955), .B2(n9860), .C1(
        P2_U3088), .C2(n15037), .ZN(P2_U3320) );
  INV_X1 U12443 ( .A(n14195), .ZN(n9864) );
  OAI222_X1 U12444 ( .A1(P1_U3086), .A2(n9864), .B1(n6656), .B2(n9863), .C1(
        n9862), .C2(n12562), .ZN(P1_U3352) );
  INV_X1 U12445 ( .A(n9947), .ZN(n9998) );
  OAI222_X1 U12446 ( .A1(P2_U3088), .A2(n9998), .B1(n13955), .B2(n9866), .C1(
        n9865), .C2(n13960), .ZN(P2_U3319) );
  INV_X1 U12447 ( .A(n10103), .ZN(n10099) );
  OAI222_X1 U12448 ( .A1(n12562), .A2(n9867), .B1(n6656), .B2(n9866), .C1(
        n10099), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U12449 ( .A(n9868), .ZN(n9869) );
  OAI222_X1 U12450 ( .A1(P3_U3151), .A2(n11572), .B1(n12584), .B2(n9870), .C1(
        n6655), .C2(n9869), .ZN(P3_U3284) );
  OAI222_X1 U12451 ( .A1(n13960), .A2(n9872), .B1(n13955), .B2(n9871), .C1(
        P2_U3088), .C2(n9935), .ZN(P2_U3325) );
  OAI222_X1 U12452 ( .A1(P2_U3088), .A2(n9911), .B1(n13955), .B2(n9874), .C1(
        n9873), .C2(n13960), .ZN(P2_U3326) );
  INV_X1 U12453 ( .A(n9875), .ZN(n9877) );
  OAI222_X1 U12454 ( .A1(n12562), .A2(n9876), .B1(n6656), .B2(n9877), .C1(
        P1_U3086), .C2(n10282), .ZN(P1_U3346) );
  OAI222_X1 U12455 ( .A1(n13960), .A2(n9878), .B1(n13955), .B2(n9877), .C1(
        P2_U3088), .C2(n10260), .ZN(P2_U3318) );
  INV_X1 U12456 ( .A(n9879), .ZN(n9880) );
  OAI222_X1 U12457 ( .A1(P3_U3151), .A2(n12073), .B1(n12584), .B2(n9881), .C1(
        n6655), .C2(n9880), .ZN(P3_U3283) );
  INV_X1 U12458 ( .A(n10335), .ZN(n9882) );
  NAND2_X1 U12459 ( .A1(n9882), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12560) );
  INV_X1 U12460 ( .A(n12560), .ZN(n9883) );
  OR2_X1 U12461 ( .A1(n10342), .A2(n9883), .ZN(n10028) );
  INV_X1 U12462 ( .A(n12501), .ZN(n11416) );
  NAND2_X1 U12463 ( .A1(n11416), .A2(n10335), .ZN(n9885) );
  NAND2_X1 U12464 ( .A1(n9885), .A2(n9884), .ZN(n10026) );
  NAND2_X1 U12465 ( .A1(n10028), .A2(n10026), .ZN(n14878) );
  INV_X1 U12466 ( .A(n14878), .ZN(n14255) );
  NOR2_X1 U12467 ( .A1(n14255), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12468 ( .A(n9886), .ZN(n9888) );
  INV_X1 U12469 ( .A(n14256), .ZN(n14252) );
  OAI222_X1 U12470 ( .A1(n12562), .A2(n9887), .B1(n6656), .B2(n9888), .C1(
        P1_U3086), .C2(n14252), .ZN(P1_U3345) );
  OAI222_X1 U12471 ( .A1(n13960), .A2(n9889), .B1(n13955), .B2(n9888), .C1(
        P2_U3088), .C2(n10375), .ZN(P2_U3317) );
  AOI21_X1 U12472 ( .B1(n9891), .B2(n9890), .A(n9120), .ZN(n9892) );
  OR2_X1 U12473 ( .A1(n9893), .A2(n9892), .ZN(n9894) );
  AND2_X1 U12474 ( .A1(n9894), .A2(n9585), .ZN(n15009) );
  AND2_X1 U12475 ( .A1(n15009), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15089) );
  INV_X1 U12476 ( .A(n15111), .ZN(n15083) );
  NOR2_X1 U12477 ( .A1(n15133), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9901) );
  NOR2_X1 U12478 ( .A1(n9585), .A2(P2_U3088), .ZN(n13952) );
  NAND2_X1 U12479 ( .A1(n9894), .A2(n13952), .ZN(n9902) );
  INV_X1 U12480 ( .A(n9902), .ZN(n9895) );
  NAND2_X1 U12481 ( .A1(n9931), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9918) );
  INV_X1 U12482 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n15225) );
  NAND2_X1 U12483 ( .A1(n13962), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9896) );
  AOI21_X1 U12484 ( .B1(n9911), .B2(n15225), .A(n9896), .ZN(n9897) );
  NAND2_X1 U12485 ( .A1(n9918), .A2(n9897), .ZN(n9919) );
  MUX2_X1 U12486 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n15225), .S(n9911), .Z(n9898) );
  OAI21_X1 U12487 ( .B1(n9974), .B2(n9907), .A(n9898), .ZN(n9899) );
  AND3_X1 U12488 ( .A1(n15085), .A2(n9919), .A3(n9899), .ZN(n9900) );
  AOI211_X1 U12489 ( .C1(n15083), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n9901), .B(
        n9900), .ZN(n9910) );
  OR2_X1 U12490 ( .A1(n9902), .A2(n13957), .ZN(n15105) );
  MUX2_X1 U12491 ( .A(n9903), .B(P2_REG2_REG_1__SCAN_IN), .S(n9911), .Z(n9905)
         );
  AND2_X1 U12492 ( .A1(n13962), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U12493 ( .A1(n9905), .A2(n9904), .ZN(n9933) );
  MUX2_X1 U12494 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9903), .S(n9911), .Z(n9906)
         );
  OAI21_X1 U12495 ( .B1(n9973), .B2(n9907), .A(n9906), .ZN(n9908) );
  NAND3_X1 U12496 ( .A1(n15091), .A2(n9933), .A3(n9908), .ZN(n9909) );
  OAI211_X1 U12497 ( .C1(n15107), .C2(n9911), .A(n9910), .B(n9909), .ZN(
        P2_U3215) );
  OAI222_X1 U12498 ( .A1(P3_U3151), .A2(n12092), .B1(n12584), .B2(n9913), .C1(
        n6655), .C2(n9912), .ZN(P3_U3282) );
  INV_X1 U12499 ( .A(n9914), .ZN(n9916) );
  INV_X1 U12500 ( .A(n10571), .ZN(n10566) );
  OAI222_X1 U12501 ( .A1(n12562), .A2(n9915), .B1(n6656), .B2(n9916), .C1(
        P1_U3086), .C2(n10566), .ZN(P1_U3344) );
  OAI222_X1 U12502 ( .A1(n13960), .A2(n9917), .B1(n13955), .B2(n9916), .C1(
        P2_U3088), .C2(n10834), .ZN(P2_U3316) );
  INV_X1 U12503 ( .A(n10260), .ZN(n9955) );
  NOR2_X1 U12504 ( .A1(n9955), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9928) );
  INV_X1 U12505 ( .A(n15010), .ZN(n9921) );
  INV_X1 U12506 ( .A(n10011), .ZN(n9920) );
  XNOR2_X1 U12507 ( .A(n9935), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n13607) );
  NAND2_X1 U12508 ( .A1(n9919), .A2(n9918), .ZN(n13608) );
  INV_X1 U12509 ( .A(n9935), .ZN(n13610) );
  AOI22_X1 U12510 ( .A1(n13607), .A2(n13608), .B1(n13610), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10002) );
  MUX2_X1 U12511 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9021), .S(n10011), .Z(
        n10001) );
  NOR2_X1 U12512 ( .A1(n10002), .A2(n10001), .ZN(n10000) );
  AOI21_X1 U12513 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n9920), .A(n10000), .ZN(
        n15017) );
  MUX2_X1 U12514 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9030), .S(n15010), .Z(
        n15016) );
  NOR2_X1 U12515 ( .A1(n15017), .A2(n15016), .ZN(n15015) );
  AOI21_X1 U12516 ( .B1(n9921), .B2(P2_REG1_REG_4__SCAN_IN), .A(n15015), .ZN(
        n15029) );
  MUX2_X1 U12517 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9922), .S(n9941), .Z(n15028) );
  NOR2_X1 U12518 ( .A1(n15029), .A2(n15028), .ZN(n15027) );
  NOR2_X1 U12519 ( .A1(n9941), .A2(n9922), .ZN(n9962) );
  MUX2_X1 U12520 ( .A(n9923), .B(P2_REG1_REG_6__SCAN_IN), .S(n9972), .Z(n9961)
         );
  OAI21_X1 U12521 ( .B1(n15027), .B2(n9962), .A(n9961), .ZN(n9960) );
  OAI21_X1 U12522 ( .B1(n9923), .B2(n9972), .A(n9960), .ZN(n15046) );
  MUX2_X1 U12523 ( .A(n9924), .B(P2_REG1_REG_7__SCAN_IN), .S(n15037), .Z(
        n15045) );
  NAND2_X1 U12524 ( .A1(n15046), .A2(n15045), .ZN(n15044) );
  OAI21_X1 U12525 ( .B1(n9924), .B2(n15037), .A(n15044), .ZN(n9989) );
  MUX2_X1 U12526 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9925), .S(n9947), .Z(n9988)
         );
  NAND2_X1 U12527 ( .A1(n9989), .A2(n9988), .ZN(n9987) );
  OAI21_X1 U12528 ( .B1(n9925), .B2(n9998), .A(n9987), .ZN(n9930) );
  MUX2_X1 U12529 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9926), .S(n10260), .Z(n9927) );
  NOR2_X1 U12530 ( .A1(n9930), .A2(n9927), .ZN(n10259) );
  AOI21_X1 U12531 ( .B1(n9928), .B2(n9930), .A(n10259), .ZN(n9959) );
  NOR2_X1 U12532 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12118), .ZN(n9929) );
  AOI21_X1 U12533 ( .B1(n15083), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n9929), .ZN(
        n9958) );
  NAND3_X1 U12534 ( .A1(n9930), .A2(n15085), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n9950) );
  INV_X1 U12535 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10899) );
  MUX2_X1 U12536 ( .A(n9934), .B(P2_REG2_REG_2__SCAN_IN), .S(n9935), .Z(n13613) );
  NAND2_X1 U12537 ( .A1(n9931), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9932) );
  NAND2_X1 U12538 ( .A1(n9933), .A2(n9932), .ZN(n13612) );
  NAND2_X1 U12539 ( .A1(n13613), .A2(n13612), .ZN(n13611) );
  OR2_X1 U12540 ( .A1(n9935), .A2(n9934), .ZN(n10005) );
  NAND2_X1 U12541 ( .A1(n13611), .A2(n10005), .ZN(n9937) );
  MUX2_X1 U12542 ( .A(n10603), .B(P2_REG2_REG_3__SCAN_IN), .S(n10011), .Z(
        n9936) );
  NAND2_X1 U12543 ( .A1(n9937), .A2(n9936), .ZN(n10008) );
  OR2_X1 U12544 ( .A1(n10011), .A2(n10603), .ZN(n9938) );
  NAND2_X1 U12545 ( .A1(n10008), .A2(n9938), .ZN(n15014) );
  MUX2_X1 U12546 ( .A(n9939), .B(P2_REG2_REG_4__SCAN_IN), .S(n15010), .Z(
        n15013) );
  NAND2_X1 U12547 ( .A1(n15014), .A2(n15013), .ZN(n15012) );
  OR2_X1 U12548 ( .A1(n15010), .A2(n9939), .ZN(n9940) );
  NAND2_X1 U12549 ( .A1(n15012), .A2(n9940), .ZN(n15033) );
  INV_X1 U12550 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10612) );
  MUX2_X1 U12551 ( .A(n10612), .B(P2_REG2_REG_5__SCAN_IN), .S(n9941), .Z(
        n15032) );
  NAND2_X1 U12552 ( .A1(n15033), .A2(n15032), .ZN(n15031) );
  INV_X1 U12553 ( .A(n9941), .ZN(n15023) );
  NAND2_X1 U12554 ( .A1(n15023), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U12555 ( .A1(n15031), .A2(n9967), .ZN(n9943) );
  INV_X1 U12556 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10642) );
  MUX2_X1 U12557 ( .A(n10642), .B(P2_REG2_REG_6__SCAN_IN), .S(n9972), .Z(n9942) );
  NAND2_X1 U12558 ( .A1(n9943), .A2(n9942), .ZN(n9969) );
  OR2_X1 U12559 ( .A1(n9972), .A2(n10642), .ZN(n9944) );
  NAND2_X1 U12560 ( .A1(n9969), .A2(n9944), .ZN(n15043) );
  MUX2_X1 U12561 ( .A(n15115), .B(P2_REG2_REG_7__SCAN_IN), .S(n15037), .Z(
        n15042) );
  NAND2_X1 U12562 ( .A1(n15043), .A2(n15042), .ZN(n15041) );
  OR2_X1 U12563 ( .A1(n15037), .A2(n15115), .ZN(n9945) );
  NAND2_X1 U12564 ( .A1(n15041), .A2(n9945), .ZN(n9992) );
  MUX2_X1 U12565 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9946), .S(n9947), .Z(n9991)
         );
  NAND2_X1 U12566 ( .A1(n9992), .A2(n9991), .ZN(n9990) );
  NAND2_X1 U12567 ( .A1(n9947), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12568 ( .A1(n9990), .A2(n9948), .ZN(n9952) );
  NAND3_X1 U12569 ( .A1(n15091), .A2(P2_REG2_REG_9__SCAN_IN), .A3(n9952), .ZN(
        n9949) );
  NAND3_X1 U12570 ( .A1(n9950), .A2(n15107), .A3(n9949), .ZN(n9956) );
  INV_X1 U12571 ( .A(n9952), .ZN(n9953) );
  NAND2_X1 U12572 ( .A1(n10260), .A2(n10899), .ZN(n10266) );
  MUX2_X1 U12573 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10899), .S(n10260), .Z(
        n9951) );
  OAI21_X1 U12574 ( .B1(n9953), .B2(n10266), .A(n10267), .ZN(n9954) );
  AOI22_X1 U12575 ( .A1(n9956), .A2(n9955), .B1(n15091), .B2(n9954), .ZN(n9957) );
  OAI211_X1 U12576 ( .C1(n9959), .C2(n15103), .A(n9958), .B(n9957), .ZN(
        P2_U3223) );
  AND2_X1 U12577 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10512) );
  INV_X1 U12578 ( .A(n9960), .ZN(n9964) );
  NOR3_X1 U12579 ( .A1(n15027), .A2(n9962), .A3(n9961), .ZN(n9963) );
  NOR3_X1 U12580 ( .A1(n15103), .A2(n9964), .A3(n9963), .ZN(n9965) );
  AOI211_X1 U12581 ( .C1(n15083), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n10512), .B(
        n9965), .ZN(n9971) );
  MUX2_X1 U12582 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10642), .S(n9972), .Z(n9966) );
  NAND3_X1 U12583 ( .A1(n15031), .A2(n9967), .A3(n9966), .ZN(n9968) );
  NAND3_X1 U12584 ( .A1(n15091), .A2(n9969), .A3(n9968), .ZN(n9970) );
  OAI211_X1 U12585 ( .C1(n15107), .C2(n9972), .A(n9971), .B(n9970), .ZN(
        P2_U3220) );
  OAI22_X1 U12586 ( .A1(n15103), .A2(n9974), .B1(n9973), .B2(n15105), .ZN(
        n9977) );
  NAND2_X1 U12587 ( .A1(n15085), .A2(n9974), .ZN(n9975) );
  OAI211_X1 U12588 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n15105), .A(n15107), .B(
        n9975), .ZN(n9976) );
  MUX2_X1 U12589 ( .A(n9977), .B(n9976), .S(n13962), .Z(n9981) );
  INV_X1 U12590 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9979) );
  OAI22_X1 U12591 ( .A1(n15111), .A2(n9979), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9978), .ZN(n9980) );
  OR2_X1 U12592 ( .A1(n9981), .A2(n9980), .ZN(P2_U3214) );
  INV_X1 U12593 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n15615) );
  NAND2_X1 U12594 ( .A1(n12874), .A2(P3_U3897), .ZN(n9982) );
  OAI21_X1 U12595 ( .B1(P3_U3897), .B2(n15615), .A(n9982), .ZN(P3_U3500) );
  INV_X1 U12596 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n15484) );
  NAND2_X1 U12597 ( .A1(n12956), .A2(P3_U3897), .ZN(n9983) );
  OAI21_X1 U12598 ( .B1(P3_U3897), .B2(n15484), .A(n9983), .ZN(P3_U3495) );
  INV_X1 U12599 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n15631) );
  NAND2_X1 U12600 ( .A1(n13015), .A2(P3_U3897), .ZN(n9984) );
  OAI21_X1 U12601 ( .B1(P3_U3897), .B2(n15631), .A(n9984), .ZN(P3_U3503) );
  INV_X1 U12602 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n15450) );
  NAND2_X1 U12603 ( .A1(n13016), .A2(P3_U3897), .ZN(n9985) );
  OAI21_X1 U12604 ( .B1(P3_U3897), .B2(n15450), .A(n9985), .ZN(P3_U3501) );
  INV_X1 U12605 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n15509) );
  NAND2_X1 U12606 ( .A1(n12652), .A2(P3_U3897), .ZN(n9986) );
  OAI21_X1 U12607 ( .B1(P3_U3897), .B2(n15509), .A(n9986), .ZN(P3_U3498) );
  OAI211_X1 U12608 ( .C1(n9989), .C2(n9988), .A(n15085), .B(n9987), .ZN(n9994)
         );
  OAI211_X1 U12609 ( .C1(n9992), .C2(n9991), .A(n15091), .B(n9990), .ZN(n9993)
         );
  NAND2_X1 U12610 ( .A1(n9994), .A2(n9993), .ZN(n9996) );
  NAND2_X1 U12611 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10933) );
  INV_X1 U12612 ( .A(n10933), .ZN(n9995) );
  AOI211_X1 U12613 ( .C1(n15083), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n9996), .B(
        n9995), .ZN(n9997) );
  OAI21_X1 U12614 ( .B1(n15107), .B2(n9998), .A(n9997), .ZN(P2_U3222) );
  INV_X1 U12615 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9999) );
  NOR2_X1 U12616 ( .A1(n15111), .A2(n9999), .ZN(n10004) );
  AOI211_X1 U12617 ( .C1(n10002), .C2(n10001), .A(n10000), .B(n15103), .ZN(
        n10003) );
  AOI211_X1 U12618 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3088), .A(n10004), 
        .B(n10003), .ZN(n10010) );
  MUX2_X1 U12619 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10603), .S(n10011), .Z(
        n10006) );
  NAND3_X1 U12620 ( .A1(n10006), .A2(n13611), .A3(n10005), .ZN(n10007) );
  NAND3_X1 U12621 ( .A1(n15091), .A2(n10008), .A3(n10007), .ZN(n10009) );
  OAI211_X1 U12622 ( .C1(n15107), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        P2_U3217) );
  INV_X1 U12623 ( .A(n10012), .ZN(n10014) );
  OAI222_X1 U12624 ( .A1(n12077), .A2(P3_U3151), .B1(n6655), .B2(n10014), .C1(
        n10013), .C2(n12584), .ZN(P3_U3281) );
  INV_X1 U12625 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n14992) );
  MUX2_X1 U12626 ( .A(n14992), .B(P1_REG1_REG_8__SCAN_IN), .S(n10103), .Z(
        n10025) );
  INV_X1 U12627 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10023) );
  INV_X1 U12628 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10020) );
  INV_X1 U12629 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10019) );
  INV_X1 U12630 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14988) );
  MUX2_X1 U12631 ( .A(n14988), .B(P1_REG1_REG_1__SCAN_IN), .S(n10035), .Z(
        n14162) );
  AND2_X1 U12632 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14161) );
  NAND2_X1 U12633 ( .A1(n14162), .A2(n14161), .ZN(n14160) );
  INV_X1 U12634 ( .A(n10035), .ZN(n14163) );
  NAND2_X1 U12635 ( .A1(n14163), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U12636 ( .A1(n14160), .A2(n10015), .ZN(n14186) );
  INV_X1 U12637 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14990) );
  MUX2_X1 U12638 ( .A(n14990), .B(P1_REG1_REG_2__SCAN_IN), .S(n14180), .Z(
        n14187) );
  NAND2_X1 U12639 ( .A1(n14186), .A2(n14187), .ZN(n14185) );
  INV_X1 U12640 ( .A(n14180), .ZN(n14179) );
  NAND2_X1 U12641 ( .A1(n14179), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U12642 ( .A1(n14185), .A2(n10016), .ZN(n14192) );
  INV_X1 U12643 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n15637) );
  MUX2_X1 U12644 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n15637), .S(n14195), .Z(
        n14193) );
  NAND2_X1 U12645 ( .A1(n14192), .A2(n14193), .ZN(n14191) );
  NAND2_X1 U12646 ( .A1(n14195), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U12647 ( .A1(n14191), .A2(n10017), .ZN(n14208) );
  MUX2_X1 U12648 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10019), .S(n14210), .Z(
        n14209) );
  NAND2_X1 U12649 ( .A1(n14208), .A2(n14209), .ZN(n14207) );
  OAI21_X1 U12650 ( .B1(n10019), .B2(n10018), .A(n14207), .ZN(n10085) );
  XNOR2_X1 U12651 ( .A(n10042), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n10086) );
  MUX2_X1 U12652 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10021), .S(n14223), .Z(
        n14226) );
  MUX2_X1 U12653 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10023), .S(n10043), .Z(
        n14240) );
  NAND2_X1 U12654 ( .A1(n14239), .A2(n14240), .ZN(n14238) );
  OAI21_X1 U12655 ( .B1(n14235), .B2(n10023), .A(n14238), .ZN(n10024) );
  NOR2_X1 U12656 ( .A1(n10024), .A2(n10025), .ZN(n10098) );
  AOI21_X1 U12657 ( .B1(n10025), .B2(n10024), .A(n10098), .ZN(n10052) );
  INV_X1 U12658 ( .A(n10026), .ZN(n10027) );
  NAND2_X1 U12659 ( .A1(n10028), .A2(n10027), .ZN(n10115) );
  INV_X1 U12660 ( .A(n10115), .ZN(n10029) );
  NAND2_X1 U12661 ( .A1(n10029), .A2(n6734), .ZN(n14295) );
  NOR2_X1 U12662 ( .A1(n10115), .A2(n14172), .ZN(n14293) );
  INV_X1 U12663 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10030) );
  NAND2_X1 U12664 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11551) );
  OAI21_X1 U12665 ( .B1(n14878), .B2(n10030), .A(n11551), .ZN(n10031) );
  AOI21_X1 U12666 ( .B1(n14293), .B2(n10103), .A(n10031), .ZN(n10051) );
  OR2_X1 U12667 ( .A1(n11968), .A2(n6734), .ZN(n10032) );
  NOR2_X2 U12668 ( .A1(n10115), .A2(n10032), .ZN(n14299) );
  INV_X1 U12669 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10033) );
  MUX2_X1 U12670 ( .A(n10033), .B(P1_REG2_REG_2__SCAN_IN), .S(n14180), .Z(
        n10037) );
  INV_X1 U12671 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10034) );
  MUX2_X1 U12672 ( .A(n10034), .B(P1_REG2_REG_1__SCAN_IN), .S(n10035), .Z(
        n14164) );
  AND2_X1 U12673 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14171) );
  NAND2_X1 U12674 ( .A1(n14164), .A2(n14171), .ZN(n14182) );
  OR2_X1 U12675 ( .A1(n10035), .A2(n10034), .ZN(n14181) );
  NAND2_X1 U12676 ( .A1(n14182), .A2(n14181), .ZN(n10036) );
  NAND2_X1 U12677 ( .A1(n10037), .A2(n10036), .ZN(n14198) );
  NAND2_X1 U12678 ( .A1(n14179), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14196) );
  NAND2_X1 U12679 ( .A1(n14198), .A2(n14196), .ZN(n10039) );
  INV_X1 U12680 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11349) );
  MUX2_X1 U12681 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11349), .S(n14195), .Z(
        n10038) );
  NAND2_X1 U12682 ( .A1(n10039), .A2(n10038), .ZN(n14213) );
  NAND2_X1 U12683 ( .A1(n14195), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14212) );
  NAND2_X1 U12684 ( .A1(n14213), .A2(n14212), .ZN(n10041) );
  INV_X1 U12685 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11329) );
  MUX2_X1 U12686 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11329), .S(n14210), .Z(
        n10040) );
  NAND2_X1 U12687 ( .A1(n10041), .A2(n10040), .ZN(n14215) );
  NAND2_X1 U12688 ( .A1(n14210), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10090) );
  INV_X1 U12689 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11405) );
  MUX2_X1 U12690 ( .A(n11405), .B(P1_REG2_REG_5__SCAN_IN), .S(n10042), .Z(
        n10091) );
  AOI21_X1 U12691 ( .B1(n14215), .B2(n10090), .A(n10091), .ZN(n14229) );
  NOR2_X1 U12692 ( .A1(n10087), .A2(n11405), .ZN(n14228) );
  MUX2_X1 U12693 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11370), .S(n14223), .Z(
        n14227) );
  OAI21_X1 U12694 ( .B1(n14229), .B2(n14228), .A(n14227), .ZN(n14243) );
  NAND2_X1 U12695 ( .A1(n14223), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14242) );
  INV_X1 U12696 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11395) );
  MUX2_X1 U12697 ( .A(n11395), .B(P1_REG2_REG_7__SCAN_IN), .S(n10043), .Z(
        n14241) );
  AOI21_X1 U12698 ( .B1(n14243), .B2(n14242), .A(n14241), .ZN(n10045) );
  NOR2_X1 U12699 ( .A1(n14235), .A2(n11395), .ZN(n10046) );
  INV_X1 U12700 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11360) );
  MUX2_X1 U12701 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11360), .S(n10103), .Z(
        n10044) );
  OAI21_X1 U12702 ( .B1(n10045), .B2(n10046), .A(n10044), .ZN(n10106) );
  INV_X1 U12703 ( .A(n10045), .ZN(n14245) );
  INV_X1 U12704 ( .A(n10046), .ZN(n10048) );
  MUX2_X1 U12705 ( .A(n11360), .B(P1_REG2_REG_8__SCAN_IN), .S(n10103), .Z(
        n10047) );
  NAND3_X1 U12706 ( .A1(n14245), .A2(n10048), .A3(n10047), .ZN(n10049) );
  NAND3_X1 U12707 ( .A1(n14299), .A2(n10106), .A3(n10049), .ZN(n10050) );
  OAI211_X1 U12708 ( .C1(n10052), .C2(n14295), .A(n10051), .B(n10050), .ZN(
        P1_U3251) );
  INV_X1 U12709 ( .A(n10053), .ZN(n10055) );
  INV_X1 U12710 ( .A(n10793), .ZN(n10788) );
  OAI222_X1 U12711 ( .A1(n12562), .A2(n10054), .B1(n6656), .B2(n10055), .C1(
        n10788), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12712 ( .A(n11436), .ZN(n10832) );
  OAI222_X1 U12713 ( .A1(n13960), .A2(n10056), .B1(n13955), .B2(n10055), .C1(
        n10832), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U12714 ( .A(n10057), .ZN(n10059) );
  OAI222_X1 U12715 ( .A1(n12060), .A2(P3_U3151), .B1(n6655), .B2(n10059), .C1(
        n10058), .C2(n12584), .ZN(P3_U3280) );
  INV_X1 U12716 ( .A(n15201), .ZN(n15146) );
  XNOR2_X1 U12717 ( .A(n10061), .B(n10060), .ZN(n10649) );
  INV_X1 U12718 ( .A(n10649), .ZN(n10071) );
  INV_X1 U12719 ( .A(n10062), .ZN(n15135) );
  AOI211_X1 U12720 ( .C1(n12047), .C2(n15135), .A(n12009), .B(n10594), .ZN(
        n10648) );
  AOI21_X1 U12721 ( .B1(n15196), .B2(n12047), .A(n10648), .ZN(n10070) );
  OAI21_X1 U12722 ( .B1(n10063), .B2(n10065), .A(n10064), .ZN(n10069) );
  NAND2_X1 U12723 ( .A1(n13605), .A2(n15128), .ZN(n10067) );
  NAND2_X1 U12724 ( .A1(n13606), .A2(n15127), .ZN(n10066) );
  AND2_X1 U12725 ( .A1(n10067), .A2(n10066), .ZN(n12045) );
  INV_X1 U12726 ( .A(n12045), .ZN(n10068) );
  AOI21_X1 U12727 ( .B1(n10069), .B2(n15131), .A(n10068), .ZN(n10652) );
  OAI211_X1 U12728 ( .C1(n15200), .C2(n10071), .A(n10070), .B(n10652), .ZN(
        n10072) );
  AOI21_X1 U12729 ( .B1(n15146), .B2(n10649), .A(n10072), .ZN(n15181) );
  NOR2_X1 U12730 ( .A1(n15162), .A2(n10073), .ZN(n10074) );
  AND2_X1 U12731 ( .A1(n10074), .A2(n15165), .ZN(n10076) );
  NAND2_X1 U12732 ( .A1(n15231), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10077) );
  OAI21_X1 U12733 ( .B1(n15181), .B2(n15231), .A(n10077), .ZN(P2_U3501) );
  INV_X1 U12734 ( .A(n10794), .ZN(n11060) );
  INV_X1 U12735 ( .A(n10078), .ZN(n10080) );
  OAI222_X1 U12736 ( .A1(P1_U3086), .A2(n11060), .B1(n6656), .B2(n10080), .C1(
        n10079), .C2(n12562), .ZN(P1_U3342) );
  INV_X1 U12737 ( .A(n15050), .ZN(n11440) );
  OAI222_X1 U12738 ( .A1(n13960), .A2(n10081), .B1(n13955), .B2(n10080), .C1(
        n11440), .C2(P2_U3088), .ZN(P2_U3314) );
  OAI222_X1 U12739 ( .A1(P3_U3151), .A2(n12083), .B1(n12584), .B2(n10083), 
        .C1(n6655), .C2(n10082), .ZN(P3_U3279) );
  AOI21_X1 U12740 ( .B1(n10086), .B2(n10085), .A(n10084), .ZN(n10096) );
  INV_X1 U12741 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n15671) );
  NOR2_X1 U12742 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15671), .ZN(n10089) );
  INV_X1 U12743 ( .A(n14293), .ZN(n14870) );
  NOR2_X1 U12744 ( .A1(n14870), .A2(n10087), .ZN(n10088) );
  AOI211_X1 U12745 ( .C1(n14255), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n10089), .B(
        n10088), .ZN(n10095) );
  INV_X1 U12746 ( .A(n14229), .ZN(n10093) );
  NAND3_X1 U12747 ( .A1(n10091), .A2(n14215), .A3(n10090), .ZN(n10092) );
  NAND3_X1 U12748 ( .A1(n14299), .A2(n10093), .A3(n10092), .ZN(n10094) );
  OAI211_X1 U12749 ( .C1(n10096), .C2(n14295), .A(n10095), .B(n10094), .ZN(
        P1_U3248) );
  INV_X1 U12750 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10097) );
  MUX2_X1 U12751 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10097), .S(n10282), .Z(
        n10101) );
  AOI21_X1 U12752 ( .B1(n14992), .B2(n10099), .A(n10098), .ZN(n10100) );
  NOR2_X1 U12753 ( .A1(n10100), .A2(n10101), .ZN(n10275) );
  AOI21_X1 U12754 ( .B1(n10101), .B2(n10100), .A(n10275), .ZN(n10111) );
  AND2_X1 U12755 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11766) );
  NOR2_X1 U12756 ( .A1(n14870), .A2(n10282), .ZN(n10102) );
  AOI211_X1 U12757 ( .C1(n14255), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n11766), .B(
        n10102), .ZN(n10110) );
  NAND2_X1 U12758 ( .A1(n10103), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10105) );
  MUX2_X1 U12759 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10281), .S(n10282), .Z(
        n10104) );
  AOI21_X1 U12760 ( .B1(n10106), .B2(n10105), .A(n10104), .ZN(n14262) );
  INV_X1 U12761 ( .A(n14262), .ZN(n10108) );
  NAND3_X1 U12762 ( .A1(n10106), .A2(n10105), .A3(n10104), .ZN(n10107) );
  NAND3_X1 U12763 ( .A1(n10108), .A2(n14299), .A3(n10107), .ZN(n10109) );
  OAI211_X1 U12764 ( .C1(n10111), .C2(n14295), .A(n10110), .B(n10109), .ZN(
        P1_U3252) );
  NOR2_X1 U12765 ( .A1(n6734), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10112) );
  NOR2_X1 U12766 ( .A1(n10112), .A2(n11968), .ZN(n14175) );
  INV_X1 U12767 ( .A(n6734), .ZN(n12556) );
  OAI21_X1 U12768 ( .B1(n12556), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14175), .ZN(
        n10113) );
  MUX2_X1 U12769 ( .A(n14175), .B(n10113), .S(n10349), .Z(n10114) );
  INV_X1 U12770 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11413) );
  OAI22_X1 U12771 ( .A1(n10115), .A2(n10114), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11413), .ZN(n10117) );
  NOR3_X1 U12772 ( .A1(n14295), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n10349), .ZN(
        n10116) );
  AOI211_X1 U12773 ( .C1(n14255), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n10117), .B(
        n10116), .ZN(n10118) );
  INV_X1 U12774 ( .A(n10118), .ZN(P1_U3243) );
  MUX2_X1 U12775 ( .A(n10120), .B(n10119), .S(n12105), .Z(n10160) );
  XNOR2_X1 U12776 ( .A(n10160), .B(n10147), .ZN(n10161) );
  MUX2_X1 U12777 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n6648), .Z(n10121) );
  MUX2_X1 U12778 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n6648), .Z(n10405) );
  NOR2_X1 U12779 ( .A1(n10405), .A2(n10404), .ZN(n10403) );
  INV_X1 U12780 ( .A(n10121), .ZN(n10122) );
  MUX2_X1 U12781 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12105), .Z(n10123) );
  XOR2_X1 U12782 ( .A(n10130), .B(n10123), .Z(n10422) );
  XOR2_X1 U12783 ( .A(n10161), .B(n10162), .Z(n10159) );
  NAND2_X1 U12784 ( .A1(P3_U3897), .A2(n12806), .ZN(n13170) );
  INV_X1 U12785 ( .A(n10671), .ZN(n10124) );
  OR2_X1 U12786 ( .A1(n10232), .A2(P3_U3151), .ZN(n12812) );
  NAND2_X1 U12787 ( .A1(n10124), .A2(n12812), .ZN(n10153) );
  NAND2_X1 U12788 ( .A1(n8227), .A2(n10232), .ZN(n10125) );
  NAND2_X1 U12789 ( .A1(n10126), .A2(n10125), .ZN(n10152) );
  INV_X1 U12790 ( .A(n10152), .ZN(n10127) );
  AND2_X1 U12791 ( .A1(n10153), .A2(n10127), .ZN(n10129) );
  MUX2_X1 U12792 ( .A(n10129), .B(P3_U3897), .S(n10128), .Z(n13166) );
  INV_X1 U12793 ( .A(n10129), .ZN(n10140) );
  INV_X1 U12794 ( .A(n13165), .ZN(n13093) );
  MUX2_X1 U12795 ( .A(n10133), .B(P3_REG1_REG_2__SCAN_IN), .S(n10130), .Z(
        n10415) );
  NAND2_X1 U12796 ( .A1(n10132), .A2(n7648), .ZN(n10190) );
  NAND2_X1 U12797 ( .A1(n10192), .A2(n7648), .ZN(n10414) );
  NAND2_X1 U12798 ( .A1(n10415), .A2(n10414), .ZN(n10413) );
  OR2_X1 U12799 ( .A1(n10130), .A2(n10133), .ZN(n10134) );
  NAND2_X1 U12800 ( .A1(n10136), .A2(n10119), .ZN(n10137) );
  NAND2_X1 U12801 ( .A1(n10168), .A2(n10137), .ZN(n10138) );
  NAND2_X1 U12802 ( .A1(n13093), .A2(n10138), .ZN(n10156) );
  INV_X1 U12803 ( .A(n13150), .ZN(n13158) );
  INV_X1 U12804 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15257) );
  NAND2_X1 U12805 ( .A1(n10404), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U12806 ( .A1(n7724), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U12807 ( .A1(n10144), .A2(n10145), .ZN(n10186) );
  INV_X1 U12808 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10185) );
  OR2_X1 U12809 ( .A1(n10186), .A2(n10185), .ZN(n10188) );
  NAND2_X1 U12810 ( .A1(n10188), .A2(n10145), .ZN(n10411) );
  OR2_X1 U12811 ( .A1(n10130), .A2(n15257), .ZN(n10146) );
  NAND2_X1 U12812 ( .A1(n10410), .A2(n10146), .ZN(n10148) );
  NAND2_X1 U12813 ( .A1(n10149), .A2(n10120), .ZN(n10150) );
  NAND2_X1 U12814 ( .A1(n10177), .A2(n10150), .ZN(n10151) );
  NAND2_X1 U12815 ( .A1(n13158), .A2(n10151), .ZN(n10155) );
  NOR2_X1 U12816 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12886), .ZN(n12884) );
  AOI21_X1 U12817 ( .B1(n15234), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n12884), .ZN(
        n10154) );
  NAND3_X1 U12818 ( .A1(n10156), .A2(n10155), .A3(n10154), .ZN(n10157) );
  AOI21_X1 U12819 ( .B1(n7213), .B2(n13166), .A(n10157), .ZN(n10158) );
  OAI21_X1 U12820 ( .B1(n10159), .B2(n13170), .A(n10158), .ZN(P3_U3185) );
  MUX2_X1 U12821 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12105), .Z(n10199) );
  XNOR2_X1 U12822 ( .A(n10199), .B(n10213), .ZN(n10200) );
  XOR2_X1 U12823 ( .A(n10200), .B(n10201), .Z(n10183) );
  INV_X1 U12824 ( .A(n10213), .ZN(n10181) );
  INV_X1 U12825 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10163) );
  XNOR2_X1 U12826 ( .A(n10213), .B(n10163), .ZN(n10165) );
  NAND2_X1 U12827 ( .A1(n10164), .A2(n10165), .ZN(n10209) );
  INV_X1 U12828 ( .A(n10165), .ZN(n10167) );
  NAND3_X1 U12829 ( .A1(n10168), .A2(n10167), .A3(n10166), .ZN(n10169) );
  AND2_X1 U12830 ( .A1(n10209), .A2(n10169), .ZN(n10171) );
  NAND2_X1 U12831 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n10699) );
  NAND2_X1 U12832 ( .A1(n15234), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10170) );
  OAI211_X1 U12833 ( .C1(n13165), .C2(n10171), .A(n10699), .B(n10170), .ZN(
        n10180) );
  XNOR2_X1 U12834 ( .A(n10213), .B(n10172), .ZN(n10174) );
  NAND2_X1 U12835 ( .A1(n10173), .A2(n10174), .ZN(n10215) );
  INV_X1 U12836 ( .A(n10174), .ZN(n10176) );
  NAND3_X1 U12837 ( .A1(n10177), .A2(n10176), .A3(n10175), .ZN(n10178) );
  AOI21_X1 U12838 ( .B1(n10215), .B2(n10178), .A(n13150), .ZN(n10179) );
  AOI211_X1 U12839 ( .C1(n13166), .C2(n10181), .A(n10180), .B(n10179), .ZN(
        n10182) );
  OAI21_X1 U12840 ( .B1(n10183), .B2(n13170), .A(n10182), .ZN(P3_U3186) );
  XOR2_X1 U12841 ( .A(n10184), .B(n10403), .Z(n10198) );
  NAND2_X1 U12842 ( .A1(n10186), .A2(n10185), .ZN(n10187) );
  NAND2_X1 U12843 ( .A1(n10188), .A2(n10187), .ZN(n10195) );
  NAND2_X1 U12844 ( .A1(n15234), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10189) );
  OAI21_X1 U12845 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n10673), .A(n10189), .ZN(
        n10194) );
  NAND2_X1 U12846 ( .A1(n10190), .A2(n7684), .ZN(n10191) );
  AOI21_X1 U12847 ( .B1(n10192), .B2(n10191), .A(n13165), .ZN(n10193) );
  AOI211_X1 U12848 ( .C1(n13158), .C2(n10195), .A(n10194), .B(n10193), .ZN(
        n10197) );
  OAI211_X1 U12849 ( .C1(n10198), .C2(n13170), .A(n10197), .B(n10196), .ZN(
        P3_U3183) );
  MUX2_X1 U12850 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n6648), .Z(n10202) );
  NAND2_X1 U12851 ( .A1(n10202), .A2(n10216), .ZN(n10205) );
  NAND2_X1 U12852 ( .A1(n10204), .A2(n10205), .ZN(n10439) );
  INV_X1 U12853 ( .A(n10439), .ZN(n10207) );
  INV_X1 U12854 ( .A(n10202), .ZN(n10203) );
  NAND2_X1 U12855 ( .A1(n10203), .A2(n10224), .ZN(n10438) );
  AOI21_X1 U12856 ( .B1(n10438), .B2(n10205), .A(n10204), .ZN(n10206) );
  AOI21_X1 U12857 ( .B1(n10207), .B2(n10438), .A(n10206), .ZN(n10226) );
  NAND2_X1 U12858 ( .A1(n10213), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U12859 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  AOI21_X1 U12860 ( .B1(n10211), .B2(n15697), .A(n10442), .ZN(n10222) );
  NOR2_X1 U12861 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10212), .ZN(n12955) );
  NAND2_X1 U12862 ( .A1(n10213), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U12863 ( .A1(n10215), .A2(n10214), .ZN(n10217) );
  AOI21_X1 U12864 ( .B1(n10218), .B2(n10923), .A(n6870), .ZN(n10219) );
  NOR2_X1 U12865 ( .A1(n13150), .A2(n10219), .ZN(n10220) );
  AOI211_X1 U12866 ( .C1(n15234), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n12955), .B(
        n10220), .ZN(n10221) );
  OAI21_X1 U12867 ( .B1(n10222), .B2(n13165), .A(n10221), .ZN(n10223) );
  AOI21_X1 U12868 ( .B1(n10224), .B2(n13166), .A(n10223), .ZN(n10225) );
  OAI21_X1 U12869 ( .B1(n10226), .B2(n13170), .A(n10225), .ZN(P3_U3187) );
  NAND2_X1 U12870 ( .A1(n13061), .A2(n10912), .ZN(n12621) );
  INV_X1 U12871 ( .A(n12621), .ZN(n10227) );
  NOR2_X1 U12872 ( .A1(n12619), .A2(n10227), .ZN(n12769) );
  NAND2_X1 U12873 ( .A1(n10231), .A2(n15295), .ZN(n10229) );
  INV_X1 U12874 ( .A(n10234), .ZN(n10228) );
  OAI22_X1 U12875 ( .A1(n10245), .A2(n10229), .B1(n10319), .B2(n10228), .ZN(
        n10230) );
  NAND2_X1 U12876 ( .A1(n10245), .A2(n10231), .ZN(n10238) );
  AND2_X1 U12877 ( .A1(n10233), .A2(n10232), .ZN(n10237) );
  NAND2_X1 U12878 ( .A1(n10319), .A2(n10234), .ZN(n10235) );
  NAND4_X1 U12879 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10239) );
  NAND2_X1 U12880 ( .A1(n10239), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10241) );
  INV_X1 U12881 ( .A(n12808), .ZN(n10317) );
  NAND2_X1 U12882 ( .A1(n10319), .A2(n10317), .ZN(n10240) );
  NAND2_X1 U12883 ( .A1(n13031), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10430) );
  NAND2_X1 U12884 ( .A1(n10430), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10250) );
  NOR2_X1 U12885 ( .A1(n12808), .A2(n10316), .ZN(n10242) );
  NAND2_X1 U12886 ( .A1(n10243), .A2(n10242), .ZN(n13028) );
  NAND2_X1 U12887 ( .A1(n10245), .A2(n12803), .ZN(n10247) );
  AND2_X1 U12888 ( .A1(n10671), .A2(n15302), .ZN(n10246) );
  AOI22_X1 U12889 ( .A1(n13037), .A2(n10244), .B1(n13044), .B2(n10248), .ZN(
        n10249) );
  OAI211_X1 U12890 ( .C1(n12769), .C2(n13046), .A(n10250), .B(n10249), .ZN(
        P3_U3172) );
  INV_X1 U12891 ( .A(n10342), .ZN(n10251) );
  NOR2_X2 U12892 ( .A1(n10252), .A2(n10251), .ZN(n14943) );
  INV_X1 U12893 ( .A(n10253), .ZN(n10254) );
  OAI22_X1 U12894 ( .A1(n14959), .A2(P1_D_REG_0__SCAN_IN), .B1(n10257), .B2(
        n10254), .ZN(n10255) );
  INV_X1 U12895 ( .A(n10255), .ZN(P1_U3445) );
  OAI22_X1 U12896 ( .A1(n14959), .A2(P1_D_REG_1__SCAN_IN), .B1(n10257), .B2(
        n10256), .ZN(n10258) );
  INV_X1 U12897 ( .A(n10258), .ZN(P1_U3446) );
  NAND2_X1 U12898 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11081)
         );
  AOI21_X1 U12899 ( .B1(n9926), .B2(n10260), .A(n10259), .ZN(n10263) );
  MUX2_X1 U12900 ( .A(n10261), .B(P2_REG1_REG_10__SCAN_IN), .S(n10375), .Z(
        n10262) );
  NAND2_X1 U12901 ( .A1(n10263), .A2(n10262), .ZN(n10374) );
  OAI211_X1 U12902 ( .C1(n10263), .C2(n10262), .A(n15085), .B(n10374), .ZN(
        n10264) );
  NAND2_X1 U12903 ( .A1(n11081), .A2(n10264), .ZN(n10265) );
  AOI21_X1 U12904 ( .B1(n15083), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10265), 
        .ZN(n10273) );
  NAND2_X1 U12905 ( .A1(n10267), .A2(n10266), .ZN(n10269) );
  INV_X1 U12906 ( .A(n10269), .ZN(n10271) );
  MUX2_X1 U12907 ( .A(n10990), .B(P2_REG2_REG_10__SCAN_IN), .S(n10375), .Z(
        n10270) );
  MUX2_X1 U12908 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10990), .S(n10375), .Z(
        n10268) );
  OAI211_X1 U12909 ( .C1(n10271), .C2(n10270), .A(n15091), .B(n10373), .ZN(
        n10272) );
  OAI211_X1 U12910 ( .C1(n15107), .C2(n10375), .A(n10273), .B(n10272), .ZN(
        P2_U3224) );
  INV_X1 U12911 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10274) );
  MUX2_X1 U12912 ( .A(n10274), .B(P1_REG1_REG_11__SCAN_IN), .S(n10571), .Z(
        n10278) );
  INV_X1 U12913 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10276) );
  MUX2_X1 U12914 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10276), .S(n14256), .Z(
        n14250) );
  AOI21_X1 U12915 ( .B1(n10278), .B2(n10277), .A(n10565), .ZN(n10292) );
  NOR2_X1 U12916 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11887), .ZN(n10280) );
  NOR2_X1 U12917 ( .A1(n14870), .A2(n10566), .ZN(n10279) );
  AOI211_X1 U12918 ( .C1(n14255), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10280), 
        .B(n10279), .ZN(n10291) );
  INV_X1 U12919 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10281) );
  NOR2_X1 U12920 ( .A1(n10282), .A2(n10281), .ZN(n14257) );
  INV_X1 U12921 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10283) );
  MUX2_X1 U12922 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10283), .S(n14256), .Z(
        n10284) );
  OAI21_X1 U12923 ( .B1(n14262), .B2(n14257), .A(n10284), .ZN(n14260) );
  NAND2_X1 U12924 ( .A1(n14256), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10287) );
  INV_X1 U12925 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10285) );
  MUX2_X1 U12926 ( .A(n10285), .B(P1_REG2_REG_11__SCAN_IN), .S(n10571), .Z(
        n10286) );
  AOI21_X1 U12927 ( .B1(n14260), .B2(n10287), .A(n10286), .ZN(n10570) );
  INV_X1 U12928 ( .A(n10570), .ZN(n10289) );
  NAND3_X1 U12929 ( .A1(n14260), .A2(n10287), .A3(n10286), .ZN(n10288) );
  NAND3_X1 U12930 ( .A1(n10289), .A2(n14299), .A3(n10288), .ZN(n10290) );
  OAI211_X1 U12931 ( .C1(n10292), .C2(n14295), .A(n10291), .B(n10290), .ZN(
        P1_U3254) );
  INV_X1 U12932 ( .A(n10293), .ZN(n10295) );
  OAI222_X1 U12933 ( .A1(n12102), .A2(P3_U3151), .B1(n6655), .B2(n10295), .C1(
        n10294), .C2(n12584), .ZN(P3_U3278) );
  NAND2_X1 U12934 ( .A1(n8837), .A2(n14908), .ZN(n12300) );
  OAI21_X1 U12935 ( .B1(n14899), .B2(n14918), .A(n7108), .ZN(n10297) );
  NAND2_X1 U12936 ( .A1(n14158), .A2(n14110), .ZN(n10358) );
  OR2_X1 U12937 ( .A1(n14908), .A2(n11414), .ZN(n10296) );
  AND2_X1 U12938 ( .A1(n10358), .A2(n10296), .ZN(n11421) );
  AND2_X1 U12939 ( .A1(n10297), .A2(n11421), .ZN(n14961) );
  NAND2_X1 U12940 ( .A1(n14991), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10298) );
  OAI21_X1 U12941 ( .B1(n14991), .B2(n14961), .A(n10298), .ZN(P1_U3528) );
  INV_X1 U12942 ( .A(n10430), .ZN(n10324) );
  INV_X1 U12943 ( .A(n12802), .ZN(n10300) );
  NAND2_X1 U12944 ( .A1(n12618), .A2(n12613), .ZN(n10301) );
  NAND2_X1 U12945 ( .A1(n10561), .A2(n10301), .ZN(n10302) );
  NAND3_X1 U12946 ( .A1(n10244), .A2(n12849), .A3(n10307), .ZN(n10308) );
  NAND2_X1 U12947 ( .A1(n10674), .A2(n12849), .ZN(n10309) );
  NAND2_X1 U12948 ( .A1(n10310), .A2(n10309), .ZN(n10311) );
  INV_X1 U12949 ( .A(n12619), .ZN(n10313) );
  NAND3_X1 U12950 ( .A1(n10313), .A2(n12772), .A3(n12903), .ZN(n10314) );
  NAND2_X1 U12951 ( .A1(n10315), .A2(n12995), .ZN(n10323) );
  NAND2_X1 U12952 ( .A1(n10317), .A2(n10316), .ZN(n10318) );
  INV_X1 U12953 ( .A(n13017), .ZN(n13041) );
  INV_X1 U12954 ( .A(n13061), .ZN(n10320) );
  OAI22_X1 U12955 ( .A1(n13041), .A2(n10320), .B1(n7745), .B2(n13028), .ZN(
        n10321) );
  AOI21_X1 U12956 ( .B1(n13044), .B2(n10307), .A(n10321), .ZN(n10322) );
  OAI211_X1 U12957 ( .C1(n10324), .C2(n10673), .A(n10323), .B(n10322), .ZN(
        P3_U3162) );
  INV_X1 U12958 ( .A(n10325), .ZN(n10327) );
  OAI222_X1 U12959 ( .A1(P2_U3088), .A2(n13627), .B1(n13955), .B2(n10327), 
        .C1(n10326), .C2(n13960), .ZN(P2_U3311) );
  INV_X1 U12960 ( .A(n11906), .ZN(n11788) );
  OAI222_X1 U12961 ( .A1(n12562), .A2(n10328), .B1(n6656), .B2(n10327), .C1(
        n11788), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12962 ( .A(n13167), .ZN(n12086) );
  OAI222_X1 U12963 ( .A1(P3_U3151), .A2(n12086), .B1(n12584), .B2(n10330), 
        .C1(n6655), .C2(n10329), .ZN(P3_U3277) );
  INV_X1 U12964 ( .A(n11302), .ZN(n10331) );
  NAND2_X1 U12965 ( .A1(n10331), .A2(n11303), .ZN(n10356) );
  INV_X1 U12966 ( .A(n10332), .ZN(n10333) );
  OAI21_X1 U12967 ( .B1(n10356), .B2(n10333), .A(n10340), .ZN(n10338) );
  AND2_X1 U12968 ( .A1(n10335), .A2(n10334), .ZN(n10336) );
  NAND2_X1 U12969 ( .A1(n10348), .A2(n10336), .ZN(n12558) );
  INV_X1 U12970 ( .A(n12558), .ZN(n10337) );
  NAND2_X1 U12971 ( .A1(n10338), .A2(n10337), .ZN(n10715) );
  OR2_X1 U12972 ( .A1(n10715), .A2(P1_U3086), .ZN(n10711) );
  INV_X1 U12973 ( .A(n10711), .ZN(n10362) );
  OR2_X1 U12974 ( .A1(n10356), .A2(n10339), .ZN(n10353) );
  INV_X1 U12975 ( .A(n10340), .ZN(n10341) );
  INV_X1 U12976 ( .A(n12502), .ZN(n10343) );
  INV_X1 U12977 ( .A(n10348), .ZN(n10344) );
  NAND2_X2 U12978 ( .A1(n12262), .A2(n6736), .ZN(n10622) );
  NOR2_X1 U12979 ( .A1(n10619), .A2(n10352), .ZN(n10621) );
  AOI21_X1 U12980 ( .B1(n10619), .B2(n10352), .A(n10621), .ZN(n14170) );
  INV_X1 U12981 ( .A(n10353), .ZN(n10355) );
  NOR2_X1 U12982 ( .A1(n14974), .A2(n11416), .ZN(n10354) );
  INV_X1 U12983 ( .A(n10356), .ZN(n10357) );
  NAND2_X1 U12984 ( .A1(n10357), .A2(n11305), .ZN(n14121) );
  OAI22_X1 U12985 ( .A1(n14170), .A2(n14103), .B1(n14121), .B2(n10358), .ZN(
        n10359) );
  AOI21_X1 U12986 ( .B1(n10360), .B2(n6638), .A(n10359), .ZN(n10361) );
  OAI21_X1 U12987 ( .B1(n10362), .B2(n11413), .A(n10361), .ZN(P1_U3232) );
  OR3_X1 U12988 ( .A1(n12769), .A2(n15302), .A3(n10363), .ZN(n10366) );
  OR2_X1 U12989 ( .A1(n10364), .A2(n13312), .ZN(n10365) );
  AND2_X1 U12990 ( .A1(n10366), .A2(n10365), .ZN(n10909) );
  MUX2_X1 U12991 ( .A(n10909), .B(n15623), .S(n15696), .Z(n10367) );
  OAI21_X1 U12992 ( .B1(n10912), .B2(n13409), .A(n10367), .ZN(P3_U3459) );
  INV_X1 U12993 ( .A(n10368), .ZN(n10370) );
  INV_X1 U12994 ( .A(n11428), .ZN(n15061) );
  OAI222_X1 U12995 ( .A1(n13960), .A2(n10369), .B1(n13955), .B2(n10370), .C1(
        n15061), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U12996 ( .A(n11063), .ZN(n11782) );
  OAI222_X1 U12997 ( .A1(n12562), .A2(n10371), .B1(n6656), .B2(n10370), .C1(
        n11782), .C2(P1_U3086), .ZN(P1_U3341) );
  NOR2_X1 U12998 ( .A1(n15105), .A2(n10386), .ZN(n10377) );
  OR2_X1 U12999 ( .A1(n10375), .A2(n10990), .ZN(n10372) );
  NAND2_X1 U13000 ( .A1(n10373), .A2(n10372), .ZN(n10388) );
  OAI21_X1 U13001 ( .B1(n10261), .B2(n10375), .A(n10374), .ZN(n10381) );
  NOR3_X1 U13002 ( .A1(n10381), .A2(P2_REG1_REG_11__SCAN_IN), .A3(n15103), 
        .ZN(n10376) );
  AOI211_X1 U13003 ( .C1(n10377), .C2(n10388), .A(n15089), .B(n10376), .ZN(
        n10392) );
  AOI21_X1 U13004 ( .B1(n10834), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10381), 
        .ZN(n10378) );
  NOR2_X1 U13005 ( .A1(n10378), .A2(n15103), .ZN(n10383) );
  MUX2_X1 U13006 ( .A(n10379), .B(P2_REG1_REG_11__SCAN_IN), .S(n10834), .Z(
        n10380) );
  NAND2_X1 U13007 ( .A1(n10381), .A2(n10380), .ZN(n10833) );
  INV_X1 U13008 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14729) );
  NAND2_X1 U13009 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11021)
         );
  OAI21_X1 U13010 ( .B1(n15111), .B2(n14729), .A(n11021), .ZN(n10382) );
  AOI21_X1 U13011 ( .B1(n10383), .B2(n10833), .A(n10382), .ZN(n10391) );
  INV_X1 U13012 ( .A(n10388), .ZN(n10385) );
  INV_X1 U13013 ( .A(n10834), .ZN(n10384) );
  NOR3_X1 U13014 ( .A1(n10385), .A2(P2_REG2_REG_11__SCAN_IN), .A3(n10384), 
        .ZN(n10389) );
  MUX2_X1 U13015 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10386), .S(n10834), .Z(
        n10387) );
  NOR2_X1 U13016 ( .A1(n10388), .A2(n10387), .ZN(n10828) );
  OAI21_X1 U13017 ( .B1(n10389), .B2(n10828), .A(n15091), .ZN(n10390) );
  OAI211_X1 U13018 ( .C1(n10392), .C2(n10834), .A(n10391), .B(n10390), .ZN(
        P2_U3225) );
  MUX2_X1 U13019 ( .A(n10909), .B(n7702), .S(n15307), .Z(n10393) );
  OAI21_X1 U13020 ( .B1(n10912), .B2(n13456), .A(n10393), .ZN(P3_U3390) );
  INV_X1 U13021 ( .A(n10394), .ZN(n10396) );
  OAI222_X1 U13022 ( .A1(n13960), .A2(n10395), .B1(n13955), .B2(n10396), .C1(
        P2_U3088), .C2(n11442), .ZN(P2_U3312) );
  OAI222_X1 U13023 ( .A1(n12562), .A2(n10397), .B1(n6656), .B2(n10396), .C1(
        P1_U3086), .C2(n6966), .ZN(P1_U3340) );
  INV_X1 U13024 ( .A(n14270), .ZN(n14276) );
  INV_X1 U13025 ( .A(n10398), .ZN(n10400) );
  OAI222_X1 U13026 ( .A1(P1_U3086), .A2(n14276), .B1(n6656), .B2(n10400), .C1(
        n10399), .C2(n12562), .ZN(P1_U3338) );
  INV_X1 U13027 ( .A(n15088), .ZN(n13628) );
  OAI222_X1 U13028 ( .A1(n13960), .A2(n10401), .B1(n13955), .B2(n10400), .C1(
        n13628), .C2(P2_U3088), .ZN(P2_U3310) );
  OAI222_X1 U13029 ( .A1(n12584), .A2(n15620), .B1(P3_U3151), .B2(n12800), 
        .C1(n6655), .C2(n10402), .ZN(P3_U3276) );
  INV_X1 U13030 ( .A(n13170), .ZN(n13132) );
  NOR3_X1 U13031 ( .A1(n13158), .A2(n13093), .A3(n13132), .ZN(n10409) );
  AOI21_X1 U13032 ( .B1(n10405), .B2(n10404), .A(n10403), .ZN(n10408) );
  AOI22_X1 U13033 ( .A1(n15234), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10407) );
  OAI211_X1 U13034 ( .C1(n10409), .C2(n10408), .A(n10407), .B(n10406), .ZN(
        P3_U3182) );
  INV_X1 U13035 ( .A(n13166), .ZN(n11582) );
  OAI21_X1 U13036 ( .B1(n10412), .B2(n10411), .A(n10410), .ZN(n10420) );
  OAI21_X1 U13037 ( .B1(n10415), .B2(n10414), .A(n10413), .ZN(n10416) );
  AND2_X1 U13038 ( .A1(n13093), .A2(n10416), .ZN(n10419) );
  INV_X1 U13039 ( .A(n15234), .ZN(n13125) );
  INV_X1 U13040 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10417) );
  OAI22_X1 U13041 ( .A1(n13125), .A2(n10417), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15239), .ZN(n10418) );
  AOI211_X1 U13042 ( .C1(n13158), .C2(n10420), .A(n10419), .B(n10418), .ZN(
        n10425) );
  XNOR2_X1 U13043 ( .A(n10422), .B(n10421), .ZN(n10423) );
  NAND2_X1 U13044 ( .A1(n10423), .A2(n13132), .ZN(n10424) );
  OAI211_X1 U13045 ( .C1(n11582), .C2(n7728), .A(n10425), .B(n10424), .ZN(
        P3_U3184) );
  NAND2_X1 U13046 ( .A1(n10427), .A2(n10426), .ZN(n10685) );
  XNOR2_X1 U13047 ( .A(n12903), .B(n7746), .ZN(n10686) );
  XNOR2_X1 U13048 ( .A(n10686), .B(n7745), .ZN(n10684) );
  XOR2_X1 U13049 ( .A(n10685), .B(n10684), .Z(n10432) );
  INV_X1 U13050 ( .A(n13044), .ZN(n13003) );
  AOI22_X1 U13051 ( .A1(n13037), .A2(n15243), .B1(n13017), .B2(n10244), .ZN(
        n10428) );
  OAI21_X1 U13052 ( .B1(n7746), .B2(n13003), .A(n10428), .ZN(n10429) );
  AOI21_X1 U13053 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10430), .A(n10429), .ZN(
        n10431) );
  OAI21_X1 U13054 ( .B1(n10432), .B2(n13046), .A(n10431), .ZN(P3_U3177) );
  INV_X1 U13055 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10446) );
  MUX2_X1 U13056 ( .A(n10446), .B(n10433), .S(n12105), .Z(n10434) );
  NAND2_X1 U13057 ( .A1(n10434), .A2(n10445), .ZN(n10462) );
  INV_X1 U13058 ( .A(n10434), .ZN(n10435) );
  NAND2_X1 U13059 ( .A1(n10435), .A2(n10477), .ZN(n10436) );
  NAND2_X1 U13060 ( .A1(n10462), .A2(n10436), .ZN(n10437) );
  AOI21_X1 U13061 ( .B1(n10439), .B2(n10438), .A(n10437), .ZN(n10496) );
  AND3_X1 U13062 ( .A1(n10439), .A2(n10438), .A3(n10437), .ZN(n10440) );
  OAI21_X1 U13063 ( .B1(n10496), .B2(n10440), .A(n13132), .ZN(n10455) );
  MUX2_X1 U13064 ( .A(n10433), .B(P3_REG1_REG_6__SCAN_IN), .S(n10445), .Z(
        n10444) );
  OAI21_X1 U13065 ( .B1(n10444), .B2(n10443), .A(n10457), .ZN(n10453) );
  MUX2_X1 U13066 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n10446), .S(n10445), .Z(
        n10447) );
  NOR2_X1 U13067 ( .A1(n10447), .A2(n10448), .ZN(n10476) );
  AOI21_X1 U13068 ( .B1(n10448), .B2(n10447), .A(n10476), .ZN(n10451) );
  NAND2_X1 U13069 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n11128) );
  INV_X1 U13070 ( .A(n11128), .ZN(n10449) );
  AOI21_X1 U13071 ( .B1(n15234), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10449), .ZN(
        n10450) );
  OAI21_X1 U13072 ( .B1(n13150), .B2(n10451), .A(n10450), .ZN(n10452) );
  AOI21_X1 U13073 ( .B1(n13093), .B2(n10453), .A(n10452), .ZN(n10454) );
  OAI211_X1 U13074 ( .C1(n11582), .C2(n10477), .A(n10455), .B(n10454), .ZN(
        P3_U3188) );
  NOR2_X1 U13075 ( .A1(n10463), .A2(n10492), .ZN(n10491) );
  NAND2_X1 U13076 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10963), .ZN(n10459) );
  OAI21_X1 U13077 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10963), .A(n10459), .ZN(
        n10460) );
  AOI21_X1 U13078 ( .B1(n10461), .B2(n10460), .A(n6869), .ZN(n10490) );
  INV_X1 U13079 ( .A(n10462), .ZN(n10495) );
  MUX2_X1 U13080 ( .A(n10464), .B(n10463), .S(n6648), .Z(n10465) );
  NAND2_X1 U13081 ( .A1(n10465), .A2(n10478), .ZN(n10474) );
  INV_X1 U13082 ( .A(n10465), .ZN(n10466) );
  NAND2_X1 U13083 ( .A1(n10466), .A2(n7305), .ZN(n10467) );
  AND2_X1 U13084 ( .A1(n10474), .A2(n10467), .ZN(n10494) );
  OAI21_X1 U13085 ( .B1(n10496), .B2(n10495), .A(n10494), .ZN(n10493) );
  MUX2_X1 U13086 ( .A(n10468), .B(n15639), .S(n12105), .Z(n10470) );
  INV_X1 U13087 ( .A(n10963), .ZN(n10469) );
  NAND2_X1 U13088 ( .A1(n10470), .A2(n10469), .ZN(n10951) );
  INV_X1 U13089 ( .A(n10470), .ZN(n10471) );
  NAND2_X1 U13090 ( .A1(n10471), .A2(n10963), .ZN(n10472) );
  NAND2_X1 U13091 ( .A1(n10951), .A2(n10472), .ZN(n10473) );
  AOI21_X1 U13092 ( .B1(n10493), .B2(n10474), .A(n10473), .ZN(n10959) );
  AND3_X1 U13093 ( .A1(n10493), .A2(n10474), .A3(n10473), .ZN(n10475) );
  OAI21_X1 U13094 ( .B1(n10959), .B2(n10475), .A(n13132), .ZN(n10489) );
  NOR2_X1 U13095 ( .A1(n10478), .A2(n10479), .ZN(n10480) );
  XNOR2_X1 U13096 ( .A(n10479), .B(n10478), .ZN(n10500) );
  NAND2_X1 U13097 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10963), .ZN(n10481) );
  OAI21_X1 U13098 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10963), .A(n10481), .ZN(
        n10482) );
  AOI21_X1 U13099 ( .B1(n10483), .B2(n10482), .A(n10962), .ZN(n10486) );
  AND2_X1 U13100 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n11246) );
  NOR2_X1 U13101 ( .A1(n11582), .A2(n10963), .ZN(n10484) );
  AOI211_X1 U13102 ( .C1(n15234), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n11246), .B(
        n10484), .ZN(n10485) );
  OAI21_X1 U13103 ( .B1(n10486), .B2(n13150), .A(n10485), .ZN(n10487) );
  INV_X1 U13104 ( .A(n10487), .ZN(n10488) );
  OAI211_X1 U13105 ( .C1(n10490), .C2(n13165), .A(n10489), .B(n10488), .ZN(
        P3_U3190) );
  AOI21_X1 U13106 ( .B1(n10463), .B2(n10492), .A(n10491), .ZN(n10508) );
  INV_X1 U13107 ( .A(n10493), .ZN(n10498) );
  NOR3_X1 U13108 ( .A1(n10496), .A2(n10495), .A3(n10494), .ZN(n10497) );
  OAI21_X1 U13109 ( .B1(n10498), .B2(n10497), .A(n13132), .ZN(n10507) );
  AOI21_X1 U13110 ( .B1(n10464), .B2(n10500), .A(n10499), .ZN(n10504) );
  NOR2_X1 U13111 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10501), .ZN(n12817) );
  NOR2_X1 U13112 ( .A1(n11582), .A2(n7305), .ZN(n10502) );
  AOI211_X1 U13113 ( .C1(n15234), .C2(P3_ADDR_REG_7__SCAN_IN), .A(n12817), .B(
        n10502), .ZN(n10503) );
  OAI21_X1 U13114 ( .B1(n10504), .B2(n13150), .A(n10503), .ZN(n10505) );
  INV_X1 U13115 ( .A(n10505), .ZN(n10506) );
  OAI211_X1 U13116 ( .C1(n10508), .C2(n13165), .A(n10507), .B(n10506), .ZN(
        P3_U3189) );
  NAND2_X1 U13117 ( .A1(n13601), .A2(n15128), .ZN(n10510) );
  NAND2_X1 U13118 ( .A1(n13603), .A2(n15127), .ZN(n10509) );
  NAND2_X1 U13119 ( .A1(n10510), .A2(n10509), .ZN(n10640) );
  NOR2_X1 U13120 ( .A1(n13539), .A2(n10636), .ZN(n10511) );
  AOI211_X1 U13121 ( .C1(n13515), .C2(n10640), .A(n10512), .B(n10511), .ZN(
        n10530) );
  XNOR2_X1 U13122 ( .A(n13543), .B(n12033), .ZN(n10767) );
  NAND2_X1 U13123 ( .A1(n13604), .A2(n9794), .ZN(n10514) );
  XNOR2_X1 U13124 ( .A(n10767), .B(n10514), .ZN(n13550) );
  AND2_X1 U13125 ( .A1(n13550), .A2(n10513), .ZN(n10546) );
  NAND2_X1 U13126 ( .A1(n13549), .A2(n10546), .ZN(n13548) );
  INV_X1 U13127 ( .A(n10767), .ZN(n10515) );
  NAND2_X1 U13128 ( .A1(n10515), .A2(n10514), .ZN(n10542) );
  NAND2_X1 U13129 ( .A1(n13548), .A2(n10542), .ZN(n10517) );
  XNOR2_X1 U13130 ( .A(n15197), .B(n12033), .ZN(n10518) );
  NAND2_X1 U13131 ( .A1(n13603), .A2(n9794), .ZN(n10519) );
  XNOR2_X1 U13132 ( .A(n10518), .B(n10519), .ZN(n10768) );
  NAND2_X1 U13133 ( .A1(n10517), .A2(n10768), .ZN(n10775) );
  INV_X1 U13134 ( .A(n10518), .ZN(n10520) );
  NAND2_X1 U13135 ( .A1(n10520), .A2(n10519), .ZN(n10527) );
  NAND2_X1 U13136 ( .A1(n10775), .A2(n10527), .ZN(n10525) );
  INV_X1 U13137 ( .A(n10523), .ZN(n10538) );
  AND2_X1 U13138 ( .A1(n13602), .A2(n13753), .ZN(n10522) );
  INV_X1 U13139 ( .A(n10522), .ZN(n10521) );
  NAND2_X1 U13140 ( .A1(n10538), .A2(n10521), .ZN(n10524) );
  NAND2_X1 U13141 ( .A1(n10523), .A2(n10522), .ZN(n10541) );
  NAND2_X1 U13142 ( .A1(n10524), .A2(n10541), .ZN(n10526) );
  AOI21_X1 U13143 ( .B1(n10525), .B2(n10526), .A(n14999), .ZN(n10528) );
  NAND2_X1 U13144 ( .A1(n10775), .A2(n10539), .ZN(n10536) );
  NAND2_X1 U13145 ( .A1(n10528), .A2(n10536), .ZN(n10529) );
  OAI211_X1 U13146 ( .C1(n15007), .C2(n10635), .A(n10530), .B(n10529), .ZN(
        P2_U3211) );
  INV_X1 U13147 ( .A(n10533), .ZN(n10930) );
  AND2_X1 U13148 ( .A1(n13601), .A2(n13753), .ZN(n10532) );
  INV_X1 U13149 ( .A(n10532), .ZN(n10531) );
  NAND2_X1 U13150 ( .A1(n10930), .A2(n10531), .ZN(n10534) );
  NAND2_X1 U13151 ( .A1(n10533), .A2(n10532), .ZN(n10929) );
  AND2_X1 U13152 ( .A1(n10534), .A2(n10929), .ZN(n10550) );
  INV_X1 U13153 ( .A(n10550), .ZN(n10535) );
  AOI21_X1 U13154 ( .B1(n10536), .B2(n10535), .A(n14999), .ZN(n10554) );
  NOR3_X1 U13155 ( .A1(n13561), .A2(n10538), .A3(n10537), .ZN(n10553) );
  INV_X1 U13156 ( .A(n10541), .ZN(n10540) );
  AND2_X1 U13157 ( .A1(n10768), .A2(n10541), .ZN(n10547) );
  INV_X1 U13158 ( .A(n10542), .ZN(n10543) );
  INV_X1 U13159 ( .A(n10545), .ZN(n10552) );
  AND2_X1 U13160 ( .A1(n10547), .A2(n10546), .ZN(n10548) );
  NAND3_X1 U13161 ( .A1(n10552), .A2(n10551), .A3(n10550), .ZN(n11006) );
  OAI21_X1 U13162 ( .B1(n10554), .B2(n10553), .A(n11006), .ZN(n10560) );
  NAND2_X1 U13163 ( .A1(n13600), .A2(n15128), .ZN(n10556) );
  NAND2_X1 U13164 ( .A1(n13602), .A2(n15127), .ZN(n10555) );
  NAND2_X1 U13165 ( .A1(n10556), .A2(n10555), .ZN(n10822) );
  NAND2_X1 U13166 ( .A1(n13515), .A2(n10822), .ZN(n10557) );
  NAND2_X1 U13167 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15038) );
  OAI211_X1 U13168 ( .C1(n15007), .C2(n15114), .A(n10557), .B(n15038), .ZN(
        n10558) );
  AOI21_X1 U13169 ( .B1(n15117), .B2(n15004), .A(n10558), .ZN(n10559) );
  NAND2_X1 U13170 ( .A1(n10560), .A2(n10559), .ZN(P2_U3185) );
  OAI222_X1 U13171 ( .A1(n6655), .A2(n10563), .B1(n12584), .B2(n10562), .C1(
        P3_U3151), .C2(n10561), .ZN(P3_U3275) );
  INV_X1 U13172 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10564) );
  MUX2_X1 U13173 ( .A(n10564), .B(P1_REG1_REG_12__SCAN_IN), .S(n10793), .Z(
        n10568) );
  AOI21_X1 U13174 ( .B1(n10274), .B2(n10566), .A(n10565), .ZN(n10567) );
  NOR2_X1 U13175 ( .A1(n10567), .A2(n10568), .ZN(n10787) );
  AOI21_X1 U13176 ( .B1(n10568), .B2(n10567), .A(n10787), .ZN(n10579) );
  INV_X1 U13177 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10569) );
  MUX2_X1 U13178 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10569), .S(n10793), .Z(
        n10573) );
  AOI21_X1 U13179 ( .B1(n10571), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10570), 
        .ZN(n10572) );
  NAND2_X1 U13180 ( .A1(n10572), .A2(n10573), .ZN(n10792) );
  OAI21_X1 U13181 ( .B1(n10573), .B2(n10572), .A(n10792), .ZN(n10577) );
  NOR2_X1 U13182 ( .A1(n10574), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14011) );
  AOI21_X1 U13183 ( .B1(n14255), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n14011), 
        .ZN(n10575) );
  OAI21_X1 U13184 ( .B1(n14870), .B2(n10788), .A(n10575), .ZN(n10576) );
  AOI21_X1 U13185 ( .B1(n10577), .B2(n14299), .A(n10576), .ZN(n10578) );
  OAI21_X1 U13186 ( .B1(n10579), .B2(n14295), .A(n10578), .ZN(P1_U3255) );
  XNOR2_X1 U13187 ( .A(n11331), .B(n14155), .ZN(n12516) );
  XOR2_X1 U13188 ( .A(n12516), .B(n10580), .Z(n11336) );
  XNOR2_X1 U13189 ( .A(n10581), .B(n12516), .ZN(n10582) );
  NOR2_X1 U13190 ( .A1(n10582), .A2(n14921), .ZN(n11327) );
  INV_X1 U13191 ( .A(n10753), .ZN(n10583) );
  AOI211_X1 U13192 ( .C1(n12327), .C2(n11337), .A(n14909), .B(n10583), .ZN(
        n11333) );
  NAND2_X1 U13193 ( .A1(n14154), .A2(n14110), .ZN(n10585) );
  NAND2_X1 U13194 ( .A1(n14156), .A2(n14111), .ZN(n10584) );
  AND2_X1 U13195 ( .A1(n10585), .A2(n10584), .ZN(n10946) );
  INV_X1 U13196 ( .A(n10946), .ZN(n11326) );
  NOR3_X1 U13197 ( .A1(n11327), .A2(n11333), .A3(n11326), .ZN(n10586) );
  OAI21_X1 U13198 ( .B1(n14895), .B2(n11336), .A(n10586), .ZN(n10591) );
  INV_X1 U13199 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10587) );
  OAI22_X1 U13200 ( .A1(n14643), .A2(n11331), .B1(n14987), .B2(n10587), .ZN(
        n10588) );
  AOI21_X1 U13201 ( .B1(n10591), .B2(n14987), .A(n10588), .ZN(n10589) );
  INV_X1 U13202 ( .A(n10589), .ZN(P1_U3471) );
  OAI22_X1 U13203 ( .A1(n14596), .A2(n11331), .B1(n14994), .B2(n10019), .ZN(
        n10590) );
  AOI21_X1 U13204 ( .B1(n10591), .B2(n14994), .A(n10590), .ZN(n10592) );
  INV_X1 U13205 ( .A(n10592), .ZN(P1_U3532) );
  XNOR2_X1 U13206 ( .A(n10593), .B(n10598), .ZN(n15186) );
  INV_X1 U13207 ( .A(n10594), .ZN(n10595) );
  AOI211_X1 U13208 ( .C1(n15183), .C2(n10595), .A(n12009), .B(n10866), .ZN(
        n15182) );
  OAI22_X1 U13209 ( .A1(n13813), .A2(n10596), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15132), .ZN(n10597) );
  AOI21_X1 U13210 ( .B1(n13835), .B2(n15182), .A(n10597), .ZN(n10605) );
  XNOR2_X1 U13211 ( .A(n10599), .B(n10598), .ZN(n10602) );
  INV_X1 U13212 ( .A(n10600), .ZN(n10601) );
  AOI21_X1 U13213 ( .B1(n10602), .B2(n15131), .A(n10601), .ZN(n15184) );
  MUX2_X1 U13214 ( .A(n10603), .B(n15184), .S(n15155), .Z(n10604) );
  OAI211_X1 U13215 ( .C1(n15139), .C2(n15186), .A(n10605), .B(n10604), .ZN(
        P2_U3262) );
  XNOR2_X1 U13216 ( .A(n10606), .B(n10607), .ZN(n15202) );
  XNOR2_X1 U13217 ( .A(n10608), .B(n10607), .ZN(n10611) );
  NAND2_X1 U13218 ( .A1(n13602), .A2(n15128), .ZN(n10610) );
  NAND2_X1 U13219 ( .A1(n13604), .A2(n15127), .ZN(n10609) );
  NAND2_X1 U13220 ( .A1(n10610), .A2(n10609), .ZN(n10765) );
  AOI21_X1 U13221 ( .B1(n10611), .B2(n15131), .A(n10765), .ZN(n15206) );
  MUX2_X1 U13222 ( .A(n10612), .B(n15206), .S(n15155), .Z(n10616) );
  NAND2_X1 U13223 ( .A1(n10865), .A2(n15197), .ZN(n10613) );
  AND3_X1 U13224 ( .A1(n10634), .A2(n15134), .A3(n10613), .ZN(n15199) );
  OAI22_X1 U13225 ( .A1(n13813), .A2(n7069), .B1(n15132), .B2(n10764), .ZN(
        n10614) );
  AOI21_X1 U13226 ( .B1(n13835), .B2(n15199), .A(n10614), .ZN(n10615) );
  OAI211_X1 U13227 ( .C1(n15139), .C2(n15202), .A(n10616), .B(n10615), .ZN(
        P2_U3260) );
  INV_X1 U13228 ( .A(n14157), .ZN(n10617) );
  AOI22_X1 U13229 ( .A1(n11281), .A2(n14157), .B1(n12262), .B2(n14969), .ZN(
        n10618) );
  XNOR2_X1 U13230 ( .A(n10618), .B(n12212), .ZN(n10717) );
  XOR2_X1 U13231 ( .A(n10718), .B(n10717), .Z(n10720) );
  OAI22_X1 U13232 ( .A1(n10622), .A2(n8436), .B1(n14964), .B2(n12274), .ZN(
        n10624) );
  XNOR2_X1 U13233 ( .A(n10623), .B(n12212), .ZN(n10625) );
  XOR2_X1 U13234 ( .A(n10624), .B(n10625), .Z(n10706) );
  NOR2_X1 U13235 ( .A1(n10707), .A2(n10706), .ZN(n10705) );
  INV_X1 U13236 ( .A(n10624), .ZN(n10626) );
  XOR2_X1 U13237 ( .A(n10720), .B(n10721), .Z(n10629) );
  INV_X1 U13238 ( .A(n6638), .ZN(n14127) );
  AOI22_X1 U13239 ( .A1(n14111), .A2(n14158), .B1(n14156), .B2(n14110), .ZN(
        n14892) );
  OAI22_X1 U13240 ( .A1(n14127), .A2(n12316), .B1(n14892), .B2(n14121), .ZN(
        n10627) );
  AOI21_X1 U13241 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10711), .A(n10627), .ZN(
        n10628) );
  OAI21_X1 U13242 ( .B1(n10629), .B2(n14103), .A(n10628), .ZN(P1_U3237) );
  INV_X1 U13243 ( .A(n10630), .ZN(n10631) );
  AOI21_X1 U13244 ( .B1(n10639), .B2(n10632), .A(n10631), .ZN(n10657) );
  INV_X1 U13245 ( .A(n10824), .ZN(n10633) );
  AOI211_X1 U13246 ( .C1(n10654), .C2(n10634), .A(n12009), .B(n10633), .ZN(
        n10653) );
  OAI22_X1 U13247 ( .A1(n13813), .A2(n10636), .B1(n15132), .B2(n10635), .ZN(
        n10637) );
  AOI21_X1 U13248 ( .B1(n10653), .B2(n13835), .A(n10637), .ZN(n10644) );
  XNOR2_X1 U13249 ( .A(n10638), .B(n10639), .ZN(n10641) );
  AOI21_X1 U13250 ( .B1(n10641), .B2(n15131), .A(n10640), .ZN(n10656) );
  MUX2_X1 U13251 ( .A(n10642), .B(n10656), .S(n15155), .Z(n10643) );
  OAI211_X1 U13252 ( .C1(n10657), .C2(n15139), .A(n10644), .B(n10643), .ZN(
        P2_U3259) );
  OAI22_X1 U13253 ( .A1(n15155), .A2(n9934), .B1(n12043), .B2(n15132), .ZN(
        n10647) );
  NOR2_X1 U13254 ( .A1(n13813), .A2(n10645), .ZN(n10646) );
  AOI211_X1 U13255 ( .C1(n10648), .C2(n13835), .A(n10647), .B(n10646), .ZN(
        n10651) );
  INV_X1 U13256 ( .A(n15139), .ZN(n15122) );
  NAND2_X1 U13257 ( .A1(n15122), .A2(n10649), .ZN(n10650) );
  OAI211_X1 U13258 ( .C1(n15157), .C2(n10652), .A(n10651), .B(n10650), .ZN(
        P2_U3263) );
  AOI21_X1 U13259 ( .B1(n15196), .B2(n10654), .A(n10653), .ZN(n10655) );
  OAI211_X1 U13260 ( .C1(n10657), .C2(n15187), .A(n10656), .B(n10655), .ZN(
        n10662) );
  NAND2_X1 U13261 ( .A1(n10662), .A2(n15233), .ZN(n10658) );
  OAI21_X1 U13262 ( .B1(n15233), .B2(n9923), .A(n10658), .ZN(P2_U3505) );
  AND3_X1 U13263 ( .A1(n15162), .A2(n15165), .A3(n10659), .ZN(n10660) );
  NAND2_X1 U13264 ( .A1(n10662), .A2(n15212), .ZN(n10663) );
  OAI21_X1 U13265 ( .B1(n15212), .B2(n9073), .A(n10663), .ZN(P2_U3448) );
  NAND2_X1 U13266 ( .A1(n13458), .A2(n10664), .ZN(n10665) );
  OAI21_X1 U13267 ( .B1(n13458), .B2(n10666), .A(n10665), .ZN(n10667) );
  INV_X1 U13268 ( .A(n10667), .ZN(n10668) );
  NAND2_X1 U13269 ( .A1(n10669), .A2(n10668), .ZN(n10745) );
  NOR2_X1 U13270 ( .A1(n15295), .A2(n12803), .ZN(n10670) );
  NAND2_X2 U13271 ( .A1(n10745), .A2(n15238), .ZN(n13344) );
  NOR2_X1 U13272 ( .A1(n12618), .A2(n12803), .ZN(n15255) );
  OR2_X1 U13273 ( .A1(n13204), .A2(n15255), .ZN(n10672) );
  NAND2_X1 U13274 ( .A1(n13344), .A2(n10672), .ZN(n13305) );
  XNOR2_X1 U13275 ( .A(n12772), .B(n12619), .ZN(n15259) );
  OAI22_X1 U13276 ( .A1(n13305), .A2(n15259), .B1(n10673), .B2(n15238), .ZN(
        n10680) );
  NAND2_X1 U13277 ( .A1(n10307), .A2(n15302), .ZN(n15261) );
  XNOR2_X1 U13278 ( .A(n12772), .B(n10674), .ZN(n10677) );
  NAND2_X1 U13279 ( .A1(n13061), .A2(n15244), .ZN(n10675) );
  OAI21_X1 U13280 ( .B1(n7745), .B2(n13312), .A(n10675), .ZN(n10676) );
  AOI21_X1 U13281 ( .B1(n10677), .B2(n15248), .A(n10676), .ZN(n15262) );
  OAI21_X1 U13282 ( .B1(n15240), .B2(n15261), .A(n15262), .ZN(n10678) );
  MUX2_X1 U13283 ( .A(P3_REG2_REG_1__SCAN_IN), .B(n10678), .S(n13344), .Z(
        n10679) );
  OR2_X1 U13284 ( .A1(n10680), .A2(n10679), .ZN(P3_U3232) );
  INV_X1 U13285 ( .A(n13631), .ZN(n15106) );
  OAI222_X1 U13286 ( .A1(P2_U3088), .A2(n15106), .B1(n13955), .B2(n10683), 
        .C1(n10681), .C2(n13960), .ZN(P2_U3309) );
  INV_X1 U13287 ( .A(n14289), .ZN(n14282) );
  OAI222_X1 U13288 ( .A1(P1_U3086), .A2(n14282), .B1(n6656), .B2(n10683), .C1(
        n10682), .C2(n12562), .ZN(P1_U3337) );
  XNOR2_X1 U13289 ( .A(n12903), .B(n10697), .ZN(n11112) );
  XNOR2_X1 U13290 ( .A(n11112), .B(n12956), .ZN(n10695) );
  NAND2_X1 U13291 ( .A1(n10685), .A2(n10684), .ZN(n10689) );
  INV_X1 U13292 ( .A(n10686), .ZN(n10687) );
  NAND2_X1 U13293 ( .A1(n10687), .A2(n7745), .ZN(n10688) );
  XNOR2_X1 U13294 ( .A(n12903), .B(n12885), .ZN(n10691) );
  XNOR2_X1 U13295 ( .A(n10691), .B(n10848), .ZN(n12880) );
  INV_X1 U13296 ( .A(n10691), .ZN(n10692) );
  NAND2_X1 U13297 ( .A1(n10692), .A2(n15243), .ZN(n10693) );
  OAI21_X1 U13298 ( .B1(n10695), .B2(n10694), .A(n11114), .ZN(n10703) );
  INV_X1 U13299 ( .A(n10845), .ZN(n10696) );
  NAND2_X1 U13300 ( .A1(n13038), .A2(n10696), .ZN(n10701) );
  AOI22_X1 U13301 ( .A1(n13044), .A2(n10697), .B1(n13017), .B2(n15243), .ZN(
        n10700) );
  NAND2_X1 U13302 ( .A1(n13037), .A2(n13059), .ZN(n10698) );
  NAND4_X1 U13303 ( .A1(n10701), .A2(n10700), .A3(n10699), .A4(n10698), .ZN(
        n10702) );
  AOI21_X1 U13304 ( .B1(n10703), .B2(n12995), .A(n10702), .ZN(n10704) );
  INV_X1 U13305 ( .A(n10704), .ZN(P3_U3170) );
  AOI21_X1 U13306 ( .B1(n10707), .B2(n10706), .A(n10705), .ZN(n10714) );
  INV_X1 U13307 ( .A(n14121), .ZN(n14830) );
  NAND2_X1 U13308 ( .A1(n8837), .A2(n14111), .ZN(n10709) );
  NAND2_X1 U13309 ( .A1(n14157), .A2(n14110), .ZN(n10708) );
  NAND2_X1 U13310 ( .A1(n10709), .A2(n10708), .ZN(n14914) );
  AOI22_X1 U13311 ( .A1(n6638), .A2(n10710), .B1(n14830), .B2(n14914), .ZN(
        n10713) );
  NAND2_X1 U13312 ( .A1(n10711), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10712) );
  OAI211_X1 U13313 ( .C1(n10714), .C2(n14103), .A(n10713), .B(n10712), .ZN(
        P1_U3222) );
  OAI22_X1 U13314 ( .A1(n12322), .A2(n12274), .B1(n12275), .B2(n11340), .ZN(
        n10716) );
  XNOR2_X1 U13315 ( .A(n10716), .B(n12212), .ZN(n10941) );
  OAI22_X1 U13316 ( .A1(n10622), .A2(n12322), .B1(n11340), .B2(n12274), .ZN(
        n10940) );
  XNOR2_X1 U13317 ( .A(n10941), .B(n10940), .ZN(n10723) );
  INV_X1 U13318 ( .A(n10717), .ZN(n10719) );
  AOI211_X1 U13319 ( .C1(n10723), .C2(n10722), .A(n14103), .B(n6863), .ZN(
        n10724) );
  INV_X1 U13320 ( .A(n10724), .ZN(n10730) );
  NAND2_X1 U13321 ( .A1(n14157), .A2(n14111), .ZN(n10726) );
  NAND2_X1 U13322 ( .A1(n14155), .A2(n14110), .ZN(n10725) );
  NAND2_X1 U13323 ( .A1(n10726), .A2(n10725), .ZN(n11347) );
  INV_X1 U13324 ( .A(n11347), .ZN(n10727) );
  INV_X1 U13325 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n15555) );
  OAI22_X1 U13326 ( .A1(n14121), .A2(n10727), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15555), .ZN(n10728) );
  AOI21_X1 U13327 ( .B1(n14975), .B2(n6638), .A(n10728), .ZN(n10729) );
  OAI211_X1 U13328 ( .C1(n14836), .C2(P1_REG3_REG_3__SCAN_IN), .A(n10730), .B(
        n10729), .ZN(P1_U3218) );
  OAI222_X1 U13329 ( .A1(P3_U3151), .A2(n12618), .B1(n12584), .B2(n10732), 
        .C1(n6655), .C2(n10731), .ZN(P3_U3274) );
  OR2_X1 U13330 ( .A1(n10734), .A2(n10733), .ZN(n10735) );
  AND2_X1 U13331 ( .A1(n10736), .A2(n10735), .ZN(n10743) );
  INV_X1 U13332 ( .A(n13204), .ZN(n15252) );
  AOI22_X1 U13333 ( .A1(n13059), .A2(n15244), .B1(n15242), .B2(n12652), .ZN(
        n10742) );
  AND2_X1 U13334 ( .A1(n10916), .A2(n10738), .ZN(n10740) );
  OAI211_X1 U13335 ( .C1(n10740), .C2(n12766), .A(n10739), .B(n15248), .ZN(
        n10741) );
  OAI211_X1 U13336 ( .C1(n10743), .C2(n15252), .A(n10742), .B(n10741), .ZN(
        n15280) );
  INV_X1 U13337 ( .A(n15280), .ZN(n10750) );
  INV_X1 U13338 ( .A(n10743), .ZN(n15282) );
  AND2_X1 U13339 ( .A1(n13344), .A2(n15255), .ZN(n13210) );
  OR2_X1 U13340 ( .A1(n15240), .A2(n15295), .ZN(n10744) );
  INV_X1 U13341 ( .A(n10746), .ZN(n11125) );
  AOI22_X1 U13342 ( .A1(n13322), .A2(n11126), .B1(n13288), .B2(n11125), .ZN(
        n10747) );
  OAI21_X1 U13343 ( .B1(n10446), .B2(n13344), .A(n10747), .ZN(n10748) );
  AOI21_X1 U13344 ( .B1(n15282), .B2(n13210), .A(n10748), .ZN(n10749) );
  OAI21_X1 U13345 ( .B1(n10750), .B2(n13328), .A(n10749), .ZN(P3_U3227) );
  OAI21_X1 U13346 ( .B1(n10752), .B2(n8497), .A(n10751), .ZN(n11402) );
  AOI211_X1 U13347 ( .C1(n12331), .C2(n10753), .A(n14909), .B(n10879), .ZN(
        n11409) );
  XOR2_X1 U13348 ( .A(n10754), .B(n12518), .Z(n10755) );
  AOI22_X1 U13349 ( .A1(n14153), .A2(n14110), .B1(n14111), .B2(n14155), .ZN(
        n11146) );
  OAI21_X1 U13350 ( .B1(n10755), .B2(n14921), .A(n11146), .ZN(n11403) );
  AOI211_X1 U13351 ( .C1(n14918), .C2(n11402), .A(n11409), .B(n11403), .ZN(
        n10761) );
  INV_X1 U13352 ( .A(n12331), .ZN(n11406) );
  INV_X1 U13353 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10756) );
  OAI22_X1 U13354 ( .A1(n14643), .A2(n11406), .B1(n14987), .B2(n10756), .ZN(
        n10757) );
  INV_X1 U13355 ( .A(n10757), .ZN(n10758) );
  OAI21_X1 U13356 ( .B1(n10761), .B2(n14985), .A(n10758), .ZN(P1_U3474) );
  OAI22_X1 U13357 ( .A1(n14596), .A2(n11406), .B1(n14994), .B2(n10020), .ZN(
        n10759) );
  INV_X1 U13358 ( .A(n10759), .ZN(n10760) );
  OAI21_X1 U13359 ( .B1(n10761), .B2(n14991), .A(n10760), .ZN(P1_U3533) );
  OAI22_X1 U13360 ( .A1(n12809), .A2(P3_U3151), .B1(SI_22_), .B2(n12584), .ZN(
        n10762) );
  AOI21_X1 U13361 ( .B1(n10763), .B2(n10995), .A(n10762), .ZN(P3_U3273) );
  INV_X1 U13362 ( .A(n10764), .ZN(n10773) );
  AND2_X1 U13363 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n15024) );
  AOI21_X1 U13364 ( .B1(n13515), .B2(n10765), .A(n15024), .ZN(n10766) );
  OAI21_X1 U13365 ( .B1(n13539), .B2(n7069), .A(n10766), .ZN(n10772) );
  INV_X1 U13366 ( .A(n13561), .ZN(n13501) );
  AOI22_X1 U13367 ( .A1(n13501), .A2(n13604), .B1(n13552), .B2(n10767), .ZN(
        n10770) );
  INV_X1 U13368 ( .A(n13548), .ZN(n10769) );
  NOR3_X1 U13369 ( .A1(n10770), .A2(n10769), .A3(n10768), .ZN(n10771) );
  AOI211_X1 U13370 ( .C1(n13546), .C2(n10773), .A(n10772), .B(n10771), .ZN(
        n10774) );
  OAI21_X1 U13371 ( .B1(n10775), .B2(n14999), .A(n10774), .ZN(P2_U3199) );
  XNOR2_X1 U13372 ( .A(n10776), .B(n12650), .ZN(n15285) );
  NAND2_X1 U13373 ( .A1(n15285), .A2(n13204), .ZN(n10781) );
  XNOR2_X1 U13374 ( .A(n10777), .B(n12650), .ZN(n10779) );
  OAI22_X1 U13375 ( .A1(n10918), .A2(n13314), .B1(n11072), .B2(n13312), .ZN(
        n10778) );
  AOI21_X1 U13376 ( .B1(n10779), .B2(n15248), .A(n10778), .ZN(n10780) );
  AND2_X1 U13377 ( .A1(n10781), .A2(n10780), .ZN(n15287) );
  INV_X1 U13378 ( .A(n10782), .ZN(n12819) );
  AOI22_X1 U13379 ( .A1(n13322), .A2(n12818), .B1(n13288), .B2(n12819), .ZN(
        n10783) );
  OAI21_X1 U13380 ( .B1(n10464), .B2(n13344), .A(n10783), .ZN(n10784) );
  AOI21_X1 U13381 ( .B1(n15285), .B2(n13210), .A(n10784), .ZN(n10785) );
  OAI21_X1 U13382 ( .B1(n15287), .B2(n15258), .A(n10785), .ZN(P3_U3226) );
  INV_X1 U13383 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n15633) );
  NAND2_X1 U13384 ( .A1(n13250), .A2(P3_U3897), .ZN(n10786) );
  OAI21_X1 U13385 ( .B1(P3_U3897), .B2(n15633), .A(n10786), .ZN(P3_U3516) );
  AOI21_X1 U13386 ( .B1(n10564), .B2(n10788), .A(n10787), .ZN(n10791) );
  INV_X1 U13387 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10789) );
  MUX2_X1 U13388 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10789), .S(n10794), .Z(
        n10790) );
  NAND2_X1 U13389 ( .A1(n10791), .A2(n10790), .ZN(n11055) );
  INV_X1 U13390 ( .A(n14295), .ZN(n14874) );
  OAI211_X1 U13391 ( .C1(n10791), .C2(n10790), .A(n11055), .B(n14874), .ZN(
        n10802) );
  OAI21_X1 U13392 ( .B1(n10793), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10792), 
        .ZN(n10796) );
  INV_X1 U13393 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11624) );
  MUX2_X1 U13394 ( .A(n11624), .B(P1_REG2_REG_13__SCAN_IN), .S(n10794), .Z(
        n10795) );
  INV_X1 U13395 ( .A(n14299), .ZN(n14871) );
  NOR2_X1 U13396 ( .A1(n10796), .A2(n10795), .ZN(n11067) );
  AOI211_X1 U13397 ( .C1(n10796), .C2(n10795), .A(n14871), .B(n11067), .ZN(
        n10800) );
  NAND2_X1 U13398 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14075)
         );
  INV_X1 U13399 ( .A(n14075), .ZN(n10797) );
  AOI21_X1 U13400 ( .B1(n14255), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10797), 
        .ZN(n10798) );
  OAI21_X1 U13401 ( .B1(n14870), .B2(n11060), .A(n10798), .ZN(n10799) );
  NOR2_X1 U13402 ( .A1(n10800), .A2(n10799), .ZN(n10801) );
  NAND2_X1 U13403 ( .A1(n10802), .A2(n10801), .ZN(P1_U3256) );
  OR2_X1 U13404 ( .A1(n10804), .A2(n10803), .ZN(n10805) );
  NAND2_X1 U13405 ( .A1(n10806), .A2(n10805), .ZN(n15269) );
  INV_X1 U13406 ( .A(n15269), .ZN(n10817) );
  INV_X1 U13407 ( .A(n13210), .ZN(n13225) );
  AOI21_X1 U13408 ( .B1(n15245), .B2(n10807), .A(n12767), .ZN(n10813) );
  NAND2_X1 U13409 ( .A1(n10808), .A2(n15248), .ZN(n10812) );
  NAND2_X1 U13410 ( .A1(n15269), .A2(n13204), .ZN(n10811) );
  AOI22_X1 U13411 ( .A1(n10809), .A2(n15244), .B1(n15242), .B2(n12956), .ZN(
        n10810) );
  OAI211_X1 U13412 ( .C1(n10813), .C2(n10812), .A(n10811), .B(n10810), .ZN(
        n15267) );
  MUX2_X1 U13413 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n15267), .S(n13344), .Z(
        n10814) );
  INV_X1 U13414 ( .A(n10814), .ZN(n10816) );
  AOI22_X1 U13415 ( .A1(n13322), .A2(n12885), .B1(n13288), .B2(n12886), .ZN(
        n10815) );
  OAI211_X1 U13416 ( .C1(n10817), .C2(n13225), .A(n10816), .B(n10815), .ZN(
        P3_U3230) );
  OAI21_X1 U13417 ( .B1(n10819), .B2(n10821), .A(n10818), .ZN(n15121) );
  INV_X1 U13418 ( .A(n15121), .ZN(n10826) );
  XOR2_X1 U13419 ( .A(n10821), .B(n10820), .Z(n10823) );
  AOI21_X1 U13420 ( .B1(n10823), .B2(n15131), .A(n10822), .ZN(n15124) );
  AOI211_X1 U13421 ( .C1(n15117), .C2(n10824), .A(n12009), .B(n11096), .ZN(
        n15113) );
  AOI21_X1 U13422 ( .B1(n15196), .B2(n15117), .A(n15113), .ZN(n10825) );
  OAI211_X1 U13423 ( .C1(n15187), .C2(n10826), .A(n15124), .B(n10825), .ZN(
        n10874) );
  NAND2_X1 U13424 ( .A1(n10874), .A2(n15233), .ZN(n10827) );
  OAI21_X1 U13425 ( .B1(n15233), .B2(n9924), .A(n10827), .ZN(P2_U3506) );
  AOI21_X1 U13426 ( .B1(n10386), .B2(n10834), .A(n10828), .ZN(n10830) );
  INV_X1 U13427 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n15546) );
  AOI22_X1 U13428 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n10832), .B1(n11436), 
        .B2(n15546), .ZN(n10829) );
  NOR2_X1 U13429 ( .A1(n10830), .A2(n10829), .ZN(n11426) );
  AOI21_X1 U13430 ( .B1(n10830), .B2(n10829), .A(n11426), .ZN(n10841) );
  INV_X1 U13431 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10831) );
  NAND2_X1 U13432 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n12572)
         );
  OAI21_X1 U13433 ( .B1(n15111), .B2(n10831), .A(n12572), .ZN(n10839) );
  AOI22_X1 U13434 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n10832), .B1(n11436), 
        .B2(n9187), .ZN(n10836) );
  OAI21_X1 U13435 ( .B1(n10834), .B2(n10379), .A(n10833), .ZN(n10835) );
  NOR2_X1 U13436 ( .A1(n10836), .A2(n10835), .ZN(n11438) );
  AOI21_X1 U13437 ( .B1(n10836), .B2(n10835), .A(n11438), .ZN(n10837) );
  NOR2_X1 U13438 ( .A1(n10837), .A2(n15103), .ZN(n10838) );
  AOI211_X1 U13439 ( .C1(n15089), .C2(n11436), .A(n10839), .B(n10838), .ZN(
        n10840) );
  OAI21_X1 U13440 ( .B1(n10841), .B2(n15105), .A(n10840), .ZN(P2_U3226) );
  OR2_X1 U13441 ( .A1(n10842), .A2(n12771), .ZN(n10843) );
  NAND2_X1 U13442 ( .A1(n10844), .A2(n10843), .ZN(n15273) );
  OAI22_X1 U13443 ( .A1(n13341), .A2(n15270), .B1(n10845), .B2(n15238), .ZN(
        n10854) );
  XNOR2_X1 U13444 ( .A(n10847), .B(n10846), .ZN(n10852) );
  NAND2_X1 U13445 ( .A1(n15273), .A2(n13204), .ZN(n10851) );
  OAI22_X1 U13446 ( .A1(n11117), .A2(n13312), .B1(n10848), .B2(n13314), .ZN(
        n10849) );
  INV_X1 U13447 ( .A(n10849), .ZN(n10850) );
  OAI211_X1 U13448 ( .C1(n10852), .C2(n13310), .A(n10851), .B(n10850), .ZN(
        n15271) );
  MUX2_X1 U13449 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15271), .S(n13344), .Z(
        n10853) );
  AOI211_X1 U13450 ( .C1(n13210), .C2(n15273), .A(n10854), .B(n10853), .ZN(
        n10855) );
  INV_X1 U13451 ( .A(n10855), .ZN(P3_U3229) );
  XNOR2_X1 U13452 ( .A(n10856), .B(n10858), .ZN(n10869) );
  OAI21_X1 U13453 ( .B1(n10859), .B2(n10858), .A(n10857), .ZN(n10863) );
  OAI22_X1 U13454 ( .A1(n10861), .A2(n13567), .B1(n10860), .B2(n15148), .ZN(
        n10862) );
  AOI21_X1 U13455 ( .B1(n10863), .B2(n15131), .A(n10862), .ZN(n10864) );
  OAI21_X1 U13456 ( .B1(n10869), .B2(n15201), .A(n10864), .ZN(n15192) );
  MUX2_X1 U13457 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n15192), .S(n15155), .Z(
        n10873) );
  INV_X1 U13458 ( .A(n13835), .ZN(n15140) );
  OAI211_X1 U13459 ( .C1(n10866), .C2(n15191), .A(n15134), .B(n10865), .ZN(
        n15190) );
  OAI22_X1 U13460 ( .A1(n13813), .A2(n15191), .B1(n13544), .B2(n15132), .ZN(
        n10867) );
  INV_X1 U13461 ( .A(n10867), .ZN(n10871) );
  INV_X1 U13462 ( .A(n6875), .ZN(n10868) );
  AND2_X1 U13463 ( .A1(n15155), .A2(n10868), .ZN(n11109) );
  INV_X1 U13464 ( .A(n10869), .ZN(n15194) );
  NAND2_X1 U13465 ( .A1(n11109), .A2(n15194), .ZN(n10870) );
  OAI211_X1 U13466 ( .C1(n15140), .C2(n15190), .A(n10871), .B(n10870), .ZN(
        n10872) );
  OR2_X1 U13467 ( .A1(n10873), .A2(n10872), .ZN(P2_U3261) );
  INV_X1 U13468 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U13469 ( .A1(n10874), .A2(n15212), .ZN(n10875) );
  OAI21_X1 U13470 ( .B1(n15212), .B2(n10876), .A(n10875), .ZN(P2_U3451) );
  OAI21_X1 U13471 ( .B1(n10878), .B2(n10881), .A(n10877), .ZN(n11367) );
  INV_X1 U13472 ( .A(n10879), .ZN(n10880) );
  AOI211_X1 U13473 ( .C1(n12343), .C2(n10880), .A(n14909), .B(n11045), .ZN(
        n11373) );
  XNOR2_X1 U13474 ( .A(n10882), .B(n10881), .ZN(n10885) );
  NAND2_X1 U13475 ( .A1(n14154), .A2(n14111), .ZN(n10884) );
  NAND2_X1 U13476 ( .A1(n14152), .A2(n14110), .ZN(n10883) );
  AND2_X1 U13477 ( .A1(n10884), .A2(n10883), .ZN(n11284) );
  OAI21_X1 U13478 ( .B1(n10885), .B2(n14921), .A(n11284), .ZN(n11368) );
  AOI211_X1 U13479 ( .C1(n14918), .C2(n11367), .A(n11373), .B(n11368), .ZN(
        n10891) );
  OAI22_X1 U13480 ( .A1(n14596), .A2(n12348), .B1(n14994), .B2(n10021), .ZN(
        n10886) );
  INV_X1 U13481 ( .A(n10886), .ZN(n10887) );
  OAI21_X1 U13482 ( .B1(n10891), .B2(n14991), .A(n10887), .ZN(P1_U3534) );
  INV_X1 U13483 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10888) );
  OAI22_X1 U13484 ( .A1(n14643), .A2(n12348), .B1(n14987), .B2(n10888), .ZN(
        n10889) );
  INV_X1 U13485 ( .A(n10889), .ZN(n10890) );
  OAI21_X1 U13486 ( .B1(n10891), .B2(n14985), .A(n10890), .ZN(P1_U3477) );
  XNOR2_X1 U13487 ( .A(n10892), .B(n10894), .ZN(n11031) );
  XNOR2_X1 U13488 ( .A(n10893), .B(n10894), .ZN(n10896) );
  AOI22_X1 U13489 ( .A1(n15127), .A2(n13600), .B1(n13597), .B2(n15128), .ZN(
        n10895) );
  OAI21_X1 U13490 ( .B1(n10896), .B2(n11793), .A(n10895), .ZN(n10897) );
  AOI21_X1 U13491 ( .B1(n15146), .B2(n11031), .A(n10897), .ZN(n11035) );
  INV_X1 U13492 ( .A(n10987), .ZN(n10898) );
  AOI211_X1 U13493 ( .C1(n11033), .C2(n11095), .A(n12009), .B(n10898), .ZN(
        n11032) );
  NOR2_X1 U13494 ( .A1(n7073), .A2(n13813), .ZN(n10901) );
  OAI22_X1 U13495 ( .A1(n15155), .A2(n10899), .B1(n12119), .B2(n15132), .ZN(
        n10900) );
  AOI211_X1 U13496 ( .C1(n11032), .C2(n13835), .A(n10901), .B(n10900), .ZN(
        n10903) );
  NAND2_X1 U13497 ( .A1(n11031), .A2(n11109), .ZN(n10902) );
  OAI211_X1 U13498 ( .C1(n11035), .C2(n15157), .A(n10903), .B(n10902), .ZN(
        P2_U3256) );
  OAI222_X1 U13499 ( .A1(n12562), .A2(n10904), .B1(n6656), .B2(n10905), .C1(
        n12498), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI222_X1 U13500 ( .A1(n13960), .A2(n10907), .B1(P2_U3088), .B2(n10906), 
        .C1(n13955), .C2(n10905), .ZN(P2_U3307) );
  MUX2_X1 U13501 ( .A(n10909), .B(n10908), .S(n15258), .Z(n10911) );
  NAND2_X1 U13502 ( .A1(n13288), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10910) );
  OAI211_X1 U13503 ( .C1(n10912), .C2(n13341), .A(n10911), .B(n10910), .ZN(
        P3_U3233) );
  XNOR2_X1 U13504 ( .A(n10913), .B(n12775), .ZN(n15275) );
  INV_X1 U13505 ( .A(n15275), .ZN(n10927) );
  NAND2_X1 U13506 ( .A1(n15275), .A2(n13204), .ZN(n10922) );
  NAND2_X1 U13507 ( .A1(n10914), .A2(n12775), .ZN(n10915) );
  NAND2_X1 U13508 ( .A1(n10916), .A2(n10915), .ZN(n10920) );
  NAND2_X1 U13509 ( .A1(n12956), .A2(n15244), .ZN(n10917) );
  OAI21_X1 U13510 ( .B1(n10918), .B2(n13312), .A(n10917), .ZN(n10919) );
  AOI21_X1 U13511 ( .B1(n10920), .B2(n15248), .A(n10919), .ZN(n10921) );
  AND2_X1 U13512 ( .A1(n10922), .A2(n10921), .ZN(n15277) );
  MUX2_X1 U13513 ( .A(n15277), .B(n10923), .S(n15258), .Z(n10926) );
  INV_X1 U13514 ( .A(n10924), .ZN(n12957) );
  AOI22_X1 U13515 ( .A1(n13322), .A2(n15274), .B1(n13288), .B2(n12957), .ZN(
        n10925) );
  OAI211_X1 U13516 ( .C1(n10927), .C2(n13225), .A(n10926), .B(n10925), .ZN(
        P3_U3228) );
  INV_X2 U13517 ( .A(n10928), .ZN(n12033) );
  NAND2_X1 U13518 ( .A1(n13600), .A2(n12009), .ZN(n11001) );
  XNOR2_X1 U13519 ( .A(n12112), .B(n11001), .ZN(n10931) );
  NAND2_X1 U13520 ( .A1(n11006), .A2(n10999), .ZN(n12117) );
  OAI21_X1 U13521 ( .B1(n10931), .B2(n11006), .A(n12117), .ZN(n10938) );
  NOR3_X1 U13522 ( .A1(n10931), .A2(n10930), .A3(n13561), .ZN(n10932) );
  AND2_X1 U13523 ( .A1(n13515), .A2(n15127), .ZN(n13541) );
  OAI21_X1 U13524 ( .B1(n10932), .B2(n13541), .A(n13601), .ZN(n10936) );
  NAND2_X1 U13525 ( .A1(n13515), .A2(n15128), .ZN(n11023) );
  INV_X1 U13526 ( .A(n11023), .ZN(n13547) );
  OAI21_X1 U13527 ( .B1(n15007), .B2(n11097), .A(n10933), .ZN(n10934) );
  AOI21_X1 U13528 ( .B1(n13547), .B2(n13598), .A(n10934), .ZN(n10935) );
  OAI211_X1 U13529 ( .C1(n15208), .C2(n13539), .A(n10936), .B(n10935), .ZN(
        n10937) );
  AOI21_X1 U13530 ( .B1(n13552), .B2(n10938), .A(n10937), .ZN(n10939) );
  INV_X1 U13531 ( .A(n10939), .ZN(P2_U3193) );
  OAI22_X1 U13532 ( .A1(n10622), .A2(n10942), .B1(n11331), .B2(n12274), .ZN(
        n11138) );
  OAI22_X1 U13533 ( .A1(n10942), .A2(n12274), .B1(n11331), .B2(n12275), .ZN(
        n10943) );
  XNOR2_X1 U13534 ( .A(n10943), .B(n12265), .ZN(n10944) );
  NAND2_X1 U13535 ( .A1(n10945), .A2(n10944), .ZN(n11141) );
  OAI211_X1 U13536 ( .C1(n10945), .C2(n10944), .A(n11141), .B(n14828), .ZN(
        n10949) );
  NAND2_X1 U13537 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14204) );
  OAI21_X1 U13538 ( .B1(n14121), .B2(n10946), .A(n14204), .ZN(n10947) );
  AOI21_X1 U13539 ( .B1(n12327), .B2(n6638), .A(n10947), .ZN(n10948) );
  OAI211_X1 U13540 ( .C1(n14836), .C2(n11330), .A(n10949), .B(n10948), .ZN(
        P1_U3230) );
  AOI21_X1 U13541 ( .B1(n10952), .B2(n10950), .A(n11209), .ZN(n10972) );
  INV_X1 U13542 ( .A(n10951), .ZN(n10958) );
  MUX2_X1 U13543 ( .A(n10953), .B(n10952), .S(n12105), .Z(n10954) );
  NAND2_X1 U13544 ( .A1(n10954), .A2(n7313), .ZN(n11230) );
  INV_X1 U13545 ( .A(n10954), .ZN(n10955) );
  NAND2_X1 U13546 ( .A1(n10955), .A2(n10964), .ZN(n10956) );
  AND2_X1 U13547 ( .A1(n11230), .A2(n10956), .ZN(n10957) );
  INV_X1 U13548 ( .A(n11231), .ZN(n10961) );
  NOR3_X1 U13549 ( .A1(n10959), .A2(n10958), .A3(n10957), .ZN(n10960) );
  OAI21_X1 U13550 ( .B1(n10961), .B2(n10960), .A(n13132), .ZN(n10971) );
  NOR2_X1 U13551 ( .A1(n10953), .A2(n10965), .ZN(n11215) );
  AOI21_X1 U13552 ( .B1(n10953), .B2(n10965), .A(n11215), .ZN(n10968) );
  NOR2_X1 U13553 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15587), .ZN(n12987) );
  AOI21_X1 U13554 ( .B1(n15234), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12987), .ZN(
        n10967) );
  NAND2_X1 U13555 ( .A1(n13166), .A2(n7313), .ZN(n10966) );
  OAI211_X1 U13556 ( .C1(n10968), .C2(n13150), .A(n10967), .B(n10966), .ZN(
        n10969) );
  INV_X1 U13557 ( .A(n10969), .ZN(n10970) );
  OAI211_X1 U13558 ( .C1(n10972), .C2(n13165), .A(n10971), .B(n10970), .ZN(
        P3_U3191) );
  INV_X1 U13559 ( .A(n10973), .ZN(n10976) );
  OAI222_X1 U13560 ( .A1(n12562), .A2(n10974), .B1(n6656), .B2(n10976), .C1(
        P1_U3086), .C2(n14301), .ZN(P1_U3336) );
  OAI222_X1 U13561 ( .A1(n13960), .A2(n10977), .B1(n13955), .B2(n10976), .C1(
        n10975), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U13562 ( .A(n10979), .B(n10978), .ZN(n15219) );
  NAND2_X1 U13563 ( .A1(n15219), .A2(n15146), .ZN(n10986) );
  XNOR2_X1 U13564 ( .A(n10980), .B(n10981), .ZN(n10984) );
  NAND2_X1 U13565 ( .A1(n13596), .A2(n15128), .ZN(n10983) );
  NAND2_X1 U13566 ( .A1(n13598), .A2(n15127), .ZN(n10982) );
  NAND2_X1 U13567 ( .A1(n10983), .A2(n10982), .ZN(n11080) );
  AOI21_X1 U13568 ( .B1(n10984), .B2(n15131), .A(n11080), .ZN(n10985) );
  AND2_X1 U13569 ( .A1(n10986), .A2(n10985), .ZN(n15221) );
  AOI21_X1 U13570 ( .B1(n15213), .B2(n10987), .A(n13753), .ZN(n10989) );
  NAND2_X1 U13571 ( .A1(n10989), .A2(n11165), .ZN(n15214) );
  INV_X1 U13572 ( .A(n13813), .ZN(n15144) );
  OAI22_X1 U13573 ( .A1(n15155), .A2(n10990), .B1(n11083), .B2(n15132), .ZN(
        n10991) );
  AOI21_X1 U13574 ( .B1(n15213), .B2(n15144), .A(n10991), .ZN(n10992) );
  OAI21_X1 U13575 ( .B1(n15214), .B2(n15140), .A(n10992), .ZN(n10993) );
  AOI21_X1 U13576 ( .B1(n15219), .B2(n11109), .A(n10993), .ZN(n10994) );
  OAI21_X1 U13577 ( .B1(n15221), .B2(n15157), .A(n10994), .ZN(P2_U3255) );
  NAND2_X1 U13578 ( .A1(n10996), .A2(n10995), .ZN(n10997) );
  OAI211_X1 U13579 ( .C1(n10998), .C2(n12584), .A(n10997), .B(n12812), .ZN(
        P3_U3272) );
  INV_X2 U13580 ( .A(n15134), .ZN(n12009) );
  NAND2_X1 U13581 ( .A1(n13598), .A2(n12009), .ZN(n11008) );
  XNOR2_X1 U13582 ( .A(n11007), .B(n11008), .ZN(n11000) );
  AND2_X1 U13583 ( .A1(n10999), .A2(n11000), .ZN(n11005) );
  INV_X1 U13584 ( .A(n11000), .ZN(n12116) );
  INV_X1 U13585 ( .A(n12112), .ZN(n11002) );
  NAND2_X1 U13586 ( .A1(n11002), .A2(n11001), .ZN(n11003) );
  AOI21_X2 U13587 ( .B1(n11006), .B2(n11005), .A(n11004), .ZN(n12126) );
  INV_X1 U13588 ( .A(n11007), .ZN(n11009) );
  NAND2_X1 U13589 ( .A1(n11009), .A2(n11008), .ZN(n11010) );
  XNOR2_X1 U13590 ( .A(n15213), .B(n12033), .ZN(n11011) );
  AND2_X1 U13591 ( .A1(n13597), .A2(n13753), .ZN(n11012) );
  NAND2_X1 U13592 ( .A1(n11011), .A2(n11012), .ZN(n11016) );
  INV_X1 U13593 ( .A(n11011), .ZN(n11025) );
  INV_X1 U13594 ( .A(n11012), .ZN(n11013) );
  NAND2_X1 U13595 ( .A1(n11025), .A2(n11013), .ZN(n11014) );
  NAND2_X1 U13596 ( .A1(n11016), .A2(n11014), .ZN(n11086) );
  INV_X1 U13597 ( .A(n11017), .ZN(n11084) );
  NAND2_X1 U13598 ( .A1(n13596), .A2(n12009), .ZN(n11490) );
  INV_X1 U13599 ( .A(n11026), .ZN(n11018) );
  INV_X1 U13600 ( .A(n11493), .ZN(n12578) );
  AOI21_X1 U13601 ( .B1(n11084), .B2(n11018), .A(n12578), .ZN(n11030) );
  INV_X1 U13602 ( .A(n11019), .ZN(n11166) );
  NAND2_X1 U13603 ( .A1(n13546), .A2(n11166), .ZN(n11020) );
  OAI211_X1 U13604 ( .C1(n11023), .C2(n11022), .A(n11021), .B(n11020), .ZN(
        n11024) );
  AOI21_X1 U13605 ( .B1(n11200), .B2(n15004), .A(n11024), .ZN(n11029) );
  NOR3_X1 U13606 ( .A1(n11026), .A2(n11025), .A3(n13561), .ZN(n11027) );
  OAI21_X1 U13607 ( .B1(n11027), .B2(n13541), .A(n13597), .ZN(n11028) );
  OAI211_X1 U13608 ( .C1(n11030), .C2(n14999), .A(n11029), .B(n11028), .ZN(
        P2_U3208) );
  INV_X1 U13609 ( .A(n11031), .ZN(n11036) );
  AOI21_X1 U13610 ( .B1(n15196), .B2(n11033), .A(n11032), .ZN(n11034) );
  OAI211_X1 U13611 ( .C1(n11036), .C2(n15200), .A(n11035), .B(n11034), .ZN(
        n11038) );
  NAND2_X1 U13612 ( .A1(n11038), .A2(n15233), .ZN(n11037) );
  OAI21_X1 U13613 ( .B1(n15233), .B2(n9926), .A(n11037), .ZN(P2_U3508) );
  NAND2_X1 U13614 ( .A1(n11038), .A2(n15212), .ZN(n11039) );
  OAI21_X1 U13615 ( .B1(n15212), .B2(n9126), .A(n11039), .ZN(P2_U3457) );
  INV_X1 U13616 ( .A(n12489), .ZN(n12510) );
  OAI222_X1 U13617 ( .A1(n12562), .A2(n11040), .B1(n6656), .B2(n11134), .C1(
        n12510), .C2(P1_U3086), .ZN(P1_U3334) );
  NAND2_X1 U13618 ( .A1(n13060), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11041) );
  OAI21_X1 U13619 ( .B1(n12608), .B2(n13060), .A(n11041), .ZN(P3_U3521) );
  NAND2_X1 U13620 ( .A1(n13060), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11042) );
  OAI21_X1 U13621 ( .B1(n12909), .B2(n13060), .A(n11042), .ZN(P3_U3520) );
  OAI21_X1 U13622 ( .B1(n11044), .B2(n12522), .A(n11043), .ZN(n11392) );
  INV_X1 U13623 ( .A(n11045), .ZN(n11046) );
  AOI211_X1 U13624 ( .C1(n12342), .C2(n11046), .A(n14909), .B(n6652), .ZN(
        n11398) );
  XNOR2_X1 U13625 ( .A(n11047), .B(n12522), .ZN(n11048) );
  AOI22_X1 U13626 ( .A1(n14153), .A2(n14111), .B1(n14110), .B2(n14151), .ZN(
        n11294) );
  OAI21_X1 U13627 ( .B1(n11048), .B2(n14921), .A(n11294), .ZN(n11393) );
  AOI211_X1 U13628 ( .C1(n14918), .C2(n11392), .A(n11398), .B(n11393), .ZN(
        n11054) );
  OAI22_X1 U13629 ( .A1(n14596), .A2(n12340), .B1(n14994), .B2(n10023), .ZN(
        n11049) );
  INV_X1 U13630 ( .A(n11049), .ZN(n11050) );
  OAI21_X1 U13631 ( .B1(n11054), .B2(n14991), .A(n11050), .ZN(P1_U3535) );
  INV_X1 U13632 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11051) );
  OAI22_X1 U13633 ( .A1(n14643), .A2(n12340), .B1(n14987), .B2(n11051), .ZN(
        n11052) );
  INV_X1 U13634 ( .A(n11052), .ZN(n11053) );
  OAI21_X1 U13635 ( .B1(n11054), .B2(n14985), .A(n11053), .ZN(P1_U3480) );
  MUX2_X1 U13636 ( .A(n11775), .B(P1_REG1_REG_14__SCAN_IN), .S(n11063), .Z(
        n11057) );
  OAI21_X1 U13637 ( .B1(n10789), .B2(n11060), .A(n11055), .ZN(n11056) );
  AOI21_X1 U13638 ( .B1(n11057), .B2(n11056), .A(n11774), .ZN(n11070) );
  NAND2_X1 U13639 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14833)
         );
  INV_X1 U13640 ( .A(n14833), .ZN(n11059) );
  NOR2_X1 U13641 ( .A1(n14870), .A2(n11782), .ZN(n11058) );
  AOI211_X1 U13642 ( .C1(n14255), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n11059), 
        .B(n11058), .ZN(n11069) );
  MUX2_X1 U13643 ( .A(n11783), .B(P1_REG2_REG_14__SCAN_IN), .S(n11063), .Z(
        n11062) );
  NOR2_X1 U13644 ( .A1(n11060), .A2(n11624), .ZN(n11065) );
  INV_X1 U13645 ( .A(n11065), .ZN(n11061) );
  NAND2_X1 U13646 ( .A1(n11062), .A2(n11061), .ZN(n11066) );
  MUX2_X1 U13647 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11783), .S(n11063), .Z(
        n11064) );
  OAI21_X1 U13648 ( .B1(n11067), .B2(n11065), .A(n11064), .ZN(n11781) );
  OAI211_X1 U13649 ( .C1(n11067), .C2(n11066), .A(n11781), .B(n14299), .ZN(
        n11068) );
  OAI211_X1 U13650 ( .C1(n11070), .C2(n14295), .A(n11069), .B(n11068), .ZN(
        P1_U3257) );
  AOI21_X1 U13651 ( .B1(n11071), .B2(n12774), .A(n13310), .ZN(n11075) );
  OAI22_X1 U13652 ( .A1(n11072), .A2(n13314), .B1(n11744), .B2(n13312), .ZN(
        n11073) );
  AOI21_X1 U13653 ( .B1(n11075), .B2(n11074), .A(n11073), .ZN(n15294) );
  OAI22_X1 U13654 ( .A1(n13341), .A2(n15296), .B1(n12989), .B2(n15238), .ZN(
        n11076) );
  AOI21_X1 U13655 ( .B1(n15258), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11076), .ZN(
        n11079) );
  XNOR2_X1 U13656 ( .A(n11077), .B(n12774), .ZN(n15299) );
  NAND2_X1 U13657 ( .A1(n15299), .A2(n13347), .ZN(n11078) );
  OAI211_X1 U13658 ( .C1(n15294), .C2(n15258), .A(n11079), .B(n11078), .ZN(
        P3_U3224) );
  NAND2_X1 U13659 ( .A1(n13515), .A2(n11080), .ZN(n11082) );
  OAI211_X1 U13660 ( .C1(n15007), .C2(n11083), .A(n11082), .B(n11081), .ZN(
        n11088) );
  AOI211_X1 U13661 ( .C1(n11086), .C2(n11085), .A(n14999), .B(n11084), .ZN(
        n11087) );
  AOI211_X1 U13662 ( .C1(n15213), .C2(n15004), .A(n11088), .B(n11087), .ZN(
        n11089) );
  INV_X1 U13663 ( .A(n11089), .ZN(P2_U3189) );
  NAND2_X1 U13664 ( .A1(n10818), .A2(n11090), .ZN(n11092) );
  NAND2_X1 U13665 ( .A1(n11092), .A2(n11091), .ZN(n11093) );
  NAND2_X1 U13666 ( .A1(n11094), .A2(n11093), .ZN(n11106) );
  INV_X1 U13667 ( .A(n11106), .ZN(n15211) );
  OAI211_X1 U13668 ( .C1(n15208), .C2(n11096), .A(n15134), .B(n11095), .ZN(
        n15207) );
  INV_X1 U13669 ( .A(n11097), .ZN(n11098) );
  AOI22_X1 U13670 ( .A1(n15144), .A2(n11099), .B1(n11098), .B2(n15154), .ZN(
        n11100) );
  OAI21_X1 U13671 ( .B1(n15207), .B2(n15140), .A(n11100), .ZN(n11108) );
  AOI22_X1 U13672 ( .A1(n15127), .A2(n13601), .B1(n13598), .B2(n15128), .ZN(
        n11105) );
  XNOR2_X1 U13673 ( .A(n11102), .B(n11101), .ZN(n11103) );
  NAND2_X1 U13674 ( .A1(n11103), .A2(n15131), .ZN(n11104) );
  OAI211_X1 U13675 ( .C1(n11106), .C2(n15201), .A(n11105), .B(n11104), .ZN(
        n15209) );
  MUX2_X1 U13676 ( .A(n15209), .B(P2_REG2_REG_8__SCAN_IN), .S(n15157), .Z(
        n11107) );
  AOI211_X1 U13677 ( .C1(n15211), .C2(n11109), .A(n11108), .B(n11107), .ZN(
        n11110) );
  INV_X1 U13678 ( .A(n11110), .ZN(P2_U3257) );
  XNOR2_X1 U13679 ( .A(n12903), .B(n15279), .ZN(n11236) );
  XNOR2_X1 U13680 ( .A(n11236), .B(n13058), .ZN(n11124) );
  NAND2_X1 U13681 ( .A1(n11112), .A2(n11111), .ZN(n11113) );
  XNOR2_X1 U13682 ( .A(n12903), .B(n11115), .ZN(n11116) );
  XNOR2_X1 U13683 ( .A(n11116), .B(n11117), .ZN(n12952) );
  NAND2_X1 U13684 ( .A1(n12953), .A2(n12952), .ZN(n11120) );
  INV_X1 U13685 ( .A(n11116), .ZN(n11118) );
  NAND2_X1 U13686 ( .A1(n11118), .A2(n11117), .ZN(n11119) );
  INV_X1 U13687 ( .A(n11238), .ZN(n11122) );
  AOI211_X1 U13688 ( .C1(n11124), .C2(n11123), .A(n13046), .B(n11122), .ZN(
        n11132) );
  NAND2_X1 U13689 ( .A1(n13038), .A2(n11125), .ZN(n11130) );
  AOI22_X1 U13690 ( .A1(n13044), .A2(n11126), .B1(n13017), .B2(n13059), .ZN(
        n11129) );
  NAND2_X1 U13691 ( .A1(n13037), .A2(n12652), .ZN(n11127) );
  NAND4_X1 U13692 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(
        n11131) );
  OR2_X1 U13693 ( .A1(n11132), .A2(n11131), .ZN(P3_U3179) );
  INV_X1 U13694 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n15571) );
  NAND2_X1 U13695 ( .A1(n6908), .A2(P3_U3897), .ZN(n11133) );
  OAI21_X1 U13696 ( .B1(P3_U3897), .B2(n15571), .A(n11133), .ZN(P3_U3519) );
  OAI222_X1 U13697 ( .A1(n13960), .A2(n11136), .B1(P2_U3088), .B2(n11135), 
        .C1(n13955), .C2(n11134), .ZN(P2_U3306) );
  INV_X1 U13698 ( .A(n11137), .ZN(n11404) );
  INV_X1 U13699 ( .A(n11138), .ZN(n11139) );
  NAND2_X1 U13700 ( .A1(n11141), .A2(n7660), .ZN(n11275) );
  INV_X1 U13701 ( .A(n11275), .ZN(n11278) );
  AOI22_X1 U13702 ( .A1(n12331), .A2(n12262), .B1(n12267), .B2(n14154), .ZN(
        n11142) );
  XOR2_X1 U13703 ( .A(n12212), .B(n11142), .Z(n11273) );
  OAI22_X1 U13704 ( .A1(n11406), .A2(n12274), .B1(n11143), .B2(n10622), .ZN(
        n11274) );
  XNOR2_X1 U13705 ( .A(n11273), .B(n11274), .ZN(n11144) );
  XNOR2_X1 U13706 ( .A(n11275), .B(n11144), .ZN(n11145) );
  NAND2_X1 U13707 ( .A1(n11145), .A2(n14828), .ZN(n11149) );
  OAI22_X1 U13708 ( .A1(n14121), .A2(n11146), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15671), .ZN(n11147) );
  AOI21_X1 U13709 ( .B1(n12331), .B2(n6638), .A(n11147), .ZN(n11148) );
  OAI211_X1 U13710 ( .C1(n14836), .C2(n11404), .A(n11149), .B(n11148), .ZN(
        P1_U3227) );
  OR2_X1 U13711 ( .A1(n11077), .A2(n11150), .ZN(n11151) );
  NAND2_X1 U13712 ( .A1(n11151), .A2(n12663), .ZN(n11152) );
  XNOR2_X1 U13713 ( .A(n11152), .B(n12776), .ZN(n15304) );
  NAND2_X1 U13714 ( .A1(n15304), .A2(n13204), .ZN(n11157) );
  INV_X1 U13715 ( .A(n12776), .ZN(n12665) );
  XNOR2_X1 U13716 ( .A(n11153), .B(n12665), .ZN(n11155) );
  OAI22_X1 U13717 ( .A1(n13012), .A2(n13312), .B1(n11740), .B2(n13314), .ZN(
        n11154) );
  AOI21_X1 U13718 ( .B1(n11155), .B2(n15248), .A(n11154), .ZN(n11156) );
  AND2_X1 U13719 ( .A1(n11157), .A2(n11156), .ZN(n15306) );
  INV_X1 U13720 ( .A(n11158), .ZN(n12875) );
  AOI22_X1 U13721 ( .A1(n13322), .A2(n15301), .B1(n13288), .B2(n12875), .ZN(
        n11159) );
  OAI21_X1 U13722 ( .B1(n11224), .B2(n13344), .A(n11159), .ZN(n11160) );
  AOI21_X1 U13723 ( .B1(n15304), .B2(n13210), .A(n11160), .ZN(n11161) );
  OAI21_X1 U13724 ( .B1(n15306), .B2(n15258), .A(n11161), .ZN(P3_U3223) );
  XNOR2_X1 U13725 ( .A(n11162), .B(n11168), .ZN(n11163) );
  AOI222_X1 U13726 ( .A1(n15131), .A2(n11163), .B1(n13595), .B2(n15128), .C1(
        n13597), .C2(n15127), .ZN(n11202) );
  INV_X1 U13727 ( .A(n11179), .ZN(n11164) );
  AOI211_X1 U13728 ( .C1(n11200), .C2(n11165), .A(n12009), .B(n11164), .ZN(
        n11199) );
  AOI22_X1 U13729 ( .A1(n15157), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11166), 
        .B2(n15154), .ZN(n11167) );
  OAI21_X1 U13730 ( .B1(n9707), .B2(n13813), .A(n11167), .ZN(n11171) );
  XNOR2_X1 U13731 ( .A(n11169), .B(n11168), .ZN(n11203) );
  NOR2_X1 U13732 ( .A1(n11203), .A2(n15139), .ZN(n11170) );
  AOI211_X1 U13733 ( .C1(n11199), .C2(n13835), .A(n11171), .B(n11170), .ZN(
        n11172) );
  OAI21_X1 U13734 ( .B1(n15157), .B2(n11202), .A(n11172), .ZN(P2_U3254) );
  XNOR2_X1 U13735 ( .A(n11173), .B(n11174), .ZN(n14820) );
  INV_X1 U13736 ( .A(n14820), .ZN(n11187) );
  AOI21_X1 U13737 ( .B1(n11175), .B2(n11174), .A(n11793), .ZN(n11178) );
  OAI22_X1 U13738 ( .A1(n12131), .A2(n15148), .B1(n11176), .B2(n13567), .ZN(
        n12571) );
  AOI21_X1 U13739 ( .B1(n11178), .B2(n11177), .A(n12571), .ZN(n14817) );
  INV_X1 U13740 ( .A(n14817), .ZN(n11185) );
  NAND2_X1 U13741 ( .A1(n14815), .A2(n11179), .ZN(n11180) );
  NAND2_X1 U13742 ( .A1(n11180), .A2(n15134), .ZN(n11181) );
  OR2_X1 U13743 ( .A1(n11267), .A2(n11181), .ZN(n14816) );
  OAI22_X1 U13744 ( .A1(n15155), .A2(n15546), .B1(n12574), .B2(n15132), .ZN(
        n11182) );
  AOI21_X1 U13745 ( .B1(n14815), .B2(n15144), .A(n11182), .ZN(n11183) );
  OAI21_X1 U13746 ( .B1(n14816), .B2(n15140), .A(n11183), .ZN(n11184) );
  AOI21_X1 U13747 ( .B1(n11185), .B2(n15155), .A(n11184), .ZN(n11186) );
  OAI21_X1 U13748 ( .B1(n15139), .B2(n11187), .A(n11186), .ZN(P2_U3253) );
  XNOR2_X1 U13749 ( .A(n11188), .B(n12782), .ZN(n11190) );
  OAI22_X1 U13750 ( .A1(n11749), .A2(n13312), .B1(n11744), .B2(n13314), .ZN(
        n11189) );
  AOI21_X1 U13751 ( .B1(n11190), .B2(n15248), .A(n11189), .ZN(n14802) );
  AND2_X1 U13752 ( .A1(n11192), .A2(n11191), .ZN(n11193) );
  XNOR2_X1 U13753 ( .A(n11193), .B(n12782), .ZN(n14798) );
  INV_X1 U13754 ( .A(n11194), .ZN(n13018) );
  AOI22_X1 U13755 ( .A1(n13322), .A2(n14799), .B1(n13018), .B2(n13288), .ZN(
        n11195) );
  OAI21_X1 U13756 ( .B1(n11196), .B2(n13344), .A(n11195), .ZN(n11197) );
  AOI21_X1 U13757 ( .B1(n14798), .B2(n13347), .A(n11197), .ZN(n11198) );
  OAI21_X1 U13758 ( .B1(n14802), .B2(n13328), .A(n11198), .ZN(P3_U3222) );
  INV_X1 U13759 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11205) );
  AOI21_X1 U13760 ( .B1(n15196), .B2(n11200), .A(n11199), .ZN(n11201) );
  OAI211_X1 U13761 ( .C1(n15187), .C2(n11203), .A(n11202), .B(n11201), .ZN(
        n11206) );
  NAND2_X1 U13762 ( .A1(n11206), .A2(n15212), .ZN(n11204) );
  OAI21_X1 U13763 ( .B1(n15212), .B2(n11205), .A(n11204), .ZN(P2_U3463) );
  NAND2_X1 U13764 ( .A1(n11206), .A2(n15233), .ZN(n11207) );
  OAI21_X1 U13765 ( .B1(n15233), .B2(n10379), .A(n11207), .ZN(P2_U3510) );
  NAND2_X1 U13766 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11464), .ZN(n11210) );
  OAI21_X1 U13767 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n11464), .A(n11210), 
        .ZN(n11211) );
  AOI21_X1 U13768 ( .B1(n11212), .B2(n11211), .A(n11465), .ZN(n11235) );
  NAND2_X1 U13769 ( .A1(n15234), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11213) );
  NAND2_X1 U13770 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n12872)
         );
  NAND2_X1 U13771 ( .A1(n11213), .A2(n12872), .ZN(n11222) );
  NOR2_X1 U13772 ( .A1(n7313), .A2(n11214), .ZN(n11216) );
  NAND2_X1 U13773 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11464), .ZN(n11217) );
  OAI21_X1 U13774 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11464), .A(n11217), 
        .ZN(n11218) );
  NOR2_X1 U13775 ( .A1(n11219), .A2(n11218), .ZN(n11453) );
  AOI21_X1 U13776 ( .B1(n11219), .B2(n11218), .A(n11453), .ZN(n11220) );
  NOR2_X1 U13777 ( .A1(n11220), .A2(n13150), .ZN(n11221) );
  AOI211_X1 U13778 ( .C1(n13166), .C2(n11225), .A(n11222), .B(n11221), .ZN(
        n11234) );
  MUX2_X1 U13779 ( .A(n11224), .B(n11223), .S(n6648), .Z(n11226) );
  NAND2_X1 U13780 ( .A1(n11226), .A2(n11225), .ZN(n11457) );
  INV_X1 U13781 ( .A(n11226), .ZN(n11227) );
  NAND2_X1 U13782 ( .A1(n11227), .A2(n11464), .ZN(n11228) );
  NAND2_X1 U13783 ( .A1(n11457), .A2(n11228), .ZN(n11229) );
  AND3_X1 U13784 ( .A1(n11231), .A2(n11230), .A3(n11229), .ZN(n11232) );
  OAI21_X1 U13785 ( .B1(n11458), .B2(n11232), .A(n13132), .ZN(n11233) );
  OAI211_X1 U13786 ( .C1(n11235), .C2(n13165), .A(n11234), .B(n11233), .ZN(
        P3_U3192) );
  NAND2_X1 U13787 ( .A1(n11236), .A2(n13058), .ZN(n11237) );
  XNOR2_X1 U13788 ( .A(n12903), .B(n15283), .ZN(n11239) );
  XNOR2_X1 U13789 ( .A(n11239), .B(n11244), .ZN(n12815) );
  NAND2_X1 U13790 ( .A1(n12816), .A2(n12815), .ZN(n12814) );
  NAND2_X1 U13791 ( .A1(n11239), .A2(n12652), .ZN(n11240) );
  NAND2_X1 U13792 ( .A1(n12814), .A2(n11240), .ZN(n11243) );
  XNOR2_X1 U13793 ( .A(n12903), .B(n11241), .ZN(n11736) );
  XNOR2_X1 U13794 ( .A(n11736), .B(n13057), .ZN(n11242) );
  OAI211_X1 U13795 ( .C1(n11243), .C2(n11242), .A(n11739), .B(n12995), .ZN(
        n11248) );
  OAI22_X1 U13796 ( .A1(n13003), .A2(n15289), .B1(n13041), .B2(n11244), .ZN(
        n11245) );
  AOI211_X1 U13797 ( .C1(n13037), .C2(n12874), .A(n11246), .B(n11245), .ZN(
        n11247) );
  OAI211_X1 U13798 ( .C1(n11250), .C2(n13031), .A(n11248), .B(n11247), .ZN(
        P3_U3161) );
  XNOR2_X1 U13799 ( .A(n11249), .B(n12770), .ZN(n15292) );
  OAI22_X1 U13800 ( .A1(n13341), .A2(n15289), .B1(n11250), .B2(n15238), .ZN(
        n11258) );
  INV_X1 U13801 ( .A(n11252), .ZN(n11253) );
  AOI21_X1 U13802 ( .B1(n12770), .B2(n11251), .A(n11253), .ZN(n11256) );
  AOI22_X1 U13803 ( .A1(n12874), .A2(n15242), .B1(n15244), .B2(n12652), .ZN(
        n11255) );
  NAND2_X1 U13804 ( .A1(n15292), .A2(n13204), .ZN(n11254) );
  OAI211_X1 U13805 ( .C1(n11256), .C2(n13310), .A(n11255), .B(n11254), .ZN(
        n15290) );
  MUX2_X1 U13806 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n15290), .S(n13344), .Z(
        n11257) );
  AOI211_X1 U13807 ( .C1(n15292), .C2(n13210), .A(n11258), .B(n11257), .ZN(
        n11259) );
  INV_X1 U13808 ( .A(n11259), .ZN(P3_U3225) );
  INV_X1 U13809 ( .A(n11260), .ZN(n11262) );
  OAI222_X1 U13810 ( .A1(n6655), .A2(n11262), .B1(n12584), .B2(n11261), .C1(
        P3_U3151), .C2(n8274), .ZN(P3_U3271) );
  XNOR2_X1 U13811 ( .A(n11263), .B(n11265), .ZN(n11264) );
  AOI22_X1 U13812 ( .A1(n13593), .A2(n15128), .B1(n13595), .B2(n15127), .ZN(
        n14996) );
  OAI21_X1 U13813 ( .B1(n11264), .B2(n11793), .A(n14996), .ZN(n14812) );
  INV_X1 U13814 ( .A(n14812), .ZN(n11272) );
  XNOR2_X1 U13815 ( .A(n11266), .B(n11265), .ZN(n14814) );
  OAI211_X1 U13816 ( .C1(n14811), .C2(n11267), .A(n15134), .B(n11592), .ZN(
        n14810) );
  OAI22_X1 U13817 ( .A1(n15155), .A2(n11424), .B1(n15008), .B2(n15132), .ZN(
        n11268) );
  AOI21_X1 U13818 ( .B1(n15005), .B2(n15144), .A(n11268), .ZN(n11269) );
  OAI21_X1 U13819 ( .B1(n14810), .B2(n15140), .A(n11269), .ZN(n11270) );
  AOI21_X1 U13820 ( .B1(n14814), .B2(n15122), .A(n11270), .ZN(n11271) );
  OAI21_X1 U13821 ( .B1(n11272), .B2(n15157), .A(n11271), .ZN(P2_U3252) );
  INV_X1 U13822 ( .A(n11274), .ZN(n11277) );
  OAI21_X2 U13823 ( .B1(n11278), .B2(n11277), .A(n11276), .ZN(n11291) );
  OR2_X1 U13824 ( .A1(n12348), .A2(n12274), .ZN(n11280) );
  NAND2_X1 U13825 ( .A1(n12268), .A2(n14153), .ZN(n11279) );
  NAND2_X1 U13826 ( .A1(n11280), .A2(n11279), .ZN(n11289) );
  OAI22_X1 U13827 ( .A1(n12348), .A2(n12275), .B1(n12344), .B2(n12274), .ZN(
        n11282) );
  XNOR2_X1 U13828 ( .A(n11282), .B(n12265), .ZN(n11288) );
  XOR2_X1 U13829 ( .A(n11289), .B(n11288), .Z(n11290) );
  XOR2_X1 U13830 ( .A(n11291), .B(n11290), .Z(n11283) );
  NAND2_X1 U13831 ( .A1(n11283), .A2(n14828), .ZN(n11287) );
  NAND2_X1 U13832 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14220) );
  OAI21_X1 U13833 ( .B1(n14121), .B2(n11284), .A(n14220), .ZN(n11285) );
  AOI21_X1 U13834 ( .B1(n12343), .B2(n6638), .A(n11285), .ZN(n11286) );
  OAI211_X1 U13835 ( .C1(n14836), .C2(n11371), .A(n11287), .B(n11286), .ZN(
        P1_U3239) );
  NOR2_X1 U13836 ( .A1(n10622), .A2(n12341), .ZN(n11292) );
  AOI21_X1 U13837 ( .B1(n12342), .B2(n12267), .A(n11292), .ZN(n11537) );
  OAI22_X1 U13838 ( .A1(n12340), .A2(n12275), .B1(n12341), .B2(n12274), .ZN(
        n11293) );
  XNOR2_X1 U13839 ( .A(n11293), .B(n12265), .ZN(n11536) );
  XNOR2_X1 U13840 ( .A(n11539), .B(n11538), .ZN(n11299) );
  INV_X1 U13841 ( .A(n14836), .ZN(n14124) );
  INV_X1 U13842 ( .A(n11394), .ZN(n11296) );
  NAND2_X1 U13843 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n14234) );
  OAI21_X1 U13844 ( .B1(n14121), .B2(n11294), .A(n14234), .ZN(n11295) );
  AOI21_X1 U13845 ( .B1(n14124), .B2(n11296), .A(n11295), .ZN(n11298) );
  NAND2_X1 U13846 ( .A1(n6638), .A2(n12342), .ZN(n11297) );
  OAI211_X1 U13847 ( .C1(n11299), .C2(n14103), .A(n11298), .B(n11297), .ZN(
        P1_U3213) );
  OAI211_X1 U13848 ( .C1(n11301), .C2(n12526), .A(n11300), .B(n14899), .ZN(
        n11381) );
  NAND2_X1 U13849 ( .A1(n14150), .A2(n14111), .ZN(n11378) );
  AND2_X1 U13850 ( .A1(n11381), .A2(n11378), .ZN(n11315) );
  NOR2_X1 U13851 ( .A1(n11303), .A2(n11302), .ZN(n11304) );
  NAND2_X1 U13852 ( .A1(n11305), .A2(n11304), .ZN(n14320) );
  INV_X1 U13853 ( .A(n11306), .ZN(n11307) );
  OAI22_X1 U13854 ( .A1(n14923), .A2(n10283), .B1(n11715), .B2(n14507), .ZN(
        n11309) );
  OAI211_X1 U13855 ( .C1(n12373), .C2(n11474), .A(n14901), .B(n11605), .ZN(
        n11379) );
  NAND2_X1 U13856 ( .A1(n14148), .A2(n14110), .ZN(n11377) );
  AOI21_X1 U13857 ( .B1(n11379), .B2(n11377), .A(n14477), .ZN(n11308) );
  AOI211_X1 U13858 ( .C1(n14900), .C2(n12372), .A(n11309), .B(n11308), .ZN(
        n11314) );
  NAND2_X1 U13859 ( .A1(n11311), .A2(n11310), .ZN(n11520) );
  OAI21_X1 U13860 ( .B1(n11311), .B2(n11310), .A(n11520), .ZN(n11383) );
  AND2_X1 U13861 ( .A1(n12212), .A2(n12501), .ZN(n11312) );
  NAND2_X1 U13862 ( .A1(n11383), .A2(n14843), .ZN(n11313) );
  OAI211_X1 U13863 ( .C1(n11315), .C2(n6653), .A(n11314), .B(n11313), .ZN(
        P1_U3283) );
  XNOR2_X1 U13864 ( .A(n11316), .B(n12781), .ZN(n11319) );
  NAND2_X1 U13865 ( .A1(n13055), .A2(n15242), .ZN(n11317) );
  OAI21_X1 U13866 ( .B1(n13012), .B2(n13314), .A(n11317), .ZN(n11318) );
  AOI21_X1 U13867 ( .B1(n11319), .B2(n15248), .A(n11318), .ZN(n14797) );
  XNOR2_X1 U13868 ( .A(n11320), .B(n12781), .ZN(n14793) );
  INV_X1 U13869 ( .A(n11321), .ZN(n12928) );
  AOI22_X1 U13870 ( .A1(n13322), .A2(n14794), .B1(n13288), .B2(n12928), .ZN(
        n11322) );
  OAI21_X1 U13871 ( .B1(n11323), .B2(n13344), .A(n11322), .ZN(n11324) );
  AOI21_X1 U13872 ( .B1(n14793), .B2(n13347), .A(n11324), .ZN(n11325) );
  OAI21_X1 U13873 ( .B1(n14797), .B2(n15258), .A(n11325), .ZN(P3_U3221) );
  NOR2_X1 U13874 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  MUX2_X1 U13875 ( .A(n11329), .B(n11328), .S(n14929), .Z(n11335) );
  OAI22_X1 U13876 ( .A1(n14925), .A2(n11331), .B1(n14507), .B2(n11330), .ZN(
        n11332) );
  AOI21_X1 U13877 ( .B1(n14911), .B2(n11333), .A(n11332), .ZN(n11334) );
  OAI211_X1 U13878 ( .C1(n14518), .C2(n11336), .A(n11335), .B(n11334), .ZN(
        P1_U3289) );
  INV_X1 U13879 ( .A(n14904), .ZN(n11339) );
  INV_X1 U13880 ( .A(n11337), .ZN(n11338) );
  AOI211_X1 U13881 ( .C1(n14975), .C2(n11339), .A(n14909), .B(n11338), .ZN(
        n14973) );
  OAI22_X1 U13882 ( .A1(n14925), .A2(n11340), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14507), .ZN(n11341) );
  AOI21_X1 U13883 ( .B1(n14911), .B2(n14973), .A(n11341), .ZN(n11351) );
  OAI21_X1 U13884 ( .B1(n11343), .B2(n12514), .A(n11342), .ZN(n11348) );
  XNOR2_X1 U13885 ( .A(n11344), .B(n12514), .ZN(n11345) );
  NOR2_X1 U13886 ( .A1(n11345), .A2(n14895), .ZN(n11346) );
  AOI211_X1 U13887 ( .C1(n14899), .C2(n11348), .A(n11347), .B(n11346), .ZN(
        n14976) );
  MUX2_X1 U13888 ( .A(n11349), .B(n14976), .S(n14929), .Z(n11350) );
  NAND2_X1 U13889 ( .A1(n11351), .A2(n11350), .ZN(P1_U3290) );
  OAI21_X1 U13890 ( .B1(n11353), .B2(n12523), .A(n11352), .ZN(n14984) );
  INV_X1 U13891 ( .A(n14984), .ZN(n11366) );
  INV_X1 U13892 ( .A(n11354), .ZN(n11355) );
  AOI21_X1 U13893 ( .B1(n11355), .B2(n12523), .A(n14921), .ZN(n11359) );
  NAND2_X1 U13894 ( .A1(n14152), .A2(n14111), .ZN(n11357) );
  NAND2_X1 U13895 ( .A1(n14150), .A2(n14110), .ZN(n11356) );
  NAND2_X1 U13896 ( .A1(n11357), .A2(n11356), .ZN(n11549) );
  AOI21_X1 U13897 ( .B1(n11359), .B2(n11358), .A(n11549), .ZN(n14981) );
  MUX2_X1 U13898 ( .A(n11360), .B(n14981), .S(n14923), .Z(n11365) );
  INV_X1 U13899 ( .A(n11475), .ZN(n11361) );
  AOI211_X1 U13900 ( .C1(n12363), .C2(n11362), .A(n14909), .B(n11361), .ZN(
        n14979) );
  OAI22_X1 U13901 ( .A1(n14925), .A2(n7192), .B1(n11552), .B2(n14507), .ZN(
        n11363) );
  AOI21_X1 U13902 ( .B1(n14979), .B2(n14911), .A(n11363), .ZN(n11364) );
  OAI211_X1 U13903 ( .C1(n11366), .C2(n14518), .A(n11365), .B(n11364), .ZN(
        P1_U3285) );
  NOR2_X1 U13904 ( .A1(n6653), .A2(n14895), .ZN(n14395) );
  INV_X1 U13905 ( .A(n14395), .ZN(n14500) );
  INV_X1 U13906 ( .A(n11367), .ZN(n11376) );
  INV_X1 U13907 ( .A(n11368), .ZN(n11369) );
  MUX2_X1 U13908 ( .A(n11370), .B(n11369), .S(n14929), .Z(n11375) );
  OAI22_X1 U13909 ( .A1(n14925), .A2(n12348), .B1(n11371), .B2(n14507), .ZN(
        n11372) );
  AOI21_X1 U13910 ( .B1(n11373), .B2(n14911), .A(n11372), .ZN(n11374) );
  OAI211_X1 U13911 ( .C1(n14500), .C2(n11376), .A(n11375), .B(n11374), .ZN(
        P1_U3287) );
  NAND2_X1 U13912 ( .A1(n11378), .A2(n11377), .ZN(n11713) );
  INV_X1 U13913 ( .A(n11713), .ZN(n11380) );
  NAND3_X1 U13914 ( .A1(n11381), .A2(n11380), .A3(n11379), .ZN(n11382) );
  AOI21_X1 U13915 ( .B1(n14918), .B2(n11383), .A(n11382), .ZN(n11388) );
  INV_X1 U13916 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11384) );
  OAI22_X1 U13917 ( .A1(n12373), .A2(n14643), .B1(n14987), .B2(n11384), .ZN(
        n11385) );
  INV_X1 U13918 ( .A(n11385), .ZN(n11386) );
  OAI21_X1 U13919 ( .B1(n11388), .B2(n14985), .A(n11386), .ZN(P1_U3489) );
  AOI22_X1 U13920 ( .A1(n14602), .A2(n12372), .B1(n14991), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11387) );
  OAI21_X1 U13921 ( .B1(n11388), .B2(n14991), .A(n11387), .ZN(P1_U3538) );
  OAI222_X1 U13922 ( .A1(n13960), .A2(n11391), .B1(P2_U3088), .B2(n11390), 
        .C1(n13955), .C2(n11389), .ZN(P2_U3305) );
  INV_X1 U13923 ( .A(n11392), .ZN(n11401) );
  NAND2_X1 U13924 ( .A1(n11393), .A2(n14929), .ZN(n11400) );
  NOR2_X1 U13925 ( .A1(n14925), .A2(n12340), .ZN(n11397) );
  OAI22_X1 U13926 ( .A1(n14923), .A2(n11395), .B1(n11394), .B2(n14507), .ZN(
        n11396) );
  AOI211_X1 U13927 ( .C1(n11398), .C2(n14911), .A(n11397), .B(n11396), .ZN(
        n11399) );
  OAI211_X1 U13928 ( .C1(n14500), .C2(n11401), .A(n11400), .B(n11399), .ZN(
        P1_U3286) );
  INV_X1 U13929 ( .A(n11402), .ZN(n11412) );
  NAND2_X1 U13930 ( .A1(n11403), .A2(n14929), .ZN(n11411) );
  OAI22_X1 U13931 ( .A1(n14923), .A2(n11405), .B1(n11404), .B2(n14507), .ZN(
        n11408) );
  NOR2_X1 U13932 ( .A1(n14925), .A2(n11406), .ZN(n11407) );
  AOI211_X1 U13933 ( .C1(n11409), .C2(n14911), .A(n11408), .B(n11407), .ZN(
        n11410) );
  OAI211_X1 U13934 ( .C1(n14500), .C2(n11412), .A(n11411), .B(n11410), .ZN(
        P1_U3288) );
  AOI21_X1 U13935 ( .B1(n12509), .B2(n14929), .A(n14911), .ZN(n11420) );
  NOR2_X1 U13936 ( .A1(n14507), .A2(n11413), .ZN(n11418) );
  INV_X1 U13937 ( .A(n11414), .ZN(n11415) );
  NOR4_X1 U13938 ( .A1(n14320), .A2(n11416), .A3(n11415), .A4(n12515), .ZN(
        n11417) );
  AOI211_X1 U13939 ( .C1(n6653), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11418), .B(
        n11417), .ZN(n11419) );
  OAI21_X1 U13940 ( .B1(n11421), .B2(n11420), .A(n11419), .ZN(P1_U3293) );
  OAI222_X1 U13941 ( .A1(n12584), .A2(n15454), .B1(P3_U3151), .B2(n11423), 
        .C1(n6655), .C2(n11422), .ZN(P3_U3270) );
  NAND2_X1 U13942 ( .A1(n15050), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11427) );
  MUX2_X1 U13943 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11424), .S(n15050), .Z(
        n15055) );
  NOR2_X1 U13944 ( .A1(n11436), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11425) );
  NOR2_X1 U13945 ( .A1(n11426), .A2(n11425), .ZN(n15056) );
  NAND2_X1 U13946 ( .A1(n15055), .A2(n15056), .ZN(n15054) );
  NAND2_X1 U13947 ( .A1(n11427), .A2(n15054), .ZN(n11429) );
  NAND2_X1 U13948 ( .A1(n11428), .A2(n11429), .ZN(n11430) );
  XNOR2_X1 U13949 ( .A(n11429), .B(n15061), .ZN(n15065) );
  NAND2_X1 U13950 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n15065), .ZN(n15064) );
  NAND2_X1 U13951 ( .A1(n11430), .A2(n15064), .ZN(n11431) );
  NAND2_X1 U13952 ( .A1(n15073), .A2(n11431), .ZN(n11432) );
  XNOR2_X1 U13953 ( .A(n11431), .B(n11442), .ZN(n15075) );
  NAND2_X1 U13954 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15075), .ZN(n15074) );
  NAND2_X1 U13955 ( .A1(n11432), .A2(n15074), .ZN(n11435) );
  INV_X1 U13956 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13620) );
  NOR2_X1 U13957 ( .A1(n13627), .A2(n13620), .ZN(n11433) );
  AOI21_X1 U13958 ( .B1(n13620), .B2(n13627), .A(n11433), .ZN(n11434) );
  NAND2_X1 U13959 ( .A1(n11434), .A2(n11435), .ZN(n13619) );
  OAI211_X1 U13960 ( .C1(n11435), .C2(n11434), .A(n15091), .B(n13619), .ZN(
        n11449) );
  NAND2_X1 U13961 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n11692)
         );
  XNOR2_X1 U13962 ( .A(n15061), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15068) );
  NOR2_X1 U13963 ( .A1(n11436), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11437) );
  NOR2_X1 U13964 ( .A1(n11438), .A2(n11437), .ZN(n15053) );
  MUX2_X1 U13965 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n11439), .S(n15050), .Z(
        n15052) );
  NAND2_X1 U13966 ( .A1(n15053), .A2(n15052), .ZN(n15051) );
  OAI21_X1 U13967 ( .B1(n11440), .B2(n11439), .A(n15051), .ZN(n15067) );
  NAND2_X1 U13968 ( .A1(n15068), .A2(n15067), .ZN(n15066) );
  OAI21_X1 U13969 ( .B1(n15061), .B2(n15541), .A(n15066), .ZN(n11441) );
  NAND2_X1 U13970 ( .A1(n15073), .A2(n11441), .ZN(n11443) );
  XNOR2_X1 U13971 ( .A(n11442), .B(n11441), .ZN(n15077) );
  NAND2_X1 U13972 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15077), .ZN(n15076) );
  NAND2_X1 U13973 ( .A1(n11443), .A2(n15076), .ZN(n11445) );
  XNOR2_X1 U13974 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13627), .ZN(n11444) );
  NAND2_X1 U13975 ( .A1(n11444), .A2(n11445), .ZN(n13625) );
  OAI211_X1 U13976 ( .C1(n11445), .C2(n11444), .A(n15085), .B(n13625), .ZN(
        n11446) );
  NAND2_X1 U13977 ( .A1(n11692), .A2(n11446), .ZN(n11447) );
  AOI21_X1 U13978 ( .B1(n15083), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11447), 
        .ZN(n11448) );
  OAI211_X1 U13979 ( .C1(n15107), .C2(n13627), .A(n11449), .B(n11448), .ZN(
        P2_U3230) );
  INV_X1 U13980 ( .A(n11472), .ZN(n11452) );
  NAND2_X1 U13981 ( .A1(n13953), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11451) );
  OAI211_X1 U13982 ( .C1(n11452), .C2(n13955), .A(n11451), .B(n11450), .ZN(
        P2_U3304) );
  AOI21_X1 U13983 ( .B1(n11196), .B2(n11454), .A(n11561), .ZN(n11470) );
  INV_X1 U13984 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14725) );
  NOR2_X1 U13985 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11455), .ZN(n13014) );
  INV_X1 U13986 ( .A(n13014), .ZN(n11456) );
  OAI21_X1 U13987 ( .B1(n13125), .B2(n14725), .A(n11456), .ZN(n11463) );
  MUX2_X1 U13988 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12105), .Z(n11573) );
  XNOR2_X1 U13989 ( .A(n11573), .B(n11572), .ZN(n11459) );
  AOI21_X1 U13990 ( .B1(n11460), .B2(n11459), .A(n11576), .ZN(n11461) );
  NOR2_X1 U13991 ( .A1(n11461), .A2(n13170), .ZN(n11462) );
  AOI211_X1 U13992 ( .C1(n13166), .C2(n11568), .A(n11463), .B(n11462), .ZN(
        n11469) );
  NOR2_X1 U13993 ( .A1(n7879), .A2(n11466), .ZN(n11570) );
  AOI21_X1 U13994 ( .B1(n7879), .B2(n11466), .A(n11570), .ZN(n11467) );
  OR2_X1 U13995 ( .A1(n11467), .A2(n13165), .ZN(n11468) );
  OAI211_X1 U13996 ( .C1(n11470), .C2(n13150), .A(n11469), .B(n11468), .ZN(
        P3_U3193) );
  NAND2_X1 U13997 ( .A1(n11472), .A2(n11471), .ZN(n11473) );
  OAI211_X1 U13998 ( .C1(n15499), .C2(n12562), .A(n11473), .B(n12560), .ZN(
        P1_U3332) );
  AOI211_X1 U13999 ( .C1(n12368), .C2(n11475), .A(n14909), .B(n11474), .ZN(
        n14880) );
  INV_X1 U14000 ( .A(n14895), .ZN(n14918) );
  OAI21_X1 U14001 ( .B1(n11477), .B2(n11481), .A(n11476), .ZN(n11485) );
  NAND2_X1 U14002 ( .A1(n14149), .A2(n14110), .ZN(n11479) );
  NAND2_X1 U14003 ( .A1(n14151), .A2(n14111), .ZN(n11478) );
  NAND2_X1 U14004 ( .A1(n11479), .A2(n11478), .ZN(n11767) );
  NAND2_X1 U14005 ( .A1(n11482), .A2(n11481), .ZN(n11483) );
  AOI21_X1 U14006 ( .B1(n11480), .B2(n11483), .A(n14921), .ZN(n11484) );
  AOI211_X1 U14007 ( .C1(n14918), .C2(n11485), .A(n11767), .B(n11484), .ZN(
        n14888) );
  INV_X1 U14008 ( .A(n14888), .ZN(n11486) );
  NOR2_X1 U14009 ( .A1(n14880), .A2(n11486), .ZN(n11489) );
  AOI22_X1 U14010 ( .A1(n14602), .A2(n12368), .B1(n14991), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11487) );
  OAI21_X1 U14011 ( .B1(n11489), .B2(n14991), .A(n11487), .ZN(P1_U3537) );
  AOI22_X1 U14012 ( .A1(n14648), .A2(n12368), .B1(n14985), .B2(
        P1_REG0_REG_9__SCAN_IN), .ZN(n11488) );
  OAI21_X1 U14013 ( .B1(n11489), .B2(n14985), .A(n11488), .ZN(P1_U3486) );
  INV_X1 U14014 ( .A(n12575), .ZN(n11491) );
  NAND2_X1 U14015 ( .A1(n11491), .A2(n11490), .ZN(n11492) );
  NAND2_X1 U14016 ( .A1(n11493), .A2(n11492), .ZN(n11495) );
  XNOR2_X1 U14017 ( .A(n14815), .B(n12033), .ZN(n11496) );
  NAND2_X1 U14018 ( .A1(n13595), .A2(n12009), .ZN(n11497) );
  XNOR2_X1 U14019 ( .A(n11496), .B(n11497), .ZN(n12576) );
  INV_X1 U14020 ( .A(n11496), .ZN(n11498) );
  NAND2_X1 U14021 ( .A1(n11498), .A2(n11497), .ZN(n11499) );
  XNOR2_X1 U14022 ( .A(n15005), .B(n12033), .ZN(n11500) );
  AND2_X1 U14023 ( .A1(n13594), .A2(n13753), .ZN(n11501) );
  NAND2_X1 U14024 ( .A1(n11500), .A2(n11501), .ZN(n11506) );
  INV_X1 U14025 ( .A(n11500), .ZN(n12132) );
  INV_X1 U14026 ( .A(n11501), .ZN(n11502) );
  NAND2_X1 U14027 ( .A1(n12132), .A2(n11502), .ZN(n11503) );
  NAND2_X1 U14028 ( .A1(n11506), .A2(n11503), .ZN(n15001) );
  NAND2_X1 U14029 ( .A1(n13593), .A2(n12009), .ZN(n11507) );
  XNOR2_X1 U14030 ( .A(n11509), .B(n11507), .ZN(n12134) );
  NAND3_X1 U14031 ( .A1(n12130), .A2(n12134), .A3(n11506), .ZN(n12139) );
  INV_X1 U14032 ( .A(n11507), .ZN(n11508) );
  NAND2_X1 U14033 ( .A1(n12139), .A2(n11510), .ZN(n11686) );
  XNOR2_X1 U14034 ( .A(n13918), .B(n11494), .ZN(n11684) );
  INV_X1 U14035 ( .A(n11688), .ZN(n11518) );
  AOI22_X1 U14036 ( .A1(n11512), .A2(n13552), .B1(n13501), .B2(n13592), .ZN(
        n11517) );
  OAI22_X1 U14037 ( .A1(n12286), .A2(n15148), .B1(n11513), .B2(n13567), .ZN(
        n11795) );
  AOI22_X1 U14038 ( .A1(n13515), .A2(n11795), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11514) );
  OAI21_X1 U14039 ( .B1(n11800), .B2(n15007), .A(n11514), .ZN(n11515) );
  AOI21_X1 U14040 ( .B1(n13918), .B2(n15004), .A(n11515), .ZN(n11516) );
  OAI21_X1 U14041 ( .B1(n11518), .B2(n11517), .A(n11516), .ZN(P2_U3213) );
  NAND2_X1 U14042 ( .A1(n11520), .A2(n11519), .ZN(n11603) );
  NAND2_X1 U14043 ( .A1(n11603), .A2(n11602), .ZN(n11601) );
  NAND2_X1 U14044 ( .A1(n11601), .A2(n11521), .ZN(n11523) );
  OAI21_X1 U14045 ( .B1(n11523), .B2(n12530), .A(n11522), .ZN(n11655) );
  INV_X1 U14046 ( .A(n11655), .ZN(n11535) );
  OAI211_X1 U14047 ( .C1(n11526), .C2(n11525), .A(n11524), .B(n14899), .ZN(
        n11530) );
  NAND2_X1 U14048 ( .A1(n14146), .A2(n14110), .ZN(n11528) );
  NAND2_X1 U14049 ( .A1(n14148), .A2(n14111), .ZN(n11527) );
  NAND2_X1 U14050 ( .A1(n11528), .A2(n11527), .ZN(n14012) );
  INV_X1 U14051 ( .A(n14012), .ZN(n11529) );
  NAND2_X1 U14052 ( .A1(n11530), .A2(n11529), .ZN(n11653) );
  NAND2_X1 U14053 ( .A1(n11653), .A2(n14929), .ZN(n11534) );
  AOI211_X1 U14054 ( .C1(n12382), .C2(n11604), .A(n14909), .B(n6649), .ZN(
        n11654) );
  NOR2_X1 U14055 ( .A1(n7204), .A2(n14925), .ZN(n11532) );
  OAI22_X1 U14056 ( .A1(n14923), .A2(n10569), .B1(n14009), .B2(n14507), .ZN(
        n11531) );
  AOI211_X1 U14057 ( .C1(n11654), .C2(n14911), .A(n11532), .B(n11531), .ZN(
        n11533) );
  OAI211_X1 U14058 ( .C1(n14500), .C2(n11535), .A(n11534), .B(n11533), .ZN(
        P1_U3281) );
  NAND2_X1 U14059 ( .A1(n12363), .A2(n12262), .ZN(n11541) );
  INV_X2 U14060 ( .A(n12274), .ZN(n12267) );
  NAND2_X1 U14061 ( .A1(n12267), .A2(n14151), .ZN(n11540) );
  NAND2_X1 U14062 ( .A1(n11541), .A2(n11540), .ZN(n11542) );
  XNOR2_X1 U14063 ( .A(n11542), .B(n6749), .ZN(n11546) );
  NOR2_X1 U14064 ( .A1(n10622), .A2(n11543), .ZN(n11544) );
  AOI21_X1 U14065 ( .B1(n12363), .B2(n12267), .A(n11544), .ZN(n11545) );
  NAND2_X1 U14066 ( .A1(n11546), .A2(n11545), .ZN(n11697) );
  OAI21_X1 U14067 ( .B1(n11546), .B2(n11545), .A(n11697), .ZN(n11547) );
  AOI21_X1 U14068 ( .B1(n11548), .B2(n11547), .A(n6861), .ZN(n11555) );
  NAND2_X1 U14069 ( .A1(n14830), .A2(n11549), .ZN(n11550) );
  OAI211_X1 U14070 ( .C1(n14836), .C2(n11552), .A(n11551), .B(n11550), .ZN(
        n11553) );
  AOI21_X1 U14071 ( .B1(n12363), .B2(n6638), .A(n11553), .ZN(n11554) );
  OAI21_X1 U14072 ( .B1(n11555), .B2(n14103), .A(n11554), .ZN(P1_U3221) );
  INV_X1 U14073 ( .A(n11556), .ZN(n11558) );
  OAI222_X1 U14074 ( .A1(P3_U3151), .A2(n11559), .B1(n6655), .B2(n11558), .C1(
        n11557), .C2(n12584), .ZN(P3_U3269) );
  NOR2_X1 U14075 ( .A1(n11568), .A2(n11560), .ZN(n11562) );
  NAND2_X1 U14076 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12073), .ZN(n11563) );
  OAI21_X1 U14077 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12073), .A(n11563), 
        .ZN(n11564) );
  NOR2_X1 U14078 ( .A1(n11565), .A2(n11564), .ZN(n12056) );
  AOI21_X1 U14079 ( .B1(n11565), .B2(n11564), .A(n12056), .ZN(n11586) );
  NOR2_X1 U14080 ( .A1(n11568), .A2(n11567), .ZN(n11569) );
  NAND2_X1 U14081 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12073), .ZN(n11571) );
  OAI21_X1 U14082 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n12073), .A(n11571), 
        .ZN(n12071) );
  XNOR2_X1 U14083 ( .A(n12072), .B(n12071), .ZN(n11584) );
  NOR2_X1 U14084 ( .A1(n11573), .A2(n11572), .ZN(n11575) );
  MUX2_X1 U14085 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6648), .Z(n12089) );
  XNOR2_X1 U14086 ( .A(n12089), .B(n12073), .ZN(n11574) );
  NOR3_X1 U14087 ( .A1(n11576), .A2(n11575), .A3(n11574), .ZN(n13067) );
  INV_X1 U14088 ( .A(n13067), .ZN(n11578) );
  OAI21_X1 U14089 ( .B1(n11576), .B2(n11575), .A(n11574), .ZN(n11577) );
  NAND3_X1 U14090 ( .A1(n11578), .A2(n13132), .A3(n11577), .ZN(n11581) );
  NOR2_X1 U14091 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11579), .ZN(n12927) );
  AOI21_X1 U14092 ( .B1(n15234), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12927), 
        .ZN(n11580) );
  OAI211_X1 U14093 ( .C1(n11582), .C2(n12073), .A(n11581), .B(n11580), .ZN(
        n11583) );
  AOI21_X1 U14094 ( .B1(n13093), .B2(n11584), .A(n11583), .ZN(n11585) );
  OAI21_X1 U14095 ( .B1(n11586), .B2(n13150), .A(n11585), .ZN(P3_U3194) );
  XNOR2_X1 U14096 ( .A(n11587), .B(n11597), .ZN(n11590) );
  NAND2_X1 U14097 ( .A1(n13592), .A2(n15128), .ZN(n11589) );
  NAND2_X1 U14098 ( .A1(n13594), .A2(n15127), .ZN(n11588) );
  NAND2_X1 U14099 ( .A1(n11589), .A2(n11588), .ZN(n12127) );
  AOI21_X1 U14100 ( .B1(n11590), .B2(n15131), .A(n12127), .ZN(n13923) );
  INV_X1 U14101 ( .A(n11591), .ZN(n11799) );
  AOI211_X1 U14102 ( .C1(n11505), .C2(n11592), .A(n12009), .B(n11591), .ZN(
        n13922) );
  INV_X1 U14103 ( .A(n11505), .ZN(n11595) );
  INV_X1 U14104 ( .A(n12129), .ZN(n11593) );
  AOI22_X1 U14105 ( .A1(n15157), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11593), 
        .B2(n15154), .ZN(n11594) );
  OAI21_X1 U14106 ( .B1(n11595), .B2(n13813), .A(n11594), .ZN(n11599) );
  XNOR2_X1 U14107 ( .A(n11596), .B(n11597), .ZN(n13925) );
  NOR2_X1 U14108 ( .A1(n13925), .A2(n15139), .ZN(n11598) );
  AOI211_X1 U14109 ( .C1(n13922), .C2(n13835), .A(n11599), .B(n11598), .ZN(
        n11600) );
  OAI21_X1 U14110 ( .B1(n15157), .B2(n13923), .A(n11600), .ZN(P2_U3251) );
  OAI21_X1 U14111 ( .B1(n11603), .B2(n11602), .A(n11601), .ZN(n14844) );
  AOI211_X1 U14112 ( .C1(n12377), .C2(n11605), .A(n14909), .B(n7205), .ZN(
        n14837) );
  OAI211_X1 U14113 ( .C1(n11607), .C2(n12527), .A(n11606), .B(n14899), .ZN(
        n11610) );
  NAND2_X1 U14114 ( .A1(n14149), .A2(n14111), .ZN(n11609) );
  NAND2_X1 U14115 ( .A1(n14147), .A2(n14110), .ZN(n11608) );
  AND2_X1 U14116 ( .A1(n11609), .A2(n11608), .ZN(n11888) );
  AND2_X1 U14117 ( .A1(n11610), .A2(n11888), .ZN(n14846) );
  INV_X1 U14118 ( .A(n14846), .ZN(n11611) );
  AOI211_X1 U14119 ( .C1(n14918), .C2(n14844), .A(n14837), .B(n11611), .ZN(
        n11616) );
  INV_X1 U14120 ( .A(n12377), .ZN(n14841) );
  INV_X1 U14121 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11612) );
  OAI22_X1 U14122 ( .A1(n14841), .A2(n14643), .B1(n14987), .B2(n11612), .ZN(
        n11613) );
  INV_X1 U14123 ( .A(n11613), .ZN(n11614) );
  OAI21_X1 U14124 ( .B1(n11616), .B2(n14985), .A(n11614), .ZN(P1_U3492) );
  AOI22_X1 U14125 ( .A1(n12377), .A2(n14602), .B1(n14991), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11615) );
  OAI21_X1 U14126 ( .B1(n11616), .B2(n14991), .A(n11615), .ZN(P1_U3539) );
  OAI21_X1 U14127 ( .B1(n11618), .B2(n12529), .A(n11617), .ZN(n11727) );
  INV_X1 U14128 ( .A(n11727), .ZN(n11629) );
  OAI211_X1 U14129 ( .C1(n11621), .C2(n11620), .A(n11619), .B(n14899), .ZN(
        n11622) );
  AOI22_X1 U14130 ( .A1(n14145), .A2(n14110), .B1(n14111), .B2(n14147), .ZN(
        n14076) );
  NAND2_X1 U14131 ( .A1(n11622), .A2(n14076), .ZN(n11725) );
  NAND2_X1 U14132 ( .A1(n11725), .A2(n14929), .ZN(n11628) );
  AOI211_X1 U14133 ( .C1(n12387), .C2(n11623), .A(n14909), .B(n7203), .ZN(
        n11726) );
  INV_X1 U14134 ( .A(n12387), .ZN(n14081) );
  NOR2_X1 U14135 ( .A1(n14081), .A2(n14925), .ZN(n11626) );
  OAI22_X1 U14136 ( .A1(n14929), .A2(n11624), .B1(n14074), .B2(n14507), .ZN(
        n11625) );
  AOI211_X1 U14137 ( .C1(n11726), .C2(n14911), .A(n11626), .B(n11625), .ZN(
        n11627) );
  OAI211_X1 U14138 ( .C1(n11629), .C2(n14518), .A(n11628), .B(n11627), .ZN(
        P1_U3280) );
  INV_X1 U14139 ( .A(n11630), .ZN(n11635) );
  OAI222_X1 U14140 ( .A1(n11632), .A2(P2_U3088), .B1(n13955), .B2(n11635), 
        .C1(n11631), .C2(n13960), .ZN(P2_U3303) );
  INV_X1 U14141 ( .A(n11633), .ZN(n11636) );
  OAI222_X1 U14142 ( .A1(P1_U3086), .A2(n11636), .B1(n6656), .B2(n11635), .C1(
        n11634), .C2(n12562), .ZN(P1_U3331) );
  INV_X1 U14143 ( .A(n11637), .ZN(n11639) );
  OAI222_X1 U14144 ( .A1(P3_U3151), .A2(n6648), .B1(n6655), .B2(n11639), .C1(
        n11638), .C2(n12584), .ZN(P3_U3268) );
  NAND2_X1 U14145 ( .A1(n11640), .A2(n15248), .ZN(n11645) );
  AOI21_X1 U14146 ( .B1(n11677), .B2(n11642), .A(n12785), .ZN(n11644) );
  AOI22_X1 U14147 ( .A1(n15244), .A2(n13055), .B1(n13053), .B2(n15242), .ZN(
        n11643) );
  OAI21_X1 U14148 ( .B1(n11645), .B2(n11644), .A(n11643), .ZN(n14785) );
  INV_X1 U14149 ( .A(n14785), .ZN(n11652) );
  OAI21_X1 U14150 ( .B1(n11647), .B2(n8239), .A(n11646), .ZN(n14787) );
  INV_X1 U14151 ( .A(n11858), .ZN(n14784) );
  INV_X1 U14152 ( .A(n11861), .ZN(n11648) );
  AOI22_X1 U14153 ( .A1(n13328), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n13288), 
        .B2(n11648), .ZN(n11649) );
  OAI21_X1 U14154 ( .B1(n14784), .B2(n13341), .A(n11649), .ZN(n11650) );
  AOI21_X1 U14155 ( .B1(n14787), .B2(n13347), .A(n11650), .ZN(n11651) );
  OAI21_X1 U14156 ( .B1(n15258), .B2(n11652), .A(n11651), .ZN(P3_U3219) );
  AOI211_X1 U14157 ( .C1(n14918), .C2(n11655), .A(n11654), .B(n11653), .ZN(
        n11660) );
  INV_X1 U14158 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11656) );
  OAI22_X1 U14159 ( .A1(n7204), .A2(n14643), .B1(n14987), .B2(n11656), .ZN(
        n11657) );
  INV_X1 U14160 ( .A(n11657), .ZN(n11658) );
  OAI21_X1 U14161 ( .B1(n11660), .B2(n14985), .A(n11658), .ZN(P1_U3495) );
  AOI22_X1 U14162 ( .A1(n12382), .A2(n14602), .B1(n14991), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11659) );
  OAI21_X1 U14163 ( .B1(n11660), .B2(n14991), .A(n11659), .ZN(P1_U3540) );
  NAND2_X1 U14164 ( .A1(n11661), .A2(n12402), .ZN(n11662) );
  NAND2_X1 U14165 ( .A1(n11831), .A2(n11662), .ZN(n11866) );
  OAI211_X1 U14166 ( .C1(n11664), .C2(n12402), .A(n11663), .B(n14899), .ZN(
        n11668) );
  NAND2_X1 U14167 ( .A1(n14146), .A2(n14111), .ZN(n11665) );
  OAI21_X1 U14168 ( .B1(n11666), .B2(n14095), .A(n11665), .ZN(n14831) );
  INV_X1 U14169 ( .A(n14831), .ZN(n11667) );
  NAND2_X1 U14170 ( .A1(n11668), .A2(n11667), .ZN(n11868) );
  NAND2_X1 U14171 ( .A1(n11868), .A2(n14929), .ZN(n11674) );
  AOI21_X1 U14172 ( .B1(n14832), .B2(n11669), .A(n14909), .ZN(n11670) );
  AND2_X1 U14173 ( .A1(n11670), .A2(n11837), .ZN(n11867) );
  OAI22_X1 U14174 ( .A1(n14929), .A2(n11783), .B1(n14835), .B2(n14507), .ZN(
        n11672) );
  NOR2_X1 U14175 ( .A1(n7202), .A2(n14925), .ZN(n11671) );
  AOI211_X1 U14176 ( .C1(n11867), .C2(n14911), .A(n11672), .B(n11671), .ZN(
        n11673) );
  OAI211_X1 U14177 ( .C1(n11866), .C2(n14518), .A(n11674), .B(n11673), .ZN(
        P1_U3279) );
  XNOR2_X1 U14178 ( .A(n11675), .B(n12783), .ZN(n14792) );
  INV_X1 U14179 ( .A(n14792), .ZN(n11683) );
  INV_X1 U14180 ( .A(n11677), .ZN(n11678) );
  AOI21_X1 U14181 ( .B1(n12783), .B2(n11676), .A(n11678), .ZN(n11679) );
  OAI222_X1 U14182 ( .A1(n13312), .A2(n11941), .B1(n13314), .B2(n11749), .C1(
        n13310), .C2(n11679), .ZN(n14790) );
  NOR2_X1 U14183 ( .A1(n13341), .A2(n14789), .ZN(n11681) );
  OAI22_X1 U14184 ( .A1(n13344), .A2(n7929), .B1(n11757), .B2(n15238), .ZN(
        n11680) );
  AOI211_X1 U14185 ( .C1(n14790), .C2(n13344), .A(n11681), .B(n11680), .ZN(
        n11682) );
  OAI21_X1 U14186 ( .B1(n13305), .B2(n11683), .A(n11682), .ZN(P3_U3220) );
  NAND2_X1 U14187 ( .A1(n13591), .A2(n12009), .ZN(n11977) );
  XNOR2_X1 U14188 ( .A(n13911), .B(n11494), .ZN(n12288) );
  XOR2_X1 U14189 ( .A(n11977), .B(n12288), .Z(n11690) );
  INV_X1 U14190 ( .A(n11684), .ZN(n11685) );
  AOI21_X1 U14191 ( .B1(n11690), .B2(n11689), .A(n12291), .ZN(n11696) );
  OAI22_X1 U14192 ( .A1(n13568), .A2(n15148), .B1(n11691), .B2(n13567), .ZN(
        n11809) );
  NAND2_X1 U14193 ( .A1(n13515), .A2(n11809), .ZN(n11693) );
  OAI211_X1 U14194 ( .C1(n15007), .C2(n11811), .A(n11693), .B(n11692), .ZN(
        n11694) );
  AOI21_X1 U14195 ( .B1(n13911), .B2(n15004), .A(n11694), .ZN(n11695) );
  OAI21_X1 U14196 ( .B1(n11696), .B2(n14999), .A(n11695), .ZN(P2_U3198) );
  NOR2_X1 U14197 ( .A1(n10622), .A2(n12369), .ZN(n11698) );
  AOI21_X1 U14198 ( .B1(n12368), .B2(n12267), .A(n11698), .ZN(n11701) );
  INV_X1 U14199 ( .A(n12368), .ZN(n14885) );
  OAI22_X1 U14200 ( .A1(n14885), .A2(n12275), .B1(n12369), .B2(n12274), .ZN(
        n11699) );
  XOR2_X1 U14201 ( .A(n12212), .B(n11699), .Z(n11764) );
  INV_X1 U14202 ( .A(n11701), .ZN(n11702) );
  NAND2_X1 U14203 ( .A1(n12372), .A2(n12262), .ZN(n11706) );
  NAND2_X1 U14204 ( .A1(n12267), .A2(n14149), .ZN(n11705) );
  NAND2_X1 U14205 ( .A1(n11706), .A2(n11705), .ZN(n11707) );
  XNOR2_X1 U14206 ( .A(n11707), .B(n6749), .ZN(n11710) );
  NOR2_X1 U14207 ( .A1(n10622), .A2(n12374), .ZN(n11708) );
  AOI21_X1 U14208 ( .B1(n12372), .B2(n12267), .A(n11708), .ZN(n11709) );
  NOR2_X1 U14209 ( .A1(n11710), .A2(n11709), .ZN(n11880) );
  NAND2_X1 U14210 ( .A1(n11710), .A2(n11709), .ZN(n11881) );
  INV_X1 U14211 ( .A(n11881), .ZN(n11711) );
  NOR2_X1 U14212 ( .A1(n11880), .A2(n11711), .ZN(n11712) );
  XNOR2_X1 U14213 ( .A(n11882), .B(n11712), .ZN(n11718) );
  AOI22_X1 U14214 ( .A1(n14830), .A2(n11713), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11714) );
  OAI21_X1 U14215 ( .B1(n11715), .B2(n14836), .A(n11714), .ZN(n11716) );
  AOI21_X1 U14216 ( .B1(n12372), .B2(n6638), .A(n11716), .ZN(n11717) );
  OAI21_X1 U14217 ( .B1(n11718), .B2(n14103), .A(n11717), .ZN(P1_U3217) );
  INV_X1 U14218 ( .A(n11719), .ZN(n11723) );
  OAI222_X1 U14219 ( .A1(n12562), .A2(n11721), .B1(n6656), .B2(n11723), .C1(
        P1_U3086), .C2(n11720), .ZN(P1_U3330) );
  OAI222_X1 U14220 ( .A1(n13960), .A2(n11724), .B1(n13955), .B2(n11723), .C1(
        n11722), .C2(P2_U3088), .ZN(P2_U3302) );
  AOI211_X1 U14221 ( .C1(n14918), .C2(n11727), .A(n11726), .B(n11725), .ZN(
        n11732) );
  AOI22_X1 U14222 ( .A1(n12387), .A2(n14602), .B1(n14991), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n11728) );
  OAI21_X1 U14223 ( .B1(n11732), .B2(n14991), .A(n11728), .ZN(P1_U3541) );
  INV_X1 U14224 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11729) );
  OAI22_X1 U14225 ( .A1(n14081), .A2(n14643), .B1(n14987), .B2(n11729), .ZN(
        n11730) );
  INV_X1 U14226 ( .A(n11730), .ZN(n11731) );
  OAI21_X1 U14227 ( .B1(n11732), .B2(n14985), .A(n11731), .ZN(P1_U3498) );
  XNOR2_X1 U14228 ( .A(n14789), .B(n12849), .ZN(n11735) );
  INV_X1 U14229 ( .A(n11735), .ZN(n11733) );
  NAND2_X1 U14230 ( .A1(n11733), .A2(n13055), .ZN(n11856) );
  NAND2_X1 U14231 ( .A1(n11735), .A2(n11734), .ZN(n11854) );
  NAND2_X1 U14232 ( .A1(n11856), .A2(n11854), .ZN(n11756) );
  INV_X1 U14233 ( .A(n11736), .ZN(n11737) );
  NAND2_X1 U14234 ( .A1(n11737), .A2(n13057), .ZN(n11738) );
  XNOR2_X1 U14235 ( .A(n12903), .B(n12988), .ZN(n11741) );
  XNOR2_X1 U14236 ( .A(n11741), .B(n11740), .ZN(n12985) );
  NAND2_X1 U14237 ( .A1(n11741), .A2(n11740), .ZN(n11742) );
  XNOR2_X1 U14238 ( .A(n12903), .B(n11743), .ZN(n11745) );
  XNOR2_X1 U14239 ( .A(n11745), .B(n11744), .ZN(n12870) );
  NAND2_X1 U14240 ( .A1(n11745), .A2(n13016), .ZN(n11746) );
  NAND2_X1 U14241 ( .A1(n12869), .A2(n11746), .ZN(n12920) );
  XNOR2_X1 U14242 ( .A(n12903), .B(n14794), .ZN(n12923) );
  XNOR2_X1 U14243 ( .A(n12903), .B(n14799), .ZN(n11748) );
  AOI22_X1 U14244 ( .A1(n11749), .A2(n12923), .B1(n11748), .B2(n13012), .ZN(
        n11747) );
  NAND2_X1 U14245 ( .A1(n12920), .A2(n11747), .ZN(n11755) );
  INV_X1 U14246 ( .A(n12923), .ZN(n11753) );
  INV_X1 U14247 ( .A(n11748), .ZN(n12922) );
  NAND2_X1 U14248 ( .A1(n12922), .A2(n13056), .ZN(n11750) );
  NAND2_X1 U14249 ( .A1(n11750), .A2(n11749), .ZN(n11752) );
  INV_X1 U14250 ( .A(n11750), .ZN(n11751) );
  AOI22_X1 U14251 ( .A1(n11753), .A2(n11752), .B1(n11751), .B2(n13015), .ZN(
        n11754) );
  NAND2_X1 U14252 ( .A1(n11755), .A2(n11754), .ZN(n11855) );
  XOR2_X1 U14253 ( .A(n11756), .B(n11855), .Z(n11763) );
  INV_X1 U14254 ( .A(n11757), .ZN(n11761) );
  NAND2_X1 U14255 ( .A1(n13017), .A2(n13015), .ZN(n11758) );
  NAND2_X1 U14256 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13064)
         );
  OAI211_X1 U14257 ( .C1(n13028), .C2(n11941), .A(n11758), .B(n13064), .ZN(
        n11760) );
  NOR2_X1 U14258 ( .A1(n13003), .A2(n14789), .ZN(n11759) );
  AOI211_X1 U14259 ( .C1(n11761), .C2(n13038), .A(n11760), .B(n11759), .ZN(
        n11762) );
  OAI21_X1 U14260 ( .B1(n11763), .B2(n13046), .A(n11762), .ZN(P3_U3174) );
  XOR2_X1 U14261 ( .A(n11765), .B(n11764), .Z(n11771) );
  AOI21_X1 U14262 ( .B1(n14830), .B2(n11767), .A(n11766), .ZN(n11769) );
  NAND2_X1 U14263 ( .A1(n6638), .A2(n12368), .ZN(n11768) );
  OAI211_X1 U14264 ( .C1(n14836), .C2(n14881), .A(n11769), .B(n11768), .ZN(
        n11770) );
  AOI21_X1 U14265 ( .B1(n11771), .B2(n14828), .A(n11770), .ZN(n11772) );
  INV_X1 U14266 ( .A(n11772), .ZN(P1_U3231) );
  INV_X1 U14267 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n11773) );
  NAND2_X1 U14268 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14035)
         );
  OAI21_X1 U14269 ( .B1(n14878), .B2(n11773), .A(n14035), .ZN(n11780) );
  OAI21_X1 U14270 ( .B1(n11776), .B2(n11785), .A(n14865), .ZN(n11778) );
  XNOR2_X1 U14271 ( .A(n11906), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11777) );
  NOR2_X1 U14272 ( .A1(n11777), .A2(n11778), .ZN(n11905) );
  AOI211_X1 U14273 ( .C1(n11778), .C2(n11777), .A(n11905), .B(n14295), .ZN(
        n11779) );
  AOI211_X1 U14274 ( .C1(n14293), .C2(n11906), .A(n11780), .B(n11779), .ZN(
        n11792) );
  OAI21_X1 U14275 ( .B1(n11783), .B2(n11782), .A(n11781), .ZN(n11784) );
  NOR2_X1 U14276 ( .A1(n11785), .A2(n11784), .ZN(n11786) );
  XNOR2_X1 U14277 ( .A(n11785), .B(n11784), .ZN(n14869) );
  NOR2_X1 U14278 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14869), .ZN(n14868) );
  NOR2_X1 U14279 ( .A1(n11786), .A2(n14868), .ZN(n11790) );
  NAND2_X1 U14280 ( .A1(n11906), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11900) );
  INV_X1 U14281 ( .A(n11900), .ZN(n11787) );
  AOI21_X1 U14282 ( .B1(n8673), .B2(n11788), .A(n11787), .ZN(n11789) );
  NAND2_X1 U14283 ( .A1(n11789), .A2(n11790), .ZN(n11899) );
  OAI211_X1 U14284 ( .C1(n11790), .C2(n11789), .A(n14299), .B(n11899), .ZN(
        n11791) );
  NAND2_X1 U14285 ( .A1(n11792), .A2(n11791), .ZN(P1_U3259) );
  AOI21_X1 U14286 ( .B1(n11794), .B2(n11804), .A(n11793), .ZN(n11797) );
  AOI21_X1 U14287 ( .B1(n11797), .B2(n11796), .A(n11795), .ZN(n13919) );
  INV_X1 U14288 ( .A(n11812), .ZN(n11798) );
  AOI211_X1 U14289 ( .C1(n13918), .C2(n11799), .A(n12009), .B(n11798), .ZN(
        n13917) );
  INV_X1 U14290 ( .A(n11800), .ZN(n11801) );
  AOI22_X1 U14291 ( .A1(n15157), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11801), 
        .B2(n15154), .ZN(n11802) );
  OAI21_X1 U14292 ( .B1(n9708), .B2(n13813), .A(n11802), .ZN(n11806) );
  XOR2_X1 U14293 ( .A(n11804), .B(n11803), .Z(n13921) );
  NOR2_X1 U14294 ( .A1(n13921), .A2(n15139), .ZN(n11805) );
  AOI211_X1 U14295 ( .C1(n13917), .C2(n13835), .A(n11806), .B(n11805), .ZN(
        n11807) );
  OAI21_X1 U14296 ( .B1(n15157), .B2(n13919), .A(n11807), .ZN(P2_U3250) );
  XNOR2_X1 U14297 ( .A(n11808), .B(n11816), .ZN(n11810) );
  AOI21_X1 U14298 ( .B1(n11810), .B2(n15131), .A(n11809), .ZN(n13915) );
  OAI22_X1 U14299 ( .A1(n15155), .A2(n13620), .B1(n11811), .B2(n15132), .ZN(
        n11815) );
  AOI21_X1 U14300 ( .B1(n11812), .B2(n13911), .A(n13753), .ZN(n11813) );
  NAND2_X1 U14301 ( .A1(n11813), .A2(n13831), .ZN(n13913) );
  NOR2_X1 U14302 ( .A1(n13913), .A2(n15140), .ZN(n11814) );
  AOI211_X1 U14303 ( .C1(n15144), .C2(n13911), .A(n11815), .B(n11814), .ZN(
        n11821) );
  NOR2_X1 U14304 ( .A1(n11817), .A2(n11816), .ZN(n11818) );
  OR2_X1 U14305 ( .A1(n11819), .A2(n11818), .ZN(n13916) );
  OR2_X1 U14306 ( .A1(n13916), .A2(n15139), .ZN(n11820) );
  OAI211_X1 U14307 ( .C1(n13915), .C2(n15157), .A(n11821), .B(n11820), .ZN(
        P2_U3249) );
  XNOR2_X1 U14308 ( .A(n11822), .B(n12689), .ZN(n11893) );
  INV_X1 U14309 ( .A(n11893), .ZN(n11829) );
  INV_X1 U14310 ( .A(n12689), .ZN(n12786) );
  XNOR2_X1 U14311 ( .A(n11823), .B(n12786), .ZN(n11824) );
  OAI222_X1 U14312 ( .A1(n13312), .A2(n12940), .B1(n13314), .B2(n11941), .C1(
        n11824), .C2(n13310), .ZN(n11892) );
  INV_X1 U14313 ( .A(n11946), .ZN(n11898) );
  INV_X1 U14314 ( .A(n11944), .ZN(n11825) );
  AOI22_X1 U14315 ( .A1(n13328), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n13288), 
        .B2(n11825), .ZN(n11826) );
  OAI21_X1 U14316 ( .B1(n11898), .B2(n13341), .A(n11826), .ZN(n11827) );
  AOI21_X1 U14317 ( .B1(n11892), .B2(n13344), .A(n11827), .ZN(n11828) );
  OAI21_X1 U14318 ( .B1(n13305), .B2(n11829), .A(n11828), .ZN(P3_U3218) );
  NAND2_X1 U14319 ( .A1(n11831), .A2(n11830), .ZN(n11832) );
  XNOR2_X1 U14320 ( .A(n11832), .B(n11834), .ZN(n14597) );
  INV_X1 U14321 ( .A(n14597), .ZN(n11844) );
  OAI211_X1 U14322 ( .C1(n11835), .C2(n11834), .A(n11833), .B(n14899), .ZN(
        n11836) );
  AOI22_X1 U14323 ( .A1(n14145), .A2(n14111), .B1(n14110), .B2(n14143), .ZN(
        n14120) );
  NAND2_X1 U14324 ( .A1(n11836), .A2(n14120), .ZN(n14598) );
  INV_X1 U14325 ( .A(n14647), .ZN(n14128) );
  AOI21_X1 U14326 ( .B1(n14647), .B2(n11837), .A(n14909), .ZN(n11838) );
  AND2_X1 U14327 ( .A1(n11838), .A2(n11917), .ZN(n14599) );
  NAND2_X1 U14328 ( .A1(n14599), .A2(n14911), .ZN(n11841) );
  INV_X1 U14329 ( .A(n11839), .ZN(n14123) );
  INV_X1 U14330 ( .A(n14507), .ZN(n14910) );
  AOI22_X1 U14331 ( .A1(n6653), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14123), 
        .B2(n14910), .ZN(n11840) );
  OAI211_X1 U14332 ( .C1(n14128), .C2(n14925), .A(n11841), .B(n11840), .ZN(
        n11842) );
  AOI21_X1 U14333 ( .B1(n14598), .B2(n14923), .A(n11842), .ZN(n11843) );
  OAI21_X1 U14334 ( .B1(n14518), .B2(n11844), .A(n11843), .ZN(P1_U3278) );
  INV_X1 U14335 ( .A(n11848), .ZN(n12787) );
  XNOR2_X1 U14336 ( .A(n11845), .B(n12787), .ZN(n11846) );
  OAI222_X1 U14337 ( .A1(n13314), .A2(n12824), .B1(n13312), .B2(n12944), .C1(
        n11846), .C2(n13310), .ZN(n13406) );
  INV_X1 U14338 ( .A(n13406), .ZN(n11853) );
  OAI21_X1 U14339 ( .B1(n11849), .B2(n11848), .A(n11847), .ZN(n13407) );
  NOR2_X1 U14340 ( .A1(n13457), .A2(n13341), .ZN(n11851) );
  OAI22_X1 U14341 ( .A1(n13344), .A2(n12100), .B1(n12947), .B2(n15238), .ZN(
        n11850) );
  AOI211_X1 U14342 ( .C1(n13407), .C2(n13347), .A(n11851), .B(n11850), .ZN(
        n11852) );
  OAI21_X1 U14343 ( .B1(n11853), .B2(n15258), .A(n11852), .ZN(P3_U3217) );
  NAND2_X1 U14344 ( .A1(n11855), .A2(n11854), .ZN(n11857) );
  NAND2_X1 U14345 ( .A1(n11857), .A2(n11856), .ZN(n11859) );
  XNOR2_X1 U14346 ( .A(n11858), .B(n12903), .ZN(n11932) );
  XNOR2_X1 U14347 ( .A(n11932), .B(n13054), .ZN(n11860) );
  NAND2_X1 U14348 ( .A1(n11859), .A2(n11860), .ZN(n11935) );
  OAI211_X1 U14349 ( .C1(n11859), .C2(n11860), .A(n11935), .B(n12995), .ZN(
        n11865) );
  NAND2_X1 U14350 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13084)
         );
  OAI21_X1 U14351 ( .B1(n13028), .B2(n12824), .A(n13084), .ZN(n11863) );
  NOR2_X1 U14352 ( .A1(n13031), .A2(n11861), .ZN(n11862) );
  AOI211_X1 U14353 ( .C1(n13017), .C2(n13055), .A(n11863), .B(n11862), .ZN(
        n11864) );
  OAI211_X1 U14354 ( .C1(n14784), .C2(n13003), .A(n11865), .B(n11864), .ZN(
        P3_U3155) );
  NOR2_X1 U14355 ( .A1(n11866), .A2(n14895), .ZN(n11869) );
  NOR3_X1 U14356 ( .A1(n11869), .A2(n11868), .A3(n11867), .ZN(n11872) );
  INV_X1 U14357 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11870) );
  MUX2_X1 U14358 ( .A(n11872), .B(n11870), .S(n14985), .Z(n11871) );
  OAI21_X1 U14359 ( .B1(n7202), .B2(n14643), .A(n11871), .ZN(P1_U3501) );
  MUX2_X1 U14360 ( .A(n11872), .B(n11775), .S(n14991), .Z(n11873) );
  OAI21_X1 U14361 ( .B1(n7202), .B2(n14596), .A(n11873), .ZN(P1_U3542) );
  INV_X1 U14362 ( .A(n11874), .ZN(n11877) );
  OAI222_X1 U14363 ( .A1(P1_U3086), .A2(n11875), .B1(n6656), .B2(n11877), .C1(
        n15601), .C2(n12562), .ZN(P1_U3329) );
  OAI222_X1 U14364 ( .A1(n11878), .A2(P2_U3088), .B1(n13955), .B2(n11877), 
        .C1(n11876), .C2(n13960), .ZN(P2_U3301) );
  AOI22_X1 U14365 ( .A1(n12377), .A2(n12267), .B1(n12268), .B2(n14148), .ZN(
        n12141) );
  AOI22_X1 U14366 ( .A1(n12377), .A2(n12262), .B1(n12267), .B2(n14148), .ZN(
        n11879) );
  XNOR2_X1 U14367 ( .A(n11879), .B(n12265), .ZN(n12140) );
  XOR2_X1 U14368 ( .A(n12141), .B(n12140), .Z(n11884) );
  AOI21_X1 U14369 ( .B1(n11882), .B2(n11881), .A(n11880), .ZN(n11883) );
  NAND2_X1 U14370 ( .A1(n11883), .A2(n11884), .ZN(n12143) );
  OAI21_X1 U14371 ( .B1(n11884), .B2(n11883), .A(n12143), .ZN(n11885) );
  NAND2_X1 U14372 ( .A1(n11885), .A2(n14828), .ZN(n11891) );
  INV_X1 U14373 ( .A(n11886), .ZN(n14838) );
  OAI22_X1 U14374 ( .A1(n14121), .A2(n11888), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11887), .ZN(n11889) );
  AOI21_X1 U14375 ( .B1(n14124), .B2(n14838), .A(n11889), .ZN(n11890) );
  OAI211_X1 U14376 ( .C1(n14841), .C2(n14127), .A(n11891), .B(n11890), .ZN(
        P1_U3236) );
  INV_X1 U14377 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n11894) );
  AOI21_X1 U14378 ( .B1(n11893), .B2(n15298), .A(n11892), .ZN(n11896) );
  MUX2_X1 U14379 ( .A(n11894), .B(n11896), .S(n15309), .Z(n11895) );
  OAI21_X1 U14380 ( .B1(n11898), .B2(n13456), .A(n11895), .ZN(P3_U3435) );
  MUX2_X1 U14381 ( .A(n13110), .B(n11896), .S(n15699), .Z(n11897) );
  OAI21_X1 U14382 ( .B1(n11898), .B2(n13409), .A(n11897), .ZN(P3_U3474) );
  NAND2_X1 U14383 ( .A1(n11900), .A2(n11899), .ZN(n11903) );
  INV_X1 U14384 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14277) );
  NOR2_X1 U14385 ( .A1(n14276), .A2(n14277), .ZN(n11901) );
  AOI21_X1 U14386 ( .B1(n14277), .B2(n14276), .A(n11901), .ZN(n11902) );
  NAND2_X1 U14387 ( .A1(n11902), .A2(n11903), .ZN(n14275) );
  OAI211_X1 U14388 ( .C1(n11903), .C2(n11902), .A(n14299), .B(n14275), .ZN(
        n11912) );
  INV_X1 U14389 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n11904) );
  NAND2_X1 U14390 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14049)
         );
  OAI21_X1 U14391 ( .B1(n14878), .B2(n11904), .A(n14049), .ZN(n11910) );
  AOI21_X1 U14392 ( .B1(n11906), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11905), 
        .ZN(n11908) );
  XNOR2_X1 U14393 ( .A(n14270), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11907) );
  NOR2_X1 U14394 ( .A1(n11908), .A2(n11907), .ZN(n14269) );
  AOI211_X1 U14395 ( .C1(n11908), .C2(n11907), .A(n14269), .B(n14295), .ZN(
        n11909) );
  AOI211_X1 U14396 ( .C1(n14293), .C2(n14270), .A(n11910), .B(n11909), .ZN(
        n11911) );
  NAND2_X1 U14397 ( .A1(n11912), .A2(n11911), .ZN(P1_U3260) );
  XOR2_X1 U14398 ( .A(n11913), .B(n12531), .Z(n11914) );
  AOI22_X1 U14399 ( .A1(n14111), .A2(n14144), .B1(n14142), .B2(n14110), .ZN(
        n14037) );
  OAI21_X1 U14400 ( .B1(n11914), .B2(n14921), .A(n14037), .ZN(n14591) );
  INV_X1 U14401 ( .A(n14591), .ZN(n11922) );
  OAI21_X1 U14402 ( .B1(n11916), .B2(n12531), .A(n11915), .ZN(n14593) );
  INV_X1 U14403 ( .A(n14039), .ZN(n14644) );
  AOI211_X1 U14404 ( .C1(n14039), .C2(n11917), .A(n14909), .B(n14510), .ZN(
        n14592) );
  NAND2_X1 U14405 ( .A1(n14592), .A2(n14911), .ZN(n11919) );
  AOI22_X1 U14406 ( .A1(n6653), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n14034), 
        .B2(n14910), .ZN(n11918) );
  OAI211_X1 U14407 ( .C1(n14644), .C2(n14925), .A(n11919), .B(n11918), .ZN(
        n11920) );
  AOI21_X1 U14408 ( .B1(n14593), .B2(n14843), .A(n11920), .ZN(n11921) );
  OAI21_X1 U14409 ( .B1(n11922), .B2(n6653), .A(n11921), .ZN(P1_U3277) );
  XNOR2_X1 U14410 ( .A(n11923), .B(n12789), .ZN(n13403) );
  INV_X1 U14411 ( .A(n13403), .ZN(n11931) );
  OAI211_X1 U14412 ( .C1(n11924), .C2(n8016), .A(n15248), .B(n13330), .ZN(
        n11926) );
  AOI22_X1 U14413 ( .A1(n13051), .A2(n15242), .B1(n15244), .B2(n13052), .ZN(
        n11925) );
  NAND2_X1 U14414 ( .A1(n11926), .A2(n11925), .ZN(n13402) );
  INV_X1 U14415 ( .A(n12968), .ZN(n13452) );
  INV_X1 U14416 ( .A(n12966), .ZN(n11927) );
  AOI22_X1 U14417 ( .A1(n13328), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13288), 
        .B2(n11927), .ZN(n11928) );
  OAI21_X1 U14418 ( .B1(n13452), .B2(n13341), .A(n11928), .ZN(n11929) );
  AOI21_X1 U14419 ( .B1(n13402), .B2(n13344), .A(n11929), .ZN(n11930) );
  OAI21_X1 U14420 ( .B1(n11931), .B2(n13305), .A(n11930), .ZN(P3_U3216) );
  XNOR2_X1 U14421 ( .A(n11946), .B(n12856), .ZN(n12825) );
  XNOR2_X1 U14422 ( .A(n12825), .B(n12824), .ZN(n11940) );
  INV_X1 U14423 ( .A(n11932), .ZN(n11933) );
  NAND2_X1 U14424 ( .A1(n11933), .A2(n13054), .ZN(n11934) );
  NAND2_X1 U14425 ( .A1(n11935), .A2(n11934), .ZN(n11939) );
  INV_X1 U14426 ( .A(n11939), .ZN(n11937) );
  INV_X1 U14427 ( .A(n11940), .ZN(n11936) );
  NAND2_X1 U14428 ( .A1(n11937), .A2(n11936), .ZN(n12827) );
  INV_X1 U14429 ( .A(n12827), .ZN(n11938) );
  AOI21_X1 U14430 ( .B1(n11940), .B2(n11939), .A(n11938), .ZN(n11948) );
  NAND2_X1 U14431 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13100)
         );
  OAI21_X1 U14432 ( .B1(n13041), .B2(n11941), .A(n13100), .ZN(n11942) );
  AOI21_X1 U14433 ( .B1(n13037), .B2(n13052), .A(n11942), .ZN(n11943) );
  OAI21_X1 U14434 ( .B1(n11944), .B2(n13031), .A(n11943), .ZN(n11945) );
  AOI21_X1 U14435 ( .B1(n13044), .B2(n11946), .A(n11945), .ZN(n11947) );
  OAI21_X1 U14436 ( .B1(n11948), .B2(n13046), .A(n11947), .ZN(P3_U3181) );
  AND2_X1 U14437 ( .A1(n11951), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U14438 ( .A1(n11951), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U14439 ( .A1(n11951), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U14440 ( .A1(n11951), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U14441 ( .A1(n11951), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U14442 ( .A1(n11951), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U14443 ( .A1(n11951), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U14444 ( .A1(n11951), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U14445 ( .A1(n11951), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U14446 ( .A1(n11951), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U14447 ( .A1(n11951), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U14448 ( .A1(n11951), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U14449 ( .A1(n11951), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U14450 ( .A1(n11951), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U14451 ( .A1(n11951), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U14452 ( .A1(n11951), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U14453 ( .A1(n11951), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U14454 ( .A1(n11951), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U14455 ( .A1(n11951), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U14456 ( .A1(n11951), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U14457 ( .A1(n11951), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U14458 ( .A1(n11951), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U14459 ( .A1(n11951), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U14460 ( .A1(n11951), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U14461 ( .A1(n11951), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U14462 ( .A1(n11951), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U14463 ( .A1(n11951), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U14464 ( .A1(n11951), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U14465 ( .A1(n11951), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U14466 ( .A1(n11951), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  INV_X1 U14467 ( .A(n11952), .ZN(n11953) );
  NAND2_X1 U14468 ( .A1(n11954), .A2(n11953), .ZN(n11956) );
  NAND2_X1 U14469 ( .A1(n14656), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11955) );
  INV_X1 U14470 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12055) );
  XNOR2_X1 U14471 ( .A(n12055), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11957) );
  XNOR2_X1 U14472 ( .A(n12598), .B(n11957), .ZN(n12586) );
  INV_X1 U14473 ( .A(n12586), .ZN(n11958) );
  OAI222_X1 U14474 ( .A1(n11960), .A2(P3_U3151), .B1(n12584), .B2(n11959), 
        .C1(n6655), .C2(n11958), .ZN(P3_U3265) );
  INV_X1 U14475 ( .A(n11961), .ZN(n11964) );
  OAI222_X1 U14476 ( .A1(n6655), .A2(n11964), .B1(P3_U3151), .B2(n11963), .C1(
        n11962), .C2(n12584), .ZN(P3_U3266) );
  INV_X1 U14477 ( .A(n11965), .ZN(n13958) );
  OAI222_X1 U14478 ( .A1(n12562), .A2(n11966), .B1(n6656), .B2(n13958), .C1(
        P1_U3086), .C2(n6734), .ZN(P1_U3328) );
  INV_X1 U14479 ( .A(n11967), .ZN(n13956) );
  OAI222_X1 U14480 ( .A1(n12562), .A2(n11969), .B1(n6656), .B2(n13956), .C1(
        n11968), .C2(P1_U3086), .ZN(P1_U3327) );
  NAND2_X1 U14481 ( .A1(n11971), .A2(n11970), .ZN(n13498) );
  AOI22_X1 U14482 ( .A1(n13547), .A2(n13606), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13498), .ZN(n11975) );
  AOI21_X1 U14483 ( .B1(n13753), .B2(n11972), .A(n14999), .ZN(n11973) );
  OAI21_X1 U14484 ( .B1(n11973), .B2(n15004), .A(n9661), .ZN(n11974) );
  OAI211_X1 U14485 ( .C1(n11976), .C2(n13561), .A(n11975), .B(n11974), .ZN(
        P2_U3204) );
  XNOR2_X1 U14486 ( .A(n13886), .B(n11494), .ZN(n11989) );
  INV_X1 U14487 ( .A(n11989), .ZN(n11991) );
  NAND2_X1 U14488 ( .A1(n13586), .A2(n12009), .ZN(n11990) );
  XNOR2_X1 U14489 ( .A(n13891), .B(n11494), .ZN(n11986) );
  INV_X1 U14490 ( .A(n11986), .ZN(n11988) );
  NOR2_X1 U14491 ( .A1(n13513), .A2(n15134), .ZN(n11985) );
  INV_X1 U14492 ( .A(n11985), .ZN(n11987) );
  XNOR2_X1 U14493 ( .A(n13896), .B(n12029), .ZN(n13562) );
  NAND2_X1 U14494 ( .A1(n13588), .A2(n12009), .ZN(n11984) );
  NOR2_X1 U14495 ( .A1(n13568), .A2(n15134), .ZN(n11980) );
  XNOR2_X1 U14496 ( .A(n13907), .B(n11494), .ZN(n11979) );
  INV_X1 U14497 ( .A(n11977), .ZN(n11978) );
  XOR2_X1 U14498 ( .A(n11980), .B(n11979), .Z(n12289) );
  OAI21_X1 U14499 ( .B1(n11980), .B2(n11979), .A(n12295), .ZN(n13573) );
  XNOR2_X1 U14500 ( .A(n13814), .B(n12029), .ZN(n13491) );
  NOR2_X1 U14501 ( .A1(n13488), .A2(n15134), .ZN(n11981) );
  NAND2_X1 U14502 ( .A1(n13491), .A2(n11981), .ZN(n11982) );
  OAI21_X1 U14503 ( .B1(n13491), .B2(n11981), .A(n11982), .ZN(n13572) );
  NOR2_X2 U14504 ( .A1(n13573), .A2(n13572), .ZN(n13571) );
  INV_X1 U14505 ( .A(n11982), .ZN(n11983) );
  XNOR2_X1 U14506 ( .A(n13562), .B(n11984), .ZN(n13494) );
  XNOR2_X1 U14507 ( .A(n11986), .B(n11985), .ZN(n13564) );
  XNOR2_X1 U14508 ( .A(n11989), .B(n11990), .ZN(n13511) );
  XNOR2_X1 U14509 ( .A(n13881), .B(n11494), .ZN(n11993) );
  XNOR2_X1 U14510 ( .A(n11994), .B(n11993), .ZN(n12564) );
  INV_X1 U14511 ( .A(n13585), .ZN(n13514) );
  NAND2_X1 U14512 ( .A1(n13585), .A2(n12009), .ZN(n11992) );
  NOR2_X1 U14513 ( .A1(n12564), .A2(n11992), .ZN(n12570) );
  AND2_X1 U14514 ( .A1(n11994), .A2(n11993), .ZN(n11995) );
  XNOR2_X1 U14515 ( .A(n13876), .B(n11494), .ZN(n11998) );
  XNOR2_X1 U14516 ( .A(n13871), .B(n12029), .ZN(n13520) );
  NAND2_X1 U14517 ( .A1(n13583), .A2(n12009), .ZN(n12001) );
  NOR2_X1 U14518 ( .A1(n13520), .A2(n12001), .ZN(n12002) );
  AOI21_X1 U14519 ( .B1(n13520), .B2(n12001), .A(n12002), .ZN(n13532) );
  INV_X1 U14520 ( .A(n12002), .ZN(n12007) );
  XNOR2_X1 U14521 ( .A(n13866), .B(n11494), .ZN(n12003) );
  AND2_X1 U14522 ( .A1(n13582), .A2(n13753), .ZN(n12004) );
  NAND2_X1 U14523 ( .A1(n12003), .A2(n12004), .ZN(n12008) );
  INV_X1 U14524 ( .A(n12003), .ZN(n12012) );
  INV_X1 U14525 ( .A(n12004), .ZN(n12005) );
  NAND2_X1 U14526 ( .A1(n12012), .A2(n12005), .ZN(n12006) );
  NAND2_X1 U14527 ( .A1(n12008), .A2(n12006), .ZN(n13522) );
  INV_X1 U14528 ( .A(n12008), .ZN(n12010) );
  XNOR2_X1 U14529 ( .A(n13694), .B(n11494), .ZN(n12025) );
  NAND2_X1 U14530 ( .A1(n13581), .A2(n12009), .ZN(n12024) );
  XNOR2_X1 U14531 ( .A(n12025), .B(n12024), .ZN(n12013) );
  NOR2_X1 U14532 ( .A1(n6754), .A2(n14999), .ZN(n12015) );
  NOR3_X1 U14533 ( .A1(n12012), .A2(n12011), .A3(n13561), .ZN(n12014) );
  OAI21_X1 U14534 ( .B1(n12015), .B2(n12014), .A(n12013), .ZN(n12023) );
  OR2_X1 U14535 ( .A1(n12036), .A2(n15148), .ZN(n12017) );
  NAND2_X1 U14536 ( .A1(n13582), .A2(n15127), .ZN(n12016) );
  NAND2_X1 U14537 ( .A1(n12017), .A2(n12016), .ZN(n13688) );
  INV_X1 U14538 ( .A(n13692), .ZN(n12019) );
  OAI22_X1 U14539 ( .A1(n12019), .A2(n15007), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12018), .ZN(n12021) );
  NOR2_X1 U14540 ( .A1(n13694), .A2(n13539), .ZN(n12020) );
  AOI211_X1 U14541 ( .C1(n13515), .C2(n13688), .A(n12021), .B(n12020), .ZN(
        n12022) );
  OAI211_X1 U14542 ( .C1(n14999), .C2(n12026), .A(n12023), .B(n12022), .ZN(
        P2_U3212) );
  INV_X1 U14543 ( .A(n12024), .ZN(n12028) );
  INV_X1 U14544 ( .A(n12025), .ZN(n12027) );
  XNOR2_X1 U14545 ( .A(n13678), .B(n12029), .ZN(n12031) );
  NOR2_X1 U14546 ( .A1(n12036), .A2(n15134), .ZN(n12030) );
  NAND2_X1 U14547 ( .A1(n12031), .A2(n12030), .ZN(n12032) );
  OAI21_X1 U14548 ( .B1(n12031), .B2(n12030), .A(n12032), .ZN(n13469) );
  NOR2_X1 U14549 ( .A1(n13473), .A2(n15134), .ZN(n12034) );
  XNOR2_X1 U14550 ( .A(n12034), .B(n11494), .ZN(n12035) );
  OR2_X1 U14551 ( .A1(n12036), .A2(n13567), .ZN(n12037) );
  OAI21_X1 U14552 ( .B1(n12038), .B2(n15148), .A(n12037), .ZN(n13668) );
  OAI22_X1 U14553 ( .A1(n13661), .A2(n15007), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12039), .ZN(n12041) );
  NOR2_X1 U14554 ( .A1(n13851), .A2(n13539), .ZN(n12040) );
  AOI211_X1 U14555 ( .C1(n13515), .C2(n13668), .A(n12041), .B(n12040), .ZN(
        n12042) );
  INV_X1 U14556 ( .A(n13498), .ZN(n12044) );
  OAI22_X1 U14557 ( .A1(n14997), .A2(n12045), .B1(n12044), .B2(n12043), .ZN(
        n12046) );
  AOI21_X1 U14558 ( .B1(n12047), .B2(n15004), .A(n12046), .ZN(n12053) );
  OAI22_X1 U14559 ( .A1(n13561), .A2(n9542), .B1(n12048), .B2(n14999), .ZN(
        n12051) );
  INV_X1 U14560 ( .A(n12049), .ZN(n12050) );
  NAND3_X1 U14561 ( .A1(n12051), .A2(n12050), .A3(n13502), .ZN(n12052) );
  OAI211_X1 U14562 ( .C1(n14999), .C2(n12054), .A(n12053), .B(n12052), .ZN(
        P2_U3209) );
  INV_X1 U14563 ( .A(n12484), .ZN(n12563) );
  OAI222_X1 U14564 ( .A1(n13955), .A2(n12563), .B1(P2_U3088), .B2(n8943), .C1(
        n12055), .C2(n13960), .ZN(P2_U3297) );
  NOR2_X1 U14565 ( .A1(n13072), .A2(n12057), .ZN(n12058) );
  NAND2_X1 U14566 ( .A1(n12077), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12094) );
  OAI21_X1 U14567 ( .B1(n12077), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12094), 
        .ZN(n13080) );
  NOR2_X1 U14568 ( .A1(n13081), .A2(n13080), .ZN(n13079) );
  INV_X1 U14569 ( .A(n13079), .ZN(n12059) );
  AND2_X1 U14570 ( .A1(n12060), .A2(n12061), .ZN(n12062) );
  NAND2_X1 U14571 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12083), .ZN(n12063) );
  OAI21_X1 U14572 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12083), .A(n12063), 
        .ZN(n13116) );
  INV_X1 U14573 ( .A(n12065), .ZN(n12066) );
  OR2_X1 U14574 ( .A1(n12066), .A2(n13148), .ZN(n13156) );
  OR2_X1 U14575 ( .A1(n13167), .A2(n13343), .ZN(n12068) );
  NAND2_X1 U14576 ( .A1(n13167), .A2(n13343), .ZN(n12067) );
  NAND2_X1 U14577 ( .A1(n12068), .A2(n12067), .ZN(n13155) );
  INV_X1 U14578 ( .A(n12068), .ZN(n12069) );
  NOR2_X1 U14579 ( .A1(n13160), .A2(n12069), .ZN(n12070) );
  XNOR2_X1 U14580 ( .A(n12800), .B(n13320), .ZN(n12107) );
  XNOR2_X1 U14581 ( .A(n12070), .B(n12107), .ZN(n12111) );
  INV_X1 U14582 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15669) );
  AND2_X1 U14583 ( .A1(n12073), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12074) );
  NOR2_X1 U14584 ( .A1(n13072), .A2(n12075), .ZN(n12076) );
  NAND2_X1 U14585 ( .A1(n12077), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12078) );
  OAI21_X1 U14586 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n12077), .A(n12078), 
        .ZN(n13082) );
  INV_X1 U14587 ( .A(n12078), .ZN(n12095) );
  NOR2_X1 U14588 ( .A1(n12079), .A2(n12095), .ZN(n12080) );
  NOR2_X1 U14589 ( .A1(n13107), .A2(n12080), .ZN(n12081) );
  NAND2_X1 U14590 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12083), .ZN(n12082) );
  OAI21_X1 U14591 ( .B1(n12083), .B2(P3_REG1_REG_16__SCAN_IN), .A(n12082), 
        .ZN(n13127) );
  NOR2_X1 U14592 ( .A1(n12085), .A2(n13138), .ZN(n13162) );
  NAND2_X1 U14593 ( .A1(n12086), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12087) );
  OAI21_X1 U14594 ( .B1(n12086), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12087), 
        .ZN(n13161) );
  INV_X1 U14595 ( .A(n12087), .ZN(n12088) );
  XNOR2_X1 U14596 ( .A(n12800), .B(n13395), .ZN(n12106) );
  NAND2_X1 U14597 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12894)
         );
  MUX2_X1 U14598 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6648), .Z(n12103) );
  INV_X1 U14599 ( .A(n12089), .ZN(n12091) );
  NOR2_X1 U14600 ( .A1(n12091), .A2(n12090), .ZN(n13066) );
  MUX2_X1 U14601 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12105), .Z(n12093) );
  XNOR2_X1 U14602 ( .A(n12093), .B(n12092), .ZN(n13065) );
  NOR2_X1 U14603 ( .A1(n12093), .A2(n12092), .ZN(n13086) );
  MUX2_X1 U14604 ( .A(n13080), .B(n13082), .S(n12105), .Z(n13090) );
  INV_X1 U14605 ( .A(n12094), .ZN(n12096) );
  MUX2_X1 U14606 ( .A(n12096), .B(n12095), .S(n12105), .Z(n12097) );
  XNOR2_X1 U14607 ( .A(n12098), .B(n12060), .ZN(n13103) );
  MUX2_X1 U14608 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6648), .Z(n13102) );
  NOR2_X1 U14609 ( .A1(n13103), .A2(n13102), .ZN(n13101) );
  AOI21_X1 U14610 ( .B1(n12099), .B2(n13107), .A(n13101), .ZN(n13121) );
  MUX2_X1 U14611 ( .A(n12100), .B(n15443), .S(n12105), .Z(n12101) );
  NOR2_X1 U14612 ( .A1(n12101), .A2(n13122), .ZN(n13117) );
  NAND2_X1 U14613 ( .A1(n12101), .A2(n13122), .ZN(n13118) );
  OAI21_X1 U14614 ( .B1(n13121), .B2(n13117), .A(n13118), .ZN(n13144) );
  XNOR2_X1 U14615 ( .A(n12103), .B(n12102), .ZN(n13145) );
  NOR2_X1 U14616 ( .A1(n13144), .A2(n13145), .ZN(n13143) );
  AOI21_X1 U14617 ( .B1(n12103), .B2(n12102), .A(n13143), .ZN(n12104) );
  XNOR2_X1 U14618 ( .A(n12104), .B(n13167), .ZN(n13153) );
  MUX2_X1 U14619 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6648), .Z(n13154) );
  NOR2_X1 U14620 ( .A1(n13153), .A2(n13154), .ZN(n13152) );
  MUX2_X1 U14621 ( .A(n12107), .B(n12106), .S(n12105), .Z(n12108) );
  OAI21_X1 U14622 ( .B1(n12111), .B2(n13150), .A(n12110), .ZN(P3_U3201) );
  NAND2_X1 U14623 ( .A1(n13552), .A2(n12112), .ZN(n12113) );
  OAI21_X1 U14624 ( .B1(n13561), .B2(n12114), .A(n12113), .ZN(n12115) );
  NAND3_X1 U14625 ( .A1(n12117), .A2(n12116), .A3(n12115), .ZN(n12124) );
  OAI22_X1 U14626 ( .A1(n15007), .A2(n12119), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12118), .ZN(n12120) );
  INV_X1 U14627 ( .A(n12120), .ZN(n12123) );
  AOI22_X1 U14628 ( .A1(n13547), .A2(n13597), .B1(n13541), .B2(n13600), .ZN(
        n12122) );
  OR2_X1 U14629 ( .A1(n13539), .A2(n7073), .ZN(n12121) );
  AND4_X1 U14630 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12125) );
  OAI21_X1 U14631 ( .B1(n12126), .B2(n14999), .A(n12125), .ZN(P2_U3203) );
  AOI22_X1 U14632 ( .A1(n13515), .A2(n12127), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12128) );
  OAI21_X1 U14633 ( .B1(n12129), .B2(n15007), .A(n12128), .ZN(n12137) );
  INV_X1 U14634 ( .A(n12130), .ZN(n14998) );
  NOR3_X1 U14635 ( .A1(n12132), .A2(n12131), .A3(n13561), .ZN(n12133) );
  AOI21_X1 U14636 ( .B1(n14998), .B2(n13552), .A(n12133), .ZN(n12135) );
  NOR2_X1 U14637 ( .A1(n12135), .A2(n12134), .ZN(n12136) );
  AOI211_X1 U14638 ( .C1(n11505), .C2(n15004), .A(n12137), .B(n12136), .ZN(
        n12138) );
  OAI21_X1 U14639 ( .B1(n12139), .B2(n14999), .A(n12138), .ZN(P2_U3187) );
  NAND2_X1 U14640 ( .A1(n12140), .A2(n12141), .ZN(n12142) );
  NAND2_X1 U14641 ( .A1(n12143), .A2(n12142), .ZN(n14006) );
  NOR2_X1 U14642 ( .A1(n10622), .A2(n12144), .ZN(n12145) );
  AOI21_X1 U14643 ( .B1(n12382), .B2(n12267), .A(n12145), .ZN(n12150) );
  NAND2_X1 U14644 ( .A1(n12382), .A2(n12262), .ZN(n12147) );
  NAND2_X1 U14645 ( .A1(n12267), .A2(n14147), .ZN(n12146) );
  NAND2_X1 U14646 ( .A1(n12147), .A2(n12146), .ZN(n12148) );
  XNOR2_X1 U14647 ( .A(n12148), .B(n12265), .ZN(n12149) );
  XOR2_X1 U14648 ( .A(n12150), .B(n12149), .Z(n14005) );
  INV_X1 U14649 ( .A(n12149), .ZN(n12151) );
  OAI22_X1 U14650 ( .A1(n14081), .A2(n12275), .B1(n12389), .B2(n12274), .ZN(
        n12152) );
  XNOR2_X1 U14651 ( .A(n12152), .B(n12265), .ZN(n12159) );
  NOR2_X1 U14652 ( .A1(n10622), .A2(n12389), .ZN(n12153) );
  AOI21_X1 U14653 ( .B1(n12387), .B2(n12267), .A(n12153), .ZN(n12160) );
  XNOR2_X1 U14654 ( .A(n12159), .B(n12160), .ZN(n14072) );
  NAND2_X1 U14655 ( .A1(n14832), .A2(n12262), .ZN(n12155) );
  NAND2_X1 U14656 ( .A1(n14145), .A2(n12267), .ZN(n12154) );
  NAND2_X1 U14657 ( .A1(n12155), .A2(n12154), .ZN(n12156) );
  XNOR2_X1 U14658 ( .A(n12156), .B(n12265), .ZN(n12163) );
  NOR2_X1 U14659 ( .A1(n10622), .A2(n12157), .ZN(n12158) );
  AOI21_X1 U14660 ( .B1(n14832), .B2(n12267), .A(n12158), .ZN(n12164) );
  XNOR2_X1 U14661 ( .A(n12163), .B(n12164), .ZN(n14826) );
  INV_X1 U14662 ( .A(n12159), .ZN(n12161) );
  OR2_X1 U14663 ( .A1(n12161), .A2(n12160), .ZN(n14824) );
  INV_X1 U14664 ( .A(n12163), .ZN(n12165) );
  NAND2_X1 U14665 ( .A1(n14647), .A2(n12262), .ZN(n12167) );
  NAND2_X1 U14666 ( .A1(n14144), .A2(n12267), .ZN(n12166) );
  NAND2_X1 U14667 ( .A1(n12167), .A2(n12166), .ZN(n12168) );
  XNOR2_X1 U14668 ( .A(n12168), .B(n12265), .ZN(n14028) );
  NAND2_X1 U14669 ( .A1(n14647), .A2(n12267), .ZN(n12170) );
  NAND2_X1 U14670 ( .A1(n12268), .A2(n14144), .ZN(n12169) );
  NAND2_X1 U14671 ( .A1(n12170), .A2(n12169), .ZN(n14118) );
  NAND2_X1 U14672 ( .A1(n14039), .A2(n12262), .ZN(n12172) );
  NAND2_X1 U14673 ( .A1(n12267), .A2(n14143), .ZN(n12171) );
  NAND2_X1 U14674 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  XNOR2_X1 U14675 ( .A(n12173), .B(n12265), .ZN(n14030) );
  NAND2_X1 U14676 ( .A1(n14039), .A2(n12267), .ZN(n12175) );
  NAND2_X1 U14677 ( .A1(n12268), .A2(n14143), .ZN(n12174) );
  NAND2_X1 U14678 ( .A1(n12175), .A2(n12174), .ZN(n14031) );
  AND2_X1 U14679 ( .A1(n14030), .A2(n14031), .ZN(n12176) );
  AOI21_X1 U14680 ( .B1(n14028), .B2(n14118), .A(n12176), .ZN(n12181) );
  INV_X1 U14681 ( .A(n12176), .ZN(n12178) );
  INV_X1 U14682 ( .A(n14118), .ZN(n12177) );
  NAND2_X1 U14683 ( .A1(n12178), .A2(n12177), .ZN(n12179) );
  OAI22_X1 U14684 ( .A1(n14028), .A2(n12179), .B1(n14031), .B2(n14030), .ZN(
        n12180) );
  OAI22_X1 U14685 ( .A1(n14514), .A2(n12275), .B1(n12406), .B2(n12274), .ZN(
        n12182) );
  XNOR2_X1 U14686 ( .A(n12182), .B(n6749), .ZN(n14044) );
  OR2_X1 U14687 ( .A1(n14514), .A2(n12274), .ZN(n12184) );
  NAND2_X1 U14688 ( .A1(n12268), .A2(n14142), .ZN(n12183) );
  AND2_X1 U14689 ( .A1(n12184), .A2(n12183), .ZN(n12186) );
  NAND2_X1 U14690 ( .A1(n14044), .A2(n12186), .ZN(n12185) );
  INV_X1 U14691 ( .A(n14044), .ZN(n12187) );
  INV_X1 U14692 ( .A(n12186), .ZN(n14043) );
  NAND2_X1 U14693 ( .A1(n12187), .A2(n14043), .ZN(n12188) );
  AOI22_X1 U14694 ( .A1(n14583), .A2(n12262), .B1(n12267), .B2(n14141), .ZN(
        n12189) );
  XNOR2_X1 U14695 ( .A(n12189), .B(n12265), .ZN(n12195) );
  AOI22_X1 U14696 ( .A1(n14583), .A2(n12267), .B1(n12268), .B2(n14141), .ZN(
        n12196) );
  XNOR2_X1 U14697 ( .A(n12195), .B(n12196), .ZN(n14094) );
  INV_X1 U14698 ( .A(n14094), .ZN(n12190) );
  NAND2_X1 U14699 ( .A1(n14637), .A2(n12262), .ZN(n12192) );
  OR2_X1 U14700 ( .A1(n14096), .A2(n12274), .ZN(n12191) );
  NAND2_X1 U14701 ( .A1(n12192), .A2(n12191), .ZN(n12193) );
  XNOR2_X1 U14702 ( .A(n12193), .B(n6749), .ZN(n12201) );
  NOR2_X1 U14703 ( .A1(n14096), .A2(n10622), .ZN(n12194) );
  AOI21_X1 U14704 ( .B1(n14637), .B2(n12267), .A(n12194), .ZN(n12200) );
  XNOR2_X1 U14705 ( .A(n12201), .B(n12200), .ZN(n13989) );
  INV_X1 U14706 ( .A(n12195), .ZN(n12198) );
  INV_X1 U14707 ( .A(n12196), .ZN(n12197) );
  NOR2_X1 U14708 ( .A1(n12198), .A2(n12197), .ZN(n13990) );
  NOR2_X1 U14709 ( .A1(n13989), .A2(n13990), .ZN(n12199) );
  NAND2_X1 U14710 ( .A1(n13988), .A2(n12199), .ZN(n13991) );
  OR2_X1 U14711 ( .A1(n12201), .A2(n12200), .ZN(n12202) );
  NAND2_X1 U14712 ( .A1(n13991), .A2(n12202), .ZN(n14064) );
  OAI22_X1 U14713 ( .A1(n12204), .A2(n12274), .B1(n12203), .B2(n10622), .ZN(
        n12208) );
  NAND2_X1 U14714 ( .A1(n14570), .A2(n12262), .ZN(n12206) );
  NAND2_X1 U14715 ( .A1(n14139), .A2(n12267), .ZN(n12205) );
  NAND2_X1 U14716 ( .A1(n12206), .A2(n12205), .ZN(n12207) );
  XNOR2_X1 U14717 ( .A(n12207), .B(n12265), .ZN(n12209) );
  XOR2_X1 U14718 ( .A(n12208), .B(n12209), .Z(n14063) );
  NAND2_X1 U14719 ( .A1(n12209), .A2(n12208), .ZN(n12210) );
  OAI22_X1 U14720 ( .A1(n14446), .A2(n12275), .B1(n14066), .B2(n12274), .ZN(
        n12211) );
  XOR2_X1 U14721 ( .A(n12212), .B(n12211), .Z(n12214) );
  AOI22_X1 U14722 ( .A1(n14632), .A2(n12267), .B1(n12268), .B2(n14138), .ZN(
        n12213) );
  NAND2_X1 U14723 ( .A1(n12214), .A2(n12213), .ZN(n14082) );
  OAI21_X1 U14724 ( .B1(n12214), .B2(n12213), .A(n14082), .ZN(n13999) );
  NAND2_X1 U14725 ( .A1(n14628), .A2(n12262), .ZN(n12216) );
  NAND2_X1 U14726 ( .A1(n14137), .A2(n12267), .ZN(n12215) );
  NAND2_X1 U14727 ( .A1(n12216), .A2(n12215), .ZN(n12217) );
  XNOR2_X1 U14728 ( .A(n12217), .B(n6749), .ZN(n12219) );
  AND2_X1 U14729 ( .A1(n14137), .A2(n12268), .ZN(n12218) );
  AOI21_X1 U14730 ( .B1(n14628), .B2(n12267), .A(n12218), .ZN(n12220) );
  NAND2_X1 U14731 ( .A1(n12219), .A2(n12220), .ZN(n13983) );
  INV_X1 U14732 ( .A(n12219), .ZN(n12222) );
  INV_X1 U14733 ( .A(n12220), .ZN(n12221) );
  NAND2_X1 U14734 ( .A1(n12222), .A2(n12221), .ZN(n12223) );
  NAND2_X1 U14735 ( .A1(n14553), .A2(n12262), .ZN(n12225) );
  NAND2_X1 U14736 ( .A1(n12267), .A2(n14136), .ZN(n12224) );
  NAND2_X1 U14737 ( .A1(n12225), .A2(n12224), .ZN(n12226) );
  XNOR2_X1 U14738 ( .A(n12226), .B(n6749), .ZN(n12229) );
  NOR2_X1 U14739 ( .A1(n10622), .A2(n12227), .ZN(n12228) );
  AOI21_X1 U14740 ( .B1(n14553), .B2(n12267), .A(n12228), .ZN(n12230) );
  NAND2_X1 U14741 ( .A1(n12229), .A2(n12230), .ZN(n14058) );
  INV_X1 U14742 ( .A(n12229), .ZN(n12232) );
  INV_X1 U14743 ( .A(n12230), .ZN(n12231) );
  NAND2_X1 U14744 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  NAND2_X1 U14745 ( .A1(n14623), .A2(n12262), .ZN(n12235) );
  NAND2_X1 U14746 ( .A1(n12267), .A2(n14135), .ZN(n12234) );
  NAND2_X1 U14747 ( .A1(n12235), .A2(n12234), .ZN(n12236) );
  XNOR2_X1 U14748 ( .A(n12236), .B(n6749), .ZN(n12238) );
  NOR2_X1 U14749 ( .A1(n10622), .A2(n13977), .ZN(n12237) );
  AOI21_X1 U14750 ( .B1(n14623), .B2(n12267), .A(n12237), .ZN(n12239) );
  NAND2_X1 U14751 ( .A1(n12238), .A2(n12239), .ZN(n14021) );
  INV_X1 U14752 ( .A(n12238), .ZN(n12241) );
  INV_X1 U14753 ( .A(n12239), .ZN(n12240) );
  NAND2_X1 U14754 ( .A1(n12241), .A2(n12240), .ZN(n12242) );
  NAND2_X1 U14755 ( .A1(n14018), .A2(n14021), .ZN(n12253) );
  NAND2_X1 U14756 ( .A1(n14619), .A2(n12262), .ZN(n12244) );
  NAND2_X1 U14757 ( .A1(n12267), .A2(n14134), .ZN(n12243) );
  NAND2_X1 U14758 ( .A1(n12244), .A2(n12243), .ZN(n12245) );
  XNOR2_X1 U14759 ( .A(n12245), .B(n6749), .ZN(n12248) );
  NOR2_X1 U14760 ( .A1(n10622), .A2(n12246), .ZN(n12247) );
  AOI21_X1 U14761 ( .B1(n14619), .B2(n12267), .A(n12247), .ZN(n12249) );
  NAND2_X1 U14762 ( .A1(n12248), .A2(n12249), .ZN(n12254) );
  INV_X1 U14763 ( .A(n12248), .ZN(n12251) );
  INV_X1 U14764 ( .A(n12249), .ZN(n12250) );
  NAND2_X1 U14765 ( .A1(n12251), .A2(n12250), .ZN(n12252) );
  NAND2_X1 U14766 ( .A1(n12253), .A2(n14019), .ZN(n14023) );
  NAND2_X1 U14767 ( .A1(n14023), .A2(n12254), .ZN(n14106) );
  OAI22_X1 U14768 ( .A1(n14616), .A2(n12275), .B1(n13969), .B2(n12274), .ZN(
        n12255) );
  XNOR2_X1 U14769 ( .A(n12255), .B(n12265), .ZN(n12259) );
  NAND2_X1 U14770 ( .A1(n12268), .A2(n14133), .ZN(n12256) );
  NAND2_X1 U14771 ( .A1(n12257), .A2(n12256), .ZN(n12258) );
  NOR2_X1 U14772 ( .A1(n12259), .A2(n12258), .ZN(n12260) );
  AOI21_X1 U14773 ( .B1(n12259), .B2(n12258), .A(n12260), .ZN(n14107) );
  INV_X1 U14774 ( .A(n12260), .ZN(n12261) );
  NAND2_X1 U14775 ( .A1(n14351), .A2(n12262), .ZN(n12264) );
  NAND2_X1 U14776 ( .A1(n12267), .A2(n14132), .ZN(n12263) );
  NAND2_X1 U14777 ( .A1(n12264), .A2(n12263), .ZN(n12266) );
  XNOR2_X1 U14778 ( .A(n12266), .B(n12265), .ZN(n12272) );
  NAND2_X1 U14779 ( .A1(n14351), .A2(n12267), .ZN(n12270) );
  NAND2_X1 U14780 ( .A1(n12268), .A2(n14132), .ZN(n12269) );
  NAND2_X1 U14781 ( .A1(n12270), .A2(n12269), .ZN(n12271) );
  NOR2_X1 U14782 ( .A1(n12272), .A2(n12271), .ZN(n12273) );
  AOI21_X1 U14783 ( .B1(n12272), .B2(n12271), .A(n12273), .ZN(n13966) );
  OAI22_X1 U14784 ( .A1(n12467), .A2(n12275), .B1(n13968), .B2(n12274), .ZN(
        n12276) );
  XNOR2_X1 U14785 ( .A(n12276), .B(n12265), .ZN(n12278) );
  OAI22_X1 U14786 ( .A1(n12467), .A2(n12274), .B1(n13968), .B2(n10622), .ZN(
        n12277) );
  XNOR2_X1 U14787 ( .A(n12278), .B(n12277), .ZN(n12279) );
  XNOR2_X1 U14788 ( .A(n12280), .B(n12279), .ZN(n12285) );
  NOR2_X1 U14789 ( .A1(n14836), .A2(n14329), .ZN(n12283) );
  OAI22_X1 U14790 ( .A1(n14121), .A2(n12281), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15462), .ZN(n12282) );
  AOI211_X1 U14791 ( .C1(n14332), .C2(n6638), .A(n12283), .B(n12282), .ZN(
        n12284) );
  OAI21_X1 U14792 ( .B1(n12285), .B2(n14103), .A(n12284), .ZN(P1_U3220) );
  OAI22_X1 U14793 ( .A1(n13488), .A2(n15148), .B1(n12286), .B2(n13567), .ZN(
        n13822) );
  AOI22_X1 U14794 ( .A1(n13515), .A2(n13822), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12287) );
  OAI21_X1 U14795 ( .B1(n13828), .B2(n15007), .A(n12287), .ZN(n12293) );
  AOI22_X1 U14796 ( .A1(n12288), .A2(n13552), .B1(n13501), .B2(n13591), .ZN(
        n12290) );
  NOR3_X1 U14797 ( .A1(n12291), .A2(n12290), .A3(n12289), .ZN(n12292) );
  AOI211_X1 U14798 ( .C1(n13907), .C2(n15004), .A(n12293), .B(n12292), .ZN(
        n12294) );
  OAI21_X1 U14799 ( .B1(n12295), .B2(n14999), .A(n12294), .ZN(P2_U3200) );
  NAND2_X1 U14800 ( .A1(n12488), .A2(n12509), .ZN(n12298) );
  MUX2_X1 U14801 ( .A(n13969), .B(n14616), .S(n12506), .Z(n12460) );
  OAI211_X1 U14802 ( .C1(n12303), .C2(n12491), .A(n12302), .B(n12305), .ZN(
        n12310) );
  NAND2_X1 U14803 ( .A1(n12310), .A2(n12309), .ZN(n12318) );
  OR2_X1 U14804 ( .A1(n14157), .A2(n12304), .ZN(n12312) );
  MUX2_X1 U14805 ( .A(n14969), .B(n14157), .S(n12304), .Z(n12313) );
  INV_X1 U14806 ( .A(n12313), .ZN(n12314) );
  NOR2_X1 U14807 ( .A1(n12317), .A2(n12316), .ZN(n12319) );
  NAND2_X1 U14808 ( .A1(n12319), .A2(n12318), .ZN(n12320) );
  NAND3_X1 U14809 ( .A1(n12321), .A2(n12320), .A3(n12514), .ZN(n12326) );
  NAND2_X1 U14810 ( .A1(n7430), .A2(n14156), .ZN(n12324) );
  NAND2_X1 U14811 ( .A1(n12322), .A2(n12491), .ZN(n12323) );
  MUX2_X1 U14812 ( .A(n12324), .B(n12323), .S(n14975), .Z(n12325) );
  MUX2_X1 U14813 ( .A(n12327), .B(n14155), .S(n12506), .Z(n12329) );
  MUX2_X1 U14814 ( .A(n14155), .B(n12327), .S(n12506), .Z(n12328) );
  INV_X1 U14815 ( .A(n12329), .ZN(n12330) );
  MUX2_X1 U14816 ( .A(n14154), .B(n12331), .S(n7430), .Z(n12335) );
  NAND2_X1 U14817 ( .A1(n12334), .A2(n12335), .ZN(n12333) );
  MUX2_X1 U14818 ( .A(n14154), .B(n12331), .S(n12491), .Z(n12332) );
  NAND2_X1 U14819 ( .A1(n12333), .A2(n12332), .ZN(n12339) );
  INV_X1 U14820 ( .A(n12334), .ZN(n12337) );
  INV_X1 U14821 ( .A(n12335), .ZN(n12336) );
  NAND2_X1 U14822 ( .A1(n12337), .A2(n12336), .ZN(n12338) );
  NAND2_X1 U14823 ( .A1(n12339), .A2(n12338), .ZN(n12362) );
  INV_X1 U14824 ( .A(n12352), .ZN(n12345) );
  NAND2_X1 U14825 ( .A1(n12342), .A2(n14152), .ZN(n12359) );
  MUX2_X1 U14826 ( .A(n14153), .B(n12343), .S(n12506), .Z(n12350) );
  MUX2_X1 U14827 ( .A(n12344), .B(n12348), .S(n12491), .Z(n12351) );
  AOI22_X1 U14828 ( .A1(n12345), .A2(n12359), .B1(n12350), .B2(n12351), .ZN(
        n12361) );
  INV_X1 U14829 ( .A(n12351), .ZN(n12347) );
  NAND2_X1 U14830 ( .A1(n12491), .A2(n14153), .ZN(n12346) );
  OAI211_X1 U14831 ( .C1(n12348), .C2(n12491), .A(n12347), .B(n12346), .ZN(
        n12358) );
  OAI21_X1 U14832 ( .B1(n12351), .B2(n12350), .A(n12349), .ZN(n12353) );
  NAND2_X1 U14833 ( .A1(n12353), .A2(n12352), .ZN(n12357) );
  NAND2_X1 U14834 ( .A1(n12363), .A2(n14151), .ZN(n12354) );
  NAND2_X1 U14835 ( .A1(n12355), .A2(n12354), .ZN(n12356) );
  OAI211_X1 U14836 ( .C1(n12359), .C2(n12358), .A(n12357), .B(n12356), .ZN(
        n12360) );
  AOI21_X1 U14837 ( .B1(n12362), .B2(n12361), .A(n12360), .ZN(n12367) );
  AND2_X1 U14838 ( .A1(n12491), .A2(n14151), .ZN(n12365) );
  NOR2_X1 U14839 ( .A1(n12491), .A2(n14151), .ZN(n12364) );
  MUX2_X1 U14840 ( .A(n12365), .B(n12364), .S(n12363), .Z(n12366) );
  MUX2_X1 U14841 ( .A(n14150), .B(n12368), .S(n7430), .Z(n12371) );
  MUX2_X1 U14842 ( .A(n12369), .B(n14885), .S(n12491), .Z(n12370) );
  MUX2_X1 U14843 ( .A(n14149), .B(n12372), .S(n12491), .Z(n12376) );
  MUX2_X1 U14844 ( .A(n12374), .B(n12373), .S(n7430), .Z(n12375) );
  MUX2_X1 U14845 ( .A(n14148), .B(n12377), .S(n7430), .Z(n12380) );
  MUX2_X1 U14846 ( .A(n14148), .B(n12377), .S(n12491), .Z(n12378) );
  INV_X1 U14847 ( .A(n12380), .ZN(n12381) );
  MUX2_X1 U14848 ( .A(n14147), .B(n12382), .S(n12491), .Z(n12385) );
  MUX2_X1 U14849 ( .A(n14147), .B(n12382), .S(n7430), .Z(n12383) );
  INV_X1 U14850 ( .A(n12385), .ZN(n12386) );
  MUX2_X1 U14851 ( .A(n14146), .B(n12387), .S(n7430), .Z(n12401) );
  INV_X1 U14852 ( .A(n12401), .ZN(n12388) );
  INV_X1 U14853 ( .A(n12412), .ZN(n12393) );
  NOR2_X1 U14854 ( .A1(n12393), .A2(n12392), .ZN(n12394) );
  NAND2_X1 U14855 ( .A1(n12395), .A2(n12394), .ZN(n12396) );
  NAND2_X1 U14856 ( .A1(n12396), .A2(n12506), .ZN(n12399) );
  NAND2_X1 U14857 ( .A1(n12411), .A2(n12397), .ZN(n12398) );
  NAND3_X1 U14858 ( .A1(n12400), .A2(n14081), .A3(n12491), .ZN(n12403) );
  MUX2_X1 U14859 ( .A(n14143), .B(n14039), .S(n12506), .Z(n12425) );
  AND2_X1 U14860 ( .A1(n14046), .A2(n7430), .ZN(n12424) );
  AOI21_X1 U14861 ( .B1(n12425), .B2(n14142), .A(n12424), .ZN(n12410) );
  AND2_X1 U14862 ( .A1(n14142), .A2(n12491), .ZN(n12418) );
  INV_X1 U14863 ( .A(n12424), .ZN(n12404) );
  NOR2_X1 U14864 ( .A1(n12404), .A2(n14142), .ZN(n12405) );
  AOI21_X1 U14865 ( .B1(n14644), .B2(n12418), .A(n12405), .ZN(n12421) );
  NAND2_X1 U14866 ( .A1(n12425), .A2(n12406), .ZN(n12407) );
  OR2_X1 U14867 ( .A1(n14039), .A2(n7430), .ZN(n12416) );
  NAND2_X1 U14868 ( .A1(n12407), .A2(n12416), .ZN(n12408) );
  NAND2_X1 U14869 ( .A1(n12408), .A2(n14514), .ZN(n12409) );
  OAI211_X1 U14870 ( .C1(n12410), .C2(n14514), .A(n12421), .B(n12409), .ZN(
        n12414) );
  MUX2_X1 U14871 ( .A(n12412), .B(n12411), .S(n7430), .Z(n12413) );
  INV_X1 U14872 ( .A(n12416), .ZN(n12417) );
  NAND2_X1 U14873 ( .A1(n12425), .A2(n12417), .ZN(n12420) );
  INV_X1 U14874 ( .A(n12418), .ZN(n12419) );
  NAND2_X1 U14875 ( .A1(n12420), .A2(n12419), .ZN(n12423) );
  INV_X1 U14876 ( .A(n12421), .ZN(n12422) );
  AOI22_X1 U14877 ( .A1(n12423), .A2(n14514), .B1(n12425), .B2(n12422), .ZN(
        n12429) );
  NAND2_X1 U14878 ( .A1(n12425), .A2(n12424), .ZN(n12426) );
  OAI21_X1 U14879 ( .B1(n12491), .B2(n14142), .A(n12426), .ZN(n12427) );
  NAND2_X1 U14880 ( .A1(n12427), .A2(n14587), .ZN(n12428) );
  MUX2_X1 U14881 ( .A(n12430), .B(n14479), .S(n12491), .Z(n12432) );
  AND2_X1 U14882 ( .A1(n12432), .A2(n12434), .ZN(n12433) );
  MUX2_X1 U14883 ( .A(n14139), .B(n14570), .S(n12506), .Z(n12438) );
  MUX2_X1 U14884 ( .A(n14139), .B(n14570), .S(n12491), .Z(n12435) );
  INV_X1 U14885 ( .A(n12438), .ZN(n12439) );
  MUX2_X1 U14886 ( .A(n14138), .B(n14632), .S(n12491), .Z(n12442) );
  MUX2_X1 U14887 ( .A(n14138), .B(n14632), .S(n7430), .Z(n12440) );
  NAND2_X1 U14888 ( .A1(n12441), .A2(n12440), .ZN(n12443) );
  MUX2_X1 U14889 ( .A(n14137), .B(n14628), .S(n12506), .Z(n12446) );
  MUX2_X1 U14890 ( .A(n14137), .B(n14628), .S(n12491), .Z(n12444) );
  INV_X1 U14891 ( .A(n12446), .ZN(n12447) );
  MUX2_X1 U14892 ( .A(n14136), .B(n14553), .S(n12491), .Z(n12449) );
  MUX2_X1 U14893 ( .A(n14136), .B(n14553), .S(n7430), .Z(n12448) );
  INV_X1 U14894 ( .A(n12449), .ZN(n12450) );
  MUX2_X1 U14895 ( .A(n14135), .B(n14623), .S(n12506), .Z(n12454) );
  MUX2_X1 U14896 ( .A(n14135), .B(n14623), .S(n12491), .Z(n12453) );
  INV_X1 U14897 ( .A(n12454), .ZN(n12455) );
  MUX2_X1 U14898 ( .A(n14134), .B(n14619), .S(n12491), .Z(n12458) );
  MUX2_X1 U14899 ( .A(n14134), .B(n14619), .S(n12506), .Z(n12456) );
  MUX2_X1 U14900 ( .A(n14133), .B(n14358), .S(n12491), .Z(n12459) );
  MUX2_X1 U14901 ( .A(n14132), .B(n14351), .S(n12491), .Z(n12462) );
  MUX2_X1 U14902 ( .A(n14351), .B(n14132), .S(n12491), .Z(n12465) );
  INV_X1 U14903 ( .A(n12462), .ZN(n12463) );
  MUX2_X1 U14904 ( .A(n12467), .B(n13968), .S(n12491), .Z(n12470) );
  MUX2_X1 U14905 ( .A(n14131), .B(n14332), .S(n12491), .Z(n12468) );
  NAND2_X1 U14906 ( .A1(n12471), .A2(n12470), .ZN(n12473) );
  INV_X1 U14907 ( .A(n14130), .ZN(n12474) );
  AOI21_X1 U14908 ( .B1(n12474), .B2(n12506), .A(n14321), .ZN(n12477) );
  AOI21_X1 U14909 ( .B1(n14130), .B2(n12491), .A(n12475), .ZN(n12476) );
  INV_X1 U14910 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14605) );
  NAND2_X1 U14911 ( .A1(n6645), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12480) );
  NAND2_X1 U14912 ( .A1(n12478), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12479) );
  OAI211_X1 U14913 ( .C1(n12481), .C2(n14605), .A(n12480), .B(n12479), .ZN(
        n14308) );
  OAI21_X1 U14914 ( .B1(n14308), .B2(n12482), .A(n14129), .ZN(n12483) );
  INV_X1 U14915 ( .A(n12483), .ZN(n12487) );
  NAND2_X1 U14916 ( .A1(n12484), .A2(n6643), .ZN(n12486) );
  INV_X1 U14917 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12596) );
  OR2_X1 U14918 ( .A1(n12495), .A2(n12596), .ZN(n12485) );
  MUX2_X1 U14919 ( .A(n12487), .B(n14313), .S(n12506), .Z(n12493) );
  NAND2_X1 U14920 ( .A1(n12506), .A2(n14308), .ZN(n12507) );
  OAI21_X1 U14921 ( .B1(n12489), .B2(n12488), .A(n12507), .ZN(n12490) );
  AOI22_X1 U14922 ( .A1(n14313), .A2(n12491), .B1(n14129), .B2(n12490), .ZN(
        n12492) );
  INV_X1 U14923 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12494) );
  NOR2_X1 U14924 ( .A1(n12495), .A2(n12494), .ZN(n12496) );
  AOI21_X2 U14925 ( .B1(n13944), .B2(n6643), .A(n12496), .ZN(n12505) );
  XNOR2_X1 U14926 ( .A(n12505), .B(n14308), .ZN(n12512) );
  INV_X1 U14927 ( .A(n12297), .ZN(n12499) );
  NAND2_X1 U14928 ( .A1(n12499), .A2(n12498), .ZN(n12500) );
  NAND2_X1 U14929 ( .A1(n12501), .A2(n12500), .ZN(n12504) );
  OR2_X1 U14930 ( .A1(n12502), .A2(n14301), .ZN(n12503) );
  NAND2_X1 U14931 ( .A1(n12504), .A2(n12503), .ZN(n12547) );
  MUX2_X1 U14932 ( .A(n12506), .B(n14308), .S(n12505), .Z(n12508) );
  NAND2_X1 U14933 ( .A1(n12510), .A2(n12509), .ZN(n12545) );
  NAND2_X1 U14934 ( .A1(n12547), .A2(n12545), .ZN(n12548) );
  INV_X1 U14935 ( .A(n12512), .ZN(n12549) );
  INV_X1 U14936 ( .A(n14129), .ZN(n12513) );
  XNOR2_X1 U14937 ( .A(n14313), .B(n12513), .ZN(n12541) );
  INV_X1 U14938 ( .A(n14490), .ZN(n14488) );
  NAND4_X1 U14939 ( .A1(n14917), .A2(n12515), .A3(n12514), .A4(n14890), .ZN(
        n12517) );
  NOR2_X1 U14940 ( .A1(n12517), .A2(n12516), .ZN(n12519) );
  NAND3_X1 U14941 ( .A1(n12520), .A2(n12519), .A3(n12518), .ZN(n12521) );
  NOR3_X1 U14942 ( .A1(n12523), .A2(n12522), .A3(n12521), .ZN(n12525) );
  NAND4_X1 U14943 ( .A1(n12527), .A2(n12526), .A3(n12525), .A4(n12524), .ZN(
        n12528) );
  OR4_X1 U14944 ( .A1(n12531), .A2(n12530), .A3(n12529), .A4(n12528), .ZN(
        n12532) );
  OR3_X1 U14945 ( .A1(n14488), .A2(n8637), .A3(n12532), .ZN(n12534) );
  OR4_X1 U14946 ( .A1(n12534), .A2(n14502), .A3(n14456), .A4(n12533), .ZN(
        n12535) );
  OR4_X1 U14947 ( .A1(n14430), .A2(n14440), .A3(n7432), .A4(n12535), .ZN(
        n12536) );
  NOR2_X1 U14948 ( .A1(n14385), .A2(n12536), .ZN(n12538) );
  NAND4_X1 U14949 ( .A1(n14361), .A2(n12538), .A3(n12537), .A4(n14410), .ZN(
        n12539) );
  NOR4_X1 U14950 ( .A1(n12541), .A2(n14339), .A3(n12540), .A4(n12539), .ZN(
        n12543) );
  NAND3_X1 U14951 ( .A1(n12549), .A2(n12543), .A3(n12542), .ZN(n12544) );
  XNOR2_X1 U14952 ( .A(n12544), .B(n14301), .ZN(n12546) );
  NOR2_X1 U14953 ( .A1(n12546), .A2(n12545), .ZN(n12555) );
  INV_X1 U14954 ( .A(n12547), .ZN(n12553) );
  NOR2_X1 U14955 ( .A1(n12549), .A2(n12548), .ZN(n12552) );
  INV_X1 U14956 ( .A(n12550), .ZN(n12551) );
  MUX2_X1 U14957 ( .A(n12553), .B(n12552), .S(n12551), .Z(n12554) );
  NAND2_X1 U14958 ( .A1(n12556), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12557) );
  OAI21_X1 U14959 ( .B1(n12560), .B2(n12297), .A(P1_B_REG_SCAN_IN), .ZN(n12559) );
  OAI222_X1 U14960 ( .A1(n6656), .A2(n12563), .B1(P1_U3086), .B2(n12561), .C1(
        n12596), .C2(n12562), .ZN(P1_U3325) );
  INV_X1 U14961 ( .A(n12564), .ZN(n12565) );
  AOI22_X1 U14962 ( .A1(n12565), .A2(n13552), .B1(n13501), .B2(n13585), .ZN(
        n12569) );
  OAI22_X1 U14963 ( .A1(n13480), .A2(n15148), .B1(n13558), .B2(n13567), .ZN(
        n13744) );
  AOI22_X1 U14964 ( .A1(n13744), .A2(n13515), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12566) );
  OAI21_X1 U14965 ( .B1(n13750), .B2(n15007), .A(n12566), .ZN(n12567) );
  AOI21_X1 U14966 ( .B1(n13881), .B2(n15004), .A(n12567), .ZN(n12568) );
  OAI21_X1 U14967 ( .B1(n12570), .B2(n12569), .A(n12568), .ZN(P2_U3207) );
  NAND2_X1 U14968 ( .A1(n13515), .A2(n12571), .ZN(n12573) );
  OAI211_X1 U14969 ( .C1(n15007), .C2(n12574), .A(n12573), .B(n12572), .ZN(
        n12580) );
  AOI22_X1 U14970 ( .A1(n12575), .A2(n13552), .B1(n13501), .B2(n13596), .ZN(
        n12577) );
  NOR3_X1 U14971 ( .A1(n12578), .A2(n12577), .A3(n12576), .ZN(n12579) );
  AOI211_X1 U14972 ( .C1(n14815), .C2(n15004), .A(n12580), .B(n12579), .ZN(
        n12581) );
  OAI21_X1 U14973 ( .B1(n12582), .B2(n14999), .A(n12581), .ZN(P2_U3196) );
  INV_X1 U14974 ( .A(SI_28_), .ZN(n12583) );
  OAI222_X1 U14975 ( .A1(n6655), .A2(n12585), .B1(n12584), .B2(n12583), .C1(
        P3_U3151), .C2(n12806), .ZN(P3_U3267) );
  NAND2_X1 U14976 ( .A1(n12586), .A2(n12601), .ZN(n12588) );
  NAND2_X1 U14977 ( .A1(n12602), .A2(SI_30_), .ZN(n12587) );
  INV_X1 U14978 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12592) );
  NAND2_X1 U14979 ( .A1(n8131), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12591) );
  INV_X1 U14980 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12589) );
  OR2_X1 U14981 ( .A1(n7754), .A2(n12589), .ZN(n12590) );
  OAI211_X1 U14982 ( .C1(n7767), .C2(n12592), .A(n12591), .B(n12590), .ZN(
        n12593) );
  INV_X1 U14983 ( .A(n12593), .ZN(n12594) );
  INV_X1 U14984 ( .A(n13173), .ZN(n13048) );
  NOR2_X1 U14985 ( .A1(n13417), .A2(n13048), .ZN(n12606) );
  AND2_X1 U14986 ( .A1(n12596), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12597) );
  OAI22_X1 U14987 ( .A1(n12598), .A2(n12597), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n12596), .ZN(n12600) );
  XNOR2_X1 U14988 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12599) );
  XNOR2_X1 U14989 ( .A(n12600), .B(n12599), .ZN(n13461) );
  NAND2_X1 U14990 ( .A1(n13461), .A2(n12601), .ZN(n12604) );
  NAND2_X1 U14991 ( .A1(n12602), .A2(SI_31_), .ZN(n12603) );
  OR2_X1 U14992 ( .A1(n13411), .A2(n13173), .ZN(n12760) );
  NAND2_X1 U14993 ( .A1(n12609), .A2(n12608), .ZN(n12757) );
  AND2_X1 U14994 ( .A1(n12757), .A2(n12754), .ZN(n12605) );
  NAND2_X1 U14995 ( .A1(n12760), .A2(n12605), .ZN(n12762) );
  AOI211_X1 U14996 ( .C1(n12607), .C2(n12763), .A(n12606), .B(n12762), .ZN(
        n12612) );
  NOR2_X1 U14997 ( .A1(n12609), .A2(n12608), .ZN(n12758) );
  NAND2_X1 U14998 ( .A1(n12758), .A2(n13411), .ZN(n12610) );
  NAND2_X1 U14999 ( .A1(n6853), .A2(n12610), .ZN(n12611) );
  INV_X1 U15000 ( .A(n12615), .ZN(n12804) );
  AND2_X1 U15001 ( .A1(n12621), .A2(n12617), .ZN(n12620) );
  MUX2_X1 U15002 ( .A(n12620), .B(n12619), .S(n12618), .Z(n12628) );
  NAND2_X1 U15003 ( .A1(n12625), .A2(n12621), .ZN(n12622) );
  NAND2_X1 U15004 ( .A1(n12622), .A2(n8227), .ZN(n12623) );
  NAND2_X1 U15005 ( .A1(n12623), .A2(n12624), .ZN(n12627) );
  MUX2_X1 U15006 ( .A(n12625), .B(n12624), .S(n8227), .Z(n12626) );
  OAI211_X1 U15007 ( .C1(n12628), .C2(n12627), .A(n15236), .B(n12626), .ZN(
        n12632) );
  NAND2_X1 U15008 ( .A1(n8232), .A2(n12629), .ZN(n12630) );
  NAND2_X1 U15009 ( .A1(n12630), .A2(n12746), .ZN(n12631) );
  NAND2_X1 U15010 ( .A1(n12632), .A2(n12631), .ZN(n12636) );
  AOI21_X1 U15011 ( .B1(n12635), .B2(n12633), .A(n12746), .ZN(n12634) );
  AOI21_X1 U15012 ( .B1(n12636), .B2(n12635), .A(n12634), .ZN(n12641) );
  OAI21_X1 U15013 ( .B1(n12746), .B2(n8232), .A(n12771), .ZN(n12640) );
  NAND2_X1 U15014 ( .A1(n12956), .A2(n15270), .ZN(n12638) );
  MUX2_X1 U15015 ( .A(n12638), .B(n12637), .S(n12746), .Z(n12639) );
  OAI211_X1 U15016 ( .C1(n12641), .C2(n12640), .A(n12775), .B(n12639), .ZN(
        n12645) );
  NAND2_X1 U15017 ( .A1(n12651), .A2(n12642), .ZN(n12643) );
  NAND2_X1 U15018 ( .A1(n12643), .A2(n8227), .ZN(n12644) );
  NAND2_X1 U15019 ( .A1(n12645), .A2(n12644), .ZN(n12649) );
  AOI21_X1 U15020 ( .B1(n12646), .B2(n12648), .A(n8227), .ZN(n12647) );
  AOI21_X1 U15021 ( .B1(n12649), .B2(n12648), .A(n12647), .ZN(n12657) );
  OAI21_X1 U15022 ( .B1(n8227), .B2(n12651), .A(n12650), .ZN(n12656) );
  NAND2_X1 U15023 ( .A1(n12652), .A2(n15283), .ZN(n12654) );
  MUX2_X1 U15024 ( .A(n12654), .B(n12653), .S(n8227), .Z(n12655) );
  OAI211_X1 U15025 ( .C1(n12657), .C2(n12656), .A(n12770), .B(n12655), .ZN(
        n12661) );
  MUX2_X1 U15026 ( .A(n12659), .B(n12658), .S(n12746), .Z(n12660) );
  NAND3_X1 U15027 ( .A1(n12661), .A2(n12774), .A3(n12660), .ZN(n12666) );
  MUX2_X1 U15028 ( .A(n12663), .B(n12662), .S(n8227), .Z(n12664) );
  NAND3_X1 U15029 ( .A1(n12666), .A2(n12665), .A3(n12664), .ZN(n12671) );
  MUX2_X1 U15030 ( .A(n12668), .B(n12667), .S(n8227), .Z(n12670) );
  AOI21_X1 U15031 ( .B1(n12671), .B2(n12670), .A(n12669), .ZN(n12674) );
  AOI21_X1 U15032 ( .B1(n12679), .B2(n12672), .A(n8227), .ZN(n12673) );
  OR2_X1 U15033 ( .A1(n12674), .A2(n12673), .ZN(n12678) );
  AOI21_X1 U15034 ( .B1(n12677), .B2(n12675), .A(n12746), .ZN(n12676) );
  AOI21_X1 U15035 ( .B1(n12678), .B2(n12677), .A(n12676), .ZN(n12684) );
  OAI21_X1 U15036 ( .B1(n12746), .B2(n12679), .A(n12783), .ZN(n12683) );
  MUX2_X1 U15037 ( .A(n12681), .B(n12680), .S(n8227), .Z(n12682) );
  OAI21_X1 U15038 ( .B1(n12684), .B2(n12683), .A(n12682), .ZN(n12685) );
  NAND2_X1 U15039 ( .A1(n12685), .A2(n8239), .ZN(n12690) );
  MUX2_X1 U15040 ( .A(n12687), .B(n12686), .S(n12746), .Z(n12688) );
  NAND3_X1 U15041 ( .A1(n12690), .A2(n12689), .A3(n12688), .ZN(n12695) );
  NAND2_X1 U15042 ( .A1(n12698), .A2(n12691), .ZN(n12692) );
  NAND2_X1 U15043 ( .A1(n12692), .A2(n12746), .ZN(n12694) );
  INV_X1 U15044 ( .A(n12697), .ZN(n12693) );
  AOI21_X1 U15045 ( .B1(n12695), .B2(n12694), .A(n12693), .ZN(n12700) );
  AOI21_X1 U15046 ( .B1(n12697), .B2(n12696), .A(n12746), .ZN(n12699) );
  OAI22_X1 U15047 ( .A1(n12700), .A2(n12699), .B1(n12746), .B2(n12698), .ZN(
        n12707) );
  INV_X1 U15048 ( .A(n12701), .ZN(n12706) );
  INV_X1 U15049 ( .A(n12708), .ZN(n12705) );
  AND2_X1 U15050 ( .A1(n12702), .A2(n8227), .ZN(n12703) );
  OAI211_X1 U15051 ( .C1(n12705), .C2(n12704), .A(n12714), .B(n12703), .ZN(
        n12710) );
  AOI22_X1 U15052 ( .A1(n12707), .A2(n12789), .B1(n12706), .B2(n12710), .ZN(
        n12712) );
  NAND3_X1 U15053 ( .A1(n12713), .A2(n12746), .A3(n12708), .ZN(n12709) );
  NAND2_X1 U15054 ( .A1(n12710), .A2(n12709), .ZN(n12711) );
  OAI21_X1 U15055 ( .B1(n12712), .B2(n13339), .A(n12711), .ZN(n12716) );
  MUX2_X1 U15056 ( .A(n12714), .B(n12713), .S(n8227), .Z(n12715) );
  NAND3_X1 U15057 ( .A1(n12716), .A2(n8243), .A3(n12715), .ZN(n12720) );
  XNOR2_X1 U15058 ( .A(n13286), .B(n13295), .ZN(n12765) );
  NAND2_X1 U15059 ( .A1(n13308), .A2(n13313), .ZN(n12717) );
  MUX2_X1 U15060 ( .A(n12718), .B(n12717), .S(n12746), .Z(n12719) );
  NAND3_X1 U15061 ( .A1(n12720), .A2(n12765), .A3(n12719), .ZN(n12724) );
  MUX2_X1 U15062 ( .A(n12722), .B(n12721), .S(n12746), .Z(n12723) );
  NAND3_X1 U15063 ( .A1(n12724), .A2(n12764), .A3(n12723), .ZN(n12728) );
  MUX2_X1 U15064 ( .A(n12726), .B(n12725), .S(n8227), .Z(n12727) );
  NAND3_X1 U15065 ( .A1(n12728), .A2(n13263), .A3(n12727), .ZN(n12732) );
  MUX2_X1 U15066 ( .A(n12730), .B(n12729), .S(n8227), .Z(n12731) );
  AOI21_X1 U15067 ( .B1(n12732), .B2(n12731), .A(n13247), .ZN(n12740) );
  OR2_X1 U15068 ( .A1(n13372), .A2(n13256), .ZN(n12734) );
  MUX2_X1 U15069 ( .A(n12734), .B(n12733), .S(n8227), .Z(n12735) );
  NAND2_X1 U15070 ( .A1(n12792), .A2(n12735), .ZN(n12739) );
  MUX2_X1 U15071 ( .A(n12737), .B(n12736), .S(n8227), .Z(n12738) );
  NAND2_X1 U15072 ( .A1(n13361), .A2(n13197), .ZN(n12741) );
  NAND2_X1 U15073 ( .A1(n12742), .A2(n12741), .ZN(n12744) );
  OR2_X1 U15074 ( .A1(n13358), .A2(n12900), .ZN(n12743) );
  NAND2_X1 U15075 ( .A1(n12744), .A2(n12743), .ZN(n12747) );
  NAND2_X1 U15076 ( .A1(n12747), .A2(n12746), .ZN(n12745) );
  OR2_X1 U15077 ( .A1(n12747), .A2(n12746), .ZN(n12748) );
  INV_X1 U15078 ( .A(n12749), .ZN(n12753) );
  MUX2_X1 U15079 ( .A(n12751), .B(n12750), .S(n8227), .Z(n12752) );
  NAND2_X1 U15080 ( .A1(n12755), .A2(n12754), .ZN(n12756) );
  INV_X1 U15081 ( .A(n12757), .ZN(n12759) );
  INV_X1 U15082 ( .A(n12758), .ZN(n12797) );
  INV_X1 U15083 ( .A(n12762), .ZN(n12799) );
  INV_X1 U15084 ( .A(n12763), .ZN(n12796) );
  INV_X1 U15085 ( .A(n12765), .ZN(n13282) );
  NOR2_X1 U15086 ( .A1(n12767), .A2(n12766), .ZN(n12768) );
  NAND4_X1 U15087 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n12768), .ZN(
        n12779) );
  INV_X1 U15088 ( .A(n12772), .ZN(n12773) );
  NAND4_X1 U15089 ( .A1(n15236), .A2(n12775), .A3(n12774), .A4(n12773), .ZN(
        n12778) );
  NOR4_X1 U15090 ( .A1(n12779), .A2(n12778), .A3(n12777), .A4(n12776), .ZN(
        n12780) );
  NAND4_X1 U15091 ( .A1(n12783), .A2(n12782), .A3(n12781), .A4(n12780), .ZN(
        n12784) );
  NOR4_X1 U15092 ( .A1(n12787), .A2(n12786), .A3(n12785), .A4(n12784), .ZN(
        n12788) );
  NAND4_X1 U15093 ( .A1(n13325), .A2(n8241), .A3(n12789), .A4(n12788), .ZN(
        n12790) );
  NOR4_X1 U15094 ( .A1(n13270), .A2(n13301), .A3(n13282), .A4(n12790), .ZN(
        n12791) );
  NAND4_X1 U15095 ( .A1(n12792), .A2(n13263), .A3(n12791), .A4(n8246), .ZN(
        n12793) );
  NOR4_X1 U15096 ( .A1(n12796), .A2(n12795), .A3(n12794), .A4(n12793), .ZN(
        n12798) );
  NAND4_X1 U15097 ( .A1(n12799), .A2(n12798), .A3(n6853), .A4(n12797), .ZN(
        n12801) );
  NOR3_X1 U15098 ( .A1(n12808), .A2(n12807), .A3(n12806), .ZN(n12811) );
  OAI21_X1 U15099 ( .B1(n12812), .B2(n12809), .A(P3_B_REG_SCAN_IN), .ZN(n12810) );
  OAI22_X1 U15100 ( .A1(n12813), .A2(n12812), .B1(n12811), .B2(n12810), .ZN(
        P3_U3296) );
  OAI211_X1 U15101 ( .C1(n12816), .C2(n12815), .A(n12814), .B(n12995), .ZN(
        n12823) );
  AOI21_X1 U15102 ( .B1(n13037), .B2(n13057), .A(n12817), .ZN(n12822) );
  AOI22_X1 U15103 ( .A1(n13044), .A2(n12818), .B1(n13017), .B2(n13058), .ZN(
        n12821) );
  NAND2_X1 U15104 ( .A1(n13038), .A2(n12819), .ZN(n12820) );
  NAND4_X1 U15105 ( .A1(n12823), .A2(n12822), .A3(n12821), .A4(n12820), .ZN(
        P3_U3153) );
  XNOR2_X1 U15106 ( .A(n13358), .B(n12856), .ZN(n12899) );
  XNOR2_X1 U15107 ( .A(n12899), .B(n13216), .ZN(n12901) );
  NAND2_X1 U15108 ( .A1(n12825), .A2(n12824), .ZN(n12826) );
  XNOR2_X1 U15109 ( .A(n12949), .B(n12856), .ZN(n12941) );
  AND2_X1 U15110 ( .A1(n12941), .A2(n12940), .ZN(n12828) );
  INV_X1 U15111 ( .A(n12941), .ZN(n12829) );
  NAND2_X1 U15112 ( .A1(n12829), .A2(n13052), .ZN(n12830) );
  XNOR2_X1 U15113 ( .A(n12968), .B(n12856), .ZN(n12831) );
  XNOR2_X1 U15114 ( .A(n12831), .B(n13333), .ZN(n12962) );
  INV_X1 U15115 ( .A(n12831), .ZN(n12832) );
  NAND2_X1 U15116 ( .A1(n12832), .A2(n13333), .ZN(n12833) );
  NAND2_X1 U15117 ( .A1(n12834), .A2(n12833), .ZN(n13025) );
  XNOR2_X1 U15118 ( .A(n13340), .B(n12856), .ZN(n12835) );
  NAND2_X1 U15119 ( .A1(n12835), .A2(n13315), .ZN(n13023) );
  NAND2_X1 U15120 ( .A1(n13025), .A2(n13023), .ZN(n12837) );
  INV_X1 U15121 ( .A(n12835), .ZN(n12836) );
  NAND2_X1 U15122 ( .A1(n12836), .A2(n13051), .ZN(n13024) );
  NAND2_X1 U15123 ( .A1(n12837), .A2(n13024), .ZN(n12893) );
  XNOR2_X1 U15124 ( .A(n13323), .B(n12856), .ZN(n12838) );
  XNOR2_X1 U15125 ( .A(n12838), .B(n13334), .ZN(n12892) );
  INV_X1 U15126 ( .A(n12838), .ZN(n12839) );
  NAND2_X1 U15127 ( .A1(n12839), .A2(n13334), .ZN(n12840) );
  XNOR2_X1 U15128 ( .A(n13308), .B(n12856), .ZN(n12841) );
  XNOR2_X1 U15129 ( .A(n12841), .B(n13050), .ZN(n12997) );
  INV_X1 U15130 ( .A(n12841), .ZN(n12842) );
  NAND2_X1 U15131 ( .A1(n12842), .A2(n13050), .ZN(n12843) );
  XNOR2_X1 U15132 ( .A(n13286), .B(n12856), .ZN(n12844) );
  XNOR2_X1 U15133 ( .A(n12844), .B(n13274), .ZN(n12914) );
  XNOR2_X1 U15134 ( .A(n13275), .B(n12849), .ZN(n12845) );
  INV_X1 U15135 ( .A(n12845), .ZN(n12846) );
  AND2_X1 U15136 ( .A1(n12847), .A2(n12846), .ZN(n12848) );
  XNOR2_X1 U15137 ( .A(n13372), .B(n12856), .ZN(n12974) );
  XNOR2_X1 U15138 ( .A(n13375), .B(n12849), .ZN(n12971) );
  INV_X1 U15139 ( .A(n12971), .ZN(n12850) );
  OAI22_X1 U15140 ( .A1(n12974), .A2(n13256), .B1(n13273), .B2(n12850), .ZN(
        n12854) );
  OAI21_X1 U15141 ( .B1(n12971), .B2(n13249), .A(n13232), .ZN(n12852) );
  NOR2_X1 U15142 ( .A1(n13232), .A2(n13249), .ZN(n12851) );
  AOI22_X1 U15143 ( .A1(n12974), .A2(n12852), .B1(n12851), .B2(n12850), .ZN(
        n12853) );
  XNOR2_X1 U15144 ( .A(n13368), .B(n12856), .ZN(n12855) );
  XNOR2_X1 U15145 ( .A(n12855), .B(n13250), .ZN(n12934) );
  XNOR2_X1 U15146 ( .A(n13361), .B(n12856), .ZN(n12857) );
  XNOR2_X1 U15147 ( .A(n12857), .B(n13197), .ZN(n13036) );
  INV_X1 U15148 ( .A(n12857), .ZN(n12858) );
  XOR2_X1 U15149 ( .A(n12901), .B(n12902), .Z(n12863) );
  AOI22_X1 U15150 ( .A1(n13233), .A2(n13017), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12860) );
  NAND2_X1 U15151 ( .A1(n13207), .A2(n13038), .ZN(n12859) );
  OAI211_X1 U15152 ( .C1(n13198), .C2(n13028), .A(n12860), .B(n12859), .ZN(
        n12861) );
  AOI21_X1 U15153 ( .B1(n13358), .B2(n13044), .A(n12861), .ZN(n12862) );
  OAI21_X1 U15154 ( .B1(n12863), .B2(n13046), .A(n12862), .ZN(P3_U3154) );
  XNOR2_X1 U15155 ( .A(n12973), .B(n13273), .ZN(n12868) );
  AOI22_X1 U15156 ( .A1(n13232), .A2(n13037), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12865) );
  NAND2_X1 U15157 ( .A1(n13038), .A2(n13260), .ZN(n12864) );
  OAI211_X1 U15158 ( .C1(n13285), .C2(n13041), .A(n12865), .B(n12864), .ZN(
        n12866) );
  AOI21_X1 U15159 ( .B1(n13375), .B2(n13044), .A(n12866), .ZN(n12867) );
  OAI21_X1 U15160 ( .B1(n12868), .B2(n13046), .A(n12867), .ZN(P3_U3156) );
  OAI211_X1 U15161 ( .C1(n12871), .C2(n12870), .A(n12869), .B(n12995), .ZN(
        n12879) );
  OAI21_X1 U15162 ( .B1(n13028), .B2(n13012), .A(n12872), .ZN(n12873) );
  INV_X1 U15163 ( .A(n12873), .ZN(n12878) );
  AOI22_X1 U15164 ( .A1(n13044), .A2(n15301), .B1(n13017), .B2(n12874), .ZN(
        n12877) );
  NAND2_X1 U15165 ( .A1(n13038), .A2(n12875), .ZN(n12876) );
  NAND4_X1 U15166 ( .A1(n12879), .A2(n12878), .A3(n12877), .A4(n12876), .ZN(
        P3_U3157) );
  AOI21_X1 U15167 ( .B1(n12881), .B2(n12880), .A(n13046), .ZN(n12883) );
  NAND2_X1 U15168 ( .A1(n12883), .A2(n12882), .ZN(n12890) );
  AOI21_X1 U15169 ( .B1(n13037), .B2(n12956), .A(n12884), .ZN(n12889) );
  AOI22_X1 U15170 ( .A1(n13044), .A2(n12885), .B1(n13017), .B2(n10809), .ZN(
        n12888) );
  NAND2_X1 U15171 ( .A1(n13038), .A2(n12886), .ZN(n12887) );
  NAND4_X1 U15172 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n12887), .ZN(
        P3_U3158) );
  INV_X1 U15173 ( .A(n13323), .ZN(n13444) );
  OAI211_X1 U15174 ( .C1(n12893), .C2(n12892), .A(n12891), .B(n12995), .ZN(
        n12898) );
  OAI21_X1 U15175 ( .B1(n13028), .B2(n13313), .A(n12894), .ZN(n12896) );
  NOR2_X1 U15176 ( .A1(n13031), .A2(n13319), .ZN(n12895) );
  AOI211_X1 U15177 ( .C1(n13017), .C2(n13051), .A(n12896), .B(n12895), .ZN(
        n12897) );
  OAI211_X1 U15178 ( .C1(n13444), .C2(n13003), .A(n12898), .B(n12897), .ZN(
        P3_U3159) );
  AOI22_X1 U15179 ( .A1(n12902), .A2(n12901), .B1(n12900), .B2(n12899), .ZN(
        n12906) );
  XNOR2_X1 U15180 ( .A(n12904), .B(n12903), .ZN(n12905) );
  XNOR2_X1 U15181 ( .A(n12906), .B(n12905), .ZN(n12912) );
  AOI22_X1 U15182 ( .A1(n13216), .A2(n13017), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12908) );
  NAND2_X1 U15183 ( .A1(n13185), .A2(n13038), .ZN(n12907) );
  OAI211_X1 U15184 ( .C1(n12909), .C2(n13028), .A(n12908), .B(n12907), .ZN(
        n12910) );
  AOI21_X1 U15185 ( .B1(n13353), .B2(n13044), .A(n12910), .ZN(n12911) );
  OAI21_X1 U15186 ( .B1(n12912), .B2(n13046), .A(n12911), .ZN(P3_U3160) );
  AOI21_X1 U15187 ( .B1(n12914), .B2(n12913), .A(n6781), .ZN(n12919) );
  NAND2_X1 U15188 ( .A1(n13038), .A2(n13287), .ZN(n12916) );
  AOI22_X1 U15189 ( .A1(n13017), .A2(n13050), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12915) );
  OAI211_X1 U15190 ( .C1(n13285), .C2(n13028), .A(n12916), .B(n12915), .ZN(
        n12917) );
  AOI21_X1 U15191 ( .B1(n13286), .B2(n13044), .A(n12917), .ZN(n12918) );
  OAI21_X1 U15192 ( .B1(n12919), .B2(n13046), .A(n12918), .ZN(P3_U3163) );
  XNOR2_X1 U15193 ( .A(n12921), .B(n12922), .ZN(n13011) );
  NOR2_X1 U15194 ( .A1(n13011), .A2(n13012), .ZN(n13010) );
  AOI21_X1 U15195 ( .B1(n12922), .B2(n12921), .A(n13010), .ZN(n12925) );
  XNOR2_X1 U15196 ( .A(n12923), .B(n13015), .ZN(n12924) );
  XNOR2_X1 U15197 ( .A(n12925), .B(n12924), .ZN(n12926) );
  NAND2_X1 U15198 ( .A1(n12926), .A2(n12995), .ZN(n12932) );
  AOI21_X1 U15199 ( .B1(n13037), .B2(n13055), .A(n12927), .ZN(n12931) );
  AOI22_X1 U15200 ( .A1(n13044), .A2(n14794), .B1(n13017), .B2(n13056), .ZN(
        n12930) );
  NAND2_X1 U15201 ( .A1(n13038), .A2(n12928), .ZN(n12929) );
  NAND4_X1 U15202 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        P3_U3164) );
  XOR2_X1 U15203 ( .A(n12934), .B(n12933), .Z(n12939) );
  AOI22_X1 U15204 ( .A1(n13233), .A2(n13037), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12936) );
  NAND2_X1 U15205 ( .A1(n13038), .A2(n13236), .ZN(n12935) );
  OAI211_X1 U15206 ( .C1(n13256), .C2(n13041), .A(n12936), .B(n12935), .ZN(
        n12937) );
  AOI21_X1 U15207 ( .B1(n13368), .B2(n13044), .A(n12937), .ZN(n12938) );
  OAI21_X1 U15208 ( .B1(n12939), .B2(n13046), .A(n12938), .ZN(P3_U3165) );
  XNOR2_X1 U15209 ( .A(n12941), .B(n12940), .ZN(n12942) );
  XNOR2_X1 U15210 ( .A(n12943), .B(n12942), .ZN(n12951) );
  NAND2_X1 U15211 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13123)
         );
  OAI21_X1 U15212 ( .B1(n13028), .B2(n12944), .A(n13123), .ZN(n12945) );
  AOI21_X1 U15213 ( .B1(n13017), .B2(n13053), .A(n12945), .ZN(n12946) );
  OAI21_X1 U15214 ( .B1(n12947), .B2(n13031), .A(n12946), .ZN(n12948) );
  AOI21_X1 U15215 ( .B1(n12949), .B2(n13044), .A(n12948), .ZN(n12950) );
  OAI21_X1 U15216 ( .B1(n12951), .B2(n13046), .A(n12950), .ZN(P3_U3166) );
  XNOR2_X1 U15217 ( .A(n12953), .B(n12952), .ZN(n12954) );
  NAND2_X1 U15218 ( .A1(n12954), .A2(n12995), .ZN(n12961) );
  AOI21_X1 U15219 ( .B1(n13037), .B2(n13058), .A(n12955), .ZN(n12960) );
  AOI22_X1 U15220 ( .A1(n13044), .A2(n15274), .B1(n13017), .B2(n12956), .ZN(
        n12959) );
  NAND2_X1 U15221 ( .A1(n13038), .A2(n12957), .ZN(n12958) );
  NAND4_X1 U15222 ( .A1(n12961), .A2(n12960), .A3(n12959), .A4(n12958), .ZN(
        P3_U3167) );
  XNOR2_X1 U15223 ( .A(n12963), .B(n12962), .ZN(n12970) );
  INV_X1 U15224 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15548) );
  NOR2_X1 U15225 ( .A1(n15548), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13140) );
  NOR2_X1 U15226 ( .A1(n13028), .A2(n13315), .ZN(n12964) );
  AOI211_X1 U15227 ( .C1(n13017), .C2(n13052), .A(n13140), .B(n12964), .ZN(
        n12965) );
  OAI21_X1 U15228 ( .B1(n12966), .B2(n13031), .A(n12965), .ZN(n12967) );
  AOI21_X1 U15229 ( .B1(n12968), .B2(n13044), .A(n12967), .ZN(n12969) );
  OAI21_X1 U15230 ( .B1(n12970), .B2(n13046), .A(n12969), .ZN(P3_U3168) );
  OAI22_X1 U15231 ( .A1(n12973), .A2(n13249), .B1(n12972), .B2(n12971), .ZN(
        n12976) );
  XNOR2_X1 U15232 ( .A(n12974), .B(n13256), .ZN(n12975) );
  XNOR2_X1 U15233 ( .A(n12976), .B(n12975), .ZN(n12981) );
  AOI22_X1 U15234 ( .A1(n13250), .A2(n13037), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12978) );
  NAND2_X1 U15235 ( .A1(n13038), .A2(n13242), .ZN(n12977) );
  OAI211_X1 U15236 ( .C1(n13273), .C2(n13041), .A(n12978), .B(n12977), .ZN(
        n12979) );
  AOI21_X1 U15237 ( .B1(n13372), .B2(n13044), .A(n12979), .ZN(n12980) );
  OAI21_X1 U15238 ( .B1(n12981), .B2(n13046), .A(n12980), .ZN(P3_U3169) );
  INV_X1 U15239 ( .A(n12982), .ZN(n12983) );
  AOI21_X1 U15240 ( .B1(n12985), .B2(n12984), .A(n12983), .ZN(n12986) );
  OR2_X1 U15241 ( .A1(n12986), .A2(n13046), .ZN(n12994) );
  AOI21_X1 U15242 ( .B1(n13037), .B2(n13016), .A(n12987), .ZN(n12993) );
  AOI22_X1 U15243 ( .A1(n13044), .A2(n12988), .B1(n13017), .B2(n13057), .ZN(
        n12992) );
  INV_X1 U15244 ( .A(n12989), .ZN(n12990) );
  NAND2_X1 U15245 ( .A1(n13038), .A2(n12990), .ZN(n12991) );
  NAND4_X1 U15246 ( .A1(n12994), .A2(n12993), .A3(n12992), .A4(n12991), .ZN(
        P3_U3171) );
  INV_X1 U15247 ( .A(n13308), .ZN(n13440) );
  OAI211_X1 U15248 ( .C1(n12998), .C2(n12997), .A(n12996), .B(n12995), .ZN(
        n13002) );
  AOI22_X1 U15249 ( .A1(n13037), .A2(n13295), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12999) );
  OAI21_X1 U15250 ( .B1(n13027), .B2(n13041), .A(n12999), .ZN(n13000) );
  AOI21_X1 U15251 ( .B1(n13298), .B2(n13038), .A(n13000), .ZN(n13001) );
  OAI211_X1 U15252 ( .C1(n13440), .C2(n13003), .A(n13002), .B(n13001), .ZN(
        P3_U3173) );
  XNOR2_X1 U15253 ( .A(n13004), .B(n13049), .ZN(n13009) );
  NAND2_X1 U15254 ( .A1(n13038), .A2(n13276), .ZN(n13006) );
  AOI22_X1 U15255 ( .A1(n13017), .A2(n13295), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13005) );
  OAI211_X1 U15256 ( .C1(n13273), .C2(n13028), .A(n13006), .B(n13005), .ZN(
        n13007) );
  AOI21_X1 U15257 ( .B1(n13275), .B2(n13044), .A(n13007), .ZN(n13008) );
  OAI21_X1 U15258 ( .B1(n13009), .B2(n13046), .A(n13008), .ZN(P3_U3175) );
  AOI211_X1 U15259 ( .C1(n13012), .C2(n13011), .A(n13046), .B(n13010), .ZN(
        n13013) );
  INV_X1 U15260 ( .A(n13013), .ZN(n13022) );
  AOI21_X1 U15261 ( .B1(n13037), .B2(n13015), .A(n13014), .ZN(n13021) );
  AOI22_X1 U15262 ( .A1(n13044), .A2(n14799), .B1(n13017), .B2(n13016), .ZN(
        n13020) );
  NAND2_X1 U15263 ( .A1(n13038), .A2(n13018), .ZN(n13019) );
  NAND4_X1 U15264 ( .A1(n13022), .A2(n13021), .A3(n13020), .A4(n13019), .ZN(
        P3_U3176) );
  NAND2_X1 U15265 ( .A1(n13024), .A2(n13023), .ZN(n13026) );
  XOR2_X1 U15266 ( .A(n13026), .B(n13025), .Z(n13034) );
  NAND2_X1 U15267 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13164)
         );
  OAI21_X1 U15268 ( .B1(n13028), .B2(n13027), .A(n13164), .ZN(n13029) );
  AOI21_X1 U15269 ( .B1(n13017), .B2(n13333), .A(n13029), .ZN(n13030) );
  OAI21_X1 U15270 ( .B1(n13342), .B2(n13031), .A(n13030), .ZN(n13032) );
  AOI21_X1 U15271 ( .B1(n13340), .B2(n13044), .A(n13032), .ZN(n13033) );
  OAI21_X1 U15272 ( .B1(n13034), .B2(n13046), .A(n13033), .ZN(P3_U3178) );
  XOR2_X1 U15273 ( .A(n13036), .B(n13035), .Z(n13047) );
  AOI22_X1 U15274 ( .A1(n13216), .A2(n13037), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13040) );
  NAND2_X1 U15275 ( .A1(n13222), .A2(n13038), .ZN(n13039) );
  OAI211_X1 U15276 ( .C1(n13042), .C2(n13041), .A(n13040), .B(n13039), .ZN(
        n13043) );
  AOI21_X1 U15277 ( .B1(n13361), .B2(n13044), .A(n13043), .ZN(n13045) );
  OAI21_X1 U15278 ( .B1(n13047), .B2(n13046), .A(n13045), .ZN(P3_U3180) );
  MUX2_X1 U15279 ( .A(n13048), .B(P3_DATAO_REG_31__SCAN_IN), .S(n13060), .Z(
        P3_U3522) );
  MUX2_X1 U15280 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13216), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15281 ( .A(n13233), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13060), .Z(
        P3_U3517) );
  MUX2_X1 U15282 ( .A(n13232), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13060), .Z(
        P3_U3515) );
  MUX2_X1 U15283 ( .A(n13249), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13060), .Z(
        P3_U3514) );
  MUX2_X1 U15284 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13049), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15285 ( .A(n13295), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13060), .Z(
        P3_U3512) );
  MUX2_X1 U15286 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13050), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15287 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13334), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15288 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13051), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15289 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13333), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15290 ( .A(n13052), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13060), .Z(
        P3_U3507) );
  MUX2_X1 U15291 ( .A(n13053), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13060), .Z(
        P3_U3506) );
  MUX2_X1 U15292 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13054), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15293 ( .A(n13055), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13060), .Z(
        P3_U3504) );
  MUX2_X1 U15294 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13056), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15295 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13057), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15296 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13058), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15297 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13059), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15298 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15243), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15299 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n10809), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15300 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n10244), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15301 ( .A(n13061), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13060), .Z(
        P3_U3491) );
  AOI21_X1 U15302 ( .B1(n7929), .B2(n13063), .A(n13062), .ZN(n13078) );
  INV_X1 U15303 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15460) );
  OAI21_X1 U15304 ( .B1(n13125), .B2(n15460), .A(n13064), .ZN(n13071) );
  INV_X1 U15305 ( .A(n13087), .ZN(n13069) );
  OAI21_X1 U15306 ( .B1(n13067), .B2(n13066), .A(n13065), .ZN(n13068) );
  AOI21_X1 U15307 ( .B1(n13069), .B2(n13068), .A(n13170), .ZN(n13070) );
  AOI211_X1 U15308 ( .C1(n13166), .C2(n13072), .A(n13071), .B(n13070), .ZN(
        n13077) );
  AOI21_X1 U15309 ( .B1(n15669), .B2(n13074), .A(n13073), .ZN(n13075) );
  OR2_X1 U15310 ( .A1(n13075), .A2(n13165), .ZN(n13076) );
  OAI211_X1 U15311 ( .C1(n13078), .C2(n13150), .A(n13077), .B(n13076), .ZN(
        P3_U3195) );
  AOI21_X1 U15312 ( .B1(n13081), .B2(n13080), .A(n13079), .ZN(n13096) );
  XNOR2_X1 U15313 ( .A(n6856), .B(n13082), .ZN(n13094) );
  INV_X1 U15314 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14739) );
  NAND2_X1 U15315 ( .A1(n13166), .A2(n13083), .ZN(n13085) );
  OAI211_X1 U15316 ( .C1(n14739), .C2(n13125), .A(n13085), .B(n13084), .ZN(
        n13092) );
  OR2_X1 U15317 ( .A1(n13087), .A2(n13086), .ZN(n13089) );
  AOI211_X1 U15318 ( .C1(n13090), .C2(n13089), .A(n13170), .B(n13088), .ZN(
        n13091) );
  AOI211_X1 U15319 ( .C1(n13094), .C2(n13093), .A(n13092), .B(n13091), .ZN(
        n13095) );
  OAI21_X1 U15320 ( .B1(n13096), .B2(n13150), .A(n13095), .ZN(P3_U3196) );
  AOI21_X1 U15321 ( .B1(n13099), .B2(n13098), .A(n13097), .ZN(n13114) );
  INV_X1 U15322 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14743) );
  OAI21_X1 U15323 ( .B1(n13125), .B2(n14743), .A(n13100), .ZN(n13106) );
  AOI21_X1 U15324 ( .B1(n13103), .B2(n13102), .A(n13101), .ZN(n13104) );
  NOR2_X1 U15325 ( .A1(n13104), .A2(n13170), .ZN(n13105) );
  AOI211_X1 U15326 ( .C1(n13166), .C2(n13107), .A(n13106), .B(n13105), .ZN(
        n13113) );
  AOI21_X1 U15327 ( .B1(n13110), .B2(n13109), .A(n13108), .ZN(n13111) );
  OR2_X1 U15328 ( .A1(n13111), .A2(n13165), .ZN(n13112) );
  OAI211_X1 U15329 ( .C1(n13114), .C2(n13150), .A(n13113), .B(n13112), .ZN(
        P3_U3197) );
  AOI21_X1 U15330 ( .B1(n6777), .B2(n13116), .A(n13115), .ZN(n13134) );
  INV_X1 U15331 ( .A(n13117), .ZN(n13119) );
  NAND2_X1 U15332 ( .A1(n13119), .A2(n13118), .ZN(n13120) );
  XNOR2_X1 U15333 ( .A(n13121), .B(n13120), .ZN(n13131) );
  INV_X1 U15334 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14750) );
  NAND2_X1 U15335 ( .A1(n13166), .A2(n13122), .ZN(n13124) );
  OAI211_X1 U15336 ( .C1(n14750), .C2(n13125), .A(n13124), .B(n13123), .ZN(
        n13130) );
  AOI21_X1 U15337 ( .B1(n6849), .B2(n13127), .A(n13126), .ZN(n13128) );
  NOR2_X1 U15338 ( .A1(n13128), .A2(n13165), .ZN(n13129) );
  AOI211_X1 U15339 ( .C1(n13132), .C2(n13131), .A(n13130), .B(n13129), .ZN(
        n13133) );
  OAI21_X1 U15340 ( .B1(n13134), .B2(n13150), .A(n13133), .ZN(P3_U3198) );
  AOI21_X1 U15341 ( .B1(n13137), .B2(n13136), .A(n13135), .ZN(n13151) );
  AOI21_X1 U15342 ( .B1(n13139), .B2(n13404), .A(n13138), .ZN(n13142) );
  AOI21_X1 U15343 ( .B1(n15234), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13140), 
        .ZN(n13141) );
  OAI21_X1 U15344 ( .B1(n13142), .B2(n13165), .A(n13141), .ZN(n13147) );
  AOI211_X1 U15345 ( .C1(n13145), .C2(n13144), .A(n13170), .B(n13143), .ZN(
        n13146) );
  AOI211_X1 U15346 ( .C1(n13166), .C2(n13148), .A(n13147), .B(n13146), .ZN(
        n13149) );
  OAI21_X1 U15347 ( .B1(n13151), .B2(n13150), .A(n13149), .ZN(P3_U3199) );
  AOI21_X1 U15348 ( .B1(n13154), .B2(n13153), .A(n13152), .ZN(n13171) );
  AND3_X1 U15349 ( .A1(n13157), .A2(n13156), .A3(n13155), .ZN(n13159) );
  OAI21_X1 U15350 ( .B1(n13160), .B2(n13159), .A(n13158), .ZN(n13169) );
  NAND2_X1 U15351 ( .A1(n15234), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13163) );
  OAI211_X1 U15352 ( .C1(n13171), .C2(n13170), .A(n13169), .B(n13168), .ZN(
        P3_U3200) );
  INV_X1 U15353 ( .A(n13411), .ZN(n13350) );
  INV_X1 U15354 ( .A(n13174), .ZN(n13175) );
  NAND2_X1 U15355 ( .A1(n13175), .A2(n13288), .ZN(n13180) );
  OAI21_X1 U15356 ( .B1(n15258), .B2(n13412), .A(n13180), .ZN(n13177) );
  AOI21_X1 U15357 ( .B1(n15258), .B2(P3_REG2_REG_31__SCAN_IN), .A(n13177), 
        .ZN(n13176) );
  OAI21_X1 U15358 ( .B1(n13350), .B2(n13341), .A(n13176), .ZN(P3_U3202) );
  AOI21_X1 U15359 ( .B1(n15258), .B2(P3_REG2_REG_30__SCAN_IN), .A(n13177), 
        .ZN(n13178) );
  OAI21_X1 U15360 ( .B1(n13417), .B2(n13341), .A(n13178), .ZN(P3_U3203) );
  NAND2_X1 U15361 ( .A1(n15258), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n13179) );
  OAI211_X1 U15362 ( .C1(n13181), .C2(n13341), .A(n13180), .B(n13179), .ZN(
        n13182) );
  OAI21_X1 U15363 ( .B1(n7657), .B2(n13305), .A(n13184), .ZN(P3_U3204) );
  INV_X1 U15364 ( .A(n13185), .ZN(n13187) );
  INV_X1 U15365 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n13186) );
  OAI22_X1 U15366 ( .A1(n13187), .A2(n15238), .B1(n13344), .B2(n13186), .ZN(
        n13188) );
  AOI21_X1 U15367 ( .B1(n13353), .B2(n13322), .A(n13188), .ZN(n13191) );
  NAND2_X1 U15368 ( .A1(n13189), .A2(n13347), .ZN(n13190) );
  OAI211_X1 U15369 ( .C1(n13192), .C2(n13328), .A(n13191), .B(n13190), .ZN(
        P3_U3205) );
  NAND2_X1 U15370 ( .A1(n13194), .A2(n13195), .ZN(n13196) );
  NAND2_X1 U15371 ( .A1(n13193), .A2(n13196), .ZN(n13200) );
  OAI22_X1 U15372 ( .A1(n13198), .A2(n13312), .B1(n13197), .B2(n13314), .ZN(
        n13199) );
  AOI21_X1 U15373 ( .B1(n13200), .B2(n15248), .A(n13199), .ZN(n13206) );
  NAND2_X1 U15374 ( .A1(n13202), .A2(n13201), .ZN(n13203) );
  NAND2_X1 U15375 ( .A1(n6798), .A2(n13203), .ZN(n13355) );
  NAND2_X1 U15376 ( .A1(n13355), .A2(n13204), .ZN(n13205) );
  INV_X1 U15377 ( .A(n13358), .ZN(n13421) );
  AOI22_X1 U15378 ( .A1(n13207), .A2(n13288), .B1(n15258), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13208) );
  OAI21_X1 U15379 ( .B1(n13421), .B2(n13341), .A(n13208), .ZN(n13209) );
  AOI21_X1 U15380 ( .B1(n13355), .B2(n13210), .A(n13209), .ZN(n13211) );
  OAI21_X1 U15381 ( .B1(n13357), .B2(n15258), .A(n13211), .ZN(P3_U3206) );
  NAND2_X1 U15382 ( .A1(n13213), .A2(n13212), .ZN(n13214) );
  NAND2_X1 U15383 ( .A1(n13215), .A2(n13214), .ZN(n13362) );
  AOI22_X1 U15384 ( .A1(n13216), .A2(n15242), .B1(n13250), .B2(n15244), .ZN(
        n13221) );
  XNOR2_X1 U15385 ( .A(n13218), .B(n13217), .ZN(n13219) );
  NAND2_X1 U15386 ( .A1(n13219), .A2(n15248), .ZN(n13220) );
  OAI211_X1 U15387 ( .C1(n13362), .C2(n15252), .A(n13221), .B(n13220), .ZN(
        n13363) );
  AOI22_X1 U15388 ( .A1(n13328), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n13222), 
        .B2(n13288), .ZN(n13224) );
  NAND2_X1 U15389 ( .A1(n13361), .A2(n13322), .ZN(n13223) );
  OAI211_X1 U15390 ( .C1(n13362), .C2(n13225), .A(n13224), .B(n13223), .ZN(
        n13226) );
  AOI21_X1 U15391 ( .B1(n13363), .B2(n13344), .A(n13226), .ZN(n13227) );
  INV_X1 U15392 ( .A(n13227), .ZN(P3_U3207) );
  XNOR2_X1 U15393 ( .A(n13228), .B(n13230), .ZN(n13370) );
  OAI211_X1 U15394 ( .C1(n13231), .C2(n13230), .A(n13229), .B(n15248), .ZN(
        n13235) );
  AOI22_X1 U15395 ( .A1(n13233), .A2(n15242), .B1(n15244), .B2(n13232), .ZN(
        n13234) );
  NAND2_X1 U15396 ( .A1(n13235), .A2(n13234), .ZN(n13367) );
  INV_X1 U15397 ( .A(n13368), .ZN(n13238) );
  AOI22_X1 U15398 ( .A1(n13328), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n13288), 
        .B2(n13236), .ZN(n13237) );
  OAI21_X1 U15399 ( .B1(n13238), .B2(n13341), .A(n13237), .ZN(n13239) );
  AOI21_X1 U15400 ( .B1(n13367), .B2(n13344), .A(n13239), .ZN(n13240) );
  OAI21_X1 U15401 ( .B1(n13305), .B2(n13370), .A(n13240), .ZN(P3_U3208) );
  AOI21_X1 U15402 ( .B1(n13247), .B2(n13241), .A(n6788), .ZN(n13374) );
  INV_X1 U15403 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13244) );
  INV_X1 U15404 ( .A(n13242), .ZN(n13243) );
  OAI22_X1 U15405 ( .A1(n13344), .A2(n13244), .B1(n13243), .B2(n15238), .ZN(
        n13245) );
  AOI21_X1 U15406 ( .B1(n13372), .B2(n13322), .A(n13245), .ZN(n13254) );
  OAI211_X1 U15407 ( .C1(n13248), .C2(n13247), .A(n13246), .B(n15248), .ZN(
        n13252) );
  AOI22_X1 U15408 ( .A1(n13250), .A2(n15242), .B1(n15244), .B2(n13249), .ZN(
        n13251) );
  NAND2_X1 U15409 ( .A1(n13252), .A2(n13251), .ZN(n13371) );
  NAND2_X1 U15410 ( .A1(n13371), .A2(n13344), .ZN(n13253) );
  OAI211_X1 U15411 ( .C1(n13374), .C2(n13305), .A(n13254), .B(n13253), .ZN(
        P3_U3209) );
  AOI21_X1 U15412 ( .B1(n13255), .B2(n13263), .A(n13310), .ZN(n13259) );
  OAI22_X1 U15413 ( .A1(n13256), .A2(n13312), .B1(n13285), .B2(n13314), .ZN(
        n13257) );
  AOI21_X1 U15414 ( .B1(n13259), .B2(n13258), .A(n13257), .ZN(n13377) );
  INV_X1 U15415 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n15614) );
  INV_X1 U15416 ( .A(n13260), .ZN(n13261) );
  OAI22_X1 U15417 ( .A1(n13344), .A2(n15614), .B1(n13261), .B2(n15238), .ZN(
        n13262) );
  AOI21_X1 U15418 ( .B1(n13375), .B2(n13322), .A(n13262), .ZN(n13268) );
  OR2_X1 U15419 ( .A1(n13264), .A2(n13263), .ZN(n13265) );
  NAND2_X1 U15420 ( .A1(n13266), .A2(n13265), .ZN(n13378) );
  OR2_X1 U15421 ( .A1(n13378), .A2(n13305), .ZN(n13267) );
  OAI211_X1 U15422 ( .C1(n13377), .C2(n13328), .A(n13268), .B(n13267), .ZN(
        P3_U3210) );
  XNOR2_X1 U15423 ( .A(n13269), .B(n13270), .ZN(n13380) );
  INV_X1 U15424 ( .A(n13380), .ZN(n13280) );
  XNOR2_X1 U15425 ( .A(n6882), .B(n13270), .ZN(n13272) );
  OAI222_X1 U15426 ( .A1(n13314), .A2(n13274), .B1(n13312), .B2(n13273), .C1(
        n13272), .C2(n13310), .ZN(n13379) );
  INV_X1 U15427 ( .A(n13275), .ZN(n13432) );
  AOI22_X1 U15428 ( .A1(n13328), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n13288), 
        .B2(n13276), .ZN(n13277) );
  OAI21_X1 U15429 ( .B1(n13432), .B2(n13341), .A(n13277), .ZN(n13278) );
  AOI21_X1 U15430 ( .B1(n13379), .B2(n13344), .A(n13278), .ZN(n13279) );
  OAI21_X1 U15431 ( .B1(n13280), .B2(n13305), .A(n13279), .ZN(P3_U3211) );
  XNOR2_X1 U15432 ( .A(n13281), .B(n13282), .ZN(n13384) );
  INV_X1 U15433 ( .A(n13384), .ZN(n13292) );
  XNOR2_X1 U15434 ( .A(n13283), .B(n13282), .ZN(n13284) );
  OAI222_X1 U15435 ( .A1(n13312), .A2(n13285), .B1(n13314), .B2(n13313), .C1(
        n13310), .C2(n13284), .ZN(n13383) );
  INV_X1 U15436 ( .A(n13286), .ZN(n13436) );
  AOI22_X1 U15437 ( .A1(n13328), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13288), 
        .B2(n13287), .ZN(n13289) );
  OAI21_X1 U15438 ( .B1(n13436), .B2(n13341), .A(n13289), .ZN(n13290) );
  AOI21_X1 U15439 ( .B1(n13383), .B2(n13344), .A(n13290), .ZN(n13291) );
  OAI21_X1 U15440 ( .B1(n13305), .B2(n13292), .A(n13291), .ZN(P3_U3212) );
  OAI211_X1 U15441 ( .C1(n13294), .C2(n13301), .A(n13293), .B(n15248), .ZN(
        n13297) );
  AOI22_X1 U15442 ( .A1(n13334), .A2(n15244), .B1(n15242), .B2(n13295), .ZN(
        n13296) );
  AND2_X1 U15443 ( .A1(n13297), .A2(n13296), .ZN(n13389) );
  INV_X1 U15444 ( .A(n13298), .ZN(n13299) );
  OAI22_X1 U15445 ( .A1(n13344), .A2(n13300), .B1(n13299), .B2(n15238), .ZN(
        n13307) );
  NAND2_X1 U15446 ( .A1(n13302), .A2(n13301), .ZN(n13303) );
  NAND2_X1 U15447 ( .A1(n13304), .A2(n13303), .ZN(n13387) );
  NOR2_X1 U15448 ( .A1(n13387), .A2(n13305), .ZN(n13306) );
  AOI211_X1 U15449 ( .C1(n13322), .C2(n13308), .A(n13307), .B(n13306), .ZN(
        n13309) );
  OAI21_X1 U15450 ( .B1(n15258), .B2(n13389), .A(n13309), .ZN(P3_U3213) );
  AOI21_X1 U15451 ( .B1(n13311), .B2(n13325), .A(n13310), .ZN(n13318) );
  OAI22_X1 U15452 ( .A1(n13315), .A2(n13314), .B1(n13313), .B2(n13312), .ZN(
        n13316) );
  AOI21_X1 U15453 ( .B1(n13318), .B2(n13317), .A(n13316), .ZN(n13393) );
  OAI22_X1 U15454 ( .A1(n13344), .A2(n13320), .B1(n13319), .B2(n15238), .ZN(
        n13321) );
  AOI21_X1 U15455 ( .B1(n13323), .B2(n13322), .A(n13321), .ZN(n13327) );
  XNOR2_X1 U15456 ( .A(n13324), .B(n8061), .ZN(n13392) );
  NAND2_X1 U15457 ( .A1(n13392), .A2(n13347), .ZN(n13326) );
  OAI211_X1 U15458 ( .C1(n13393), .C2(n13328), .A(n13327), .B(n13326), .ZN(
        P3_U3214) );
  AND2_X1 U15459 ( .A1(n13330), .A2(n13329), .ZN(n13332) );
  OAI21_X1 U15460 ( .B1(n13332), .B2(n13339), .A(n13331), .ZN(n13335) );
  AOI222_X1 U15461 ( .A1(n15248), .A2(n13335), .B1(n13334), .B2(n15242), .C1(
        n13333), .C2(n15244), .ZN(n13397) );
  INV_X1 U15462 ( .A(n13336), .ZN(n13337) );
  AOI21_X1 U15463 ( .B1(n13339), .B2(n13338), .A(n13337), .ZN(n13399) );
  INV_X1 U15464 ( .A(n13340), .ZN(n13448) );
  NOR2_X1 U15465 ( .A1(n13448), .A2(n13341), .ZN(n13346) );
  OAI22_X1 U15466 ( .A1(n13344), .A2(n13343), .B1(n13342), .B2(n15238), .ZN(
        n13345) );
  AOI211_X1 U15467 ( .C1(n13399), .C2(n13347), .A(n13346), .B(n13345), .ZN(
        n13348) );
  OAI21_X1 U15468 ( .B1(n13397), .B2(n15258), .A(n13348), .ZN(P3_U3215) );
  NOR2_X1 U15469 ( .A1(n13412), .A2(n15696), .ZN(n13351) );
  AOI21_X1 U15470 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15696), .A(n13351), 
        .ZN(n13349) );
  OAI21_X1 U15471 ( .B1(n13350), .B2(n13409), .A(n13349), .ZN(P3_U3490) );
  AOI21_X1 U15472 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15696), .A(n13351), 
        .ZN(n13352) );
  OAI21_X1 U15473 ( .B1(n13417), .B2(n13409), .A(n13352), .ZN(P3_U3489) );
  INV_X1 U15474 ( .A(n13409), .ZN(n13359) );
  INV_X1 U15475 ( .A(n13354), .ZN(P3_U3487) );
  NAND2_X1 U15476 ( .A1(n13355), .A2(n15303), .ZN(n13356) );
  INV_X1 U15477 ( .A(n13360), .ZN(P3_U3486) );
  INV_X1 U15478 ( .A(n13361), .ZN(n13425) );
  INV_X1 U15479 ( .A(n13362), .ZN(n13364) );
  AOI21_X1 U15480 ( .B1(n15303), .B2(n13364), .A(n13363), .ZN(n13422) );
  MUX2_X1 U15481 ( .A(n13365), .B(n13422), .S(n15699), .Z(n13366) );
  OAI21_X1 U15482 ( .B1(n13425), .B2(n13409), .A(n13366), .ZN(P3_U3485) );
  AOI21_X1 U15483 ( .B1(n15302), .B2(n13368), .A(n13367), .ZN(n13369) );
  OAI21_X1 U15484 ( .B1(n9740), .B2(n13370), .A(n13369), .ZN(n13426) );
  MUX2_X1 U15485 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13426), .S(n15699), .Z(
        P3_U3484) );
  AOI21_X1 U15486 ( .B1(n15302), .B2(n13372), .A(n13371), .ZN(n13373) );
  OAI21_X1 U15487 ( .B1(n13374), .B2(n9740), .A(n13373), .ZN(n13427) );
  MUX2_X1 U15488 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13427), .S(n15699), .Z(
        P3_U3483) );
  NAND2_X1 U15489 ( .A1(n13375), .A2(n15302), .ZN(n13376) );
  OAI211_X1 U15490 ( .C1(n9740), .C2(n13378), .A(n13377), .B(n13376), .ZN(
        n13428) );
  MUX2_X1 U15491 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13428), .S(n15699), .Z(
        P3_U3482) );
  INV_X1 U15492 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13381) );
  AOI21_X1 U15493 ( .B1(n15298), .B2(n13380), .A(n13379), .ZN(n13429) );
  MUX2_X1 U15494 ( .A(n13381), .B(n13429), .S(n15699), .Z(n13382) );
  OAI21_X1 U15495 ( .B1(n13432), .B2(n13409), .A(n13382), .ZN(P3_U3481) );
  AOI21_X1 U15496 ( .B1(n13384), .B2(n15298), .A(n13383), .ZN(n13433) );
  MUX2_X1 U15497 ( .A(n13385), .B(n13433), .S(n15699), .Z(n13386) );
  OAI21_X1 U15498 ( .B1(n13436), .B2(n13409), .A(n13386), .ZN(P3_U3480) );
  OR2_X1 U15499 ( .A1(n13387), .A2(n9740), .ZN(n13388) );
  MUX2_X1 U15500 ( .A(n13390), .B(n13438), .S(n15699), .Z(n13391) );
  OAI21_X1 U15501 ( .B1(n13440), .B2(n13409), .A(n13391), .ZN(P3_U3479) );
  NAND2_X1 U15502 ( .A1(n13392), .A2(n15298), .ZN(n13394) );
  AND2_X1 U15503 ( .A1(n13394), .A2(n13393), .ZN(n13442) );
  MUX2_X1 U15504 ( .A(n13395), .B(n13442), .S(n15699), .Z(n13396) );
  OAI21_X1 U15505 ( .B1(n13444), .B2(n13409), .A(n13396), .ZN(P3_U3478) );
  INV_X1 U15506 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13400) );
  INV_X1 U15507 ( .A(n13397), .ZN(n13398) );
  AOI21_X1 U15508 ( .B1(n13399), .B2(n15298), .A(n13398), .ZN(n13445) );
  MUX2_X1 U15509 ( .A(n13400), .B(n13445), .S(n15699), .Z(n13401) );
  OAI21_X1 U15510 ( .B1(n13448), .B2(n13409), .A(n13401), .ZN(P3_U3477) );
  AOI21_X1 U15511 ( .B1(n13403), .B2(n15298), .A(n13402), .ZN(n13449) );
  MUX2_X1 U15512 ( .A(n13404), .B(n13449), .S(n15699), .Z(n13405) );
  OAI21_X1 U15513 ( .B1(n13452), .B2(n13409), .A(n13405), .ZN(P3_U3476) );
  AOI21_X1 U15514 ( .B1(n15298), .B2(n13407), .A(n13406), .ZN(n13453) );
  MUX2_X1 U15515 ( .A(n15443), .B(n13453), .S(n15699), .Z(n13408) );
  OAI21_X1 U15516 ( .B1(n13457), .B2(n13409), .A(n13408), .ZN(P3_U3475) );
  NAND2_X1 U15517 ( .A1(n13411), .A2(n13410), .ZN(n13414) );
  INV_X1 U15518 ( .A(n13412), .ZN(n13413) );
  NAND2_X1 U15519 ( .A1(n13413), .A2(n15309), .ZN(n13416) );
  OAI211_X1 U15520 ( .C1(n12589), .C2(n15309), .A(n13414), .B(n13416), .ZN(
        P3_U3458) );
  NAND2_X1 U15521 ( .A1(n15307), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13415) );
  OAI211_X1 U15522 ( .C1(n13417), .C2(n13456), .A(n13416), .B(n13415), .ZN(
        P3_U3457) );
  INV_X1 U15523 ( .A(n13418), .ZN(n13419) );
  MUX2_X1 U15524 ( .A(n13419), .B(n15474), .S(n15307), .Z(n13420) );
  OAI21_X1 U15525 ( .B1(n13421), .B2(n13456), .A(n13420), .ZN(P3_U3454) );
  INV_X1 U15526 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13423) );
  MUX2_X1 U15527 ( .A(n13423), .B(n13422), .S(n15309), .Z(n13424) );
  OAI21_X1 U15528 ( .B1(n13425), .B2(n13456), .A(n13424), .ZN(P3_U3453) );
  MUX2_X1 U15529 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13426), .S(n15309), .Z(
        P3_U3452) );
  MUX2_X1 U15530 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13427), .S(n15309), .Z(
        P3_U3451) );
  MUX2_X1 U15531 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13428), .S(n15309), .Z(
        P3_U3450) );
  INV_X1 U15532 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13430) );
  MUX2_X1 U15533 ( .A(n13430), .B(n13429), .S(n15309), .Z(n13431) );
  OAI21_X1 U15534 ( .B1(n13432), .B2(n13456), .A(n13431), .ZN(P3_U3449) );
  INV_X1 U15535 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13434) );
  MUX2_X1 U15536 ( .A(n13434), .B(n13433), .S(n15309), .Z(n13435) );
  OAI21_X1 U15537 ( .B1(n13436), .B2(n13456), .A(n13435), .ZN(P3_U3448) );
  MUX2_X1 U15538 ( .A(n13438), .B(n13437), .S(n15307), .Z(n13439) );
  OAI21_X1 U15539 ( .B1(n13440), .B2(n13456), .A(n13439), .ZN(P3_U3447) );
  INV_X1 U15540 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13441) );
  MUX2_X1 U15541 ( .A(n13442), .B(n13441), .S(n15307), .Z(n13443) );
  OAI21_X1 U15542 ( .B1(n13444), .B2(n13456), .A(n13443), .ZN(P3_U3446) );
  MUX2_X1 U15543 ( .A(n13446), .B(n13445), .S(n15309), .Z(n13447) );
  OAI21_X1 U15544 ( .B1(n13448), .B2(n13456), .A(n13447), .ZN(P3_U3444) );
  INV_X1 U15545 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13450) );
  MUX2_X1 U15546 ( .A(n13450), .B(n13449), .S(n15309), .Z(n13451) );
  OAI21_X1 U15547 ( .B1(n13452), .B2(n13456), .A(n13451), .ZN(P3_U3441) );
  INV_X1 U15548 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13454) );
  MUX2_X1 U15549 ( .A(n13454), .B(n13453), .S(n15309), .Z(n13455) );
  OAI21_X1 U15550 ( .B1(n13457), .B2(n13456), .A(n13455), .ZN(P3_U3438) );
  MUX2_X1 U15551 ( .A(P3_D_REG_1__SCAN_IN), .B(n13458), .S(n13459), .Z(
        P3_U3377) );
  MUX2_X1 U15552 ( .A(P3_D_REG_0__SCAN_IN), .B(n13460), .S(n13459), .Z(
        P3_U3376) );
  INV_X1 U15553 ( .A(n13461), .ZN(n13467) );
  NOR4_X1 U15554 ( .A1(n13463), .A2(P3_IR_REG_30__SCAN_IN), .A3(n13462), .A4(
        P3_U3151), .ZN(n13464) );
  AOI21_X1 U15555 ( .B1(n13465), .B2(SI_31_), .A(n13464), .ZN(n13466) );
  OAI21_X1 U15556 ( .B1(n13467), .B2(n6655), .A(n13466), .ZN(P3_U3264) );
  AOI21_X1 U15557 ( .B1(n13470), .B2(n13469), .A(n14999), .ZN(n13472) );
  NAND2_X1 U15558 ( .A1(n13472), .A2(n13471), .ZN(n13478) );
  OAI22_X1 U15559 ( .A1(n13473), .A2(n15148), .B1(n13526), .B2(n13567), .ZN(
        n13682) );
  INV_X1 U15560 ( .A(n13676), .ZN(n13475) );
  OAI22_X1 U15561 ( .A1(n13475), .A2(n15007), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13474), .ZN(n13476) );
  AOI21_X1 U15562 ( .B1(n13682), .B2(n13515), .A(n13476), .ZN(n13477) );
  OAI211_X1 U15563 ( .C1(n13678), .C2(n13539), .A(n13478), .B(n13477), .ZN(
        P2_U3186) );
  INV_X1 U15564 ( .A(n13479), .ZN(n13481) );
  OAI22_X1 U15565 ( .A1(n13481), .A2(n14999), .B1(n13480), .B2(n13561), .ZN(
        n13483) );
  NAND2_X1 U15566 ( .A1(n13483), .A2(n13482), .ZN(n13487) );
  AOI22_X1 U15567 ( .A1(n13583), .A2(n15128), .B1(n15127), .B2(n13585), .ZN(
        n13730) );
  OAI22_X1 U15568 ( .A1(n13730), .A2(n14997), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13484), .ZN(n13485) );
  AOI21_X1 U15569 ( .B1(n13736), .B2(n13546), .A(n13485), .ZN(n13486) );
  OAI211_X1 U15570 ( .C1(n13739), .C2(n13539), .A(n13487), .B(n13486), .ZN(
        P2_U3188) );
  OAI22_X1 U15571 ( .A1(n13513), .A2(n15148), .B1(n13488), .B2(n13567), .ZN(
        n13792) );
  AOI22_X1 U15572 ( .A1(n13515), .A2(n13792), .B1(P2_REG3_REG_19__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13489) );
  OAI21_X1 U15573 ( .B1(n13796), .B2(n15007), .A(n13489), .ZN(n13490) );
  AOI21_X1 U15574 ( .B1(n13896), .B2(n15004), .A(n13490), .ZN(n13497) );
  INV_X1 U15575 ( .A(n13571), .ZN(n13493) );
  NAND3_X1 U15576 ( .A1(n13491), .A2(n13501), .A3(n13589), .ZN(n13492) );
  OAI21_X1 U15577 ( .B1(n13493), .B2(n14999), .A(n13492), .ZN(n13495) );
  NAND2_X1 U15578 ( .A1(n13495), .A2(n13494), .ZN(n13496) );
  OAI211_X1 U15579 ( .C1(n6838), .C2(n14999), .A(n13497), .B(n13496), .ZN(
        P2_U3191) );
  AOI22_X1 U15580 ( .A1(n13547), .A2(n15129), .B1(n13541), .B2(n11972), .ZN(
        n13509) );
  AOI22_X1 U15581 ( .A1(n15004), .A2(n15143), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13498), .ZN(n13508) );
  NAND3_X1 U15582 ( .A1(n13501), .A2(n13500), .A3(n13499), .ZN(n13507) );
  OAI21_X1 U15583 ( .B1(n13504), .B2(n13503), .A(n13502), .ZN(n13505) );
  NAND2_X1 U15584 ( .A1(n13552), .A2(n13505), .ZN(n13506) );
  NAND4_X1 U15585 ( .A1(n13509), .A2(n13508), .A3(n13507), .A4(n13506), .ZN(
        P2_U3194) );
  OAI211_X1 U15586 ( .C1(n13512), .C2(n13511), .A(n13510), .B(n13552), .ZN(
        n13519) );
  OAI22_X1 U15587 ( .A1(n13514), .A2(n15148), .B1(n13513), .B2(n13567), .ZN(
        n13762) );
  AOI22_X1 U15588 ( .A1(n13762), .A2(n13515), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13518) );
  NAND2_X1 U15589 ( .A1(n13886), .A2(n15004), .ZN(n13517) );
  NAND2_X1 U15590 ( .A1(n13546), .A2(n13766), .ZN(n13516) );
  NAND4_X1 U15591 ( .A1(n13519), .A2(n13518), .A3(n13517), .A4(n13516), .ZN(
        P2_U3195) );
  INV_X1 U15592 ( .A(n13583), .ZN(n13525) );
  NOR3_X1 U15593 ( .A1(n13520), .A2(n13525), .A3(n13561), .ZN(n13524) );
  AOI21_X1 U15594 ( .B1(n13521), .B2(n13522), .A(n14999), .ZN(n13523) );
  OAI21_X1 U15595 ( .B1(n13524), .B2(n13523), .A(n6754), .ZN(n13531) );
  OAI22_X1 U15596 ( .A1(n13526), .A2(n15148), .B1(n13525), .B2(n13567), .ZN(
        n13701) );
  INV_X1 U15597 ( .A(n13708), .ZN(n13528) );
  OAI22_X1 U15598 ( .A1(n13528), .A2(n15007), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13527), .ZN(n13529) );
  AOI21_X1 U15599 ( .B1(n13701), .B2(n13515), .A(n13529), .ZN(n13530) );
  OAI211_X1 U15600 ( .C1(n13711), .C2(n13539), .A(n13531), .B(n13530), .ZN(
        P2_U3197) );
  OAI211_X1 U15601 ( .C1(n13533), .C2(n13532), .A(n13521), .B(n13552), .ZN(
        n13538) );
  INV_X1 U15602 ( .A(n13534), .ZN(n13722) );
  AOI22_X1 U15603 ( .A1(n13582), .A2(n15128), .B1(n15127), .B2(n13584), .ZN(
        n13716) );
  OAI22_X1 U15604 ( .A1(n13716), .A2(n14997), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13535), .ZN(n13536) );
  AOI21_X1 U15605 ( .B1(n13722), .B2(n13546), .A(n13536), .ZN(n13537) );
  OAI211_X1 U15606 ( .C1(n13725), .C2(n13539), .A(n13538), .B(n13537), .ZN(
        P2_U3201) );
  NOR3_X1 U15607 ( .A1(n13561), .A2(n13540), .A3(n13550), .ZN(n13542) );
  OAI21_X1 U15608 ( .B1(n13542), .B2(n13541), .A(n13605), .ZN(n13556) );
  AOI22_X1 U15609 ( .A1(n15004), .A2(n13543), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13555) );
  INV_X1 U15610 ( .A(n13544), .ZN(n13545) );
  AOI22_X1 U15611 ( .A1(n13547), .A2(n13603), .B1(n13546), .B2(n13545), .ZN(
        n13554) );
  OAI21_X1 U15612 ( .B1(n13550), .B2(n13549), .A(n13548), .ZN(n13551) );
  NAND2_X1 U15613 ( .A1(n13552), .A2(n13551), .ZN(n13553) );
  NAND4_X1 U15614 ( .A1(n13556), .A2(n13555), .A3(n13554), .A4(n13553), .ZN(
        P2_U3202) );
  INV_X1 U15615 ( .A(n13557), .ZN(n13780) );
  OAI22_X1 U15616 ( .A1(n13558), .A2(n15148), .B1(n13569), .B2(n13567), .ZN(
        n13776) );
  AOI22_X1 U15617 ( .A1(n13776), .A2(n13515), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13559) );
  OAI21_X1 U15618 ( .B1(n13780), .B2(n15007), .A(n13559), .ZN(n13560) );
  AOI21_X1 U15619 ( .B1(n13891), .B2(n15004), .A(n13560), .ZN(n13566) );
  OAI22_X1 U15620 ( .A1(n13562), .A2(n14999), .B1(n13569), .B2(n13561), .ZN(
        n13563) );
  NAND3_X1 U15621 ( .A1(n6838), .A2(n13564), .A3(n13563), .ZN(n13565) );
  OAI211_X1 U15622 ( .C1(n6855), .C2(n14999), .A(n13566), .B(n13565), .ZN(
        P2_U3205) );
  OAI22_X1 U15623 ( .A1(n13569), .A2(n15148), .B1(n13568), .B2(n13567), .ZN(
        n13806) );
  NAND2_X1 U15624 ( .A1(n13515), .A2(n13806), .ZN(n13570) );
  NAND2_X1 U15625 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15109)
         );
  OAI211_X1 U15626 ( .C1(n15007), .C2(n13815), .A(n13570), .B(n15109), .ZN(
        n13575) );
  AOI211_X1 U15627 ( .C1(n13573), .C2(n13572), .A(n14999), .B(n13571), .ZN(
        n13574) );
  AOI211_X1 U15628 ( .C1(n13902), .C2(n15004), .A(n13575), .B(n13574), .ZN(
        n13576) );
  INV_X1 U15629 ( .A(n13576), .ZN(P2_U3210) );
  INV_X2 U15630 ( .A(P2_U3947), .ZN(n13599) );
  MUX2_X1 U15631 ( .A(n13646), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13599), .Z(
        P2_U3562) );
  MUX2_X1 U15632 ( .A(n13577), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13599), .Z(
        P2_U3561) );
  MUX2_X1 U15633 ( .A(n13578), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13599), .Z(
        P2_U3560) );
  MUX2_X1 U15634 ( .A(n13579), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13599), .Z(
        P2_U3559) );
  MUX2_X1 U15635 ( .A(n13580), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13599), .Z(
        P2_U3558) );
  MUX2_X1 U15636 ( .A(n13581), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13599), .Z(
        P2_U3557) );
  MUX2_X1 U15637 ( .A(n13582), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13599), .Z(
        P2_U3556) );
  MUX2_X1 U15638 ( .A(n13583), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13599), .Z(
        P2_U3555) );
  MUX2_X1 U15639 ( .A(n13584), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13599), .Z(
        P2_U3554) );
  MUX2_X1 U15640 ( .A(n13585), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13599), .Z(
        P2_U3553) );
  MUX2_X1 U15641 ( .A(n13586), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13599), .Z(
        P2_U3552) );
  MUX2_X1 U15642 ( .A(n13587), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13599), .Z(
        P2_U3551) );
  MUX2_X1 U15643 ( .A(n13588), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13599), .Z(
        P2_U3550) );
  MUX2_X1 U15644 ( .A(n13589), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13599), .Z(
        P2_U3549) );
  MUX2_X1 U15645 ( .A(n13590), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13599), .Z(
        P2_U3548) );
  MUX2_X1 U15646 ( .A(n13591), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13599), .Z(
        P2_U3547) );
  MUX2_X1 U15647 ( .A(n13592), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13599), .Z(
        P2_U3546) );
  MUX2_X1 U15648 ( .A(n13593), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13599), .Z(
        P2_U3545) );
  MUX2_X1 U15649 ( .A(n13594), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13599), .Z(
        P2_U3544) );
  MUX2_X1 U15650 ( .A(n13595), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13599), .Z(
        P2_U3543) );
  MUX2_X1 U15651 ( .A(n13596), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13599), .Z(
        P2_U3542) );
  MUX2_X1 U15652 ( .A(n13597), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13599), .Z(
        P2_U3541) );
  MUX2_X1 U15653 ( .A(n13598), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13599), .Z(
        P2_U3540) );
  MUX2_X1 U15654 ( .A(n13600), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13599), .Z(
        P2_U3539) );
  MUX2_X1 U15655 ( .A(n13601), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13599), .Z(
        P2_U3538) );
  MUX2_X1 U15656 ( .A(n13602), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13599), .Z(
        P2_U3537) );
  MUX2_X1 U15657 ( .A(n13603), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13599), .Z(
        P2_U3536) );
  MUX2_X1 U15658 ( .A(n13604), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13599), .Z(
        P2_U3535) );
  MUX2_X1 U15659 ( .A(n13605), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13599), .Z(
        P2_U3534) );
  MUX2_X1 U15660 ( .A(n15129), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13599), .Z(
        P2_U3533) );
  MUX2_X1 U15661 ( .A(n13606), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13599), .Z(
        P2_U3532) );
  MUX2_X1 U15662 ( .A(n11972), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13599), .Z(
        P2_U3531) );
  XOR2_X1 U15663 ( .A(n13608), .B(n13607), .Z(n13609) );
  AOI22_X1 U15664 ( .A1(n13610), .A2(n15089), .B1(n15085), .B2(n13609), .ZN(
        n13617) );
  OAI211_X1 U15665 ( .C1(n13613), .C2(n13612), .A(n15091), .B(n13611), .ZN(
        n13616) );
  NAND2_X1 U15666 ( .A1(n15083), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n13615) );
  NAND2_X1 U15667 ( .A1(P2_U3088), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n13614) );
  NAND4_X1 U15668 ( .A1(n13617), .A2(n13616), .A3(n13615), .A4(n13614), .ZN(
        P2_U3216) );
  INV_X1 U15669 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n15529) );
  NAND2_X1 U15670 ( .A1(n15088), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13621) );
  INV_X1 U15671 ( .A(n13621), .ZN(n13618) );
  AOI21_X1 U15672 ( .B1(n13829), .B2(n13628), .A(n13618), .ZN(n15093) );
  OAI21_X1 U15673 ( .B1(n13627), .B2(n13620), .A(n13619), .ZN(n15092) );
  NAND2_X1 U15674 ( .A1(n15093), .A2(n15092), .ZN(n15090) );
  NAND2_X1 U15675 ( .A1(n13621), .A2(n15090), .ZN(n13622) );
  NOR2_X1 U15676 ( .A1(n13631), .A2(n13622), .ZN(n13623) );
  XNOR2_X1 U15677 ( .A(n13631), .B(n13622), .ZN(n15099) );
  NOR2_X1 U15678 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n15099), .ZN(n15098) );
  NOR2_X1 U15679 ( .A1(n13623), .A2(n15098), .ZN(n13624) );
  XOR2_X1 U15680 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13624), .Z(n13635) );
  XNOR2_X1 U15681 ( .A(n13628), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15087) );
  INV_X1 U15682 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13626) );
  OAI21_X1 U15683 ( .B1(n13627), .B2(n13626), .A(n13625), .ZN(n15086) );
  NAND2_X1 U15684 ( .A1(n15087), .A2(n15086), .ZN(n15084) );
  OAI21_X1 U15685 ( .B1(n13629), .B2(n13628), .A(n15084), .ZN(n13630) );
  NAND2_X1 U15686 ( .A1(n13631), .A2(n13630), .ZN(n13632) );
  XOR2_X1 U15687 ( .A(n13631), .B(n13630), .Z(n15101) );
  NAND2_X1 U15688 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n15101), .ZN(n15100) );
  NAND2_X1 U15689 ( .A1(n13632), .A2(n15100), .ZN(n13633) );
  XOR2_X1 U15690 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13633), .Z(n13634) );
  AOI22_X1 U15691 ( .A1(n13635), .A2(n15091), .B1(n15085), .B2(n13634), .ZN(
        n13640) );
  INV_X1 U15692 ( .A(n13634), .ZN(n13637) );
  NOR2_X1 U15693 ( .A1(n13635), .A2(n15105), .ZN(n13636) );
  AOI211_X1 U15694 ( .C1(n15085), .C2(n13637), .A(n15089), .B(n13636), .ZN(
        n13639) );
  MUX2_X1 U15695 ( .A(n13640), .B(n13639), .S(n13638), .Z(n13642) );
  NAND2_X1 U15696 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n13641)
         );
  OAI211_X1 U15697 ( .C1(n15529), .C2(n15111), .A(n13642), .B(n13641), .ZN(
        P2_U3233) );
  NAND2_X1 U15698 ( .A1(n13652), .A2(n13843), .ZN(n13651) );
  NAND2_X1 U15699 ( .A1(n13647), .A2(n13646), .ZN(n13841) );
  NOR2_X1 U15700 ( .A1(n15157), .A2(n13841), .ZN(n13654) );
  NOR2_X1 U15701 ( .A1(n13644), .A2(n13813), .ZN(n13649) );
  AOI211_X1 U15702 ( .C1(n15157), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13654), 
        .B(n13649), .ZN(n13650) );
  OAI21_X1 U15703 ( .B1(n13840), .B2(n15140), .A(n13650), .ZN(P2_U3234) );
  OAI211_X1 U15704 ( .C1(n13652), .C2(n13843), .A(n15134), .B(n13651), .ZN(
        n13842) );
  NOR2_X1 U15705 ( .A1(n13843), .A2(n13813), .ZN(n13653) );
  AOI211_X1 U15706 ( .C1(n15157), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13654), 
        .B(n13653), .ZN(n13655) );
  OAI21_X1 U15707 ( .B1(n13842), .B2(n15140), .A(n13655), .ZN(P2_U3235) );
  XNOR2_X1 U15708 ( .A(n13657), .B(n13656), .ZN(n13853) );
  OR2_X1 U15709 ( .A1(n13851), .A2(n13675), .ZN(n13658) );
  INV_X1 U15710 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13660) );
  OAI22_X1 U15711 ( .A1(n13661), .A2(n15132), .B1(n13660), .B2(n15155), .ZN(
        n13662) );
  INV_X1 U15712 ( .A(n13662), .ZN(n13663) );
  OAI21_X1 U15713 ( .B1(n13851), .B2(n13813), .A(n13663), .ZN(n13664) );
  AOI21_X1 U15714 ( .B1(n13850), .B2(n13835), .A(n13664), .ZN(n13673) );
  NAND2_X1 U15715 ( .A1(n13665), .A2(n15131), .ZN(n13671) );
  AOI21_X1 U15716 ( .B1(n13679), .B2(n13667), .A(n13666), .ZN(n13670) );
  INV_X1 U15717 ( .A(n13668), .ZN(n13669) );
  OAI21_X1 U15718 ( .B1(n13671), .B2(n13670), .A(n13669), .ZN(n13849) );
  NAND2_X1 U15719 ( .A1(n13849), .A2(n15155), .ZN(n13672) );
  OAI211_X1 U15720 ( .C1(n13853), .C2(n15139), .A(n13673), .B(n13672), .ZN(
        P2_U3237) );
  NOR2_X1 U15721 ( .A1(n13678), .A2(n13691), .ZN(n13674) );
  AOI22_X1 U15722 ( .A1(n13676), .A2(n15154), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15157), .ZN(n13677) );
  OAI21_X1 U15723 ( .B1(n13678), .B2(n13813), .A(n13677), .ZN(n13685) );
  OAI21_X1 U15724 ( .B1(n13681), .B2(n13680), .A(n13679), .ZN(n13683) );
  NOR2_X1 U15725 ( .A1(n13859), .A2(n15157), .ZN(n13684) );
  AOI211_X1 U15726 ( .C1(n7659), .C2(n13835), .A(n13685), .B(n13684), .ZN(
        n13686) );
  OAI21_X1 U15727 ( .B1(n13860), .B2(n15139), .A(n13686), .ZN(P2_U3238) );
  XNOR2_X1 U15728 ( .A(n13687), .B(n13696), .ZN(n13689) );
  AOI21_X1 U15729 ( .B1(n13689), .B2(n15131), .A(n13688), .ZN(n13863) );
  NOR2_X1 U15730 ( .A1(n13694), .A2(n13707), .ZN(n13690) );
  AOI22_X1 U15731 ( .A1(n13692), .A2(n15154), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15157), .ZN(n13693) );
  OAI21_X1 U15732 ( .B1(n13694), .B2(n13813), .A(n13693), .ZN(n13698) );
  XOR2_X1 U15733 ( .A(n13696), .B(n13695), .Z(n13864) );
  NOR2_X1 U15734 ( .A1(n13864), .A2(n15139), .ZN(n13697) );
  AOI211_X1 U15735 ( .C1(n7647), .C2(n13835), .A(n13698), .B(n13697), .ZN(
        n13699) );
  OAI21_X1 U15736 ( .B1(n15157), .B2(n13863), .A(n13699), .ZN(P2_U3239) );
  XNOR2_X1 U15737 ( .A(n13700), .B(n13703), .ZN(n13702) );
  AOI21_X1 U15738 ( .B1(n13702), .B2(n15131), .A(n13701), .ZN(n13868) );
  XNOR2_X1 U15739 ( .A(n13704), .B(n13703), .ZN(n13869) );
  INV_X1 U15740 ( .A(n13869), .ZN(n13713) );
  NAND2_X1 U15741 ( .A1(n13866), .A2(n6804), .ZN(n13705) );
  NAND2_X1 U15742 ( .A1(n13705), .A2(n15134), .ZN(n13706) );
  NOR2_X1 U15743 ( .A1(n13707), .A2(n13706), .ZN(n13865) );
  NAND2_X1 U15744 ( .A1(n13865), .A2(n13835), .ZN(n13710) );
  AOI22_X1 U15745 ( .A1(n13708), .A2(n15154), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n15157), .ZN(n13709) );
  OAI211_X1 U15746 ( .C1(n13711), .C2(n13813), .A(n13710), .B(n13709), .ZN(
        n13712) );
  AOI21_X1 U15747 ( .B1(n13713), .B2(n15122), .A(n13712), .ZN(n13714) );
  OAI21_X1 U15748 ( .B1(n15157), .B2(n13868), .A(n13714), .ZN(P2_U3240) );
  XNOR2_X1 U15749 ( .A(n13715), .B(n13719), .ZN(n13718) );
  INV_X1 U15750 ( .A(n13716), .ZN(n13717) );
  AOI21_X1 U15751 ( .B1(n13718), .B2(n15131), .A(n13717), .ZN(n13873) );
  XNOR2_X1 U15752 ( .A(n13720), .B(n13719), .ZN(n13874) );
  INV_X1 U15753 ( .A(n13874), .ZN(n13727) );
  AOI21_X1 U15754 ( .B1(n13871), .B2(n6761), .A(n13753), .ZN(n13721) );
  AND2_X1 U15755 ( .A1(n13721), .A2(n6804), .ZN(n13870) );
  NAND2_X1 U15756 ( .A1(n13870), .A2(n13835), .ZN(n13724) );
  AOI22_X1 U15757 ( .A1(n13722), .A2(n15154), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n15157), .ZN(n13723) );
  OAI211_X1 U15758 ( .C1(n13725), .C2(n13813), .A(n13724), .B(n13723), .ZN(
        n13726) );
  AOI21_X1 U15759 ( .B1(n13727), .B2(n15122), .A(n13726), .ZN(n13728) );
  OAI21_X1 U15760 ( .B1(n15157), .B2(n13873), .A(n13728), .ZN(P2_U3241) );
  XNOR2_X1 U15761 ( .A(n13729), .B(n13733), .ZN(n13732) );
  INV_X1 U15762 ( .A(n13730), .ZN(n13731) );
  AOI21_X1 U15763 ( .B1(n13732), .B2(n15131), .A(n13731), .ZN(n13878) );
  XNOR2_X1 U15764 ( .A(n13734), .B(n13733), .ZN(n13879) );
  INV_X1 U15765 ( .A(n13879), .ZN(n13741) );
  AOI21_X1 U15766 ( .B1(n13876), .B2(n13754), .A(n13753), .ZN(n13735) );
  AND2_X1 U15767 ( .A1(n13735), .A2(n6761), .ZN(n13875) );
  NAND2_X1 U15768 ( .A1(n13875), .A2(n13835), .ZN(n13738) );
  AOI22_X1 U15769 ( .A1(n15157), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n13736), 
        .B2(n15154), .ZN(n13737) );
  OAI211_X1 U15770 ( .C1(n13739), .C2(n13813), .A(n13738), .B(n13737), .ZN(
        n13740) );
  AOI21_X1 U15771 ( .B1(n13741), .B2(n15122), .A(n13740), .ZN(n13742) );
  OAI21_X1 U15772 ( .B1(n15157), .B2(n13878), .A(n13742), .ZN(P2_U3242) );
  XOR2_X1 U15773 ( .A(n13748), .B(n13743), .Z(n13745) );
  AOI21_X1 U15774 ( .B1(n13745), .B2(n15131), .A(n13744), .ZN(n13883) );
  AOI21_X1 U15775 ( .B1(n13748), .B2(n13747), .A(n13746), .ZN(n13749) );
  INV_X1 U15776 ( .A(n13749), .ZN(n13884) );
  OAI22_X1 U15777 ( .A1(n15155), .A2(n13751), .B1(n13750), .B2(n15132), .ZN(
        n13752) );
  AOI21_X1 U15778 ( .B1(n13881), .B2(n15144), .A(n13752), .ZN(n13757) );
  AOI21_X1 U15779 ( .B1(n13881), .B2(n13765), .A(n13753), .ZN(n13755) );
  AND2_X1 U15780 ( .A1(n13755), .A2(n13754), .ZN(n13880) );
  NAND2_X1 U15781 ( .A1(n13880), .A2(n13835), .ZN(n13756) );
  OAI211_X1 U15782 ( .C1(n13884), .C2(n15139), .A(n13757), .B(n13756), .ZN(
        n13758) );
  INV_X1 U15783 ( .A(n13758), .ZN(n13759) );
  OAI21_X1 U15784 ( .B1(n15157), .B2(n13883), .A(n13759), .ZN(P2_U3243) );
  XNOR2_X1 U15785 ( .A(n13761), .B(n13760), .ZN(n13763) );
  AOI21_X1 U15786 ( .B1(n13763), .B2(n15131), .A(n13762), .ZN(n13888) );
  OR2_X1 U15787 ( .A1(n7485), .A2(n13785), .ZN(n13764) );
  AND3_X1 U15788 ( .A1(n13765), .A2(n13764), .A3(n15134), .ZN(n13885) );
  NAND2_X1 U15789 ( .A1(n13886), .A2(n15144), .ZN(n13768) );
  NAND2_X1 U15790 ( .A1(n13766), .A2(n15154), .ZN(n13767) );
  OAI211_X1 U15791 ( .C1(n15155), .C2(n13769), .A(n13768), .B(n13767), .ZN(
        n13773) );
  XNOR2_X1 U15792 ( .A(n13771), .B(n13770), .ZN(n13889) );
  NOR2_X1 U15793 ( .A1(n13889), .A2(n15139), .ZN(n13772) );
  AOI211_X1 U15794 ( .C1(n13885), .C2(n13835), .A(n13773), .B(n13772), .ZN(
        n13774) );
  OAI21_X1 U15795 ( .B1(n15157), .B2(n13888), .A(n13774), .ZN(P2_U3244) );
  XNOR2_X1 U15796 ( .A(n13775), .B(n13778), .ZN(n13777) );
  AOI21_X1 U15797 ( .B1(n13777), .B2(n15131), .A(n13776), .ZN(n13893) );
  XNOR2_X1 U15798 ( .A(n13779), .B(n13778), .ZN(n13894) );
  INV_X1 U15799 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13781) );
  OAI22_X1 U15800 ( .A1(n15155), .A2(n13781), .B1(n13780), .B2(n15132), .ZN(
        n13782) );
  AOI21_X1 U15801 ( .B1(n13891), .B2(n15144), .A(n13782), .ZN(n13787) );
  NAND2_X1 U15802 ( .A1(n13794), .A2(n13891), .ZN(n13783) );
  NAND2_X1 U15803 ( .A1(n13783), .A2(n15134), .ZN(n13784) );
  NOR2_X1 U15804 ( .A1(n13785), .A2(n13784), .ZN(n13890) );
  NAND2_X1 U15805 ( .A1(n13890), .A2(n13835), .ZN(n13786) );
  OAI211_X1 U15806 ( .C1(n13894), .C2(n15139), .A(n13787), .B(n13786), .ZN(
        n13788) );
  INV_X1 U15807 ( .A(n13788), .ZN(n13789) );
  OAI21_X1 U15808 ( .B1(n13893), .B2(n15157), .A(n13789), .ZN(P2_U3245) );
  XNOR2_X1 U15809 ( .A(n13791), .B(n13800), .ZN(n13793) );
  AOI21_X1 U15810 ( .B1(n13793), .B2(n15131), .A(n13792), .ZN(n13898) );
  INV_X1 U15811 ( .A(n13794), .ZN(n13795) );
  AOI211_X1 U15812 ( .C1(n13896), .C2(n13811), .A(n12009), .B(n13795), .ZN(
        n13895) );
  INV_X1 U15813 ( .A(n13796), .ZN(n13797) );
  AOI22_X1 U15814 ( .A1(n15157), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13797), 
        .B2(n15154), .ZN(n13798) );
  OAI21_X1 U15815 ( .B1(n13799), .B2(n13813), .A(n13798), .ZN(n13803) );
  XOR2_X1 U15816 ( .A(n13801), .B(n13800), .Z(n13899) );
  NOR2_X1 U15817 ( .A1(n13899), .A2(n15139), .ZN(n13802) );
  AOI211_X1 U15818 ( .C1(n13895), .C2(n13835), .A(n13803), .B(n13802), .ZN(
        n13804) );
  OAI21_X1 U15819 ( .B1(n15157), .B2(n13898), .A(n13804), .ZN(P2_U3246) );
  XNOR2_X1 U15820 ( .A(n13805), .B(n13809), .ZN(n13807) );
  AOI21_X1 U15821 ( .B1(n13807), .B2(n15131), .A(n13806), .ZN(n13904) );
  OAI21_X1 U15822 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(n13900) );
  NAND2_X1 U15823 ( .A1(n13900), .A2(n15122), .ZN(n13820) );
  INV_X1 U15824 ( .A(n13811), .ZN(n13812) );
  AOI211_X1 U15825 ( .C1(n13902), .C2(n7078), .A(n12009), .B(n13812), .ZN(
        n13901) );
  NOR2_X1 U15826 ( .A1(n13814), .A2(n13813), .ZN(n13818) );
  OAI22_X1 U15827 ( .A1(n15155), .A2(n13816), .B1(n13815), .B2(n15132), .ZN(
        n13817) );
  AOI211_X1 U15828 ( .C1(n13901), .C2(n13835), .A(n13818), .B(n13817), .ZN(
        n13819) );
  OAI211_X1 U15829 ( .C1(n15157), .C2(n13904), .A(n13820), .B(n13819), .ZN(
        P2_U3247) );
  XNOR2_X1 U15830 ( .A(n13821), .B(n13825), .ZN(n13823) );
  AOI21_X1 U15831 ( .B1(n13823), .B2(n15131), .A(n13822), .ZN(n13909) );
  AOI21_X1 U15832 ( .B1(n13826), .B2(n13825), .A(n13824), .ZN(n13827) );
  INV_X1 U15833 ( .A(n13827), .ZN(n13910) );
  OAI22_X1 U15834 ( .A1(n15155), .A2(n13829), .B1(n13828), .B2(n15132), .ZN(
        n13830) );
  AOI21_X1 U15835 ( .B1(n13907), .B2(n15144), .A(n13830), .ZN(n13837) );
  NAND2_X1 U15836 ( .A1(n13831), .A2(n13907), .ZN(n13832) );
  NAND2_X1 U15837 ( .A1(n13832), .A2(n15134), .ZN(n13833) );
  NOR2_X1 U15838 ( .A1(n13834), .A2(n13833), .ZN(n13906) );
  NAND2_X1 U15839 ( .A1(n13906), .A2(n13835), .ZN(n13836) );
  OAI211_X1 U15840 ( .C1(n13910), .C2(n15139), .A(n13837), .B(n13836), .ZN(
        n13838) );
  INV_X1 U15841 ( .A(n13838), .ZN(n13839) );
  OAI21_X1 U15842 ( .B1(n15157), .B2(n13909), .A(n13839), .ZN(P2_U3248) );
  OAI211_X1 U15843 ( .C1(n13644), .C2(n15215), .A(n13840), .B(n13841), .ZN(
        n13926) );
  MUX2_X1 U15844 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13926), .S(n15233), .Z(
        P2_U3530) );
  OAI211_X1 U15845 ( .C1(n13843), .C2(n15215), .A(n13842), .B(n13841), .ZN(
        n13927) );
  MUX2_X1 U15846 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13927), .S(n15233), .Z(
        P2_U3529) );
  INV_X1 U15847 ( .A(n13849), .ZN(n13856) );
  INV_X1 U15848 ( .A(n13850), .ZN(n13852) );
  NAND3_X1 U15849 ( .A1(n13856), .A2(n13855), .A3(n13854), .ZN(n13929) );
  MUX2_X1 U15850 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13929), .S(n15233), .Z(
        P2_U3527) );
  AOI21_X1 U15851 ( .B1(n15196), .B2(n13857), .A(n7659), .ZN(n13858) );
  OAI211_X1 U15852 ( .C1(n13860), .C2(n15187), .A(n13859), .B(n13858), .ZN(
        n13930) );
  MUX2_X1 U15853 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13930), .S(n15233), .Z(
        P2_U3526) );
  AOI21_X1 U15854 ( .B1(n15196), .B2(n13861), .A(n7647), .ZN(n13862) );
  OAI211_X1 U15855 ( .C1(n13864), .C2(n15187), .A(n13863), .B(n13862), .ZN(
        n13931) );
  MUX2_X1 U15856 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13931), .S(n15233), .Z(
        P2_U3525) );
  AOI21_X1 U15857 ( .B1(n15196), .B2(n13866), .A(n13865), .ZN(n13867) );
  OAI211_X1 U15858 ( .C1(n13869), .C2(n15187), .A(n13868), .B(n13867), .ZN(
        n13932) );
  MUX2_X1 U15859 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13932), .S(n15233), .Z(
        P2_U3524) );
  AOI21_X1 U15860 ( .B1(n15196), .B2(n13871), .A(n13870), .ZN(n13872) );
  OAI211_X1 U15861 ( .C1(n13874), .C2(n15187), .A(n13873), .B(n13872), .ZN(
        n13933) );
  MUX2_X1 U15862 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13933), .S(n15233), .Z(
        P2_U3523) );
  AOI21_X1 U15863 ( .B1(n15196), .B2(n13876), .A(n13875), .ZN(n13877) );
  OAI211_X1 U15864 ( .C1(n13879), .C2(n15187), .A(n13878), .B(n13877), .ZN(
        n13934) );
  MUX2_X1 U15865 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13934), .S(n15233), .Z(
        P2_U3522) );
  AOI21_X1 U15866 ( .B1(n15196), .B2(n13881), .A(n13880), .ZN(n13882) );
  OAI211_X1 U15867 ( .C1(n13884), .C2(n15187), .A(n13883), .B(n13882), .ZN(
        n13935) );
  MUX2_X1 U15868 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13935), .S(n15233), .Z(
        P2_U3521) );
  AOI21_X1 U15869 ( .B1(n15196), .B2(n13886), .A(n13885), .ZN(n13887) );
  OAI211_X1 U15870 ( .C1(n13889), .C2(n15187), .A(n13888), .B(n13887), .ZN(
        n13936) );
  MUX2_X1 U15871 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13936), .S(n15233), .Z(
        P2_U3520) );
  AOI21_X1 U15872 ( .B1(n15196), .B2(n13891), .A(n13890), .ZN(n13892) );
  OAI211_X1 U15873 ( .C1(n15187), .C2(n13894), .A(n13893), .B(n13892), .ZN(
        n13937) );
  MUX2_X1 U15874 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13937), .S(n15233), .Z(
        P2_U3519) );
  AOI21_X1 U15875 ( .B1(n15196), .B2(n13896), .A(n13895), .ZN(n13897) );
  OAI211_X1 U15876 ( .C1(n13899), .C2(n15187), .A(n13898), .B(n13897), .ZN(
        n13938) );
  MUX2_X1 U15877 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13938), .S(n15233), .Z(
        P2_U3518) );
  INV_X1 U15878 ( .A(n13900), .ZN(n13905) );
  AOI21_X1 U15879 ( .B1(n15196), .B2(n13902), .A(n13901), .ZN(n13903) );
  OAI211_X1 U15880 ( .C1(n13905), .C2(n15187), .A(n13904), .B(n13903), .ZN(
        n13939) );
  MUX2_X1 U15881 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13939), .S(n15233), .Z(
        P2_U3517) );
  AOI21_X1 U15882 ( .B1(n15196), .B2(n13907), .A(n13906), .ZN(n13908) );
  OAI211_X1 U15883 ( .C1(n13910), .C2(n15187), .A(n13909), .B(n13908), .ZN(
        n13940) );
  MUX2_X1 U15884 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13940), .S(n15233), .Z(
        P2_U3516) );
  NAND2_X1 U15885 ( .A1(n13911), .A2(n15196), .ZN(n13912) );
  AND2_X1 U15886 ( .A1(n13913), .A2(n13912), .ZN(n13914) );
  OAI211_X1 U15887 ( .C1(n15187), .C2(n13916), .A(n13915), .B(n13914), .ZN(
        n13941) );
  MUX2_X1 U15888 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13941), .S(n15233), .Z(
        P2_U3515) );
  AOI21_X1 U15889 ( .B1(n15196), .B2(n13918), .A(n13917), .ZN(n13920) );
  OAI211_X1 U15890 ( .C1(n15187), .C2(n13921), .A(n13920), .B(n13919), .ZN(
        n13942) );
  MUX2_X1 U15891 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13942), .S(n15233), .Z(
        P2_U3514) );
  AOI21_X1 U15892 ( .B1(n15196), .B2(n11505), .A(n13922), .ZN(n13924) );
  OAI211_X1 U15893 ( .C1(n15187), .C2(n13925), .A(n13924), .B(n13923), .ZN(
        n13943) );
  MUX2_X1 U15894 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13943), .S(n15233), .Z(
        P2_U3513) );
  INV_X2 U15895 ( .A(n15222), .ZN(n15212) );
  MUX2_X1 U15896 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13926), .S(n15212), .Z(
        P2_U3498) );
  MUX2_X1 U15897 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13927), .S(n15212), .Z(
        P2_U3497) );
  MUX2_X1 U15898 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13928), .S(n15212), .Z(
        P2_U3496) );
  MUX2_X1 U15899 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13929), .S(n15212), .Z(
        P2_U3495) );
  MUX2_X1 U15900 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13930), .S(n15212), .Z(
        P2_U3494) );
  MUX2_X1 U15901 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13931), .S(n15212), .Z(
        P2_U3493) );
  MUX2_X1 U15902 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13932), .S(n15212), .Z(
        P2_U3492) );
  MUX2_X1 U15903 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13933), .S(n15212), .Z(
        P2_U3491) );
  MUX2_X1 U15904 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13934), .S(n15212), .Z(
        P2_U3490) );
  MUX2_X1 U15905 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13935), .S(n15212), .Z(
        P2_U3489) );
  MUX2_X1 U15906 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13936), .S(n15212), .Z(
        P2_U3488) );
  MUX2_X1 U15907 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13937), .S(n15212), .Z(
        P2_U3487) );
  MUX2_X1 U15908 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13938), .S(n15212), .Z(
        P2_U3486) );
  MUX2_X1 U15909 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13939), .S(n15212), .Z(
        P2_U3484) );
  MUX2_X1 U15910 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13940), .S(n15212), .Z(
        P2_U3481) );
  MUX2_X1 U15911 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13941), .S(n15212), .Z(
        P2_U3478) );
  MUX2_X1 U15912 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13942), .S(n15212), .Z(
        P2_U3475) );
  MUX2_X1 U15913 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13943), .S(n15212), .Z(
        P2_U3472) );
  INV_X1 U15914 ( .A(n13944), .ZN(n14653) );
  NOR4_X1 U15915 ( .A1(n13946), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13945), .A4(
        P2_U3088), .ZN(n13947) );
  AOI21_X1 U15916 ( .B1(n13953), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13947), 
        .ZN(n13948) );
  OAI21_X1 U15917 ( .B1(n14653), .B2(n13955), .A(n13948), .ZN(P2_U3296) );
  INV_X1 U15918 ( .A(n13949), .ZN(n14654) );
  OAI222_X1 U15919 ( .A1(n13955), .A2(n14654), .B1(P2_U3088), .B2(n13951), 
        .C1(n13950), .C2(n13960), .ZN(P2_U3298) );
  AOI21_X1 U15920 ( .B1(n13953), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13952), 
        .ZN(n13954) );
  OAI21_X1 U15921 ( .B1(n13956), .B2(n13955), .A(n13954), .ZN(P2_U3299) );
  OAI222_X1 U15922 ( .A1(n13960), .A2(n13959), .B1(n13955), .B2(n13958), .C1(
        P2_U3088), .C2(n13957), .ZN(P2_U3300) );
  INV_X1 U15923 ( .A(n13961), .ZN(n13963) );
  MUX2_X1 U15924 ( .A(n13963), .B(n13962), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  OAI21_X1 U15925 ( .B1(n13966), .B2(n13965), .A(n13964), .ZN(n13967) );
  NAND2_X1 U15926 ( .A1(n13967), .A2(n14828), .ZN(n13976) );
  INV_X1 U15927 ( .A(n14348), .ZN(n13974) );
  NOR2_X1 U15928 ( .A1(n13968), .A2(n14095), .ZN(n13971) );
  NOR2_X1 U15929 ( .A1(n13969), .A2(n14065), .ZN(n13970) );
  OR2_X1 U15930 ( .A1(n13971), .A2(n13970), .ZN(n14341) );
  INV_X1 U15931 ( .A(n14341), .ZN(n13972) );
  OAI22_X1 U15932 ( .A1(n14121), .A2(n13972), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15574), .ZN(n13973) );
  AOI21_X1 U15933 ( .B1(n14124), .B2(n13974), .A(n13973), .ZN(n13975) );
  OAI211_X1 U15934 ( .C1(n8823), .C2(n14127), .A(n13976), .B(n13975), .ZN(
        P1_U3214) );
  OAI22_X1 U15935 ( .A1(n13978), .A2(n14065), .B1(n13977), .B2(n14095), .ZN(
        n14406) );
  AOI22_X1 U15936 ( .A1(n14406), .A2(n14830), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13979) );
  OAI21_X1 U15937 ( .B1(n14408), .B2(n14836), .A(n13979), .ZN(n13986) );
  NAND3_X1 U15938 ( .A1(n13981), .A2(n13983), .A3(n7505), .ZN(n13984) );
  AOI21_X1 U15939 ( .B1(n13980), .B2(n13984), .A(n14103), .ZN(n13985) );
  AOI211_X1 U15940 ( .C1(n14553), .C2(n6638), .A(n13986), .B(n13985), .ZN(
        n13987) );
  INV_X1 U15941 ( .A(n13987), .ZN(P1_U3216) );
  INV_X1 U15942 ( .A(n14637), .ZN(n14472) );
  INV_X1 U15943 ( .A(n13988), .ZN(n14092) );
  OAI21_X1 U15944 ( .B1(n14092), .B2(n13990), .A(n13989), .ZN(n13992) );
  NAND3_X1 U15945 ( .A1(n13992), .A2(n14828), .A3(n13991), .ZN(n13996) );
  NOR2_X1 U15946 ( .A1(n14047), .A2(n14065), .ZN(n13993) );
  AOI21_X1 U15947 ( .B1(n14139), .B2(n14110), .A(n13993), .ZN(n14576) );
  NAND2_X1 U15948 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14304)
         );
  OAI21_X1 U15949 ( .B1(n14121), .B2(n14576), .A(n14304), .ZN(n13994) );
  AOI21_X1 U15950 ( .B1(n14124), .B2(n14474), .A(n13994), .ZN(n13995) );
  OAI211_X1 U15951 ( .C1(n14472), .C2(n14127), .A(n13996), .B(n13995), .ZN(
        P1_U3219) );
  INV_X1 U15952 ( .A(n13998), .ZN(n14084) );
  AOI21_X1 U15953 ( .B1(n13997), .B2(n13999), .A(n14084), .ZN(n14004) );
  NOR2_X1 U15954 ( .A1(n14836), .A2(n14447), .ZN(n14002) );
  AND2_X1 U15955 ( .A1(n14139), .A2(n14111), .ZN(n14000) );
  AOI21_X1 U15956 ( .B1(n14137), .B2(n14110), .A(n14000), .ZN(n14443) );
  INV_X1 U15957 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15545) );
  OAI22_X1 U15958 ( .A1(n14443), .A2(n14121), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15545), .ZN(n14001) );
  AOI211_X1 U15959 ( .C1(n14632), .C2(n6638), .A(n14002), .B(n14001), .ZN(
        n14003) );
  OAI21_X1 U15960 ( .B1(n14004), .B2(n14103), .A(n14003), .ZN(P1_U3223) );
  AOI21_X1 U15961 ( .B1(n14006), .B2(n14005), .A(n14103), .ZN(n14008) );
  NAND2_X1 U15962 ( .A1(n14008), .A2(n14007), .ZN(n14014) );
  NOR2_X1 U15963 ( .A1(n14836), .A2(n14009), .ZN(n14010) );
  AOI211_X1 U15964 ( .C1(n14830), .C2(n14012), .A(n14011), .B(n14010), .ZN(
        n14013) );
  OAI211_X1 U15965 ( .C1(n7204), .C2(n14127), .A(n14014), .B(n14013), .ZN(
        P1_U3224) );
  AND2_X1 U15966 ( .A1(n14135), .A2(n14111), .ZN(n14015) );
  AOI21_X1 U15967 ( .B1(n14133), .B2(n14110), .A(n14015), .ZN(n14540) );
  INV_X1 U15968 ( .A(n14540), .ZN(n14016) );
  AOI22_X1 U15969 ( .A1(n14830), .A2(n14016), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14017) );
  OAI21_X1 U15970 ( .B1(n14372), .B2(n14836), .A(n14017), .ZN(n14025) );
  INV_X1 U15971 ( .A(n14019), .ZN(n14020) );
  NAND3_X1 U15972 ( .A1(n14018), .A2(n14021), .A3(n14020), .ZN(n14022) );
  AOI21_X1 U15973 ( .B1(n14023), .B2(n14022), .A(n14103), .ZN(n14024) );
  AOI211_X1 U15974 ( .C1(n14619), .C2(n6638), .A(n14025), .B(n14024), .ZN(
        n14026) );
  INV_X1 U15975 ( .A(n14026), .ZN(P1_U3225) );
  INV_X1 U15976 ( .A(n14028), .ZN(n14029) );
  XNOR2_X1 U15977 ( .A(n14027), .B(n14028), .ZN(n14119) );
  NAND2_X1 U15978 ( .A1(n14119), .A2(n14118), .ZN(n14117) );
  OAI21_X1 U15979 ( .B1(n14029), .B2(n14027), .A(n14117), .ZN(n14033) );
  XOR2_X1 U15980 ( .A(n14031), .B(n14030), .Z(n14032) );
  XNOR2_X1 U15981 ( .A(n14033), .B(n14032), .ZN(n14041) );
  NAND2_X1 U15982 ( .A1(n14124), .A2(n14034), .ZN(n14036) );
  OAI211_X1 U15983 ( .C1(n14037), .C2(n14121), .A(n14036), .B(n14035), .ZN(
        n14038) );
  AOI21_X1 U15984 ( .B1(n14039), .B2(n6638), .A(n14038), .ZN(n14040) );
  OAI21_X1 U15985 ( .B1(n14041), .B2(n14103), .A(n14040), .ZN(P1_U3226) );
  XNOR2_X1 U15986 ( .A(n14044), .B(n14043), .ZN(n14045) );
  XNOR2_X1 U15987 ( .A(n14042), .B(n14045), .ZN(n14052) );
  OAI22_X1 U15988 ( .A1(n14047), .A2(n14095), .B1(n14046), .B2(n14065), .ZN(
        n14504) );
  NAND2_X1 U15989 ( .A1(n14830), .A2(n14504), .ZN(n14048) );
  OAI211_X1 U15990 ( .C1(n14836), .C2(n14508), .A(n14049), .B(n14048), .ZN(
        n14050) );
  AOI21_X1 U15991 ( .B1(n14587), .B2(n6638), .A(n14050), .ZN(n14051) );
  OAI21_X1 U15992 ( .B1(n14052), .B2(n14103), .A(n14051), .ZN(P1_U3228) );
  NAND2_X1 U15993 ( .A1(n14136), .A2(n14111), .ZN(n14054) );
  NAND2_X1 U15994 ( .A1(n14134), .A2(n14110), .ZN(n14053) );
  NAND2_X1 U15995 ( .A1(n14054), .A2(n14053), .ZN(n14389) );
  AOI22_X1 U15996 ( .A1(n14830), .A2(n14389), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14055) );
  OAI21_X1 U15997 ( .B1(n14398), .B2(n14836), .A(n14055), .ZN(n14061) );
  INV_X1 U15998 ( .A(n14056), .ZN(n14057) );
  NAND3_X1 U15999 ( .A1(n13980), .A2(n14058), .A3(n14057), .ZN(n14059) );
  AOI21_X1 U16000 ( .B1(n14018), .B2(n14059), .A(n14103), .ZN(n14060) );
  AOI211_X1 U16001 ( .C1(n14623), .C2(n6638), .A(n14061), .B(n14060), .ZN(
        n14062) );
  INV_X1 U16002 ( .A(n14062), .ZN(P1_U3229) );
  XNOR2_X1 U16003 ( .A(n14064), .B(n14063), .ZN(n14070) );
  OAI22_X1 U16004 ( .A1(n14066), .A2(n14095), .B1(n14096), .B2(n14065), .ZN(
        n14458) );
  AOI22_X1 U16005 ( .A1(n14458), .A2(n14830), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14067) );
  OAI21_X1 U16006 ( .B1(n14461), .B2(n14836), .A(n14067), .ZN(n14068) );
  AOI21_X1 U16007 ( .B1(n14570), .B2(n6638), .A(n14068), .ZN(n14069) );
  OAI21_X1 U16008 ( .B1(n14070), .B2(n14103), .A(n14069), .ZN(P1_U3233) );
  OAI211_X1 U16009 ( .C1(n14073), .C2(n14072), .A(n14071), .B(n14828), .ZN(
        n14080) );
  INV_X1 U16010 ( .A(n14074), .ZN(n14078) );
  OAI21_X1 U16011 ( .B1(n14121), .B2(n14076), .A(n14075), .ZN(n14077) );
  AOI21_X1 U16012 ( .B1(n14124), .B2(n14078), .A(n14077), .ZN(n14079) );
  OAI211_X1 U16013 ( .C1(n14081), .C2(n14127), .A(n14080), .B(n14079), .ZN(
        P1_U3234) );
  NOR3_X1 U16014 ( .A1(n14084), .A2(n6898), .A3(n14083), .ZN(n14085) );
  OAI21_X1 U16015 ( .B1(n14085), .B2(n6895), .A(n14828), .ZN(n14090) );
  AND2_X1 U16016 ( .A1(n14136), .A2(n14110), .ZN(n14086) );
  AOI21_X1 U16017 ( .B1(n14138), .B2(n14111), .A(n14086), .ZN(n14425) );
  INV_X1 U16018 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14087) );
  OAI22_X1 U16019 ( .A1(n14425), .A2(n14121), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14087), .ZN(n14088) );
  AOI21_X1 U16020 ( .B1(n14429), .B2(n14124), .A(n14088), .ZN(n14089) );
  OAI211_X1 U16021 ( .C1(n14127), .C2(n14091), .A(n14090), .B(n14089), .ZN(
        P1_U3235) );
  AOI21_X1 U16022 ( .B1(n14094), .B2(n14093), .A(n14092), .ZN(n14104) );
  OR2_X1 U16023 ( .A1(n14096), .A2(n14095), .ZN(n14098) );
  NAND2_X1 U16024 ( .A1(n14142), .A2(n14111), .ZN(n14097) );
  AND2_X1 U16025 ( .A1(n14098), .A2(n14097), .ZN(n14491) );
  NAND2_X1 U16026 ( .A1(n14124), .A2(n14494), .ZN(n14099) );
  NAND2_X1 U16027 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14266)
         );
  OAI211_X1 U16028 ( .C1(n14491), .C2(n14121), .A(n14099), .B(n14266), .ZN(
        n14100) );
  AOI21_X1 U16029 ( .B1(n14583), .B2(n6638), .A(n14100), .ZN(n14102) );
  OAI21_X1 U16030 ( .B1(n14104), .B2(n14103), .A(n14102), .ZN(P1_U3238) );
  OAI21_X1 U16031 ( .B1(n14107), .B2(n14106), .A(n14105), .ZN(n14108) );
  NAND2_X1 U16032 ( .A1(n14108), .A2(n14828), .ZN(n14116) );
  INV_X1 U16033 ( .A(n14109), .ZN(n14357) );
  NAND2_X1 U16034 ( .A1(n14132), .A2(n14110), .ZN(n14113) );
  NAND2_X1 U16035 ( .A1(n14134), .A2(n14111), .ZN(n14112) );
  AND2_X1 U16036 ( .A1(n14113), .A2(n14112), .ZN(n14532) );
  OAI22_X1 U16037 ( .A1(n14121), .A2(n14532), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15531), .ZN(n14114) );
  AOI21_X1 U16038 ( .B1(n14124), .B2(n14357), .A(n14114), .ZN(n14115) );
  OAI211_X1 U16039 ( .C1(n14616), .C2(n14127), .A(n14116), .B(n14115), .ZN(
        P1_U3240) );
  OAI211_X1 U16040 ( .C1(n14119), .C2(n14118), .A(n14117), .B(n14828), .ZN(
        n14126) );
  NAND2_X1 U16041 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14876)
         );
  OAI21_X1 U16042 ( .B1(n14121), .B2(n14120), .A(n14876), .ZN(n14122) );
  AOI21_X1 U16043 ( .B1(n14124), .B2(n14123), .A(n14122), .ZN(n14125) );
  OAI211_X1 U16044 ( .C1(n14128), .C2(n14127), .A(n14126), .B(n14125), .ZN(
        P1_U3241) );
  MUX2_X1 U16045 ( .A(n14308), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14159), .Z(
        P1_U3591) );
  MUX2_X1 U16046 ( .A(n14129), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14159), .Z(
        P1_U3590) );
  MUX2_X1 U16047 ( .A(n14130), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14159), .Z(
        P1_U3589) );
  MUX2_X1 U16048 ( .A(n14131), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14159), .Z(
        P1_U3588) );
  MUX2_X1 U16049 ( .A(n14132), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14159), .Z(
        P1_U3587) );
  MUX2_X1 U16050 ( .A(n14133), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14159), .Z(
        P1_U3586) );
  MUX2_X1 U16051 ( .A(n14134), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14159), .Z(
        P1_U3585) );
  MUX2_X1 U16052 ( .A(n14135), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14159), .Z(
        P1_U3584) );
  MUX2_X1 U16053 ( .A(n14136), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14159), .Z(
        P1_U3583) );
  MUX2_X1 U16054 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14137), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16055 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14138), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16056 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14139), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16057 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14140), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16058 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14141), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16059 ( .A(n14142), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14159), .Z(
        P1_U3577) );
  MUX2_X1 U16060 ( .A(n14143), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14159), .Z(
        P1_U3576) );
  MUX2_X1 U16061 ( .A(n14144), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14159), .Z(
        P1_U3575) );
  MUX2_X1 U16062 ( .A(n14145), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14159), .Z(
        P1_U3574) );
  MUX2_X1 U16063 ( .A(n14146), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14159), .Z(
        P1_U3573) );
  MUX2_X1 U16064 ( .A(n14147), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14159), .Z(
        P1_U3572) );
  MUX2_X1 U16065 ( .A(n14148), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14159), .Z(
        P1_U3571) );
  MUX2_X1 U16066 ( .A(n14149), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14159), .Z(
        P1_U3570) );
  MUX2_X1 U16067 ( .A(n14150), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14159), .Z(
        P1_U3569) );
  MUX2_X1 U16068 ( .A(n14151), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14159), .Z(
        P1_U3568) );
  MUX2_X1 U16069 ( .A(n14152), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14159), .Z(
        P1_U3567) );
  MUX2_X1 U16070 ( .A(n14153), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14159), .Z(
        P1_U3566) );
  MUX2_X1 U16071 ( .A(n14154), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14159), .Z(
        P1_U3565) );
  MUX2_X1 U16072 ( .A(n14155), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14159), .Z(
        P1_U3564) );
  MUX2_X1 U16073 ( .A(n14156), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14159), .Z(
        P1_U3563) );
  MUX2_X1 U16074 ( .A(n14157), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14159), .Z(
        P1_U3562) );
  MUX2_X1 U16075 ( .A(n14158), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14159), .Z(
        P1_U3561) );
  MUX2_X1 U16076 ( .A(n8837), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14159), .Z(
        P1_U3560) );
  OAI211_X1 U16077 ( .C1(n14162), .C2(n14161), .A(n14874), .B(n14160), .ZN(
        n14168) );
  AOI22_X1 U16078 ( .A1(n14255), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14167) );
  NAND2_X1 U16079 ( .A1(n14293), .A2(n14163), .ZN(n14166) );
  OAI211_X1 U16080 ( .C1(n14171), .C2(n14164), .A(n14299), .B(n14182), .ZN(
        n14165) );
  NAND4_X1 U16081 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        P1_U3244) );
  MUX2_X1 U16082 ( .A(n14171), .B(n14170), .S(n6734), .Z(n14173) );
  NAND2_X1 U16083 ( .A1(n14173), .A2(n14172), .ZN(n14174) );
  OAI211_X1 U16084 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14175), .A(n14174), .B(
        P1_U4016), .ZN(n14219) );
  INV_X1 U16085 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14177) );
  INV_X1 U16086 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14176) );
  OAI22_X1 U16087 ( .A1(n14878), .A2(n14177), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14176), .ZN(n14178) );
  AOI21_X1 U16088 ( .B1(n14179), .B2(n14293), .A(n14178), .ZN(n14190) );
  MUX2_X1 U16089 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10033), .S(n14180), .Z(
        n14183) );
  NAND3_X1 U16090 ( .A1(n14183), .A2(n14182), .A3(n14181), .ZN(n14184) );
  NAND3_X1 U16091 ( .A1(n14299), .A2(n14198), .A3(n14184), .ZN(n14189) );
  OAI211_X1 U16092 ( .C1(n14187), .C2(n14186), .A(n14874), .B(n14185), .ZN(
        n14188) );
  NAND4_X1 U16093 ( .A1(n14219), .A2(n14190), .A3(n14189), .A4(n14188), .ZN(
        P1_U3245) );
  OAI211_X1 U16094 ( .C1(n14193), .C2(n14192), .A(n14874), .B(n14191), .ZN(
        n14203) );
  NOR2_X1 U16095 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15555), .ZN(n14194) );
  AOI21_X1 U16096 ( .B1(n14255), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n14194), .ZN(
        n14202) );
  NAND2_X1 U16097 ( .A1(n14293), .A2(n14195), .ZN(n14201) );
  MUX2_X1 U16098 ( .A(n11349), .B(P1_REG2_REG_3__SCAN_IN), .S(n14195), .Z(
        n14197) );
  NAND3_X1 U16099 ( .A1(n14198), .A2(n14197), .A3(n14196), .ZN(n14199) );
  NAND3_X1 U16100 ( .A1(n14299), .A2(n14213), .A3(n14199), .ZN(n14200) );
  NAND4_X1 U16101 ( .A1(n14203), .A2(n14202), .A3(n14201), .A4(n14200), .ZN(
        P1_U3246) );
  INV_X1 U16102 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14205) );
  OAI21_X1 U16103 ( .B1(n14878), .B2(n14205), .A(n14204), .ZN(n14206) );
  AOI21_X1 U16104 ( .B1(n14293), .B2(n14210), .A(n14206), .ZN(n14218) );
  OAI211_X1 U16105 ( .C1(n14209), .C2(n14208), .A(n14874), .B(n14207), .ZN(
        n14217) );
  MUX2_X1 U16106 ( .A(n11329), .B(P1_REG2_REG_4__SCAN_IN), .S(n14210), .Z(
        n14211) );
  NAND3_X1 U16107 ( .A1(n14213), .A2(n14212), .A3(n14211), .ZN(n14214) );
  NAND3_X1 U16108 ( .A1(n14299), .A2(n14215), .A3(n14214), .ZN(n14216) );
  NAND4_X1 U16109 ( .A1(n14219), .A2(n14218), .A3(n14217), .A4(n14216), .ZN(
        P1_U3247) );
  INV_X1 U16110 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14221) );
  OAI21_X1 U16111 ( .B1(n14878), .B2(n14221), .A(n14220), .ZN(n14222) );
  AOI21_X1 U16112 ( .B1(n14293), .B2(n14223), .A(n14222), .ZN(n14233) );
  OAI211_X1 U16113 ( .C1(n14226), .C2(n14225), .A(n14874), .B(n14224), .ZN(
        n14232) );
  OR3_X1 U16114 ( .A1(n14229), .A2(n14228), .A3(n14227), .ZN(n14230) );
  NAND3_X1 U16115 ( .A1(n14299), .A2(n14243), .A3(n14230), .ZN(n14231) );
  NAND3_X1 U16116 ( .A1(n14233), .A2(n14232), .A3(n14231), .ZN(P1_U3249) );
  INV_X1 U16117 ( .A(n14234), .ZN(n14237) );
  NOR2_X1 U16118 ( .A1(n14870), .A2(n14235), .ZN(n14236) );
  AOI211_X1 U16119 ( .C1(n14255), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n14237), .B(
        n14236), .ZN(n14248) );
  OAI211_X1 U16120 ( .C1(n14240), .C2(n14239), .A(n14874), .B(n14238), .ZN(
        n14247) );
  NAND3_X1 U16121 ( .A1(n14243), .A2(n14242), .A3(n14241), .ZN(n14244) );
  NAND3_X1 U16122 ( .A1(n14299), .A2(n14245), .A3(n14244), .ZN(n14246) );
  NAND3_X1 U16123 ( .A1(n14248), .A2(n14247), .A3(n14246), .ZN(P1_U3250) );
  OAI211_X1 U16124 ( .C1(n14251), .C2(n14250), .A(n14249), .B(n14874), .ZN(
        n14265) );
  AND2_X1 U16125 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14254) );
  NOR2_X1 U16126 ( .A1(n14870), .A2(n14252), .ZN(n14253) );
  AOI211_X1 U16127 ( .C1(n14255), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n14254), 
        .B(n14253), .ZN(n14264) );
  MUX2_X1 U16128 ( .A(n10283), .B(P1_REG2_REG_10__SCAN_IN), .S(n14256), .Z(
        n14259) );
  INV_X1 U16129 ( .A(n14257), .ZN(n14258) );
  NAND2_X1 U16130 ( .A1(n14259), .A2(n14258), .ZN(n14261) );
  OAI211_X1 U16131 ( .C1(n14262), .C2(n14261), .A(n14260), .B(n14299), .ZN(
        n14263) );
  NAND3_X1 U16132 ( .A1(n14265), .A2(n14264), .A3(n14263), .ZN(P1_U3253) );
  INV_X1 U16133 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14267) );
  OAI21_X1 U16134 ( .B1(n14878), .B2(n14267), .A(n14266), .ZN(n14268) );
  AOI21_X1 U16135 ( .B1(n14293), .B2(n14289), .A(n14268), .ZN(n14281) );
  INV_X1 U16136 ( .A(n14271), .ZN(n14274) );
  INV_X1 U16137 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14272) );
  INV_X1 U16138 ( .A(n14285), .ZN(n14273) );
  OAI211_X1 U16139 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14274), .A(n14874), 
        .B(n14273), .ZN(n14280) );
  OAI21_X1 U16140 ( .B1(n14277), .B2(n14276), .A(n14275), .ZN(n14288) );
  XNOR2_X1 U16141 ( .A(n14282), .B(n14288), .ZN(n14278) );
  NAND2_X1 U16142 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14278), .ZN(n14291) );
  OAI211_X1 U16143 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14278), .A(n14299), 
        .B(n14291), .ZN(n14279) );
  NAND3_X1 U16144 ( .A1(n14281), .A2(n14280), .A3(n14279), .ZN(P1_U3261) );
  INV_X1 U16145 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14306) );
  NOR2_X1 U16146 ( .A1(n14283), .A2(n14282), .ZN(n14284) );
  XOR2_X1 U16147 ( .A(n14287), .B(n14286), .Z(n14300) );
  NAND2_X1 U16148 ( .A1(n14289), .A2(n14288), .ZN(n14290) );
  NAND2_X1 U16149 ( .A1(n14291), .A2(n14290), .ZN(n14292) );
  XNOR2_X1 U16150 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14292), .ZN(n14297) );
  AOI21_X1 U16151 ( .B1(n14297), .B2(n14299), .A(n14293), .ZN(n14294) );
  OAI21_X1 U16152 ( .B1(n14300), .B2(n14295), .A(n14294), .ZN(n14296) );
  INV_X1 U16153 ( .A(n14296), .ZN(n14303) );
  INV_X1 U16154 ( .A(n14297), .ZN(n14298) );
  AOI22_X1 U16155 ( .A1(n14300), .A2(n14874), .B1(n14299), .B2(n14298), .ZN(
        n14302) );
  MUX2_X1 U16156 ( .A(n14303), .B(n14302), .S(n14301), .Z(n14305) );
  OAI211_X1 U16157 ( .C1(n14306), .C2(n14878), .A(n14305), .B(n14304), .ZN(
        P1_U3262) );
  NAND2_X1 U16158 ( .A1(n14519), .A2(n14911), .ZN(n14311) );
  AND2_X1 U16159 ( .A1(n14308), .A2(n14307), .ZN(n14522) );
  INV_X1 U16160 ( .A(n14522), .ZN(n14309) );
  NOR2_X1 U16161 ( .A1(n6653), .A2(n14309), .ZN(n14315) );
  AOI21_X1 U16162 ( .B1(n6653), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14315), .ZN(
        n14310) );
  OAI211_X1 U16163 ( .C1(n12505), .C2(n14925), .A(n14311), .B(n14310), .ZN(
        P1_U3263) );
  INV_X1 U16164 ( .A(n14313), .ZN(n14610) );
  AOI211_X1 U16165 ( .C1(n14314), .C2(n14313), .A(n14909), .B(n14312), .ZN(
        n14523) );
  NAND2_X1 U16166 ( .A1(n14523), .A2(n14911), .ZN(n14317) );
  AOI21_X1 U16167 ( .B1(n6653), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14315), .ZN(
        n14316) );
  OAI211_X1 U16168 ( .C1(n14610), .C2(n14925), .A(n14317), .B(n14316), .ZN(
        P1_U3264) );
  OAI22_X1 U16169 ( .A1(n14320), .A2(n14319), .B1(n14318), .B2(n14507), .ZN(
        n14323) );
  NOR2_X1 U16170 ( .A1(n14321), .A2(n14925), .ZN(n14322) );
  AOI211_X1 U16171 ( .C1(n6653), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14323), .B(
        n14322), .ZN(n14324) );
  OAI21_X1 U16172 ( .B1(n14325), .B2(n14477), .A(n14324), .ZN(n14326) );
  AOI21_X1 U16173 ( .B1(n14327), .B2(n14843), .A(n14326), .ZN(n14328) );
  OAI21_X1 U16174 ( .B1(n6779), .B2(n6653), .A(n14328), .ZN(P1_U3356) );
  OAI22_X1 U16175 ( .A1(n14923), .A2(n14330), .B1(n14329), .B2(n14507), .ZN(
        n14331) );
  AOI21_X1 U16176 ( .B1(n14332), .B2(n14900), .A(n14331), .ZN(n14333) );
  OAI21_X1 U16177 ( .B1(n14334), .B2(n14477), .A(n14333), .ZN(n14335) );
  AOI21_X1 U16178 ( .B1(n14336), .B2(n14843), .A(n14335), .ZN(n14337) );
  OAI21_X1 U16179 ( .B1(n14338), .B2(n6653), .A(n14337), .ZN(P1_U3265) );
  XNOR2_X1 U16180 ( .A(n14340), .B(n14339), .ZN(n14342) );
  AOI21_X1 U16181 ( .B1(n14342), .B2(n14899), .A(n14341), .ZN(n14527) );
  NAND2_X1 U16182 ( .A1(n14343), .A2(n7242), .ZN(n14344) );
  NAND2_X1 U16183 ( .A1(n14345), .A2(n14344), .ZN(n14525) );
  AND2_X1 U16184 ( .A1(n14351), .A2(n14356), .ZN(n14346) );
  INV_X1 U16185 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14349) );
  OAI22_X1 U16186 ( .A1(n14929), .A2(n14349), .B1(n14348), .B2(n14507), .ZN(
        n14350) );
  AOI21_X1 U16187 ( .B1(n14351), .B2(n14900), .A(n14350), .ZN(n14352) );
  OAI21_X1 U16188 ( .B1(n14526), .B2(n14477), .A(n14352), .ZN(n14353) );
  AOI21_X1 U16189 ( .B1(n14525), .B2(n14395), .A(n14353), .ZN(n14354) );
  OAI21_X1 U16190 ( .B1(n14527), .B2(n6653), .A(n14354), .ZN(P1_U3266) );
  XNOR2_X1 U16191 ( .A(n14355), .B(n14361), .ZN(n14535) );
  OAI211_X1 U16192 ( .C1(n14616), .C2(n14371), .A(n14901), .B(n14356), .ZN(
        n14531) );
  AOI22_X1 U16193 ( .A1(n6653), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14357), 
        .B2(n14910), .ZN(n14360) );
  NAND2_X1 U16194 ( .A1(n14358), .A2(n14900), .ZN(n14359) );
  OAI211_X1 U16195 ( .C1(n14531), .C2(n14477), .A(n14360), .B(n14359), .ZN(
        n14365) );
  XNOR2_X1 U16196 ( .A(n14362), .B(n14361), .ZN(n14363) );
  NAND2_X1 U16197 ( .A1(n14363), .A2(n14899), .ZN(n14533) );
  AOI21_X1 U16198 ( .B1(n14533), .B2(n14532), .A(n6653), .ZN(n14364) );
  AOI211_X1 U16199 ( .C1(n14843), .C2(n14535), .A(n14365), .B(n14364), .ZN(
        n14366) );
  INV_X1 U16200 ( .A(n14366), .ZN(P1_U3267) );
  OAI21_X1 U16201 ( .B1(n14368), .B2(n14376), .A(n14367), .ZN(n14538) );
  INV_X1 U16202 ( .A(n14538), .ZN(n14383) );
  NAND2_X1 U16203 ( .A1(n14619), .A2(n14396), .ZN(n14369) );
  NAND2_X1 U16204 ( .A1(n14369), .A2(n14901), .ZN(n14370) );
  OR2_X1 U16205 ( .A1(n14371), .A2(n14370), .ZN(n14539) );
  INV_X1 U16206 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14373) );
  OAI22_X1 U16207 ( .A1(n14923), .A2(n14373), .B1(n14372), .B2(n14507), .ZN(
        n14374) );
  AOI21_X1 U16208 ( .B1(n14619), .B2(n14900), .A(n14374), .ZN(n14375) );
  OAI21_X1 U16209 ( .B1(n14539), .B2(n14477), .A(n14375), .ZN(n14382) );
  NAND2_X1 U16210 ( .A1(n14377), .A2(n14376), .ZN(n14378) );
  NAND2_X1 U16211 ( .A1(n14379), .A2(n14378), .ZN(n14380) );
  NAND2_X1 U16212 ( .A1(n14380), .A2(n14899), .ZN(n14541) );
  AOI21_X1 U16213 ( .B1(n14541), .B2(n14540), .A(n6653), .ZN(n14381) );
  AOI211_X1 U16214 ( .C1(n14383), .C2(n14843), .A(n14382), .B(n14381), .ZN(
        n14384) );
  INV_X1 U16215 ( .A(n14384), .ZN(P1_U3268) );
  NAND2_X1 U16216 ( .A1(n14386), .A2(n14385), .ZN(n14387) );
  NAND3_X1 U16217 ( .A1(n14388), .A2(n14899), .A3(n14387), .ZN(n14391) );
  INV_X1 U16218 ( .A(n14389), .ZN(n14390) );
  NAND2_X1 U16219 ( .A1(n14391), .A2(n14390), .ZN(n14548) );
  INV_X1 U16220 ( .A(n14548), .ZN(n14404) );
  NAND2_X1 U16221 ( .A1(n14392), .A2(n8863), .ZN(n14393) );
  NAND2_X1 U16222 ( .A1(n14394), .A2(n14393), .ZN(n14546) );
  NAND2_X1 U16223 ( .A1(n14546), .A2(n14395), .ZN(n14403) );
  AOI21_X1 U16224 ( .B1(n14623), .B2(n14413), .A(n14909), .ZN(n14397) );
  AND2_X1 U16225 ( .A1(n14397), .A2(n14396), .ZN(n14547) );
  OAI22_X1 U16226 ( .A1(n14923), .A2(n14399), .B1(n14398), .B2(n14507), .ZN(
        n14401) );
  NOR2_X1 U16227 ( .A1(n7200), .A2(n14925), .ZN(n14400) );
  AOI211_X1 U16228 ( .C1(n14547), .C2(n14911), .A(n14401), .B(n14400), .ZN(
        n14402) );
  OAI211_X1 U16229 ( .C1(n14404), .C2(n6653), .A(n14403), .B(n14402), .ZN(
        P1_U3269) );
  XNOR2_X1 U16230 ( .A(n14405), .B(n14410), .ZN(n14407) );
  AOI21_X1 U16231 ( .B1(n14407), .B2(n14899), .A(n14406), .ZN(n14556) );
  OAI21_X1 U16232 ( .B1(n14408), .B2(n14507), .A(n14556), .ZN(n14418) );
  INV_X1 U16233 ( .A(n14410), .ZN(n14412) );
  OAI21_X1 U16234 ( .B1(n14409), .B2(n14412), .A(n14411), .ZN(n14557) );
  AOI22_X1 U16235 ( .A1(n14553), .A2(n14900), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n6653), .ZN(n14416) );
  AOI21_X1 U16236 ( .B1(n14553), .B2(n14414), .A(n7201), .ZN(n14554) );
  NAND3_X1 U16237 ( .A1(n14554), .A2(n14901), .A3(n14911), .ZN(n14415) );
  OAI211_X1 U16238 ( .C1(n14557), .C2(n14518), .A(n14416), .B(n14415), .ZN(
        n14417) );
  AOI21_X1 U16239 ( .B1(n14923), .B2(n14418), .A(n14417), .ZN(n14419) );
  INV_X1 U16240 ( .A(n14419), .ZN(P1_U3270) );
  NAND2_X1 U16241 ( .A1(n14420), .A2(n14421), .ZN(n14422) );
  NAND2_X1 U16242 ( .A1(n14422), .A2(n14430), .ZN(n14424) );
  NAND2_X1 U16243 ( .A1(n14424), .A2(n14423), .ZN(n14427) );
  INV_X1 U16244 ( .A(n14425), .ZN(n14426) );
  AOI21_X1 U16245 ( .B1(n14427), .B2(n14899), .A(n14426), .ZN(n14561) );
  INV_X1 U16246 ( .A(n14561), .ZN(n14428) );
  AOI21_X1 U16247 ( .B1(n14429), .B2(n14910), .A(n14428), .ZN(n14438) );
  OR2_X1 U16248 ( .A1(n14431), .A2(n14430), .ZN(n14432) );
  NAND2_X1 U16249 ( .A1(n14433), .A2(n14432), .ZN(n14558) );
  XNOR2_X1 U16250 ( .A(n14628), .B(n6877), .ZN(n14434) );
  NAND2_X1 U16251 ( .A1(n14434), .A2(n14901), .ZN(n14560) );
  AOI22_X1 U16252 ( .A1(n14628), .A2(n14900), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n6653), .ZN(n14435) );
  OAI21_X1 U16253 ( .B1(n14560), .B2(n14477), .A(n14435), .ZN(n14436) );
  AOI21_X1 U16254 ( .B1(n14558), .B2(n14843), .A(n14436), .ZN(n14437) );
  OAI21_X1 U16255 ( .B1(n14438), .B2(n6653), .A(n14437), .ZN(P1_U3271) );
  XNOR2_X1 U16256 ( .A(n14439), .B(n14440), .ZN(n14566) );
  OAI211_X1 U16257 ( .C1(n14442), .C2(n14441), .A(n14420), .B(n14899), .ZN(
        n14444) );
  AND2_X1 U16258 ( .A1(n14444), .A2(n14443), .ZN(n14565) );
  INV_X1 U16259 ( .A(n14565), .ZN(n14452) );
  OAI211_X1 U16260 ( .C1(n14446), .C2(n14462), .A(n14901), .B(n14445), .ZN(
        n14564) );
  INV_X1 U16261 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14448) );
  OAI22_X1 U16262 ( .A1(n14929), .A2(n14448), .B1(n14447), .B2(n14507), .ZN(
        n14449) );
  AOI21_X1 U16263 ( .B1(n14632), .B2(n14900), .A(n14449), .ZN(n14450) );
  OAI21_X1 U16264 ( .B1(n14564), .B2(n14477), .A(n14450), .ZN(n14451) );
  AOI21_X1 U16265 ( .B1(n14452), .B2(n14923), .A(n14451), .ZN(n14453) );
  OAI21_X1 U16266 ( .B1(n14518), .B2(n14566), .A(n14453), .ZN(P1_U3272) );
  XNOR2_X1 U16267 ( .A(n14455), .B(n14454), .ZN(n14573) );
  AOI21_X1 U16268 ( .B1(n14457), .B2(n14456), .A(n14921), .ZN(n14460) );
  AOI21_X1 U16269 ( .B1(n14460), .B2(n14459), .A(n14458), .ZN(n14572) );
  OAI21_X1 U16270 ( .B1(n14461), .B2(n14507), .A(n14572), .ZN(n14466) );
  AOI211_X1 U16271 ( .C1(n14570), .C2(n6846), .A(n14909), .B(n14462), .ZN(
        n14569) );
  INV_X1 U16272 ( .A(n14569), .ZN(n14464) );
  AOI22_X1 U16273 ( .A1(n14570), .A2(n14900), .B1(n6653), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14463) );
  OAI21_X1 U16274 ( .B1(n14464), .B2(n14477), .A(n14463), .ZN(n14465) );
  AOI21_X1 U16275 ( .B1(n14466), .B2(n14923), .A(n14465), .ZN(n14467) );
  OAI21_X1 U16276 ( .B1(n14573), .B2(n14518), .A(n14467), .ZN(P1_U3273) );
  NAND2_X1 U16277 ( .A1(n14469), .A2(n14468), .ZN(n14470) );
  NAND2_X1 U16278 ( .A1(n14471), .A2(n14470), .ZN(n14574) );
  XNOR2_X1 U16279 ( .A(n14472), .B(n6845), .ZN(n14473) );
  NAND2_X1 U16280 ( .A1(n14473), .A2(n14901), .ZN(n14575) );
  AOI22_X1 U16281 ( .A1(n6653), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14474), 
        .B2(n14910), .ZN(n14476) );
  NAND2_X1 U16282 ( .A1(n14637), .A2(n14900), .ZN(n14475) );
  OAI211_X1 U16283 ( .C1(n14575), .C2(n14477), .A(n14476), .B(n14475), .ZN(
        n14485) );
  NAND2_X1 U16284 ( .A1(n14478), .A2(n14479), .ZN(n14480) );
  NAND2_X1 U16285 ( .A1(n14480), .A2(n7432), .ZN(n14482) );
  NAND2_X1 U16286 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  NAND2_X1 U16287 ( .A1(n14483), .A2(n14899), .ZN(n14578) );
  AOI21_X1 U16288 ( .B1(n14578), .B2(n14576), .A(n6653), .ZN(n14484) );
  AOI211_X1 U16289 ( .C1(n14843), .C2(n14574), .A(n14485), .B(n14484), .ZN(
        n14486) );
  INV_X1 U16290 ( .A(n14486), .ZN(P1_U3274) );
  XNOR2_X1 U16291 ( .A(n14487), .B(n14488), .ZN(n14585) );
  OAI211_X1 U16292 ( .C1(n14490), .C2(n14489), .A(n14478), .B(n14899), .ZN(
        n14492) );
  NAND2_X1 U16293 ( .A1(n14492), .A2(n14491), .ZN(n14581) );
  INV_X1 U16294 ( .A(n14583), .ZN(n14497) );
  AOI21_X1 U16295 ( .B1(n14511), .B2(n14583), .A(n14909), .ZN(n14493) );
  AND2_X1 U16296 ( .A1(n14493), .A2(n6845), .ZN(n14582) );
  NAND2_X1 U16297 ( .A1(n14582), .A2(n14911), .ZN(n14496) );
  AOI22_X1 U16298 ( .A1(n6653), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14494), 
        .B2(n14910), .ZN(n14495) );
  OAI211_X1 U16299 ( .C1(n14497), .C2(n14925), .A(n14496), .B(n14495), .ZN(
        n14498) );
  AOI21_X1 U16300 ( .B1(n14581), .B2(n14929), .A(n14498), .ZN(n14499) );
  OAI21_X1 U16301 ( .B1(n14500), .B2(n14585), .A(n14499), .ZN(P1_U3275) );
  XNOR2_X1 U16302 ( .A(n14501), .B(n8855), .ZN(n14590) );
  AOI21_X1 U16303 ( .B1(n14503), .B2(n14502), .A(n14921), .ZN(n14506) );
  AOI21_X1 U16304 ( .B1(n14506), .B2(n14505), .A(n14504), .ZN(n14589) );
  OAI21_X1 U16305 ( .B1(n14508), .B2(n14507), .A(n14589), .ZN(n14509) );
  NAND2_X1 U16306 ( .A1(n14509), .A2(n14929), .ZN(n14517) );
  INV_X1 U16307 ( .A(n14510), .ZN(n14513) );
  INV_X1 U16308 ( .A(n14511), .ZN(n14512) );
  AOI211_X1 U16309 ( .C1(n14587), .C2(n14513), .A(n14909), .B(n14512), .ZN(
        n14586) );
  OAI22_X1 U16310 ( .A1(n14514), .A2(n14925), .B1(n14277), .B2(n14929), .ZN(
        n14515) );
  AOI21_X1 U16311 ( .B1(n14586), .B2(n14911), .A(n14515), .ZN(n14516) );
  OAI211_X1 U16312 ( .C1(n14590), .C2(n14518), .A(n14517), .B(n14516), .ZN(
        P1_U3276) );
  INV_X1 U16313 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14520) );
  NOR2_X1 U16314 ( .A1(n14519), .A2(n14522), .ZN(n14604) );
  MUX2_X1 U16315 ( .A(n14520), .B(n14604), .S(n14994), .Z(n14521) );
  OAI21_X1 U16316 ( .B1(n12505), .B2(n14596), .A(n14521), .ZN(P1_U3559) );
  NOR2_X1 U16317 ( .A1(n14523), .A2(n14522), .ZN(n14607) );
  MUX2_X1 U16318 ( .A(n15557), .B(n14607), .S(n14994), .Z(n14524) );
  OAI21_X1 U16319 ( .B1(n14610), .B2(n14596), .A(n14524), .ZN(P1_U3558) );
  NAND2_X1 U16320 ( .A1(n14525), .A2(n14918), .ZN(n14528) );
  NAND3_X1 U16321 ( .A1(n14528), .A2(n14527), .A3(n14526), .ZN(n14611) );
  MUX2_X1 U16322 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14611), .S(n14994), .Z(
        n14529) );
  INV_X1 U16323 ( .A(n14529), .ZN(n14530) );
  OAI21_X1 U16324 ( .B1(n8823), .B2(n14596), .A(n14530), .ZN(P1_U3555) );
  NAND3_X1 U16325 ( .A1(n14533), .A2(n14532), .A3(n14531), .ZN(n14534) );
  AOI21_X1 U16326 ( .B1(n14535), .B2(n14918), .A(n14534), .ZN(n14614) );
  MUX2_X1 U16327 ( .A(n14536), .B(n14614), .S(n14994), .Z(n14537) );
  OAI21_X1 U16328 ( .B1(n14616), .B2(n14596), .A(n14537), .ZN(P1_U3554) );
  OR2_X1 U16329 ( .A1(n14538), .A2(n14895), .ZN(n14543) );
  AND3_X1 U16330 ( .A1(n14541), .A2(n14540), .A3(n14539), .ZN(n14542) );
  NAND2_X1 U16331 ( .A1(n14543), .A2(n14542), .ZN(n14617) );
  MUX2_X1 U16332 ( .A(n14617), .B(P1_REG1_REG_25__SCAN_IN), .S(n14991), .Z(
        n14544) );
  AOI21_X1 U16333 ( .B1(n14602), .B2(n14619), .A(n14544), .ZN(n14545) );
  INV_X1 U16334 ( .A(n14545), .ZN(P1_U3553) );
  NAND2_X1 U16335 ( .A1(n14546), .A2(n14918), .ZN(n14550) );
  NOR2_X1 U16336 ( .A1(n14548), .A2(n14547), .ZN(n14549) );
  NAND2_X1 U16337 ( .A1(n14550), .A2(n14549), .ZN(n14621) );
  MUX2_X1 U16338 ( .A(n14621), .B(P1_REG1_REG_24__SCAN_IN), .S(n14991), .Z(
        n14551) );
  AOI21_X1 U16339 ( .B1(n14602), .B2(n14623), .A(n14551), .ZN(n14552) );
  INV_X1 U16340 ( .A(n14552), .ZN(P1_U3552) );
  AOI22_X1 U16341 ( .A1(n14554), .A2(n14901), .B1(n14553), .B2(n14974), .ZN(
        n14555) );
  OAI211_X1 U16342 ( .C1(n14557), .C2(n14895), .A(n14556), .B(n14555), .ZN(
        n14625) );
  MUX2_X1 U16343 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14625), .S(n14994), .Z(
        P1_U3551) );
  NAND2_X1 U16344 ( .A1(n14558), .A2(n14918), .ZN(n14559) );
  NAND3_X1 U16345 ( .A1(n14561), .A2(n14560), .A3(n14559), .ZN(n14626) );
  MUX2_X1 U16346 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14626), .S(n14994), .Z(
        n14562) );
  AOI21_X1 U16347 ( .B1(n14602), .B2(n14628), .A(n14562), .ZN(n14563) );
  INV_X1 U16348 ( .A(n14563), .ZN(P1_U3550) );
  OAI211_X1 U16349 ( .C1(n14566), .C2(n14895), .A(n14565), .B(n14564), .ZN(
        n14630) );
  MUX2_X1 U16350 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14630), .S(n14994), .Z(
        n14567) );
  AOI21_X1 U16351 ( .B1(n14602), .B2(n14632), .A(n14567), .ZN(n14568) );
  INV_X1 U16352 ( .A(n14568), .ZN(P1_U3549) );
  AOI21_X1 U16353 ( .B1(n14570), .B2(n14974), .A(n14569), .ZN(n14571) );
  OAI211_X1 U16354 ( .C1(n14573), .C2(n14895), .A(n14572), .B(n14571), .ZN(
        n14634) );
  MUX2_X1 U16355 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14634), .S(n14994), .Z(
        P1_U3548) );
  NAND2_X1 U16356 ( .A1(n14574), .A2(n14918), .ZN(n14577) );
  NAND4_X1 U16357 ( .A1(n14578), .A2(n14577), .A3(n14576), .A4(n14575), .ZN(
        n14635) );
  MUX2_X1 U16358 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14635), .S(n14994), .Z(
        n14579) );
  AOI21_X1 U16359 ( .B1(n14602), .B2(n14637), .A(n14579), .ZN(n14580) );
  INV_X1 U16360 ( .A(n14580), .ZN(P1_U3547) );
  AOI211_X1 U16361 ( .C1(n14583), .C2(n14974), .A(n14582), .B(n14581), .ZN(
        n14584) );
  OAI21_X1 U16362 ( .B1(n14895), .B2(n14585), .A(n14584), .ZN(n14639) );
  MUX2_X1 U16363 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14639), .S(n14994), .Z(
        P1_U3546) );
  AOI21_X1 U16364 ( .B1(n14587), .B2(n14974), .A(n14586), .ZN(n14588) );
  OAI211_X1 U16365 ( .C1(n14895), .C2(n14590), .A(n14589), .B(n14588), .ZN(
        n14640) );
  MUX2_X1 U16366 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14640), .S(n14994), .Z(
        P1_U3545) );
  INV_X1 U16367 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14594) );
  AOI211_X1 U16368 ( .C1(n14918), .C2(n14593), .A(n14592), .B(n14591), .ZN(
        n14641) );
  MUX2_X1 U16369 ( .A(n14594), .B(n14641), .S(n14994), .Z(n14595) );
  OAI21_X1 U16370 ( .B1(n14644), .B2(n14596), .A(n14595), .ZN(P1_U3544) );
  AND2_X1 U16371 ( .A1(n14597), .A2(n14918), .ZN(n14600) );
  MUX2_X1 U16372 ( .A(n14645), .B(P1_REG1_REG_15__SCAN_IN), .S(n14991), .Z(
        n14601) );
  AOI21_X1 U16373 ( .B1(n14602), .B2(n14647), .A(n14601), .ZN(n14603) );
  INV_X1 U16374 ( .A(n14603), .ZN(P1_U3543) );
  MUX2_X1 U16375 ( .A(n14605), .B(n14604), .S(n14987), .Z(n14606) );
  OAI21_X1 U16376 ( .B1(n12505), .B2(n14643), .A(n14606), .ZN(P1_U3527) );
  INV_X1 U16377 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14608) );
  MUX2_X1 U16378 ( .A(n14608), .B(n14607), .S(n14987), .Z(n14609) );
  OAI21_X1 U16379 ( .B1(n14610), .B2(n14643), .A(n14609), .ZN(P1_U3526) );
  MUX2_X1 U16380 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14611), .S(n14987), .Z(
        n14612) );
  INV_X1 U16381 ( .A(n14612), .ZN(n14613) );
  OAI21_X1 U16382 ( .B1(n8823), .B2(n14643), .A(n14613), .ZN(P1_U3523) );
  MUX2_X1 U16383 ( .A(n15558), .B(n14614), .S(n14987), .Z(n14615) );
  OAI21_X1 U16384 ( .B1(n14616), .B2(n14643), .A(n14615), .ZN(P1_U3522) );
  MUX2_X1 U16385 ( .A(n14617), .B(P1_REG0_REG_25__SCAN_IN), .S(n14985), .Z(
        n14618) );
  AOI21_X1 U16386 ( .B1(n14648), .B2(n14619), .A(n14618), .ZN(n14620) );
  INV_X1 U16387 ( .A(n14620), .ZN(P1_U3521) );
  MUX2_X1 U16388 ( .A(n14621), .B(P1_REG0_REG_24__SCAN_IN), .S(n14985), .Z(
        n14622) );
  AOI21_X1 U16389 ( .B1(n14648), .B2(n14623), .A(n14622), .ZN(n14624) );
  INV_X1 U16390 ( .A(n14624), .ZN(P1_U3520) );
  MUX2_X1 U16391 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14625), .S(n14987), .Z(
        P1_U3519) );
  MUX2_X1 U16392 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14626), .S(n14987), .Z(
        n14627) );
  AOI21_X1 U16393 ( .B1(n14648), .B2(n14628), .A(n14627), .ZN(n14629) );
  INV_X1 U16394 ( .A(n14629), .ZN(P1_U3518) );
  MUX2_X1 U16395 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14630), .S(n14987), .Z(
        n14631) );
  AOI21_X1 U16396 ( .B1(n14648), .B2(n14632), .A(n14631), .ZN(n14633) );
  INV_X1 U16397 ( .A(n14633), .ZN(P1_U3517) );
  MUX2_X1 U16398 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14634), .S(n14987), .Z(
        P1_U3516) );
  MUX2_X1 U16399 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14635), .S(n14987), .Z(
        n14636) );
  AOI21_X1 U16400 ( .B1(n14648), .B2(n14637), .A(n14636), .ZN(n14638) );
  INV_X1 U16401 ( .A(n14638), .ZN(P1_U3515) );
  MUX2_X1 U16402 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14639), .S(n14987), .Z(
        P1_U3513) );
  MUX2_X1 U16403 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14640), .S(n14987), .Z(
        P1_U3510) );
  MUX2_X1 U16404 ( .A(n15640), .B(n14641), .S(n14987), .Z(n14642) );
  OAI21_X1 U16405 ( .B1(n14644), .B2(n14643), .A(n14642), .ZN(P1_U3507) );
  MUX2_X1 U16406 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14645), .S(n14987), .Z(
        n14646) );
  AOI21_X1 U16407 ( .B1(n14648), .B2(n14647), .A(n14646), .ZN(n14649) );
  INV_X1 U16408 ( .A(n14649), .ZN(P1_U3504) );
  NOR4_X1 U16409 ( .A1(n6697), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8411), .A4(
        P1_U3086), .ZN(n14650) );
  AOI21_X1 U16410 ( .B1(n14651), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14650), 
        .ZN(n14652) );
  OAI21_X1 U16411 ( .B1(n14653), .B2(n6656), .A(n14652), .ZN(P1_U3324) );
  OAI222_X1 U16412 ( .A1(n12562), .A2(n14656), .B1(P1_U3086), .B2(n14655), 
        .C1(n6656), .C2(n14654), .ZN(P1_U3326) );
  MUX2_X1 U16413 ( .A(n12297), .B(n14657), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16414 ( .A(n14658), .ZN(n14659) );
  MUX2_X1 U16415 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14659), .S(P1_U3086), .Z(
        P1_U3355) );
  INV_X1 U16416 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14678) );
  XOR2_X1 U16417 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(n14678), .Z(n14730) );
  AND2_X1 U16418 ( .A1(n14725), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n14676) );
  INV_X1 U16419 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14675) );
  XOR2_X1 U16420 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n14715) );
  XOR2_X1 U16421 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n10030), .Z(n14680) );
  AOI22_X1 U16422 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n10417), .B1(
        P3_ADDR_REG_2__SCAN_IN), .B2(n14177), .ZN(n14684) );
  NAND2_X1 U16423 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14663), .ZN(n14664) );
  NAND2_X1 U16424 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14665), .ZN(n14666) );
  NAND2_X1 U16425 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14667), .ZN(n14669) );
  INV_X1 U16426 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14699) );
  OR2_X1 U16427 ( .A1(n14221), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14670) );
  INV_X1 U16428 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15575) );
  NAND2_X1 U16429 ( .A1(n14671), .A2(n15575), .ZN(n14672) );
  NOR2_X1 U16430 ( .A1(n14715), .A2(n14714), .ZN(n14674) );
  NAND2_X1 U16431 ( .A1(n14730), .A2(n14731), .ZN(n14677) );
  INV_X1 U16432 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U16433 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .B1(n15483), .B2(n15460), .ZN(n14679) );
  XOR2_X1 U16434 ( .A(n14735), .B(n14679), .Z(n14853) );
  XOR2_X1 U16435 ( .A(n14681), .B(n14680), .Z(n14713) );
  XNOR2_X1 U16436 ( .A(n14205), .B(n14682), .ZN(n14695) );
  XOR2_X1 U16437 ( .A(n14695), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15703) );
  INV_X1 U16438 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14773) );
  XNOR2_X1 U16439 ( .A(n14684), .B(n14683), .ZN(n14692) );
  NAND2_X1 U16440 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14688), .ZN(n14690) );
  AOI21_X1 U16441 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14687), .A(n14686), .ZN(
        n15702) );
  NOR2_X1 U16442 ( .A1(n15702), .A2(n9979), .ZN(n15713) );
  NAND2_X1 U16443 ( .A1(n14690), .A2(n14689), .ZN(n14691) );
  NAND2_X1 U16444 ( .A1(n14692), .A2(n14691), .ZN(n14770) );
  NOR2_X1 U16445 ( .A1(n14692), .A2(n14691), .ZN(n14771) );
  AOI21_X1 U16446 ( .B1(n14773), .B2(n14770), .A(n14771), .ZN(n15710) );
  XNOR2_X1 U16447 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14693), .ZN(n15709) );
  NAND2_X1 U16448 ( .A1(n15710), .A2(n15709), .ZN(n14694) );
  NOR2_X1 U16449 ( .A1(n15710), .A2(n15709), .ZN(n15708) );
  AOI21_X1 U16450 ( .B1(n9999), .B2(n14694), .A(n15708), .ZN(n15704) );
  NAND2_X1 U16451 ( .A1(n15703), .A2(n15704), .ZN(n14697) );
  NAND2_X1 U16452 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14695), .ZN(n14696) );
  XNOR2_X1 U16453 ( .A(n14699), .B(n14698), .ZN(n14700) );
  INV_X1 U16454 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14702) );
  XOR2_X1 U16455 ( .A(n14221), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14704) );
  XNOR2_X1 U16456 ( .A(n14704), .B(n14703), .ZN(n14774) );
  NAND2_X1 U16457 ( .A1(n14775), .A2(n14774), .ZN(n14707) );
  NAND2_X1 U16458 ( .A1(n14705), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14706) );
  NAND2_X1 U16459 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14709), .ZN(n14712) );
  XOR2_X1 U16460 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14710), .Z(n15706) );
  NAND2_X1 U16461 ( .A1(n15707), .A2(n15706), .ZN(n14711) );
  XNOR2_X1 U16462 ( .A(n14715), .B(n14714), .ZN(n14716) );
  NAND2_X1 U16463 ( .A1(n14718), .A2(n14716), .ZN(n14720) );
  NAND2_X1 U16464 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n14777), .ZN(n14719) );
  NAND2_X1 U16465 ( .A1(n14722), .A2(n14721), .ZN(n14723) );
  XOR2_X1 U16466 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14723), .Z(n14724) );
  XOR2_X1 U16467 ( .A(n14725), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n14727) );
  XOR2_X1 U16468 ( .A(n14727), .B(n14726), .Z(n14849) );
  NAND2_X1 U16469 ( .A1(n14848), .A2(n14849), .ZN(n14728) );
  NOR2_X1 U16470 ( .A1(n14848), .A2(n14849), .ZN(n14847) );
  XNOR2_X1 U16471 ( .A(n14731), .B(n14730), .ZN(n14733) );
  XOR2_X1 U16472 ( .A(n14739), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n14736) );
  NAND2_X1 U16473 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15460), .ZN(n14734) );
  XOR2_X1 U16474 ( .A(n14736), .B(n14741), .Z(n14737) );
  NOR2_X1 U16475 ( .A1(n14738), .A2(n14737), .ZN(n14857) );
  OR2_X1 U16476 ( .A1(n14739), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n14740) );
  INV_X1 U16477 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14879) );
  XNOR2_X1 U16478 ( .A(n14879), .B(P3_ADDR_REG_15__SCAN_IN), .ZN(n14742) );
  XOR2_X1 U16479 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n14750), .Z(n14745) );
  XOR2_X1 U16480 ( .A(n14745), .B(n14749), .Z(n14746) );
  NOR2_X1 U16481 ( .A1(n14747), .A2(n14746), .ZN(n14863) );
  XNOR2_X1 U16482 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14752), .ZN(n14781) );
  INV_X1 U16483 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U16484 ( .A1(n14751), .A2(n11904), .ZN(n14754) );
  NAND2_X1 U16485 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14752), .ZN(n14753) );
  NAND2_X1 U16486 ( .A1(n14754), .A2(n14753), .ZN(n14757) );
  INV_X1 U16487 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14760) );
  NOR2_X1 U16488 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14760), .ZN(n14755) );
  AOI21_X1 U16489 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14760), .A(n14755), 
        .ZN(n14758) );
  XNOR2_X1 U16490 ( .A(n14757), .B(n14758), .ZN(n14756) );
  NAND2_X1 U16491 ( .A1(n14758), .A2(n14757), .ZN(n14759) );
  OAI21_X1 U16492 ( .B1(n14760), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14759), 
        .ZN(n14766) );
  INV_X1 U16493 ( .A(n14761), .ZN(n14763) );
  NAND2_X1 U16494 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14762) );
  NAND2_X1 U16495 ( .A1(n14763), .A2(n14762), .ZN(n14764) );
  XNOR2_X1 U16496 ( .A(n14764), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n14765) );
  INV_X1 U16497 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15112) );
  XOR2_X1 U16498 ( .A(n15112), .B(n14767), .Z(SUB_1596_U62) );
  AOI21_X1 U16499 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14768) );
  OAI21_X1 U16500 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14768), 
        .ZN(U28) );
  AOI21_X1 U16501 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14769) );
  OAI21_X1 U16502 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14769), 
        .ZN(U29) );
  INV_X1 U16503 ( .A(n14770), .ZN(n14772) );
  AOI222_X1 U16504 ( .A1(n14773), .A2(n14772), .B1(n14773), .B2(n14771), .C1(
        n15710), .C2(n14770), .ZN(SUB_1596_U61) );
  XOR2_X1 U16505 ( .A(n14775), .B(n14774), .Z(SUB_1596_U57) );
  XNOR2_X1 U16506 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14776), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16507 ( .A(n14777), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  XNOR2_X1 U16508 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14778), .ZN(SUB_1596_U70)
         );
  OAI21_X1 U16509 ( .B1(n14781), .B2(n14780), .A(n14779), .ZN(n14783) );
  XOR2_X1 U16510 ( .A(n14783), .B(n14782), .Z(SUB_1596_U63) );
  NOR2_X1 U16511 ( .A1(n14784), .A2(n15295), .ZN(n14786) );
  AOI211_X1 U16512 ( .C1(n15298), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        n14803) );
  AOI22_X1 U16513 ( .A1(n15699), .A2(n14803), .B1(n14788), .B2(n15696), .ZN(
        P3_U3473) );
  NOR2_X1 U16514 ( .A1(n14789), .A2(n15295), .ZN(n14791) );
  AOI211_X1 U16515 ( .C1(n14792), .C2(n15298), .A(n14791), .B(n14790), .ZN(
        n14805) );
  AOI22_X1 U16516 ( .A1(n15699), .A2(n14805), .B1(n15669), .B2(n15696), .ZN(
        P3_U3472) );
  NAND2_X1 U16517 ( .A1(n14793), .A2(n15298), .ZN(n14796) );
  NAND2_X1 U16518 ( .A1(n14794), .A2(n15302), .ZN(n14795) );
  AND3_X1 U16519 ( .A1(n14797), .A2(n14796), .A3(n14795), .ZN(n14807) );
  AOI22_X1 U16520 ( .A1(n15699), .A2(n14807), .B1(n7895), .B2(n15696), .ZN(
        P3_U3471) );
  NAND2_X1 U16521 ( .A1(n14798), .A2(n15298), .ZN(n14801) );
  NAND2_X1 U16522 ( .A1(n14799), .A2(n15302), .ZN(n14800) );
  AND3_X1 U16523 ( .A1(n14802), .A2(n14801), .A3(n14800), .ZN(n14809) );
  AOI22_X1 U16524 ( .A1(n15699), .A2(n14809), .B1(n7879), .B2(n15696), .ZN(
        P3_U3470) );
  AOI22_X1 U16525 ( .A1(n15309), .A2(n14803), .B1(n7952), .B2(n15307), .ZN(
        P3_U3432) );
  INV_X1 U16526 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14804) );
  AOI22_X1 U16527 ( .A1(n15309), .A2(n14805), .B1(n14804), .B2(n15307), .ZN(
        P3_U3429) );
  INV_X1 U16528 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14806) );
  AOI22_X1 U16529 ( .A1(n15309), .A2(n14807), .B1(n14806), .B2(n15307), .ZN(
        P3_U3426) );
  INV_X1 U16530 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14808) );
  AOI22_X1 U16531 ( .A1(n15309), .A2(n14809), .B1(n14808), .B2(n15307), .ZN(
        P3_U3423) );
  INV_X1 U16532 ( .A(n15187), .ZN(n15178) );
  OAI21_X1 U16533 ( .B1(n14811), .B2(n15215), .A(n14810), .ZN(n14813) );
  AOI211_X1 U16534 ( .C1(n15178), .C2(n14814), .A(n14813), .B(n14812), .ZN(
        n14821) );
  AOI22_X1 U16535 ( .A1(n15233), .A2(n14821), .B1(n11439), .B2(n15231), .ZN(
        P2_U3512) );
  INV_X1 U16536 ( .A(n14815), .ZN(n14818) );
  OAI211_X1 U16537 ( .C1(n14818), .C2(n15215), .A(n14817), .B(n14816), .ZN(
        n14819) );
  AOI21_X1 U16538 ( .B1(n14820), .B2(n15178), .A(n14819), .ZN(n14823) );
  AOI22_X1 U16539 ( .A1(n15233), .A2(n14823), .B1(n9187), .B2(n15231), .ZN(
        P2_U3511) );
  AOI22_X1 U16540 ( .A1(n15212), .A2(n14821), .B1(n9210), .B2(n15222), .ZN(
        P2_U3469) );
  INV_X1 U16541 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14822) );
  AOI22_X1 U16542 ( .A1(n15212), .A2(n14823), .B1(n14822), .B2(n15222), .ZN(
        P2_U3466) );
  AND2_X1 U16543 ( .A1(n14071), .A2(n14824), .ZN(n14827) );
  OAI21_X1 U16544 ( .B1(n14827), .B2(n14826), .A(n14825), .ZN(n14829) );
  AOI222_X1 U16545 ( .A1(n6638), .A2(n14832), .B1(n14831), .B2(n14830), .C1(
        n14829), .C2(n14828), .ZN(n14834) );
  OAI211_X1 U16546 ( .C1(n14836), .C2(n14835), .A(n14834), .B(n14833), .ZN(
        P1_U3215) );
  NAND2_X1 U16547 ( .A1(n14837), .A2(n14911), .ZN(n14840) );
  AOI22_X1 U16548 ( .A1(n6653), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n14838), 
        .B2(n14910), .ZN(n14839) );
  OAI211_X1 U16549 ( .C1(n14841), .C2(n14925), .A(n14840), .B(n14839), .ZN(
        n14842) );
  AOI21_X1 U16550 ( .B1(n14844), .B2(n14843), .A(n14842), .ZN(n14845) );
  OAI21_X1 U16551 ( .B1(n6653), .B2(n14846), .A(n14845), .ZN(P1_U3282) );
  AOI21_X1 U16552 ( .B1(n14849), .B2(n14848), .A(n14847), .ZN(n14850) );
  XOR2_X1 U16553 ( .A(n14850), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  XOR2_X1 U16554 ( .A(n10831), .B(n14851), .Z(SUB_1596_U68) );
  AOI21_X1 U16555 ( .B1(n14854), .B2(n14853), .A(n14852), .ZN(n14855) );
  XOR2_X1 U16556 ( .A(n14855), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  NOR2_X1 U16557 ( .A1(n14857), .A2(n14856), .ZN(n14858) );
  XOR2_X1 U16558 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n14858), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16559 ( .A1(n14860), .A2(n14859), .ZN(n14861) );
  XOR2_X1 U16560 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14861), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16561 ( .A1(n14863), .A2(n14862), .ZN(n14864) );
  XOR2_X1 U16562 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14864), .Z(SUB_1596_U64)
         );
  OAI21_X1 U16563 ( .B1(n14867), .B2(n14866), .A(n14865), .ZN(n14875) );
  AOI21_X1 U16564 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14869), .A(n14868), 
        .ZN(n14872) );
  OAI22_X1 U16565 ( .A1(n14872), .A2(n14871), .B1(n6966), .B2(n14870), .ZN(
        n14873) );
  AOI21_X1 U16566 ( .B1(n14875), .B2(n14874), .A(n14873), .ZN(n14877) );
  OAI211_X1 U16567 ( .C1(n14879), .C2(n14878), .A(n14877), .B(n14876), .ZN(
        P1_U3258) );
  NAND2_X1 U16568 ( .A1(n14880), .A2(n14911), .ZN(n14884) );
  INV_X1 U16569 ( .A(n14881), .ZN(n14882) );
  AOI22_X1 U16570 ( .A1(n6653), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n14882), .B2(
        n14910), .ZN(n14883) );
  OAI211_X1 U16571 ( .C1(n14885), .C2(n14925), .A(n14884), .B(n14883), .ZN(
        n14886) );
  INV_X1 U16572 ( .A(n14886), .ZN(n14887) );
  OAI21_X1 U16573 ( .B1(n6653), .B2(n14888), .A(n14887), .ZN(P1_U3284) );
  OAI21_X1 U16574 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n14898) );
  INV_X1 U16575 ( .A(n14892), .ZN(n14897) );
  NOR2_X1 U16576 ( .A1(n7649), .A2(n14895), .ZN(n14896) );
  AOI211_X1 U16577 ( .C1(n14899), .C2(n14898), .A(n14897), .B(n14896), .ZN(
        n14970) );
  AOI222_X1 U16578 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n6653), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14910), .C1(n14969), .C2(n14900), .ZN(
        n14906) );
  NAND2_X1 U16579 ( .A1(n14907), .A2(n14969), .ZN(n14902) );
  NAND2_X1 U16580 ( .A1(n14902), .A2(n14901), .ZN(n14903) );
  NOR2_X1 U16581 ( .A1(n14904), .A2(n14903), .ZN(n14968) );
  NAND2_X1 U16582 ( .A1(n14968), .A2(n14911), .ZN(n14905) );
  OAI211_X1 U16583 ( .C1(n6653), .C2(n14970), .A(n14906), .B(n14905), .ZN(
        P1_U3291) );
  OAI21_X1 U16584 ( .B1(n14964), .B2(n14908), .A(n14907), .ZN(n14912) );
  NOR2_X1 U16585 ( .A1(n14912), .A2(n14909), .ZN(n14962) );
  AOI22_X1 U16586 ( .A1(n14911), .A2(n14962), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14910), .ZN(n14928) );
  XNOR2_X1 U16587 ( .A(n8436), .B(n14912), .ZN(n14913) );
  MUX2_X1 U16588 ( .A(n14917), .B(n14913), .S(n8838), .Z(n14922) );
  INV_X1 U16589 ( .A(n14914), .ZN(n14920) );
  INV_X1 U16590 ( .A(n14915), .ZN(n14916) );
  NAND2_X1 U16591 ( .A1(n7643), .A2(n14918), .ZN(n14919) );
  OAI211_X1 U16592 ( .C1(n14922), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        n14965) );
  NAND2_X1 U16593 ( .A1(n14923), .A2(n14965), .ZN(n14924) );
  OAI21_X1 U16594 ( .B1(n14925), .B2(n14964), .A(n14924), .ZN(n14926) );
  INV_X1 U16595 ( .A(n14926), .ZN(n14927) );
  OAI211_X1 U16596 ( .C1(n10034), .C2(n14929), .A(n14928), .B(n14927), .ZN(
        P1_U3292) );
  INV_X1 U16597 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14930) );
  NOR2_X1 U16598 ( .A1(n14959), .A2(n14930), .ZN(P1_U3294) );
  INV_X1 U16599 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14931) );
  NOR2_X1 U16600 ( .A1(n14959), .A2(n14931), .ZN(P1_U3295) );
  INV_X1 U16601 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14932) );
  NOR2_X1 U16602 ( .A1(n14959), .A2(n14932), .ZN(P1_U3296) );
  INV_X1 U16603 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14933) );
  NOR2_X1 U16604 ( .A1(n14943), .A2(n14933), .ZN(P1_U3297) );
  INV_X1 U16605 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14934) );
  NOR2_X1 U16606 ( .A1(n14943), .A2(n14934), .ZN(P1_U3298) );
  INV_X1 U16607 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15512) );
  NOR2_X1 U16608 ( .A1(n14943), .A2(n15512), .ZN(P1_U3299) );
  INV_X1 U16609 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14935) );
  NOR2_X1 U16610 ( .A1(n14943), .A2(n14935), .ZN(P1_U3300) );
  INV_X1 U16611 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14936) );
  NOR2_X1 U16612 ( .A1(n14943), .A2(n14936), .ZN(P1_U3301) );
  INV_X1 U16613 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14937) );
  NOR2_X1 U16614 ( .A1(n14943), .A2(n14937), .ZN(P1_U3302) );
  INV_X1 U16615 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14938) );
  NOR2_X1 U16616 ( .A1(n14943), .A2(n14938), .ZN(P1_U3303) );
  INV_X1 U16617 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14939) );
  NOR2_X1 U16618 ( .A1(n14943), .A2(n14939), .ZN(P1_U3304) );
  INV_X1 U16619 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15439) );
  NOR2_X1 U16620 ( .A1(n14943), .A2(n15439), .ZN(P1_U3305) );
  INV_X1 U16621 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14940) );
  NOR2_X1 U16622 ( .A1(n14943), .A2(n14940), .ZN(P1_U3306) );
  INV_X1 U16623 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14941) );
  NOR2_X1 U16624 ( .A1(n14943), .A2(n14941), .ZN(P1_U3307) );
  INV_X1 U16625 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14942) );
  NOR2_X1 U16626 ( .A1(n14943), .A2(n14942), .ZN(P1_U3308) );
  INV_X1 U16627 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14944) );
  NOR2_X1 U16628 ( .A1(n14959), .A2(n14944), .ZN(P1_U3309) );
  INV_X1 U16629 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14945) );
  NOR2_X1 U16630 ( .A1(n14959), .A2(n14945), .ZN(P1_U3310) );
  INV_X1 U16631 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14946) );
  NOR2_X1 U16632 ( .A1(n14959), .A2(n14946), .ZN(P1_U3311) );
  INV_X1 U16633 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14947) );
  NOR2_X1 U16634 ( .A1(n14959), .A2(n14947), .ZN(P1_U3312) );
  INV_X1 U16635 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14948) );
  NOR2_X1 U16636 ( .A1(n14959), .A2(n14948), .ZN(P1_U3313) );
  INV_X1 U16637 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14949) );
  NOR2_X1 U16638 ( .A1(n14959), .A2(n14949), .ZN(P1_U3314) );
  INV_X1 U16639 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14950) );
  NOR2_X1 U16640 ( .A1(n14959), .A2(n14950), .ZN(P1_U3315) );
  INV_X1 U16641 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14951) );
  NOR2_X1 U16642 ( .A1(n14959), .A2(n14951), .ZN(P1_U3316) );
  INV_X1 U16643 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14952) );
  NOR2_X1 U16644 ( .A1(n14959), .A2(n14952), .ZN(P1_U3317) );
  INV_X1 U16645 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14953) );
  NOR2_X1 U16646 ( .A1(n14959), .A2(n14953), .ZN(P1_U3318) );
  INV_X1 U16647 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14954) );
  NOR2_X1 U16648 ( .A1(n14959), .A2(n14954), .ZN(P1_U3319) );
  INV_X1 U16649 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14955) );
  NOR2_X1 U16650 ( .A1(n14959), .A2(n14955), .ZN(P1_U3320) );
  INV_X1 U16651 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14956) );
  NOR2_X1 U16652 ( .A1(n14959), .A2(n14956), .ZN(P1_U3321) );
  INV_X1 U16653 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14957) );
  NOR2_X1 U16654 ( .A1(n14959), .A2(n14957), .ZN(P1_U3322) );
  INV_X1 U16655 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14958) );
  NOR2_X1 U16656 ( .A1(n14959), .A2(n14958), .ZN(P1_U3323) );
  INV_X1 U16657 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14960) );
  AOI22_X1 U16658 ( .A1(n14987), .A2(n14961), .B1(n14960), .B2(n14985), .ZN(
        P1_U3459) );
  INV_X1 U16659 ( .A(n14962), .ZN(n14963) );
  OAI21_X1 U16660 ( .B1(n14964), .B2(n14982), .A(n14963), .ZN(n14966) );
  NOR2_X1 U16661 ( .A1(n14966), .A2(n14965), .ZN(n14989) );
  INV_X1 U16662 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14967) );
  AOI22_X1 U16663 ( .A1(n14987), .A2(n14989), .B1(n14967), .B2(n14985), .ZN(
        P1_U3462) );
  AOI21_X1 U16664 ( .B1(n14969), .B2(n14974), .A(n14968), .ZN(n14971) );
  INV_X1 U16665 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U16666 ( .A1(n14987), .A2(n7661), .B1(n14972), .B2(n14985), .ZN(
        P1_U3465) );
  AOI21_X1 U16667 ( .B1(n14975), .B2(n14974), .A(n14973), .ZN(n14977) );
  INV_X1 U16668 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U16669 ( .A1(n14987), .A2(n7646), .B1(n14978), .B2(n14985), .ZN(
        P1_U3468) );
  INV_X1 U16670 ( .A(n14979), .ZN(n14980) );
  OAI211_X1 U16671 ( .C1(n7192), .C2(n14982), .A(n14981), .B(n14980), .ZN(
        n14983) );
  AOI21_X1 U16672 ( .B1(n14918), .B2(n14984), .A(n14983), .ZN(n14993) );
  INV_X1 U16673 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14986) );
  AOI22_X1 U16674 ( .A1(n14987), .A2(n14993), .B1(n14986), .B2(n14985), .ZN(
        P1_U3483) );
  AOI22_X1 U16675 ( .A1(n14994), .A2(n14989), .B1(n14988), .B2(n14991), .ZN(
        P1_U3529) );
  AOI22_X1 U16676 ( .A1(n14994), .A2(n7661), .B1(n14990), .B2(n14991), .ZN(
        P1_U3530) );
  AOI22_X1 U16677 ( .A1(n14994), .A2(n7646), .B1(n15637), .B2(n14991), .ZN(
        P1_U3531) );
  AOI22_X1 U16678 ( .A1(n14994), .A2(n14993), .B1(n14992), .B2(n14991), .ZN(
        P1_U3536) );
  NOR2_X1 U16679 ( .A1(n15083), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI22_X1 U16680 ( .A1(n14997), .A2(n14996), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14995), .ZN(n15003) );
  AOI211_X1 U16681 ( .C1(n15001), .C2(n15000), .A(n14999), .B(n14998), .ZN(
        n15002) );
  AOI211_X1 U16682 ( .C1(n15005), .C2(n15004), .A(n15003), .B(n15002), .ZN(
        n15006) );
  OAI21_X1 U16683 ( .B1(n15008), .B2(n15007), .A(n15006), .ZN(P2_U3206) );
  INV_X1 U16684 ( .A(n15009), .ZN(n15062) );
  OAI21_X1 U16685 ( .B1(n15062), .B2(n15010), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15011) );
  OAI21_X1 U16686 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15011), .ZN(n15022) );
  OAI211_X1 U16687 ( .C1(n15014), .C2(n15013), .A(n15091), .B(n15012), .ZN(
        n15021) );
  NAND2_X1 U16688 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15083), .ZN(n15020) );
  AOI211_X1 U16689 ( .C1(n15017), .C2(n15016), .A(n15015), .B(n15103), .ZN(
        n15018) );
  INV_X1 U16690 ( .A(n15018), .ZN(n15019) );
  NAND4_X1 U16691 ( .A1(n15022), .A2(n15021), .A3(n15020), .A4(n15019), .ZN(
        P2_U3218) );
  NAND2_X1 U16692 ( .A1(n15089), .A2(n15023), .ZN(n15026) );
  AOI21_X1 U16693 ( .B1(n15083), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n15024), .ZN(
        n15025) );
  AND2_X1 U16694 ( .A1(n15026), .A2(n15025), .ZN(n15036) );
  AOI211_X1 U16695 ( .C1(n15029), .C2(n15028), .A(n15027), .B(n15103), .ZN(
        n15030) );
  INV_X1 U16696 ( .A(n15030), .ZN(n15035) );
  OAI211_X1 U16697 ( .C1(n15033), .C2(n15032), .A(n15091), .B(n15031), .ZN(
        n15034) );
  NAND3_X1 U16698 ( .A1(n15036), .A2(n15035), .A3(n15034), .ZN(P2_U3219) );
  INV_X1 U16699 ( .A(n15037), .ZN(n15040) );
  OAI21_X1 U16700 ( .B1(n15111), .B2(n14708), .A(n15038), .ZN(n15039) );
  AOI21_X1 U16701 ( .B1(n15040), .B2(n15089), .A(n15039), .ZN(n15049) );
  OAI211_X1 U16702 ( .C1(n15043), .C2(n15042), .A(n15091), .B(n15041), .ZN(
        n15048) );
  OAI211_X1 U16703 ( .C1(n15046), .C2(n15045), .A(n15044), .B(n15085), .ZN(
        n15047) );
  NAND3_X1 U16704 ( .A1(n15049), .A2(n15048), .A3(n15047), .ZN(P2_U3221) );
  AOI22_X1 U16705 ( .A1(n15083), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n15060) );
  NAND2_X1 U16706 ( .A1(n15089), .A2(n15050), .ZN(n15059) );
  OAI211_X1 U16707 ( .C1(n15053), .C2(n15052), .A(n15085), .B(n15051), .ZN(
        n15058) );
  OAI211_X1 U16708 ( .C1(n15056), .C2(n15055), .A(n15091), .B(n15054), .ZN(
        n15057) );
  NAND4_X1 U16709 ( .A1(n15060), .A2(n15059), .A3(n15058), .A4(n15057), .ZN(
        P2_U3227) );
  OAI21_X1 U16710 ( .B1(n15062), .B2(n15061), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15063) );
  OAI21_X1 U16711 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15063), .ZN(n15072) );
  OAI211_X1 U16712 ( .C1(n15065), .C2(P2_REG2_REG_14__SCAN_IN), .A(n15091), 
        .B(n15064), .ZN(n15071) );
  NAND2_X1 U16713 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n15083), .ZN(n15070) );
  OAI211_X1 U16714 ( .C1(n15068), .C2(n15067), .A(n15085), .B(n15066), .ZN(
        n15069) );
  NAND4_X1 U16715 ( .A1(n15072), .A2(n15071), .A3(n15070), .A4(n15069), .ZN(
        P2_U3228) );
  AOI22_X1 U16716 ( .A1(n15083), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15081) );
  NAND2_X1 U16717 ( .A1(n15089), .A2(n15073), .ZN(n15080) );
  OAI211_X1 U16718 ( .C1(n15075), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15091), 
        .B(n15074), .ZN(n15079) );
  OAI211_X1 U16719 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15077), .A(n15085), 
        .B(n15076), .ZN(n15078) );
  NAND4_X1 U16720 ( .A1(n15081), .A2(n15080), .A3(n15079), .A4(n15078), .ZN(
        P2_U3229) );
  AOI22_X1 U16721 ( .A1(n15083), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n15097) );
  OAI211_X1 U16722 ( .C1(n15087), .C2(n15086), .A(n15085), .B(n15084), .ZN(
        n15096) );
  NAND2_X1 U16723 ( .A1(n15089), .A2(n15088), .ZN(n15095) );
  OAI211_X1 U16724 ( .C1(n15093), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        n15094) );
  NAND4_X1 U16725 ( .A1(n15097), .A2(n15096), .A3(n15095), .A4(n15094), .ZN(
        P2_U3231) );
  AOI21_X1 U16726 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n15099), .A(n15098), 
        .ZN(n15104) );
  OAI21_X1 U16727 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n15101), .A(n15100), 
        .ZN(n15102) );
  OAI222_X1 U16728 ( .A1(n15107), .A2(n15106), .B1(n15105), .B2(n15104), .C1(
        n15103), .C2(n15102), .ZN(n15108) );
  INV_X1 U16729 ( .A(n15108), .ZN(n15110) );
  OAI211_X1 U16730 ( .C1(n15112), .C2(n15111), .A(n15110), .B(n15109), .ZN(
        P2_U3232) );
  INV_X1 U16731 ( .A(n15113), .ZN(n15119) );
  OAI22_X1 U16732 ( .A1(n15155), .A2(n15115), .B1(n15114), .B2(n15132), .ZN(
        n15116) );
  AOI21_X1 U16733 ( .B1(n15144), .B2(n15117), .A(n15116), .ZN(n15118) );
  OAI21_X1 U16734 ( .B1(n15119), .B2(n15140), .A(n15118), .ZN(n15120) );
  AOI21_X1 U16735 ( .B1(n15122), .B2(n15121), .A(n15120), .ZN(n15123) );
  OAI21_X1 U16736 ( .B1(n15157), .B2(n15124), .A(n15123), .ZN(P2_U3258) );
  OAI21_X1 U16737 ( .B1(n15126), .B2(n15138), .A(n15125), .ZN(n15130) );
  AOI222_X1 U16738 ( .A1(n15131), .A2(n15130), .B1(n15129), .B2(n15128), .C1(
        n11972), .C2(n15127), .ZN(n15174) );
  OAI22_X1 U16739 ( .A1(n15155), .A2(n9903), .B1(n15133), .B2(n15132), .ZN(
        n15142) );
  OAI211_X1 U16740 ( .C1(n15175), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        n15173) );
  XNOR2_X1 U16741 ( .A(n15138), .B(n15137), .ZN(n15172) );
  OAI22_X1 U16742 ( .A1(n15140), .A2(n15173), .B1(n15172), .B2(n15139), .ZN(
        n15141) );
  AOI211_X1 U16743 ( .C1(n15144), .C2(n15143), .A(n15142), .B(n15141), .ZN(
        n15145) );
  OAI21_X1 U16744 ( .B1(n15157), .B2(n15174), .A(n15145), .ZN(P2_U3264) );
  OAI21_X1 U16745 ( .B1(n15146), .B2(n15131), .A(n15170), .ZN(n15147) );
  OAI21_X1 U16746 ( .B1(n9542), .B2(n15148), .A(n15147), .ZN(n15168) );
  INV_X1 U16747 ( .A(n15170), .ZN(n15152) );
  NAND2_X1 U16748 ( .A1(n15149), .A2(n9661), .ZN(n15167) );
  OAI22_X1 U16749 ( .A1(n15152), .A2(n6875), .B1(n15150), .B2(n15167), .ZN(
        n15153) );
  AOI211_X1 U16750 ( .C1(n15154), .C2(P2_REG3_REG_0__SCAN_IN), .A(n15168), .B(
        n15153), .ZN(n15156) );
  AOI22_X1 U16751 ( .A1(n15157), .A2(n9973), .B1(n15156), .B2(n15155), .ZN(
        P2_U3265) );
  NOR2_X1 U16752 ( .A1(n15163), .A2(n15158), .ZN(n15159) );
  AND2_X1 U16753 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15160), .ZN(P2_U3266) );
  AND2_X1 U16754 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15160), .ZN(P2_U3267) );
  AND2_X1 U16755 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15160), .ZN(P2_U3268) );
  AND2_X1 U16756 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15160), .ZN(P2_U3269) );
  INV_X1 U16757 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15636) );
  NOR2_X1 U16758 ( .A1(n15159), .A2(n15636), .ZN(P2_U3270) );
  AND2_X1 U16759 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15160), .ZN(P2_U3271) );
  AND2_X1 U16760 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15160), .ZN(P2_U3272) );
  AND2_X1 U16761 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15160), .ZN(P2_U3273) );
  AND2_X1 U16762 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15160), .ZN(P2_U3274) );
  AND2_X1 U16763 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15160), .ZN(P2_U3275) );
  INV_X1 U16764 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15569) );
  NOR2_X1 U16765 ( .A1(n15159), .A2(n15569), .ZN(P2_U3276) );
  AND2_X1 U16766 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15160), .ZN(P2_U3277) );
  AND2_X1 U16767 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15160), .ZN(P2_U3278) );
  AND2_X1 U16768 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15160), .ZN(P2_U3279) );
  AND2_X1 U16769 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15160), .ZN(P2_U3280) );
  AND2_X1 U16770 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15160), .ZN(P2_U3281) );
  AND2_X1 U16771 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15160), .ZN(P2_U3282) );
  AND2_X1 U16772 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15160), .ZN(P2_U3283) );
  AND2_X1 U16773 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15160), .ZN(P2_U3284) );
  AND2_X1 U16774 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15160), .ZN(P2_U3285) );
  AND2_X1 U16775 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15160), .ZN(P2_U3286) );
  AND2_X1 U16776 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15160), .ZN(P2_U3287) );
  AND2_X1 U16777 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15160), .ZN(P2_U3288) );
  AND2_X1 U16778 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15160), .ZN(P2_U3289) );
  AND2_X1 U16779 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15160), .ZN(P2_U3290) );
  AND2_X1 U16780 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15160), .ZN(P2_U3291) );
  AND2_X1 U16781 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15160), .ZN(P2_U3292) );
  AND2_X1 U16782 ( .A1(n15160), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3293) );
  AND2_X1 U16783 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15160), .ZN(P2_U3294) );
  AND2_X1 U16784 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15160), .ZN(P2_U3295) );
  AOI22_X1 U16785 ( .A1(n15166), .A2(n15162), .B1(n15161), .B2(n15163), .ZN(
        P2_U3416) );
  AOI22_X1 U16786 ( .A1(n15166), .A2(n15165), .B1(n15164), .B2(n15163), .ZN(
        P2_U3417) );
  INV_X1 U16787 ( .A(n15167), .ZN(n15169) );
  AOI211_X1 U16788 ( .C1(n15218), .C2(n15170), .A(n15169), .B(n15168), .ZN(
        n15224) );
  INV_X1 U16789 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15171) );
  AOI22_X1 U16790 ( .A1(n15212), .A2(n15224), .B1(n15171), .B2(n15222), .ZN(
        P2_U3430) );
  INV_X1 U16791 ( .A(n15172), .ZN(n15177) );
  OAI211_X1 U16792 ( .C1(n15175), .C2(n15215), .A(n15174), .B(n15173), .ZN(
        n15176) );
  AOI21_X1 U16793 ( .B1(n15178), .B2(n15177), .A(n15176), .ZN(n15226) );
  INV_X1 U16794 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15179) );
  AOI22_X1 U16795 ( .A1(n15212), .A2(n15226), .B1(n15179), .B2(n15222), .ZN(
        P2_U3433) );
  INV_X1 U16796 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15180) );
  AOI22_X1 U16797 ( .A1(n15212), .A2(n15181), .B1(n15180), .B2(n15222), .ZN(
        P2_U3436) );
  AOI21_X1 U16798 ( .B1(n15196), .B2(n15183), .A(n15182), .ZN(n15185) );
  OAI211_X1 U16799 ( .C1(n15187), .C2(n15186), .A(n15185), .B(n15184), .ZN(
        n15188) );
  INV_X1 U16800 ( .A(n15188), .ZN(n15227) );
  INV_X1 U16801 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15189) );
  AOI22_X1 U16802 ( .A1(n15212), .A2(n15227), .B1(n15189), .B2(n15222), .ZN(
        P2_U3439) );
  OAI21_X1 U16803 ( .B1(n15191), .B2(n15215), .A(n15190), .ZN(n15193) );
  AOI211_X1 U16804 ( .C1(n15218), .C2(n15194), .A(n15193), .B(n15192), .ZN(
        n15228) );
  INV_X1 U16805 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15195) );
  AOI22_X1 U16806 ( .A1(n15212), .A2(n15228), .B1(n15195), .B2(n15222), .ZN(
        P2_U3442) );
  AND2_X1 U16807 ( .A1(n15197), .A2(n15196), .ZN(n15198) );
  NOR2_X1 U16808 ( .A1(n15199), .A2(n15198), .ZN(n15205) );
  OR2_X1 U16809 ( .A1(n15202), .A2(n15200), .ZN(n15204) );
  OR2_X1 U16810 ( .A1(n15202), .A2(n15201), .ZN(n15203) );
  AND4_X1 U16811 ( .A1(n15206), .A2(n15205), .A3(n15204), .A4(n15203), .ZN(
        n15229) );
  AOI22_X1 U16812 ( .A1(n15212), .A2(n15229), .B1(n9048), .B2(n15222), .ZN(
        P2_U3445) );
  OAI21_X1 U16813 ( .B1(n15208), .B2(n15215), .A(n15207), .ZN(n15210) );
  AOI211_X1 U16814 ( .C1(n15218), .C2(n15211), .A(n15210), .B(n15209), .ZN(
        n15230) );
  INV_X1 U16815 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15592) );
  AOI22_X1 U16816 ( .A1(n15212), .A2(n15230), .B1(n15592), .B2(n15222), .ZN(
        P2_U3454) );
  INV_X1 U16817 ( .A(n15213), .ZN(n15216) );
  OAI21_X1 U16818 ( .B1(n15216), .B2(n15215), .A(n15214), .ZN(n15217) );
  AOI21_X1 U16819 ( .B1(n15219), .B2(n15218), .A(n15217), .ZN(n15220) );
  AND2_X1 U16820 ( .A1(n15221), .A2(n15220), .ZN(n15232) );
  INV_X1 U16821 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15223) );
  AOI22_X1 U16822 ( .A1(n15212), .A2(n15232), .B1(n15223), .B2(n15222), .ZN(
        P2_U3460) );
  AOI22_X1 U16823 ( .A1(n15233), .A2(n15224), .B1(n9974), .B2(n15231), .ZN(
        P2_U3499) );
  AOI22_X1 U16824 ( .A1(n15233), .A2(n15226), .B1(n15225), .B2(n15231), .ZN(
        P2_U3500) );
  AOI22_X1 U16825 ( .A1(n15233), .A2(n15227), .B1(n9021), .B2(n15231), .ZN(
        P2_U3502) );
  AOI22_X1 U16826 ( .A1(n15233), .A2(n15228), .B1(n9030), .B2(n15231), .ZN(
        P2_U3503) );
  AOI22_X1 U16827 ( .A1(n15233), .A2(n15229), .B1(n9922), .B2(n15231), .ZN(
        P2_U3504) );
  AOI22_X1 U16828 ( .A1(n15233), .A2(n15230), .B1(n9925), .B2(n15231), .ZN(
        P2_U3507) );
  AOI22_X1 U16829 ( .A1(n15233), .A2(n15232), .B1(n10261), .B2(n15231), .ZN(
        P2_U3509) );
  NOR2_X1 U16830 ( .A1(P3_U3897), .A2(n15234), .ZN(P3_U3150) );
  OAI21_X1 U16831 ( .B1(n15237), .B2(n15236), .A(n15235), .ZN(n15265) );
  NOR2_X1 U16832 ( .A1(n7746), .A2(n15295), .ZN(n15264) );
  INV_X1 U16833 ( .A(n15264), .ZN(n15241) );
  OAI22_X1 U16834 ( .A1(n15241), .A2(n15240), .B1(n15239), .B2(n15238), .ZN(
        n15254) );
  INV_X1 U16835 ( .A(n15265), .ZN(n15253) );
  AOI22_X1 U16836 ( .A1(n15244), .A2(n10244), .B1(n15243), .B2(n15242), .ZN(
        n15251) );
  OAI21_X1 U16837 ( .B1(n15247), .B2(n15246), .A(n15245), .ZN(n15249) );
  NAND2_X1 U16838 ( .A1(n15249), .A2(n15248), .ZN(n15250) );
  OAI211_X1 U16839 ( .C1(n15253), .C2(n15252), .A(n15251), .B(n15250), .ZN(
        n15263) );
  AOI211_X1 U16840 ( .C1(n15255), .C2(n15265), .A(n15254), .B(n15263), .ZN(
        n15256) );
  AOI22_X1 U16841 ( .A1(n15258), .A2(n15257), .B1(n15256), .B2(n13344), .ZN(
        P3_U3231) );
  OR2_X1 U16842 ( .A1(n15259), .A2(n9740), .ZN(n15260) );
  AND3_X1 U16843 ( .A1(n15262), .A2(n15261), .A3(n15260), .ZN(n15310) );
  AOI22_X1 U16844 ( .A1(n15309), .A2(n15310), .B1(n7683), .B2(n15307), .ZN(
        P3_U3393) );
  AOI211_X1 U16845 ( .C1(n15303), .C2(n15265), .A(n15264), .B(n15263), .ZN(
        n15311) );
  AOI22_X1 U16846 ( .A1(n15309), .A2(n15311), .B1(n7711), .B2(n15307), .ZN(
        P3_U3396) );
  NOR2_X1 U16847 ( .A1(n15266), .A2(n15295), .ZN(n15268) );
  AOI211_X1 U16848 ( .C1(n15303), .C2(n15269), .A(n15268), .B(n15267), .ZN(
        n15312) );
  AOI22_X1 U16849 ( .A1(n15309), .A2(n15312), .B1(n7730), .B2(n15307), .ZN(
        P3_U3399) );
  NOR2_X1 U16850 ( .A1(n15270), .A2(n15295), .ZN(n15272) );
  AOI211_X1 U16851 ( .C1(n15303), .C2(n15273), .A(n15272), .B(n15271), .ZN(
        n15313) );
  AOI22_X1 U16852 ( .A1(n15309), .A2(n15313), .B1(n7753), .B2(n15307), .ZN(
        P3_U3402) );
  AOI22_X1 U16853 ( .A1(n15275), .A2(n15303), .B1(n15302), .B2(n15274), .ZN(
        n15276) );
  AND2_X1 U16854 ( .A1(n15277), .A2(n15276), .ZN(n15698) );
  INV_X1 U16855 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15278) );
  AOI22_X1 U16856 ( .A1(n15309), .A2(n15698), .B1(n15278), .B2(n15307), .ZN(
        P3_U3405) );
  NOR2_X1 U16857 ( .A1(n15279), .A2(n15295), .ZN(n15281) );
  AOI211_X1 U16858 ( .C1(n15303), .C2(n15282), .A(n15281), .B(n15280), .ZN(
        n15314) );
  AOI22_X1 U16859 ( .A1(n15309), .A2(n15314), .B1(n7791), .B2(n15307), .ZN(
        P3_U3408) );
  NOR2_X1 U16860 ( .A1(n15283), .A2(n15295), .ZN(n15284) );
  AOI21_X1 U16861 ( .B1(n15285), .B2(n15303), .A(n15284), .ZN(n15286) );
  AND2_X1 U16862 ( .A1(n15287), .A2(n15286), .ZN(n15315) );
  INV_X1 U16863 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15288) );
  AOI22_X1 U16864 ( .A1(n15309), .A2(n15315), .B1(n15288), .B2(n15307), .ZN(
        P3_U3411) );
  NOR2_X1 U16865 ( .A1(n15289), .A2(n15295), .ZN(n15291) );
  AOI211_X1 U16866 ( .C1(n15292), .C2(n15303), .A(n15291), .B(n15290), .ZN(
        n15316) );
  INV_X1 U16867 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15293) );
  AOI22_X1 U16868 ( .A1(n15309), .A2(n15316), .B1(n15293), .B2(n15307), .ZN(
        P3_U3414) );
  OAI21_X1 U16869 ( .B1(n15296), .B2(n15295), .A(n15294), .ZN(n15297) );
  AOI21_X1 U16870 ( .B1(n15299), .B2(n15298), .A(n15297), .ZN(n15317) );
  INV_X1 U16871 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15300) );
  AOI22_X1 U16872 ( .A1(n15309), .A2(n15317), .B1(n15300), .B2(n15307), .ZN(
        P3_U3417) );
  AOI22_X1 U16873 ( .A1(n15304), .A2(n15303), .B1(n15302), .B2(n15301), .ZN(
        n15305) );
  AND2_X1 U16874 ( .A1(n15306), .A2(n15305), .ZN(n15318) );
  INV_X1 U16875 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15308) );
  AOI22_X1 U16876 ( .A1(n15309), .A2(n15318), .B1(n15308), .B2(n15307), .ZN(
        P3_U3420) );
  AOI22_X1 U16877 ( .A1(n15699), .A2(n15310), .B1(n7684), .B2(n15696), .ZN(
        P3_U3460) );
  AOI22_X1 U16878 ( .A1(n15699), .A2(n15311), .B1(n10133), .B2(n15696), .ZN(
        P3_U3461) );
  AOI22_X1 U16879 ( .A1(n15699), .A2(n15312), .B1(n10119), .B2(n15696), .ZN(
        P3_U3462) );
  AOI22_X1 U16880 ( .A1(n15699), .A2(n15313), .B1(n10163), .B2(n15696), .ZN(
        P3_U3463) );
  AOI22_X1 U16881 ( .A1(n15699), .A2(n15314), .B1(n10433), .B2(n15696), .ZN(
        P3_U3465) );
  AOI22_X1 U16882 ( .A1(n15699), .A2(n15315), .B1(n10463), .B2(n15696), .ZN(
        P3_U3466) );
  AOI22_X1 U16883 ( .A1(n15699), .A2(n15316), .B1(n15639), .B2(n15696), .ZN(
        P3_U3467) );
  AOI22_X1 U16884 ( .A1(n15699), .A2(n15317), .B1(n10952), .B2(n15696), .ZN(
        P3_U3468) );
  AOI22_X1 U16885 ( .A1(n15699), .A2(n15318), .B1(n11223), .B2(n15696), .ZN(
        P3_U3469) );
  OAI22_X1 U16886 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(keyinput12), .B1(
        keyinput36), .B2(P1_IR_REG_6__SCAN_IN), .ZN(n15319) );
  AOI221_X1 U16887 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(keyinput12), .C1(
        P1_IR_REG_6__SCAN_IN), .C2(keyinput36), .A(n15319), .ZN(n15326) );
  OAI22_X1 U16888 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(keyinput98), .B1(
        P1_REG0_REG_27__SCAN_IN), .B2(keyinput122), .ZN(n15320) );
  AOI221_X1 U16889 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(keyinput98), .C1(
        keyinput122), .C2(P1_REG0_REG_27__SCAN_IN), .A(n15320), .ZN(n15325) );
  OAI22_X1 U16890 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput101), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput26), .ZN(n15321) );
  AOI221_X1 U16891 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput101), .C1(
        keyinput26), .C2(P1_IR_REG_31__SCAN_IN), .A(n15321), .ZN(n15324) );
  OAI22_X1 U16892 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(keyinput40), .B1(SI_25_), .B2(keyinput13), .ZN(n15322) );
  AOI221_X1 U16893 ( .B1(P1_DATAO_REG_15__SCAN_IN), .B2(keyinput40), .C1(
        keyinput13), .C2(SI_25_), .A(n15322), .ZN(n15323) );
  NAND4_X1 U16894 ( .A1(n15326), .A2(n15325), .A3(n15324), .A4(n15323), .ZN(
        n15354) );
  OAI22_X1 U16895 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput71), .B1(
        keyinput64), .B2(P2_ADDR_REG_14__SCAN_IN), .ZN(n15327) );
  AOI221_X1 U16896 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput71), .C1(
        P2_ADDR_REG_14__SCAN_IN), .C2(keyinput64), .A(n15327), .ZN(n15334) );
  OAI22_X1 U16897 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput84), .B1(
        keyinput22), .B2(P2_D_REG_4__SCAN_IN), .ZN(n15328) );
  AOI221_X1 U16898 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput84), .C1(
        P2_D_REG_4__SCAN_IN), .C2(keyinput22), .A(n15328), .ZN(n15333) );
  OAI22_X1 U16899 ( .A1(P2_REG0_REG_6__SCAN_IN), .A2(keyinput113), .B1(
        P2_REG2_REG_30__SCAN_IN), .B2(keyinput11), .ZN(n15329) );
  AOI221_X1 U16900 ( .B1(P2_REG0_REG_6__SCAN_IN), .B2(keyinput113), .C1(
        keyinput11), .C2(P2_REG2_REG_30__SCAN_IN), .A(n15329), .ZN(n15332) );
  OAI22_X1 U16901 ( .A1(P3_REG0_REG_4__SCAN_IN), .A2(keyinput86), .B1(
        keyinput8), .B2(P1_D_REG_26__SCAN_IN), .ZN(n15330) );
  AOI221_X1 U16902 ( .B1(P3_REG0_REG_4__SCAN_IN), .B2(keyinput86), .C1(
        P1_D_REG_26__SCAN_IN), .C2(keyinput8), .A(n15330), .ZN(n15331) );
  NAND4_X1 U16903 ( .A1(n15334), .A2(n15333), .A3(n15332), .A4(n15331), .ZN(
        n15353) );
  OAI22_X1 U16904 ( .A1(P3_REG0_REG_27__SCAN_IN), .A2(keyinput69), .B1(
        P1_REG1_REG_7__SCAN_IN), .B2(keyinput124), .ZN(n15335) );
  AOI221_X1 U16905 ( .B1(P3_REG0_REG_27__SCAN_IN), .B2(keyinput69), .C1(
        keyinput124), .C2(P1_REG1_REG_7__SCAN_IN), .A(n15335), .ZN(n15342) );
  OAI22_X1 U16906 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(keyinput121), .B1(
        keyinput82), .B2(P2_REG3_REG_15__SCAN_IN), .ZN(n15336) );
  AOI221_X1 U16907 ( .B1(P2_DATAO_REG_5__SCAN_IN), .B2(keyinput121), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput82), .A(n15336), .ZN(n15341) );
  OAI22_X1 U16908 ( .A1(P1_D_REG_20__SCAN_IN), .A2(keyinput103), .B1(
        P1_ADDR_REG_5__SCAN_IN), .B2(keyinput4), .ZN(n15337) );
  AOI221_X1 U16909 ( .B1(P1_D_REG_20__SCAN_IN), .B2(keyinput103), .C1(
        keyinput4), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n15337), .ZN(n15340) );
  OAI22_X1 U16910 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput57), .B1(
        keyinput66), .B2(P1_REG3_REG_19__SCAN_IN), .ZN(n15338) );
  AOI221_X1 U16911 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput57), .C1(
        P1_REG3_REG_19__SCAN_IN), .C2(keyinput66), .A(n15338), .ZN(n15339) );
  NAND4_X1 U16912 ( .A1(n15342), .A2(n15341), .A3(n15340), .A4(n15339), .ZN(
        n15352) );
  OAI22_X1 U16913 ( .A1(P3_REG1_REG_21__SCAN_IN), .A2(keyinput102), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(keyinput35), .ZN(n15343) );
  AOI221_X1 U16914 ( .B1(P3_REG1_REG_21__SCAN_IN), .B2(keyinput102), .C1(
        keyinput35), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n15343), .ZN(n15350) );
  OAI22_X1 U16915 ( .A1(P2_REG0_REG_25__SCAN_IN), .A2(keyinput80), .B1(
        P3_DATAO_REG_4__SCAN_IN), .B2(keyinput108), .ZN(n15344) );
  AOI221_X1 U16916 ( .B1(P2_REG0_REG_25__SCAN_IN), .B2(keyinput80), .C1(
        keyinput108), .C2(P3_DATAO_REG_4__SCAN_IN), .A(n15344), .ZN(n15349) );
  OAI22_X1 U16917 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput48), .B1(
        keyinput45), .B2(P2_REG1_REG_3__SCAN_IN), .ZN(n15345) );
  AOI221_X1 U16918 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput48), .C1(
        P2_REG1_REG_3__SCAN_IN), .C2(keyinput45), .A(n15345), .ZN(n15348) );
  OAI22_X1 U16919 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(keyinput114), .B1(
        P3_ADDR_REG_8__SCAN_IN), .B2(keyinput34), .ZN(n15346) );
  AOI221_X1 U16920 ( .B1(P3_ADDR_REG_13__SCAN_IN), .B2(keyinput114), .C1(
        keyinput34), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n15346), .ZN(n15347) );
  NAND4_X1 U16921 ( .A1(n15350), .A2(n15349), .A3(n15348), .A4(n15347), .ZN(
        n15351) );
  NOR4_X1 U16922 ( .A1(n15354), .A2(n15353), .A3(n15352), .A4(n15351), .ZN(
        n15695) );
  AOI22_X1 U16923 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput251), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(keyinput142), .ZN(n15355) );
  OAI221_X1 U16924 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput251), .C1(
        P1_DATAO_REG_5__SCAN_IN), .C2(keyinput142), .A(n15355), .ZN(n15362) );
  AOI22_X1 U16925 ( .A1(P2_REG1_REG_24__SCAN_IN), .A2(keyinput151), .B1(
        P3_REG2_REG_23__SCAN_IN), .B2(keyinput217), .ZN(n15356) );
  OAI221_X1 U16926 ( .B1(P2_REG1_REG_24__SCAN_IN), .B2(keyinput151), .C1(
        P3_REG2_REG_23__SCAN_IN), .C2(keyinput217), .A(n15356), .ZN(n15361) );
  AOI22_X1 U16927 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput243), .B1(
        P1_REG1_REG_26__SCAN_IN), .B2(keyinput202), .ZN(n15357) );
  OAI221_X1 U16928 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput243), .C1(
        P1_REG1_REG_26__SCAN_IN), .C2(keyinput202), .A(n15357), .ZN(n15360) );
  AOI22_X1 U16929 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(keyinput165), .B1(
        P2_REG2_REG_22__SCAN_IN), .B2(keyinput174), .ZN(n15358) );
  OAI221_X1 U16930 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(keyinput165), .C1(
        P2_REG2_REG_22__SCAN_IN), .C2(keyinput174), .A(n15358), .ZN(n15359) );
  NOR4_X1 U16931 ( .A1(n15362), .A2(n15361), .A3(n15360), .A4(n15359), .ZN(
        n15390) );
  AOI22_X1 U16932 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(keyinput153), .B1(SI_19_), .B2(keyinput198), .ZN(n15363) );
  OAI221_X1 U16933 ( .B1(P1_REG2_REG_24__SCAN_IN), .B2(keyinput153), .C1(
        SI_19_), .C2(keyinput198), .A(n15363), .ZN(n15370) );
  AOI22_X1 U16934 ( .A1(P1_REG0_REG_16__SCAN_IN), .A2(keyinput247), .B1(SI_7_), 
        .B2(keyinput184), .ZN(n15364) );
  OAI221_X1 U16935 ( .B1(P1_REG0_REG_16__SCAN_IN), .B2(keyinput247), .C1(SI_7_), .C2(keyinput184), .A(n15364), .ZN(n15369) );
  AOI22_X1 U16936 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(keyinput252), .B1(
        P3_REG2_REG_27__SCAN_IN), .B2(keyinput227), .ZN(n15365) );
  OAI221_X1 U16937 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(keyinput252), .C1(
        P3_REG2_REG_27__SCAN_IN), .C2(keyinput227), .A(n15365), .ZN(n15368) );
  AOI22_X1 U16938 ( .A1(P1_D_REG_18__SCAN_IN), .A2(keyinput134), .B1(
        P2_ADDR_REG_19__SCAN_IN), .B2(keyinput157), .ZN(n15366) );
  OAI221_X1 U16939 ( .B1(P1_D_REG_18__SCAN_IN), .B2(keyinput134), .C1(
        P2_ADDR_REG_19__SCAN_IN), .C2(keyinput157), .A(n15366), .ZN(n15367) );
  NOR4_X1 U16940 ( .A1(n15370), .A2(n15369), .A3(n15368), .A4(n15367), .ZN(
        n15389) );
  AOI22_X1 U16941 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(keyinput200), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput164), .ZN(n15371) );
  OAI221_X1 U16942 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(keyinput200), .C1(
        P1_IR_REG_6__SCAN_IN), .C2(keyinput164), .A(n15371), .ZN(n15378) );
  AOI22_X1 U16943 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput169), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(keyinput168), .ZN(n15372) );
  OAI221_X1 U16944 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput169), .C1(
        P1_DATAO_REG_15__SCAN_IN), .C2(keyinput168), .A(n15372), .ZN(n15377)
         );
  AOI22_X1 U16945 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(keyinput162), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput246), .ZN(n15373) );
  OAI221_X1 U16946 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(keyinput162), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput246), .A(n15373), .ZN(n15376) );
  AOI22_X1 U16947 ( .A1(P3_REG1_REG_21__SCAN_IN), .A2(keyinput230), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(keyinput249), .ZN(n15374) );
  OAI221_X1 U16948 ( .B1(P3_REG1_REG_21__SCAN_IN), .B2(keyinput230), .C1(
        P2_DATAO_REG_5__SCAN_IN), .C2(keyinput249), .A(n15374), .ZN(n15375) );
  NOR4_X1 U16949 ( .A1(n15378), .A2(n15377), .A3(n15376), .A4(n15375), .ZN(
        n15388) );
  AOI22_X1 U16950 ( .A1(P3_DATAO_REG_25__SCAN_IN), .A2(keyinput172), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput175), .ZN(n15379) );
  OAI221_X1 U16951 ( .B1(P3_DATAO_REG_25__SCAN_IN), .B2(keyinput172), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput175), .A(n15379), .ZN(n15386) );
  AOI22_X1 U16952 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(keyinput193), .B1(
        P2_IR_REG_7__SCAN_IN), .B2(keyinput135), .ZN(n15380) );
  OAI221_X1 U16953 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(keyinput193), .C1(
        P2_IR_REG_7__SCAN_IN), .C2(keyinput135), .A(n15380), .ZN(n15385) );
  AOI22_X1 U16954 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(keyinput132), .B1(
        P2_IR_REG_13__SCAN_IN), .B2(keyinput238), .ZN(n15381) );
  OAI221_X1 U16955 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(keyinput132), .C1(
        P2_IR_REG_13__SCAN_IN), .C2(keyinput238), .A(n15381), .ZN(n15384) );
  AOI22_X1 U16956 ( .A1(P2_D_REG_4__SCAN_IN), .A2(keyinput150), .B1(
        P1_D_REG_13__SCAN_IN), .B2(keyinput221), .ZN(n15382) );
  OAI221_X1 U16957 ( .B1(P2_D_REG_4__SCAN_IN), .B2(keyinput150), .C1(
        P1_D_REG_13__SCAN_IN), .C2(keyinput221), .A(n15382), .ZN(n15383) );
  NOR4_X1 U16958 ( .A1(n15386), .A2(n15385), .A3(n15384), .A4(n15383), .ZN(
        n15387) );
  NAND4_X1 U16959 ( .A1(n15390), .A2(n15389), .A3(n15388), .A4(n15387), .ZN(
        n15527) );
  AOI22_X1 U16960 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(keyinput203), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(keyinput133), .ZN(n15391) );
  OAI221_X1 U16961 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(keyinput203), .C1(
        P1_DATAO_REG_9__SCAN_IN), .C2(keyinput133), .A(n15391), .ZN(n15398) );
  AOI22_X1 U16962 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(keyinput166), .B1(SI_5_), 
        .B2(keyinput156), .ZN(n15392) );
  OAI221_X1 U16963 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(keyinput166), .C1(SI_5_), 
        .C2(keyinput156), .A(n15392), .ZN(n15397) );
  AOI22_X1 U16964 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput160), .B1(
        P3_DATAO_REG_12__SCAN_IN), .B2(keyinput234), .ZN(n15393) );
  OAI221_X1 U16965 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput160), .C1(
        P3_DATAO_REG_12__SCAN_IN), .C2(keyinput234), .A(n15393), .ZN(n15396)
         );
  AOI22_X1 U16966 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(keyinput206), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(keyinput216), .ZN(n15394) );
  OAI221_X1 U16967 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(keyinput206), .C1(
        P2_IR_REG_30__SCAN_IN), .C2(keyinput216), .A(n15394), .ZN(n15395) );
  NOR4_X1 U16968 ( .A1(n15398), .A2(n15397), .A3(n15396), .A4(n15395), .ZN(
        n15426) );
  AOI22_X1 U16969 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput154), .B1(
        P3_IR_REG_30__SCAN_IN), .B2(keyinput138), .ZN(n15399) );
  OAI221_X1 U16970 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput154), .C1(
        P3_IR_REG_30__SCAN_IN), .C2(keyinput138), .A(n15399), .ZN(n15406) );
  AOI22_X1 U16971 ( .A1(P2_REG0_REG_19__SCAN_IN), .A2(keyinput235), .B1(
        P3_REG3_REG_16__SCAN_IN), .B2(keyinput195), .ZN(n15400) );
  OAI221_X1 U16972 ( .B1(P2_REG0_REG_19__SCAN_IN), .B2(keyinput235), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput195), .A(n15400), .ZN(n15405) );
  AOI22_X1 U16973 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(keyinput143), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput190), .ZN(n15401) );
  OAI221_X1 U16974 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(keyinput143), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput190), .A(n15401), .ZN(n15404) );
  AOI22_X1 U16975 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(keyinput213), .B1(
        P2_REG1_REG_3__SCAN_IN), .B2(keyinput173), .ZN(n15402) );
  OAI221_X1 U16976 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(keyinput213), .C1(
        P2_REG1_REG_3__SCAN_IN), .C2(keyinput173), .A(n15402), .ZN(n15403) );
  NOR4_X1 U16977 ( .A1(n15406), .A2(n15405), .A3(n15404), .A4(n15403), .ZN(
        n15425) );
  AOI22_X1 U16978 ( .A1(P3_D_REG_12__SCAN_IN), .A2(keyinput170), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(keyinput229), .ZN(n15407) );
  OAI221_X1 U16979 ( .B1(P3_D_REG_12__SCAN_IN), .B2(keyinput170), .C1(
        P1_DATAO_REG_0__SCAN_IN), .C2(keyinput229), .A(n15407), .ZN(n15414) );
  AOI22_X1 U16980 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(keyinput144), .B1(
        P3_D_REG_16__SCAN_IN), .B2(keyinput228), .ZN(n15408) );
  OAI221_X1 U16981 ( .B1(P2_REG2_REG_21__SCAN_IN), .B2(keyinput144), .C1(
        P3_D_REG_16__SCAN_IN), .C2(keyinput228), .A(n15408), .ZN(n15413) );
  AOI22_X1 U16982 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(keyinput152), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput210), .ZN(n15409) );
  OAI221_X1 U16983 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(keyinput152), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput210), .A(n15409), .ZN(n15412) );
  AOI22_X1 U16984 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(keyinput192), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(keyinput181), .ZN(n15410) );
  OAI221_X1 U16985 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(keyinput192), .C1(
        P1_REG3_REG_3__SCAN_IN), .C2(keyinput181), .A(n15410), .ZN(n15411) );
  NOR4_X1 U16986 ( .A1(n15414), .A2(n15413), .A3(n15412), .A4(n15411), .ZN(
        n15424) );
  AOI22_X1 U16987 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(keyinput233), .B1(
        P2_REG2_REG_14__SCAN_IN), .B2(keyinput129), .ZN(n15415) );
  OAI221_X1 U16988 ( .B1(P3_DATAO_REG_11__SCAN_IN), .B2(keyinput233), .C1(
        P2_REG2_REG_14__SCAN_IN), .C2(keyinput129), .A(n15415), .ZN(n15422) );
  AOI22_X1 U16989 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(keyinput225), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput176), .ZN(n15416) );
  OAI221_X1 U16990 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(keyinput225), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput176), .A(n15416), .ZN(n15421) );
  AOI22_X1 U16991 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(keyinput201), .B1(
        P1_D_REG_5__SCAN_IN), .B2(keyinput240), .ZN(n15417) );
  OAI221_X1 U16992 ( .B1(P3_ADDR_REG_1__SCAN_IN), .B2(keyinput201), .C1(
        P1_D_REG_5__SCAN_IN), .C2(keyinput240), .A(n15417), .ZN(n15420) );
  AOI22_X1 U16993 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(keyinput161), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput224), .ZN(n15418) );
  OAI221_X1 U16994 ( .B1(P1_REG3_REG_5__SCAN_IN), .B2(keyinput161), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput224), .A(n15418), .ZN(n15419) );
  NOR4_X1 U16995 ( .A1(n15422), .A2(n15421), .A3(n15420), .A4(n15419), .ZN(
        n15423) );
  NAND4_X1 U16996 ( .A1(n15426), .A2(n15425), .A3(n15424), .A4(n15423), .ZN(
        n15526) );
  AOI22_X1 U16997 ( .A1(n15615), .A2(keyinput167), .B1(n15636), .B2(
        keyinput196), .ZN(n15427) );
  OAI221_X1 U16998 ( .B1(n15615), .B2(keyinput167), .C1(n15636), .C2(
        keyinput196), .A(n15427), .ZN(n15435) );
  INV_X1 U16999 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15630) );
  AOI22_X1 U17000 ( .A1(n10831), .A2(keyinput223), .B1(n15630), .B2(
        keyinput187), .ZN(n15428) );
  OAI221_X1 U17001 ( .B1(n10831), .B2(keyinput223), .C1(n15630), .C2(
        keyinput187), .A(n15428), .ZN(n15434) );
  INV_X1 U17002 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n15549) );
  AOI22_X1 U17003 ( .A1(n15549), .A2(keyinput245), .B1(n15532), .B2(
        keyinput248), .ZN(n15429) );
  OAI221_X1 U17004 ( .B1(n15549), .B2(keyinput245), .C1(n15532), .C2(
        keyinput248), .A(n15429), .ZN(n15433) );
  AOI22_X1 U17005 ( .A1(n15557), .A2(keyinput211), .B1(n15431), .B2(
        keyinput208), .ZN(n15430) );
  OAI221_X1 U17006 ( .B1(n15557), .B2(keyinput211), .C1(n15431), .C2(
        keyinput208), .A(n15430), .ZN(n15432) );
  NOR4_X1 U17007 ( .A1(n15435), .A2(n15434), .A3(n15433), .A4(n15432), .ZN(
        n15473) );
  AOI22_X1 U17008 ( .A1(n15437), .A2(keyinput155), .B1(keyinput222), .B2(
        n15575), .ZN(n15436) );
  OAI221_X1 U17009 ( .B1(n15437), .B2(keyinput155), .C1(n15575), .C2(
        keyinput222), .A(n15436), .ZN(n15447) );
  AOI22_X1 U17010 ( .A1(n10463), .A2(keyinput140), .B1(keyinput231), .B2(
        n15439), .ZN(n15438) );
  OAI221_X1 U17011 ( .B1(n10463), .B2(keyinput140), .C1(n15439), .C2(
        keyinput231), .A(n15438), .ZN(n15446) );
  AOI22_X1 U17012 ( .A1(n15669), .A2(keyinput177), .B1(keyinput194), .B2(
        n15441), .ZN(n15440) );
  OAI221_X1 U17013 ( .B1(n15669), .B2(keyinput177), .C1(n15441), .C2(
        keyinput194), .A(n15440), .ZN(n15445) );
  AOI22_X1 U17014 ( .A1(n15443), .A2(keyinput215), .B1(keyinput253), .B2(
        n15574), .ZN(n15442) );
  OAI221_X1 U17015 ( .B1(n15443), .B2(keyinput215), .C1(n15574), .C2(
        keyinput253), .A(n15442), .ZN(n15444) );
  NOR4_X1 U17016 ( .A1(n15447), .A2(n15446), .A3(n15445), .A4(n15444), .ZN(
        n15472) );
  AOI22_X1 U17017 ( .A1(n15450), .A2(keyinput219), .B1(n15449), .B2(
        keyinput250), .ZN(n15448) );
  OAI221_X1 U17018 ( .B1(n15450), .B2(keyinput219), .C1(n15449), .C2(
        keyinput250), .A(n15448), .ZN(n15458) );
  AOI22_X1 U17019 ( .A1(n15601), .A2(keyinput239), .B1(keyinput214), .B2(n7753), .ZN(n15451) );
  OAI221_X1 U17020 ( .B1(n15601), .B2(keyinput239), .C1(n7753), .C2(
        keyinput214), .A(n15451), .ZN(n15457) );
  INV_X1 U17021 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n15634) );
  AOI22_X1 U17022 ( .A1(n15634), .A2(keyinput159), .B1(n15558), .B2(
        keyinput130), .ZN(n15452) );
  OAI221_X1 U17023 ( .B1(n15634), .B2(keyinput159), .C1(n15558), .C2(
        keyinput130), .A(n15452), .ZN(n15456) );
  AOI22_X1 U17024 ( .A1(n15454), .A2(keyinput141), .B1(keyinput189), .B2(
        n15592), .ZN(n15453) );
  OAI221_X1 U17025 ( .B1(n15454), .B2(keyinput141), .C1(n15592), .C2(
        keyinput189), .A(n15453), .ZN(n15455) );
  NOR4_X1 U17026 ( .A1(n15458), .A2(n15457), .A3(n15456), .A4(n15455), .ZN(
        n15471) );
  AOI22_X1 U17027 ( .A1(n15590), .A2(keyinput148), .B1(keyinput242), .B2(
        n15460), .ZN(n15459) );
  OAI221_X1 U17028 ( .B1(n15590), .B2(keyinput148), .C1(n15460), .C2(
        keyinput242), .A(n15459), .ZN(n15469) );
  AOI22_X1 U17029 ( .A1(n9073), .A2(keyinput241), .B1(n15462), .B2(keyinput137), .ZN(n15461) );
  OAI221_X1 U17030 ( .B1(n9073), .B2(keyinput241), .C1(n15462), .C2(
        keyinput137), .A(n15461), .ZN(n15468) );
  AOI22_X1 U17031 ( .A1(n15639), .A2(keyinput158), .B1(keyinput204), .B2(
        n15603), .ZN(n15463) );
  OAI221_X1 U17032 ( .B1(n15639), .B2(keyinput158), .C1(n15603), .C2(
        keyinput204), .A(n15463), .ZN(n15467) );
  XNOR2_X1 U17033 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput205), .ZN(n15465) );
  XNOR2_X1 U17034 ( .A(P1_REG3_REG_21__SCAN_IN), .B(keyinput186), .ZN(n15464)
         );
  NAND2_X1 U17035 ( .A1(n15465), .A2(n15464), .ZN(n15466) );
  NOR4_X1 U17036 ( .A1(n15469), .A2(n15468), .A3(n15467), .A4(n15466), .ZN(
        n15470) );
  NAND4_X1 U17037 ( .A1(n15473), .A2(n15472), .A3(n15471), .A4(n15470), .ZN(
        n15525) );
  XOR2_X1 U17038 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(keyinput180), .Z(n15478) );
  XNOR2_X1 U17039 ( .A(n15474), .B(keyinput197), .ZN(n15477) );
  XNOR2_X1 U17040 ( .A(n15475), .B(keyinput191), .ZN(n15476) );
  NOR3_X1 U17041 ( .A1(n15478), .A2(n15477), .A3(n15476), .ZN(n15481) );
  XNOR2_X1 U17042 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput183), .ZN(n15480)
         );
  XNOR2_X1 U17043 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput131), .ZN(n15479)
         );
  NAND3_X1 U17044 ( .A1(n15481), .A2(n15480), .A3(n15479), .ZN(n15487) );
  AOI22_X1 U17045 ( .A1(n15483), .A2(keyinput218), .B1(n15531), .B2(
        keyinput254), .ZN(n15482) );
  OAI221_X1 U17046 ( .B1(n15483), .B2(keyinput218), .C1(n15531), .C2(
        keyinput254), .A(n15482), .ZN(n15486) );
  XNOR2_X1 U17047 ( .A(n15484), .B(keyinput236), .ZN(n15485) );
  NOR3_X1 U17048 ( .A1(n15487), .A2(n15486), .A3(n15485), .ZN(n15523) );
  AOI22_X1 U17049 ( .A1(n10119), .A2(keyinput226), .B1(keyinput182), .B2(
        n10417), .ZN(n15488) );
  OAI221_X1 U17050 ( .B1(n10119), .B2(keyinput226), .C1(n10417), .C2(
        keyinput182), .A(n15488), .ZN(n15497) );
  AOI22_X1 U17051 ( .A1(n9187), .A2(keyinput232), .B1(n15569), .B2(keyinput149), .ZN(n15489) );
  OAI221_X1 U17052 ( .B1(n9187), .B2(keyinput232), .C1(n15569), .C2(
        keyinput149), .A(n15489), .ZN(n15496) );
  INV_X1 U17053 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15490) );
  XOR2_X1 U17054 ( .A(n15490), .B(keyinput163), .Z(n15494) );
  XOR2_X1 U17055 ( .A(n15546), .B(keyinput255), .Z(n15493) );
  XNOR2_X1 U17056 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput146), .ZN(n15492)
         );
  XNOR2_X1 U17057 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput185), .ZN(n15491)
         );
  NAND4_X1 U17058 ( .A1(n15494), .A2(n15493), .A3(n15492), .A4(n15491), .ZN(
        n15495) );
  NOR3_X1 U17059 ( .A1(n15497), .A2(n15496), .A3(n15495), .ZN(n15522) );
  AOI22_X1 U17060 ( .A1(n9126), .A2(keyinput237), .B1(n15499), .B2(keyinput212), .ZN(n15498) );
  OAI221_X1 U17061 ( .B1(n9126), .B2(keyinput237), .C1(n15499), .C2(
        keyinput212), .A(n15498), .ZN(n15507) );
  XNOR2_X1 U17062 ( .A(keyinput199), .B(n9111), .ZN(n15506) );
  XNOR2_X1 U17063 ( .A(keyinput209), .B(n11349), .ZN(n15505) );
  XNOR2_X1 U17064 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput179), .ZN(n15503) );
  XNOR2_X1 U17065 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput207), .ZN(n15502) );
  XNOR2_X1 U17066 ( .A(P3_REG1_REG_0__SCAN_IN), .B(keyinput171), .ZN(n15501)
         );
  XNOR2_X1 U17067 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput128), .ZN(n15500)
         );
  NAND4_X1 U17068 ( .A1(n15503), .A2(n15502), .A3(n15501), .A4(n15500), .ZN(
        n15504) );
  NOR4_X1 U17069 ( .A1(n15507), .A2(n15506), .A3(n15505), .A4(n15504), .ZN(
        n15521) );
  INV_X1 U17070 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15510) );
  AOI22_X1 U17071 ( .A1(n15510), .A2(keyinput145), .B1(keyinput178), .B2(
        n15509), .ZN(n15508) );
  OAI221_X1 U17072 ( .B1(n15510), .B2(keyinput145), .C1(n15509), .C2(
        keyinput178), .A(n15508), .ZN(n15519) );
  AOI22_X1 U17073 ( .A1(n15512), .A2(keyinput136), .B1(keyinput188), .B2(
        n15560), .ZN(n15511) );
  OAI221_X1 U17074 ( .B1(n15512), .B2(keyinput136), .C1(n15560), .C2(
        keyinput188), .A(n15511), .ZN(n15518) );
  XOR2_X1 U17075 ( .A(n9509), .B(keyinput139), .Z(n15516) );
  XNOR2_X1 U17076 ( .A(keyinput244), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n15515)
         );
  XNOR2_X1 U17077 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput220), .ZN(n15514) );
  XNOR2_X1 U17078 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput147), .ZN(n15513)
         );
  NAND4_X1 U17079 ( .A1(n15516), .A2(n15515), .A3(n15514), .A4(n15513), .ZN(
        n15517) );
  NOR3_X1 U17080 ( .A1(n15519), .A2(n15518), .A3(n15517), .ZN(n15520) );
  NAND4_X1 U17081 ( .A1(n15523), .A2(n15522), .A3(n15521), .A4(n15520), .ZN(
        n15524) );
  NOR4_X1 U17082 ( .A1(n15527), .A2(n15526), .A3(n15525), .A4(n15524), .ZN(
        n15651) );
  AOI22_X1 U17083 ( .A1(n9224), .A2(keyinput1), .B1(n15529), .B2(keyinput29), 
        .ZN(n15528) );
  OAI221_X1 U17084 ( .B1(n9224), .B2(keyinput1), .C1(n15529), .C2(keyinput29), 
        .A(n15528), .ZN(n15539) );
  AOI22_X1 U17085 ( .A1(n15532), .A2(keyinput120), .B1(keyinput126), .B2(
        n15531), .ZN(n15530) );
  OAI221_X1 U17086 ( .B1(n15532), .B2(keyinput120), .C1(n15531), .C2(
        keyinput126), .A(n15530), .ZN(n15538) );
  XNOR2_X1 U17087 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(keyinput52), .ZN(n15536)
         );
  XNOR2_X1 U17088 ( .A(SI_7_), .B(keyinput56), .ZN(n15535) );
  XNOR2_X1 U17089 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput19), .ZN(n15534)
         );
  XNOR2_X1 U17090 ( .A(keyinput116), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n15533)
         );
  NAND4_X1 U17091 ( .A1(n15536), .A2(n15535), .A3(n15534), .A4(n15533), .ZN(
        n15537) );
  NOR3_X1 U17092 ( .A1(n15539), .A2(n15538), .A3(n15537), .ZN(n15585) );
  AOI22_X1 U17093 ( .A1(n15541), .A2(keyinput78), .B1(n13769), .B2(keyinput16), 
        .ZN(n15540) );
  OAI221_X1 U17094 ( .B1(n15541), .B2(keyinput78), .C1(n13769), .C2(keyinput16), .A(n15540), .ZN(n15553) );
  AOI22_X1 U17095 ( .A1(n13751), .A2(keyinput46), .B1(n15543), .B2(keyinput47), 
        .ZN(n15542) );
  OAI221_X1 U17096 ( .B1(n13751), .B2(keyinput46), .C1(n15543), .C2(keyinput47), .A(n15542), .ZN(n15552) );
  AOI22_X1 U17097 ( .A1(n15546), .A2(keyinput127), .B1(n15545), .B2(keyinput58), .ZN(n15544) );
  OAI221_X1 U17098 ( .B1(n15546), .B2(keyinput127), .C1(n15545), .C2(
        keyinput58), .A(n15544), .ZN(n15551) );
  AOI22_X1 U17099 ( .A1(n15549), .A2(keyinput117), .B1(n15548), .B2(keyinput96), .ZN(n15547) );
  OAI221_X1 U17100 ( .B1(n15549), .B2(keyinput117), .C1(n15548), .C2(
        keyinput96), .A(n15547), .ZN(n15550) );
  NOR4_X1 U17101 ( .A1(n15553), .A2(n15552), .A3(n15551), .A4(n15550), .ZN(
        n15584) );
  AOI22_X1 U17102 ( .A1(n14399), .A2(keyinput25), .B1(n15555), .B2(keyinput53), 
        .ZN(n15554) );
  OAI221_X1 U17103 ( .B1(n14399), .B2(keyinput25), .C1(n15555), .C2(keyinput53), .A(n15554), .ZN(n15567) );
  AOI22_X1 U17104 ( .A1(n15558), .A2(keyinput2), .B1(keyinput83), .B2(n15557), 
        .ZN(n15556) );
  OAI221_X1 U17105 ( .B1(n15558), .B2(keyinput2), .C1(n15557), .C2(keyinput83), 
        .A(n15556), .ZN(n15566) );
  AOI22_X1 U17106 ( .A1(n15561), .A2(keyinput107), .B1(n15560), .B2(keyinput60), .ZN(n15559) );
  OAI221_X1 U17107 ( .B1(n15561), .B2(keyinput107), .C1(n15560), .C2(
        keyinput60), .A(n15559), .ZN(n15565) );
  XNOR2_X1 U17108 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput14), .ZN(n15563)
         );
  XNOR2_X1 U17109 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput74), .ZN(n15562)
         );
  NAND2_X1 U17110 ( .A1(n15563), .A2(n15562), .ZN(n15564) );
  NOR4_X1 U17111 ( .A1(n15567), .A2(n15566), .A3(n15565), .A4(n15564), .ZN(
        n15583) );
  AOI22_X1 U17112 ( .A1(n15569), .A2(keyinput21), .B1(keyinput109), .B2(n9126), 
        .ZN(n15568) );
  OAI221_X1 U17113 ( .B1(n15569), .B2(keyinput21), .C1(n9126), .C2(keyinput109), .A(n15568), .ZN(n15581) );
  AOI22_X1 U17114 ( .A1(n10642), .A2(keyinput38), .B1(keyinput32), .B2(n15571), 
        .ZN(n15570) );
  OAI221_X1 U17115 ( .B1(n10642), .B2(keyinput38), .C1(n15571), .C2(keyinput32), .A(n15570), .ZN(n15580) );
  INV_X1 U17116 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n15573) );
  AOI22_X1 U17117 ( .A1(n15574), .A2(keyinput125), .B1(n15573), .B2(keyinput10), .ZN(n15572) );
  OAI221_X1 U17118 ( .B1(n15574), .B2(keyinput125), .C1(n15573), .C2(
        keyinput10), .A(n15572), .ZN(n15579) );
  XOR2_X1 U17119 ( .A(n15575), .B(keyinput94), .Z(n15577) );
  XNOR2_X1 U17120 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput18), .ZN(n15576)
         );
  NAND2_X1 U17121 ( .A1(n15577), .A2(n15576), .ZN(n15578) );
  NOR4_X1 U17122 ( .A1(n15581), .A2(n15580), .A3(n15579), .A4(n15578), .ZN(
        n15582) );
  NAND4_X1 U17123 ( .A1(n15585), .A2(n15584), .A3(n15583), .A4(n15582), .ZN(
        n15650) );
  AOI22_X1 U17124 ( .A1(n10831), .A2(keyinput95), .B1(n15587), .B2(keyinput55), 
        .ZN(n15586) );
  OAI221_X1 U17125 ( .B1(n10831), .B2(keyinput95), .C1(n15587), .C2(keyinput55), .A(n15586), .ZN(n15599) );
  AOI22_X1 U17126 ( .A1(n15590), .A2(keyinput20), .B1(keyinput23), .B2(n15589), 
        .ZN(n15588) );
  OAI221_X1 U17127 ( .B1(n15590), .B2(keyinput20), .C1(n15589), .C2(keyinput23), .A(n15588), .ZN(n15598) );
  INV_X1 U17128 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15591) );
  XNOR2_X1 U17129 ( .A(n15591), .B(keyinput42), .ZN(n15597) );
  XOR2_X1 U17130 ( .A(n15592), .B(keyinput61), .Z(n15595) );
  XNOR2_X1 U17131 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput62), .ZN(n15594) );
  XNOR2_X1 U17132 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput92), .ZN(n15593) );
  NAND3_X1 U17133 ( .A1(n15595), .A2(n15594), .A3(n15593), .ZN(n15596) );
  NOR4_X1 U17134 ( .A1(n15599), .A2(n15598), .A3(n15597), .A4(n15596), .ZN(
        n15648) );
  AOI22_X1 U17135 ( .A1(n15601), .A2(keyinput111), .B1(keyinput97), .B2(n9030), 
        .ZN(n15600) );
  OAI221_X1 U17136 ( .B1(n15601), .B2(keyinput111), .C1(n9030), .C2(keyinput97), .A(n15600), .ZN(n15612) );
  INV_X1 U17137 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n15604) );
  AOI22_X1 U17138 ( .A1(n15604), .A2(keyinput100), .B1(keyinput76), .B2(n15603), .ZN(n15602) );
  OAI221_X1 U17139 ( .B1(n15604), .B2(keyinput100), .C1(n15603), .C2(
        keyinput76), .A(n15602), .ZN(n15611) );
  XOR2_X1 U17140 ( .A(n15605), .B(keyinput73), .Z(n15609) );
  XNOR2_X1 U17141 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput63), .ZN(n15608) );
  XNOR2_X1 U17142 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput0), .ZN(n15607) );
  XNOR2_X1 U17143 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput77), .ZN(n15606) );
  NAND4_X1 U17144 ( .A1(n15609), .A2(n15608), .A3(n15607), .A4(n15606), .ZN(
        n15610) );
  NOR3_X1 U17145 ( .A1(n15612), .A2(n15611), .A3(n15610), .ZN(n15647) );
  AOI22_X1 U17146 ( .A1(n15615), .A2(keyinput39), .B1(n15614), .B2(keyinput89), 
        .ZN(n15613) );
  OAI221_X1 U17147 ( .B1(n15615), .B2(keyinput39), .C1(n15614), .C2(keyinput89), .A(n15613), .ZN(n15618) );
  INV_X1 U17148 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15616) );
  XNOR2_X1 U17149 ( .A(n15616), .B(keyinput41), .ZN(n15617) );
  NOR2_X1 U17150 ( .A1(n15618), .A2(n15617), .ZN(n15628) );
  AOI22_X1 U17151 ( .A1(n14177), .A2(keyinput85), .B1(n15620), .B2(keyinput70), 
        .ZN(n15619) );
  OAI221_X1 U17152 ( .B1(n14177), .B2(keyinput85), .C1(n15620), .C2(keyinput70), .A(n15619), .ZN(n15621) );
  INV_X1 U17153 ( .A(n15621), .ZN(n15627) );
  AOI22_X1 U17154 ( .A1(n11439), .A2(keyinput65), .B1(n15623), .B2(keyinput43), 
        .ZN(n15622) );
  OAI221_X1 U17155 ( .B1(n11439), .B2(keyinput65), .C1(n15623), .C2(keyinput43), .A(n15622), .ZN(n15624) );
  INV_X1 U17156 ( .A(n15624), .ZN(n15626) );
  XNOR2_X1 U17157 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput7), .ZN(n15625) );
  AND4_X1 U17158 ( .A1(n15628), .A2(n15627), .A3(n15626), .A4(n15625), .ZN(
        n15646) );
  AOI22_X1 U17159 ( .A1(n15631), .A2(keyinput106), .B1(n15630), .B2(keyinput59), .ZN(n15629) );
  OAI221_X1 U17160 ( .B1(n15631), .B2(keyinput106), .C1(n15630), .C2(
        keyinput59), .A(n15629), .ZN(n15644) );
  AOI22_X1 U17161 ( .A1(n15634), .A2(keyinput31), .B1(keyinput44), .B2(n15633), 
        .ZN(n15632) );
  OAI221_X1 U17162 ( .B1(n15634), .B2(keyinput31), .C1(n15633), .C2(keyinput44), .A(n15632), .ZN(n15643) );
  AOI22_X1 U17163 ( .A1(n15637), .A2(keyinput75), .B1(keyinput68), .B2(n15636), 
        .ZN(n15635) );
  OAI221_X1 U17164 ( .B1(n15637), .B2(keyinput75), .C1(n15636), .C2(keyinput68), .A(n15635), .ZN(n15642) );
  AOI22_X1 U17165 ( .A1(n15640), .A2(keyinput119), .B1(n15639), .B2(keyinput30), .ZN(n15638) );
  OAI221_X1 U17166 ( .B1(n15640), .B2(keyinput119), .C1(n15639), .C2(
        keyinput30), .A(n15638), .ZN(n15641) );
  NOR4_X1 U17167 ( .A1(n15644), .A2(n15643), .A3(n15642), .A4(n15641), .ZN(
        n15645) );
  NAND4_X1 U17168 ( .A1(n15648), .A2(n15647), .A3(n15646), .A4(n15645), .ZN(
        n15649) );
  NOR3_X1 U17169 ( .A1(n15651), .A2(n15650), .A3(n15649), .ZN(n15694) );
  OAI22_X1 U17170 ( .A1(P1_REG0_REG_24__SCAN_IN), .A2(keyinput27), .B1(
        P1_ADDR_REG_6__SCAN_IN), .B2(keyinput37), .ZN(n15652) );
  AOI221_X1 U17171 ( .B1(P1_REG0_REG_24__SCAN_IN), .B2(keyinput27), .C1(
        keyinput37), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n15652), .ZN(n15659) );
  OAI22_X1 U17172 ( .A1(P3_REG2_REG_27__SCAN_IN), .A2(keyinput99), .B1(
        P3_REG1_REG_16__SCAN_IN), .B2(keyinput87), .ZN(n15653) );
  AOI221_X1 U17173 ( .B1(P3_REG2_REG_27__SCAN_IN), .B2(keyinput99), .C1(
        keyinput87), .C2(P3_REG1_REG_16__SCAN_IN), .A(n15653), .ZN(n15658) );
  OAI22_X1 U17174 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(keyinput79), .B1(
        P3_DATAO_REG_11__SCAN_IN), .B2(keyinput105), .ZN(n15654) );
  AOI221_X1 U17175 ( .B1(P2_IR_REG_22__SCAN_IN), .B2(keyinput79), .C1(
        keyinput105), .C2(P3_DATAO_REG_11__SCAN_IN), .A(n15654), .ZN(n15657)
         );
  OAI22_X1 U17176 ( .A1(P1_D_REG_13__SCAN_IN), .A2(keyinput93), .B1(keyinput17), .B2(P1_REG0_REG_9__SCAN_IN), .ZN(n15655) );
  AOI221_X1 U17177 ( .B1(P1_D_REG_13__SCAN_IN), .B2(keyinput93), .C1(
        P1_REG0_REG_9__SCAN_IN), .C2(keyinput17), .A(n15655), .ZN(n15656) );
  NAND4_X1 U17178 ( .A1(n15659), .A2(n15658), .A3(n15657), .A4(n15656), .ZN(
        n15692) );
  OAI22_X1 U17179 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(keyinput9), .B1(
        keyinput88), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n15660) );
  AOI221_X1 U17180 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(keyinput9), .C1(
        P2_IR_REG_30__SCAN_IN), .C2(keyinput88), .A(n15660), .ZN(n15667) );
  OAI22_X1 U17181 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(keyinput110), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(keyinput123), .ZN(n15661) );
  AOI221_X1 U17182 ( .B1(P2_IR_REG_13__SCAN_IN), .B2(keyinput110), .C1(
        keyinput123), .C2(P2_REG3_REG_0__SCAN_IN), .A(n15661), .ZN(n15666) );
  OAI22_X1 U17183 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(keyinput90), .B1(
        keyinput91), .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n15662) );
  AOI221_X1 U17184 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(keyinput90), .C1(
        P3_DATAO_REG_10__SCAN_IN), .C2(keyinput91), .A(n15662), .ZN(n15665) );
  OAI22_X1 U17185 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(keyinput5), .B1(
        keyinput24), .B2(P2_ADDR_REG_4__SCAN_IN), .ZN(n15663) );
  AOI221_X1 U17186 ( .B1(P1_DATAO_REG_9__SCAN_IN), .B2(keyinput5), .C1(
        P2_ADDR_REG_4__SCAN_IN), .C2(keyinput24), .A(n15663), .ZN(n15664) );
  NAND4_X1 U17187 ( .A1(n15667), .A2(n15666), .A3(n15665), .A4(n15664), .ZN(
        n15691) );
  OAI22_X1 U17188 ( .A1(n15669), .A2(keyinput49), .B1(keyinput15), .B2(
        P1_ADDR_REG_12__SCAN_IN), .ZN(n15668) );
  AOI221_X1 U17189 ( .B1(n15669), .B2(keyinput49), .C1(P1_ADDR_REG_12__SCAN_IN), .C2(keyinput15), .A(n15668), .ZN(n15680) );
  OAI22_X1 U17190 ( .A1(n15671), .A2(keyinput33), .B1(n11904), .B2(keyinput72), 
        .ZN(n15670) );
  AOI221_X1 U17191 ( .B1(n15671), .B2(keyinput33), .C1(keyinput72), .C2(n11904), .A(n15670), .ZN(n15679) );
  OAI22_X1 U17192 ( .A1(n9187), .A2(keyinput104), .B1(keyinput115), .B2(
        P2_REG3_REG_9__SCAN_IN), .ZN(n15672) );
  AOI221_X1 U17193 ( .B1(n9187), .B2(keyinput104), .C1(P2_REG3_REG_9__SCAN_IN), 
        .C2(keyinput115), .A(n15672), .ZN(n15678) );
  XNOR2_X1 U17194 ( .A(n15673), .B(keyinput28), .ZN(n15676) );
  XNOR2_X1 U17195 ( .A(n15674), .B(keyinput51), .ZN(n15675) );
  NOR2_X1 U17196 ( .A1(n15676), .A2(n15675), .ZN(n15677) );
  NAND4_X1 U17197 ( .A1(n15680), .A2(n15679), .A3(n15678), .A4(n15677), .ZN(
        n15690) );
  OAI22_X1 U17198 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(keyinput54), .B1(
        P3_DATAO_REG_7__SCAN_IN), .B2(keyinput50), .ZN(n15681) );
  AOI221_X1 U17199 ( .B1(P3_ADDR_REG_2__SCAN_IN), .B2(keyinput54), .C1(
        keyinput50), .C2(P3_DATAO_REG_7__SCAN_IN), .A(n15681), .ZN(n15688) );
  OAI22_X1 U17200 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(keyinput3), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput118), .ZN(n15682) );
  AOI221_X1 U17201 ( .B1(P1_DATAO_REG_7__SCAN_IN), .B2(keyinput3), .C1(
        keyinput118), .C2(P2_REG3_REG_14__SCAN_IN), .A(n15682), .ZN(n15687) );
  OAI22_X1 U17202 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput67), .B1(
        P1_D_REG_5__SCAN_IN), .B2(keyinput112), .ZN(n15683) );
  AOI221_X1 U17203 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput67), .C1(
        keyinput112), .C2(P1_D_REG_5__SCAN_IN), .A(n15683), .ZN(n15686) );
  OAI22_X1 U17204 ( .A1(P1_D_REG_18__SCAN_IN), .A2(keyinput6), .B1(
        P1_REG2_REG_3__SCAN_IN), .B2(keyinput81), .ZN(n15684) );
  AOI221_X1 U17205 ( .B1(P1_D_REG_18__SCAN_IN), .B2(keyinput6), .C1(keyinput81), .C2(P1_REG2_REG_3__SCAN_IN), .A(n15684), .ZN(n15685) );
  NAND4_X1 U17206 ( .A1(n15688), .A2(n15687), .A3(n15686), .A4(n15685), .ZN(
        n15689) );
  NOR4_X1 U17207 ( .A1(n15692), .A2(n15691), .A3(n15690), .A4(n15689), .ZN(
        n15693) );
  NAND3_X1 U17208 ( .A1(n15695), .A2(n15694), .A3(n15693), .ZN(n15701) );
  AOI22_X1 U17209 ( .A1(n15699), .A2(n15698), .B1(n15697), .B2(n15696), .ZN(
        n15700) );
  XNOR2_X1 U17210 ( .A(n15701), .B(n15700), .ZN(P3_U3464) );
  AOI21_X1 U17211 ( .B1(n15702), .B2(n9979), .A(n15713), .ZN(SUB_1596_U53) );
  XOR2_X1 U17212 ( .A(n15704), .B(n15703), .Z(SUB_1596_U59) );
  XNOR2_X1 U17213 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15705), .ZN(SUB_1596_U58)
         );
  XOR2_X1 U17214 ( .A(n15707), .B(n15706), .Z(SUB_1596_U56) );
  AOI21_X1 U17215 ( .B1(n15710), .B2(n15709), .A(n15708), .ZN(n15711) );
  XOR2_X1 U17216 ( .A(n15711), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  XOR2_X1 U17217 ( .A(n15713), .B(n15712), .Z(SUB_1596_U5) );
  AND3_X1 U8357 ( .A1(n7744), .A2(n7743), .A3(n7742), .ZN(n12885) );
  CLKBUF_X2 U7395 ( .A(n8050), .Z(n6642) );
  CLKBUF_X1 U7419 ( .A(n12304), .Z(n12506) );
  CLKBUF_X1 U7424 ( .A(n13271), .Z(n6882) );
  CLKBUF_X1 U7428 ( .A(n8941), .Z(n13946) );
  AOI21_X1 U7468 ( .B1(n13183), .B2(n13344), .A(n13182), .ZN(n13184) );
endmodule

