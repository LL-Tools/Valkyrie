

module b17_C_gen_AntiSAT_k_128_5 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9631, n9632, n9633, n9634, n9635, n9637, n9639, n9640, n9641, n9642,
         n9643, n9644, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9668, n9669, n9670, n9671, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18428, n18429, n18430, n18431, n18432, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258;

  AND2_X1 U11075 ( .A1(n15045), .A2(n15151), .ZN(n15010) );
  NAND2_X1 U11076 ( .A1(n11662), .A2(n16040), .ZN(n9817) );
  NOR2_X1 U11077 ( .A1(n19002), .A2(n18992), .ZN(n18382) );
  NAND4_X1 U11078 ( .A1(n10234), .A2(n14009), .A3(n10240), .A4(n10232), .ZN(
        n14107) );
  NOR2_X1 U11079 ( .A1(n11301), .A2(n18145), .ZN(n11304) );
  CLKBUF_X2 U11080 ( .A(n12742), .Z(n15224) );
  AOI21_X1 U11081 ( .B1(n16109), .B2(n16108), .A(n14174), .ZN(n16199) );
  NOR2_X2 U11082 ( .A1(n18998), .A2(n11273), .ZN(n16109) );
  CLKBUF_X3 U11083 ( .A(n13531), .Z(n9653) );
  OR2_X1 U11084 ( .A1(n11366), .A2(n11340), .ZN(n19709) );
  OR2_X1 U11085 ( .A1(n11366), .A2(n11361), .ZN(n19789) );
  OR2_X1 U11086 ( .A1(n11372), .A2(n13903), .ZN(n19895) );
  NAND2_X1 U11087 ( .A1(n9826), .A2(n11347), .ZN(n19676) );
  OR2_X1 U11088 ( .A1(n13065), .A2(n10951), .ZN(n10689) );
  AOI211_X1 U11089 ( .C1(n17450), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n11230), .B(n11229), .ZN(n11271) );
  CLKBUF_X2 U11090 ( .A(n11068), .Z(n17544) );
  CLKBUF_X2 U11091 ( .A(n11769), .Z(n12366) );
  CLKBUF_X1 U11092 ( .A(n14390), .Z(n9643) );
  CLKBUF_X2 U11094 ( .A(n12648), .Z(n9664) );
  CLKBUF_X3 U11095 ( .A(n11064), .Z(n9647) );
  CLKBUF_X1 U11096 ( .A(n14436), .Z(n9639) );
  CLKBUF_X2 U11098 ( .A(n11776), .Z(n12650) );
  CLKBUF_X1 U11099 ( .A(n14390), .Z(n9642) );
  OR3_X1 U11100 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n19020), .ZN(n11021) );
  CLKBUF_X2 U11101 ( .A(n14466), .Z(n9660) );
  NAND2_X2 U11102 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19020) );
  NAND2_X2 U11103 ( .A1(n10409), .A2(n10408), .ZN(n10486) );
  MUX2_X1 U11104 ( .A(n10396), .B(n10395), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10697) );
  NAND4_X2 U11105 ( .A1(n11734), .A2(n11733), .A3(n11732), .A4(n11731), .ZN(
        n13514) );
  AND2_X1 U11106 ( .A1(n10420), .A2(n10419), .ZN(n13116) );
  INV_X1 U11107 ( .A(n12608), .ZN(n12648) );
  NAND2_X1 U11108 ( .A1(n11726), .A2(n11719), .ZN(n12634) );
  NAND2_X1 U11109 ( .A1(n13381), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16071) );
  AND2_X1 U11110 ( .A1(n10154), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11718) );
  NOR3_X2 U11111 ( .A1(n17713), .A2(n18987), .A3(n18510), .ZN(n9631) );
  INV_X1 U11112 ( .A(n18521), .ZN(n18510) );
  OAI22_X2 U11114 ( .A1(n16781), .A2(n15341), .B1(n21231), .B2(n15340), .ZN(
        n20909) );
  NAND2_X2 U11115 ( .A1(n16286), .A2(n14263), .ZN(n15340) );
  INV_X1 U11116 ( .A(n19065), .ZN(n9632) );
  INV_X1 U11117 ( .A(n9632), .ZN(n9633) );
  INV_X1 U11118 ( .A(n9632), .ZN(n9634) );
  NAND2_X1 U11120 ( .A1(n11660), .A2(n11503), .ZN(n11655) );
  CLKBUF_X2 U11121 ( .A(n11846), .Z(n12651) );
  INV_X1 U11122 ( .A(n12603), .ZN(n12378) );
  AND2_X1 U11123 ( .A1(n13514), .A2(n13875), .ZN(n11833) );
  INV_X2 U11124 ( .A(n11744), .ZN(n12578) );
  AND2_X1 U11125 ( .A1(n10122), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11726) );
  AND2_X2 U11126 ( .A1(n10366), .A2(n13923), .ZN(n14466) );
  NAND2_X1 U11127 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10679), .ZN(
        n14440) );
  OR2_X1 U11128 ( .A1(n13271), .A2(n9675), .ZN(n11366) );
  AND2_X1 U11129 ( .A1(n11932), .A2(n13514), .ZN(n12788) );
  BUF_X4 U11130 ( .A(n14466), .Z(n9661) );
  INV_X2 U11132 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10680) );
  XNOR2_X1 U11133 ( .A(n11469), .B(n10179), .ZN(n11654) );
  AND2_X1 U11134 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13380) );
  NOR2_X1 U11136 ( .A1(n15418), .A2(n14527), .ZN(n14552) );
  NOR2_X1 U11137 ( .A1(n13849), .A2(n13848), .ZN(n13851) );
  NAND2_X1 U11138 ( .A1(n11661), .A2(n15724), .ZN(n11663) );
  OR2_X1 U11139 ( .A1(n11654), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14136) );
  NAND2_X1 U11140 ( .A1(n13023), .A2(n10463), .ZN(n10508) );
  NAND2_X1 U11141 ( .A1(n13379), .A2(n11353), .ZN(n11446) );
  NAND2_X1 U11142 ( .A1(n11355), .A2(n13379), .ZN(n11450) );
  CLKBUF_X3 U11143 ( .A(n17539), .Z(n9649) );
  INV_X1 U11144 ( .A(n17500), .ZN(n17545) );
  NAND2_X1 U11145 ( .A1(n11017), .A2(n19185), .ZN(n17247) );
  NAND2_X1 U11146 ( .A1(n13958), .A2(n13954), .ZN(n14093) );
  NAND2_X2 U11147 ( .A1(n14318), .A2(n14093), .ZN(n14656) );
  INV_X1 U11148 ( .A(n14721), .ZN(n12542) );
  NOR2_X1 U11149 ( .A1(n15045), .A2(n14999), .ZN(n15021) );
  INV_X1 U11150 ( .A(n12742), .ZN(n15018) );
  AND2_X1 U11151 ( .A1(n13296), .A2(n13293), .ZN(n13517) );
  BUF_X2 U11152 ( .A(n10532), .Z(n10652) );
  BUF_X1 U11154 ( .A(n19379), .Z(n9658) );
  INV_X1 U11155 ( .A(n19015), .ZN(n18400) );
  AND2_X1 U11156 ( .A1(n14099), .A2(n13686), .ZN(n20349) );
  NAND4_X1 U11157 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n13875) );
  NAND2_X1 U11158 ( .A1(n15460), .A2(n9790), .ZN(n14457) );
  AND2_X1 U11159 ( .A1(n11334), .A2(n11332), .ZN(n13050) );
  NOR2_X1 U11160 ( .A1(n15585), .A2(n15584), .ZN(n15789) );
  BUF_X1 U11161 ( .A(n13174), .Z(n9644) );
  INV_X1 U11162 ( .A(n14116), .ZN(n14611) );
  INV_X1 U11163 ( .A(n11607), .ZN(n15376) );
  INV_X1 U11164 ( .A(n10314), .ZN(n17394) );
  NOR4_X2 U11165 ( .A1(n19212), .A2(n17195), .A3(n16199), .A4(n19044), .ZN(
        n17581) );
  INV_X1 U11166 ( .A(n9647), .ZN(n17557) );
  INV_X1 U11167 ( .A(n11241), .ZN(n17539) );
  NAND2_X1 U11168 ( .A1(n9741), .A2(n9972), .ZN(n11284) );
  NOR3_X2 U11169 ( .A1(n11427), .A2(n11504), .A3(n10111), .ZN(n10109) );
  AND2_X1 U11170 ( .A1(n11718), .A2(n11726), .ZN(n11846) );
  INV_X1 U11171 ( .A(n9906), .ZN(n9635) );
  INV_X2 U11173 ( .A(n9635), .ZN(n9637) );
  AND2_X1 U11174 ( .A1(n11726), .A2(n11724), .ZN(n11776) );
  NOR2_X4 U11175 ( .A1(n10471), .A2(n10470), .ZN(n13023) );
  NAND2_X2 U11176 ( .A1(n10443), .A2(n10442), .ZN(n10691) );
  NOR2_X4 U11177 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16072) );
  XNOR2_X2 U11178 ( .A(n11935), .B(n11934), .ZN(n12098) );
  OAI22_X2 U11179 ( .A1(n13569), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12687), 
        .B2(n12007), .ZN(n11935) );
  AND2_X1 U11181 ( .A1(n10397), .A2(n10680), .ZN(n14436) );
  AOI211_X4 U11182 ( .C1(n17520), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n11245), .B(n11244), .ZN(n12869) );
  BUF_X8 U11183 ( .A(n17394), .Z(n9641) );
  NOR2_X2 U11184 ( .A1(n10355), .A2(n13983), .ZN(n10356) );
  BUF_X8 U11185 ( .A(n10444), .Z(n14577) );
  AOI21_X2 U11186 ( .B1(n11995), .B2(n21045), .A(n10310), .ZN(n12673) );
  INV_X2 U11187 ( .A(n15296), .ZN(n11995) );
  AND2_X1 U11188 ( .A1(n10397), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14390) );
  XNOR2_X1 U11189 ( .A(n11351), .B(n11335), .ZN(n13174) );
  NOR2_X2 U11190 ( .A1(n18130), .A2(n11132), .ZN(n11136) );
  INV_X4 U11191 ( .A(n10648), .ZN(n10642) );
  NOR2_X1 U11194 ( .A1(n17247), .A2(n11022), .ZN(n11064) );
  NAND2_X2 U11195 ( .A1(n13056), .A2(n10792), .ZN(n10951) );
  AND2_X1 U11196 ( .A1(n11725), .A2(n11724), .ZN(n9650) );
  AND2_X1 U11197 ( .A1(n11725), .A2(n11724), .ZN(n12586) );
  INV_X2 U11198 ( .A(n11062), .ZN(n9651) );
  INV_X1 U11199 ( .A(n9651), .ZN(n9652) );
  OR2_X1 U11200 ( .A1(n19167), .A2(n11026), .ZN(n11062) );
  AOI211_X2 U11201 ( .C1(n15147), .C2(n15144), .A(n15143), .B(n15145), .ZN(
        n16195) );
  AOI211_X1 U11202 ( .C1(n16589), .C2(n16455), .A(n15621), .B(n15620), .ZN(
        n15622) );
  NAND2_X1 U11203 ( .A1(n12542), .A2(n12541), .ZN(n14707) );
  OAI21_X1 U11204 ( .B1(n12845), .B2(n15224), .A(n12847), .ZN(n14992) );
  AOI21_X1 U11205 ( .B1(n9838), .B2(n9837), .A(n9907), .ZN(n9836) );
  AND2_X1 U11206 ( .A1(n10175), .A2(n9784), .ZN(n16115) );
  XNOR2_X1 U11207 ( .A(n14107), .B(n12204), .ZN(n14912) );
  OR2_X1 U11208 ( .A1(n9732), .A2(n9908), .ZN(n9907) );
  NOR2_X1 U11209 ( .A1(n15413), .A2(n15405), .ZN(n15406) );
  NOR2_X1 U11210 ( .A1(n17881), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17880) );
  NOR2_X1 U11211 ( .A1(n15091), .A2(n15093), .ZN(n15080) );
  NAND2_X1 U11212 ( .A1(n11654), .A2(n11667), .ZN(n10178) );
  OR2_X1 U11213 ( .A1(n17910), .A2(n9883), .ZN(n17903) );
  OR2_X1 U11214 ( .A1(n18108), .A2(n9885), .ZN(n11139) );
  OR2_X1 U11215 ( .A1(n13540), .A2(n13519), .ZN(n20453) );
  NAND2_X1 U11216 ( .A1(n13512), .A2(n13511), .ZN(n13540) );
  AND2_X1 U11217 ( .A1(n14099), .A2(n13672), .ZN(n13683) );
  NOR3_X1 U11218 ( .A1(n19296), .A2(n11667), .A3(n15958), .ZN(n15654) );
  NAND2_X1 U11219 ( .A1(n16054), .A2(n10296), .ZN(n13619) );
  NOR2_X1 U11220 ( .A1(n17464), .A2(n17460), .ZN(n17444) );
  NOR2_X1 U11221 ( .A1(n18147), .A2(n18146), .ZN(n18145) );
  NAND2_X1 U11222 ( .A1(n20547), .A2(n11991), .ZN(n11994) );
  NAND2_X1 U11223 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17482), .ZN(n17460) );
  AND2_X1 U11224 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17465), .ZN(n17482) );
  NOR2_X1 U11225 ( .A1(n11299), .A2(n18159), .ZN(n18147) );
  INV_X2 U11226 ( .A(n15449), .ZN(n15448) );
  AND2_X1 U11227 ( .A1(n10543), .A2(n10542), .ZN(n10547) );
  OR3_X1 U11228 ( .A1(n10094), .A2(n10096), .A3(n14160), .ZN(n10093) );
  CLKBUF_X2 U11229 ( .A(n10533), .Z(n10606) );
  OR2_X1 U11230 ( .A1(n10672), .A2(n20258), .ZN(n10512) );
  OR2_X1 U11231 ( .A1(n11272), .A2(n18997), .ZN(n14173) );
  INV_X1 U11232 ( .A(n13246), .ZN(n21043) );
  AOI211_X1 U11234 ( .C1(n9651), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n11190), .B(n11189), .ZN(n11259) );
  OR2_X1 U11235 ( .A1(n11789), .A2(n11788), .ZN(n11834) );
  BUF_X1 U11236 ( .A(n10476), .Z(n19603) );
  OR2_X1 U11237 ( .A1(n11775), .A2(n11774), .ZN(n13308) );
  INV_X4 U11238 ( .A(n10481), .ZN(n10457) );
  OR2_X2 U11239 ( .A1(n11832), .A2(n11831), .ZN(n13954) );
  NOR2_X1 U11240 ( .A1(n10358), .A2(n15705), .ZN(n10361) );
  NOR2_X1 U11241 ( .A1(n11758), .A2(n11757), .ZN(n11759) );
  AOI211_X1 U11242 ( .C1(n17544), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n11196), .B(n11195), .ZN(n11197) );
  INV_X2 U11243 ( .A(n11744), .ZN(n12647) );
  INV_X1 U11244 ( .A(n12492), .ZN(n9665) );
  INV_X4 U11245 ( .A(n11822), .ZN(n12580) );
  INV_X4 U11246 ( .A(n17547), .ZN(n17526) );
  INV_X4 U11247 ( .A(n9710), .ZN(n17497) );
  NAND2_X1 U11248 ( .A1(n11025), .A2(n11024), .ZN(n17468) );
  INV_X4 U11249 ( .A(n17388), .ZN(n17501) );
  INV_X1 U11250 ( .A(n9668), .ZN(n9654) );
  INV_X4 U11251 ( .A(n11180), .ZN(n17546) );
  INV_X8 U11252 ( .A(n11021), .ZN(n17541) );
  INV_X2 U11253 ( .A(n9709), .ZN(n9655) );
  INV_X2 U11254 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11017) );
  AND2_X1 U11255 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11724) );
  AND2_X1 U11256 ( .A1(n15760), .A2(n15761), .ZN(n10016) );
  NOR2_X1 U11257 ( .A1(n12819), .A2(n12818), .ZN(n12820) );
  AND2_X1 U11258 ( .A1(n9968), .A2(n9966), .ZN(n15956) );
  OAI21_X1 U11259 ( .B1(n14992), .B2(n12850), .A(n12849), .ZN(n12851) );
  NAND2_X1 U11260 ( .A1(n9836), .A2(n11610), .ZN(n15582) );
  AOI21_X1 U11261 ( .B1(n10269), .B2(n9924), .A(n15689), .ZN(n9923) );
  NAND2_X1 U11262 ( .A1(n15021), .A2(n9925), .ZN(n9928) );
  CLKBUF_X1 U11263 ( .A(n14720), .Z(n14735) );
  AND2_X1 U11264 ( .A1(n15009), .A2(n9926), .ZN(n9925) );
  NAND2_X1 U11265 ( .A1(n15019), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15009) );
  OR2_X1 U11266 ( .A1(n16164), .A2(n15230), .ZN(n16189) );
  NAND2_X1 U11267 ( .A1(n12754), .A2(n15052), .ZN(n15045) );
  NAND3_X1 U11268 ( .A1(n11663), .A2(n9817), .A3(n11669), .ZN(n16572) );
  NAND2_X1 U11269 ( .A1(n15063), .A2(n15062), .ZN(n15061) );
  AND2_X1 U11270 ( .A1(n9896), .A2(n9894), .ZN(n16757) );
  NOR3_X1 U11271 ( .A1(n11153), .A2(n11152), .A3(n12887), .ZN(n11156) );
  CLKBUF_X1 U11272 ( .A(n14807), .Z(n14849) );
  NOR2_X1 U11273 ( .A1(n15417), .A2(n15419), .ZN(n15418) );
  OAI21_X1 U11274 ( .B1(n17855), .B2(n16752), .A(n16751), .ZN(n9897) );
  NAND2_X1 U11275 ( .A1(n16062), .A2(n11659), .ZN(n10193) );
  XNOR2_X1 U11276 ( .A(n14526), .B(n10297), .ZN(n15417) );
  AND2_X1 U11277 ( .A1(n14526), .A2(n10297), .ZN(n14527) );
  AND2_X1 U11278 ( .A1(n9983), .A2(n9982), .ZN(n17855) );
  NAND2_X1 U11279 ( .A1(n9985), .A2(n9984), .ZN(n9983) );
  NAND2_X1 U11280 ( .A1(n14912), .A2(n14911), .ZN(n14850) );
  NAND2_X1 U11281 ( .A1(n10176), .A2(n10177), .ZN(n10175) );
  AND2_X1 U11282 ( .A1(n16173), .A2(n16745), .ZN(n11150) );
  AND2_X1 U11283 ( .A1(n15406), .A2(n15400), .ZN(n15399) );
  INV_X1 U11284 ( .A(n14016), .ZN(n10234) );
  NAND3_X1 U11285 ( .A1(n10201), .A2(n9788), .A3(n10200), .ZN(n14505) );
  NAND2_X1 U11286 ( .A1(n10140), .A2(n16292), .ZN(n15126) );
  AND2_X1 U11287 ( .A1(n10035), .A2(n15614), .ZN(n10034) );
  OR2_X1 U11288 ( .A1(n15415), .A2(n15416), .ZN(n15413) );
  XNOR2_X1 U11289 ( .A(n12829), .B(n10990), .ZN(n19435) );
  NAND2_X1 U11290 ( .A1(n9948), .A2(n15080), .ZN(n15071) );
  OR2_X1 U11291 ( .A1(n15439), .A2(n10202), .ZN(n10200) );
  OAI21_X1 U11292 ( .B1(n17904), .B2(n17905), .A(n9877), .ZN(n17881) );
  AOI21_X1 U11293 ( .B1(n10029), .B2(n10033), .A(n9761), .ZN(n10028) );
  XNOR2_X1 U11294 ( .A(n11606), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15614) );
  NAND2_X1 U11295 ( .A1(n16453), .A2(n11618), .ZN(n11606) );
  AOI21_X1 U11296 ( .B1(n10178), .B2(n19376), .A(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9916) );
  AND2_X1 U11297 ( .A1(n15227), .A2(n12744), .ZN(n15091) );
  AND2_X1 U11298 ( .A1(n17903), .A2(n9789), .ZN(n9877) );
  AND2_X1 U11299 ( .A1(n10031), .A2(n10030), .ZN(n10029) );
  NAND2_X1 U11300 ( .A1(n12070), .A2(n12069), .ZN(n12668) );
  NOR2_X1 U11301 ( .A1(n11597), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10112) );
  OAI22_X1 U11302 ( .A1(n15320), .A2(n12697), .B1(n13246), .B2(n12696), .ZN(
        n12698) );
  NOR3_X2 U11303 ( .A1(n15905), .A2(n15525), .A3(n10098), .ZN(n15527) );
  NAND2_X1 U11304 ( .A1(n11597), .A2(n11595), .ZN(n12957) );
  NAND2_X1 U11305 ( .A1(n18004), .A2(n18109), .ZN(n17971) );
  NOR3_X2 U11306 ( .A1(n11597), .A2(P2_EBX_REG_25__SCAN_IN), .A3(
        P2_EBX_REG_24__SCAN_IN), .ZN(n16454) );
  INV_X1 U11307 ( .A(n11468), .ZN(n10179) );
  OR2_X2 U11308 ( .A1(n11594), .A2(n11593), .ZN(n11597) );
  OR2_X1 U11309 ( .A1(n15379), .A2(n15555), .ZN(n15905) );
  AND2_X1 U11310 ( .A1(n11463), .A2(n11462), .ZN(n11468) );
  INV_X1 U11311 ( .A(n12149), .ZN(n12070) );
  NOR2_X1 U11312 ( .A1(n15987), .A2(n10093), .ZN(n15381) );
  CLKBUF_X1 U11313 ( .A(n14268), .Z(n14970) );
  OAI211_X1 U11314 ( .C1(n9884), .C2(n9885), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n9882), .ZN(n10169) );
  NAND2_X2 U11315 ( .A1(n12121), .A2(n12099), .ZN(n20582) );
  CLKBUF_X1 U11316 ( .A(n13595), .Z(n21021) );
  OAI22_X1 U11317 ( .A1(n11363), .A2(n13760), .B1(n19676), .B2(n11362), .ZN(
        n11370) );
  NOR2_X1 U11318 ( .A1(n18345), .A2(n18344), .ZN(n18343) );
  AND2_X1 U11319 ( .A1(n13374), .A2(n13285), .ZN(n13286) );
  OR2_X1 U11320 ( .A1(n13540), .A2(n13525), .ZN(n16371) );
  OR2_X1 U11321 ( .A1(n13540), .A2(n13524), .ZN(n15149) );
  OR2_X1 U11322 ( .A1(n13284), .A2(n13283), .ZN(n13373) );
  OR2_X1 U11323 ( .A1(n11137), .A2(n11318), .ZN(n18432) );
  OAI21_X1 U11324 ( .B1(n13282), .B2(n13281), .A(n10298), .ZN(n13375) );
  AND2_X1 U11325 ( .A1(n11136), .A2(n18442), .ZN(n11137) );
  INV_X1 U11326 ( .A(n18196), .ZN(n18211) );
  AND2_X1 U11327 ( .A1(n13248), .A2(n13200), .ZN(n21047) );
  AND2_X1 U11328 ( .A1(n13903), .A2(n11347), .ZN(n11348) );
  NAND2_X1 U11329 ( .A1(n11972), .A2(n11971), .ZN(n11998) );
  NAND2_X1 U11330 ( .A1(n13619), .A2(n10101), .ZN(n16622) );
  NOR2_X2 U11331 ( .A1(n19212), .A2(n16865), .ZN(n18199) );
  NAND2_X1 U11332 ( .A1(n11569), .A2(n11568), .ZN(n11571) );
  NAND2_X1 U11333 ( .A1(n9832), .A2(n10182), .ZN(n11327) );
  NOR2_X1 U11334 ( .A1(n19393), .A2(n19269), .ZN(n19261) );
  NAND2_X1 U11335 ( .A1(n11994), .A2(n11917), .ZN(n9937) );
  AND2_X1 U11336 ( .A1(n10049), .A2(n10048), .ZN(n19269) );
  NAND2_X1 U11337 ( .A1(n9690), .A2(n9770), .ZN(n9936) );
  CLKBUF_X1 U11338 ( .A(n12115), .Z(n20546) );
  NOR2_X1 U11339 ( .A1(n17711), .A2(n16202), .ZN(n17738) );
  AND2_X1 U11340 ( .A1(n11938), .A2(n11936), .ZN(n11991) );
  NAND2_X1 U11341 ( .A1(n11127), .A2(n11126), .ZN(n18148) );
  NAND2_X1 U11342 ( .A1(n11898), .A2(n11897), .ZN(n11938) );
  NOR2_X1 U11343 ( .A1(n14116), .A2(n19559), .ZN(n19607) );
  NAND2_X1 U11344 ( .A1(n11528), .A2(n9767), .ZN(n11562) );
  NOR2_X1 U11345 ( .A1(n14611), .A2(n19559), .ZN(n19608) );
  OR2_X1 U11346 ( .A1(n18164), .A2(n10159), .ZN(n10158) );
  NAND2_X1 U11347 ( .A1(n11602), .A2(n11532), .ZN(n11528) );
  AND2_X1 U11348 ( .A1(n10539), .A2(n10538), .ZN(n13189) );
  OR2_X1 U11349 ( .A1(n10652), .A2(n15732), .ZN(n10543) );
  NAND2_X2 U11350 ( .A1(n11129), .A2(n16746), .ZN(n18109) );
  NOR2_X1 U11351 ( .A1(n18173), .A2(n18172), .ZN(n18171) );
  XNOR2_X1 U11352 ( .A(n11121), .B(n18490), .ZN(n18173) );
  NAND2_X1 U11353 ( .A1(n9815), .A2(n10514), .ZN(n10530) );
  CLKBUF_X1 U11354 ( .A(n17840), .Z(n17849) );
  AND2_X1 U11355 ( .A1(n10156), .A2(n9746), .ZN(n11121) );
  NOR2_X1 U11356 ( .A1(n19212), .A2(n17848), .ZN(n17840) );
  AND2_X1 U11357 ( .A1(n9863), .A2(n9862), .ZN(n18984) );
  CLKBUF_X1 U11358 ( .A(n17581), .Z(n9669) );
  NAND2_X1 U11359 ( .A1(n13517), .A2(n11878), .ZN(n11879) );
  OR2_X1 U11360 ( .A1(n18186), .A2(n18185), .ZN(n10156) );
  NAND2_X1 U11361 ( .A1(n9861), .A2(n11275), .ZN(n9863) );
  OAI21_X1 U11362 ( .B1(n11254), .B2(n11250), .A(n12871), .ZN(n11262) );
  OR3_X1 U11363 ( .A1(n12793), .A2(n12792), .A3(n12789), .ZN(n12790) );
  OR2_X1 U11364 ( .A1(n13024), .A2(n20263), .ZN(n10514) );
  NOR2_X1 U11365 ( .A1(n12776), .A2(n13498), .ZN(n12795) );
  OR2_X1 U11366 ( .A1(n17785), .A2(n12870), .ZN(n9861) );
  NOR2_X1 U11367 ( .A1(n17735), .A2(n17744), .ZN(n11120) );
  AND2_X1 U11368 ( .A1(n11884), .A2(n13520), .ZN(n13349) );
  INV_X2 U11369 ( .A(n10512), .ZN(n10648) );
  NOR2_X1 U11370 ( .A1(n10512), .A2(n10535), .ZN(n10536) );
  CLKBUF_X1 U11371 ( .A(n13059), .Z(n13384) );
  NAND2_X1 U11372 ( .A1(n11418), .A2(n11417), .ZN(n11426) );
  NAND2_X1 U11373 ( .A1(n12788), .A2(n13303), .ZN(n12806) );
  AND2_X1 U11374 ( .A1(n10458), .A2(n10498), .ZN(n13117) );
  MUX2_X1 U11375 ( .A(P2_EBX_REG_4__SCAN_IN), .B(n11005), .S(n10792), .Z(
        n11427) );
  AND2_X1 U11376 ( .A1(n11874), .A2(n13954), .ZN(n13209) );
  NAND2_X1 U11377 ( .A1(n11900), .A2(n14265), .ZN(n10225) );
  NOR2_X1 U11378 ( .A1(n10480), .A2(n10472), .ZN(n13329) );
  INV_X1 U11379 ( .A(n9663), .ZN(n18578) );
  NAND2_X1 U11380 ( .A1(n10498), .A2(n10497), .ZN(n16662) );
  AND2_X1 U11381 ( .A1(n9888), .A2(n9887), .ZN(n17725) );
  AND3_X1 U11382 ( .A1(n10486), .A2(n10499), .A3(n10457), .ZN(n10498) );
  INV_X1 U11383 ( .A(n11833), .ZN(n11875) );
  NAND2_X1 U11384 ( .A1(n13875), .A2(n11834), .ZN(n14267) );
  CLKBUF_X1 U11385 ( .A(n11834), .Z(n13967) );
  INV_X1 U11386 ( .A(n10476), .ZN(n13054) );
  OR2_X1 U11387 ( .A1(n10754), .A2(n10753), .ZN(n11380) );
  OR2_X1 U11388 ( .A1(n10733), .A2(n10732), .ZN(n10999) );
  NAND2_X1 U11389 ( .A1(n11117), .A2(n11116), .ZN(n18205) );
  AND2_X1 U11390 ( .A1(n11061), .A2(n10308), .ZN(n17735) );
  OAI211_X1 U11391 ( .C1(n14198), .C2(n14190), .A(n11082), .B(n11081), .ZN(
        n17729) );
  OR2_X2 U11392 ( .A1(n10825), .A2(n10824), .ZN(n11618) );
  INV_X1 U11393 ( .A(n13514), .ZN(n15338) );
  OR2_X1 U11394 ( .A1(n10791), .A2(n10790), .ZN(n11460) );
  NAND2_X2 U11395 ( .A1(n10319), .A2(n11759), .ZN(n14265) );
  NOR2_X1 U11396 ( .A1(n10084), .A2(n10320), .ZN(n10126) );
  OR2_X1 U11397 ( .A1(n11859), .A2(n10085), .ZN(n10084) );
  INV_X2 U11398 ( .A(n13116), .ZN(n10499) );
  NAND2_X1 U11399 ( .A1(n9819), .A2(n9818), .ZN(n10476) );
  AOI211_X1 U11400 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n11090), .B(n11089), .ZN(n11091) );
  AND4_X1 U11401 ( .A1(n9726), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n11852) );
  NAND2_X2 U11402 ( .A1(n9821), .A2(n9820), .ZN(n10477) );
  AND4_X1 U11403 ( .A1(n11804), .A2(n11803), .A3(n11802), .A4(n11801), .ZN(
        n11815) );
  NAND2_X1 U11404 ( .A1(n11756), .A2(n9714), .ZN(n11757) );
  OR2_X2 U11405 ( .A1(n16814), .A2(n16760), .ZN(n16817) );
  NAND2_X1 U11406 ( .A1(n10429), .A2(n10680), .ZN(n10430) );
  AND4_X1 U11407 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11733) );
  AND4_X1 U11408 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11756) );
  AND4_X1 U11409 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11872) );
  AND4_X1 U11410 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11873) );
  AND4_X1 U11411 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .ZN(
        n10429) );
  NAND2_X1 U11412 ( .A1(n18905), .A2(n18853), .ZN(n18776) );
  INV_X1 U11413 ( .A(n17468), .ZN(n9670) );
  AND2_X1 U11414 ( .A1(n10403), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10404) );
  AND3_X1 U11415 ( .A1(n10411), .A2(n10680), .A3(n10410), .ZN(n10414) );
  AND2_X2 U11416 ( .A1(n9660), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14406) );
  INV_X2 U11417 ( .A(n17468), .ZN(n17450) );
  NAND2_X2 U11418 ( .A1(n19151), .A2(n19081), .ZN(n19140) );
  INV_X2 U11419 ( .A(n12634), .ZN(n12365) );
  INV_X2 U11420 ( .A(n9709), .ZN(n17540) );
  BUF_X2 U11421 ( .A(n14466), .Z(n9659) );
  INV_X1 U11422 ( .A(n10316), .ZN(n9662) );
  INV_X1 U11423 ( .A(n12637), .ZN(n12615) );
  NAND2_X2 U11424 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20274), .ZN(n20173) );
  INV_X1 U11425 ( .A(n19156), .ZN(n19065) );
  NAND2_X2 U11426 ( .A1(n20274), .A2(n20133), .ZN(n20176) );
  NOR2_X1 U11427 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18544), .ZN(n18905) );
  INV_X2 U11428 ( .A(n16850), .ZN(U215) );
  INV_X1 U11429 ( .A(n12492), .ZN(n12616) );
  INV_X4 U11430 ( .A(n11036), .ZN(n17433) );
  INV_X1 U11431 ( .A(n11023), .ZN(n11025) );
  INV_X2 U11432 ( .A(n21053), .ZN(n21013) );
  OR2_X2 U11434 ( .A1(n11018), .A2(n19020), .ZN(n17388) );
  OR3_X2 U11435 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n17247), .ZN(n11241) );
  AND2_X1 U11436 ( .A1(n11725), .A2(n11719), .ZN(n11769) );
  OR2_X2 U11437 ( .A1(n11023), .A2(n11018), .ZN(n10316) );
  AND2_X2 U11438 ( .A1(n14601), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14398) );
  AND2_X2 U11439 ( .A1(n14594), .A2(n10680), .ZN(n10765) );
  NAND2_X1 U11440 ( .A1(n10303), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11036) );
  OR2_X1 U11441 ( .A1(n11022), .A2(n11023), .ZN(n9710) );
  INV_X2 U11442 ( .A(n19220), .ZN(n19151) );
  INV_X1 U11443 ( .A(n12544), .ZN(n12643) );
  AND3_X1 U11444 ( .A1(n10356), .A2(n10069), .A3(n10067), .ZN(n10352) );
  INV_X2 U11445 ( .A(n16853), .ZN(n16855) );
  OR3_X2 U11446 ( .A1(n17247), .A2(n19177), .A3(n19167), .ZN(n9709) );
  INV_X1 U11447 ( .A(n12544), .ZN(n9657) );
  NAND2_X1 U11448 ( .A1(n19167), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11018) );
  AND2_X1 U11449 ( .A1(n10226), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13362) );
  AND2_X2 U11450 ( .A1(n13381), .A2(n13923), .ZN(n14601) );
  NOR2_X2 U11451 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13584) );
  AND2_X1 U11452 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13358) );
  AND2_X1 U11453 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U11454 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U11455 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19026) );
  INV_X2 U11456 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19167) );
  NAND2_X1 U11457 ( .A1(n13379), .A2(n11348), .ZN(n11447) );
  NAND2_X1 U11458 ( .A1(n13379), .A2(n11346), .ZN(n19920) );
  NAND2_X2 U11459 ( .A1(n11469), .A2(n11468), .ZN(n11502) );
  NOR2_X2 U11460 ( .A1(n17357), .A2(n17384), .ZN(n17372) );
  OAI22_X1 U11461 ( .A1(n11700), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n20256), 
        .B2(n10651), .ZN(n19379) );
  AND2_X1 U11462 ( .A1(n16024), .A2(n15941), .ZN(n16508) );
  OR2_X1 U11463 ( .A1(n15694), .A2(n9822), .ZN(n15869) );
  BUF_X2 U11464 ( .A(n11352), .Z(n9675) );
  XNOR2_X1 U11465 ( .A(n11329), .B(n11328), .ZN(n11352) );
  NOR2_X4 U11466 ( .A1(n13749), .A2(n13750), .ZN(n16403) );
  OR2_X2 U11467 ( .A1(n13735), .A2(n13734), .ZN(n13749) );
  INV_X2 U11468 ( .A(n16071), .ZN(n14602) );
  INV_X2 U11469 ( .A(n16071), .ZN(n9676) );
  NAND2_X1 U11470 ( .A1(n10691), .A2(n10468), .ZN(n9906) );
  INV_X4 U11471 ( .A(n10468), .ZN(n16663) );
  INV_X1 U11472 ( .A(n12492), .ZN(n9666) );
  NAND2_X1 U11473 ( .A1(n11726), .A2(n13362), .ZN(n12637) );
  NAND2_X2 U11474 ( .A1(n11501), .A2(n11500), .ZN(n11660) );
  INV_X2 U11475 ( .A(n12544), .ZN(n9668) );
  NAND2_X1 U11476 ( .A1(n13584), .A2(n11724), .ZN(n12544) );
  NAND2_X1 U11477 ( .A1(n13958), .A2(n13499), .ZN(n13531) );
  NOR2_X2 U11478 ( .A1(n11136), .A2(n18442), .ZN(n11318) );
  NAND2_X2 U11479 ( .A1(n10484), .A2(n16663), .ZN(n10673) );
  AND2_X2 U11480 ( .A1(n13381), .A2(n13923), .ZN(n9671) );
  AND2_X1 U11482 ( .A1(n10365), .A2(n16653), .ZN(n9673) );
  AND2_X1 U11483 ( .A1(n10365), .A2(n16653), .ZN(n9674) );
  AND2_X4 U11484 ( .A1(n10366), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10397) );
  INV_X1 U11485 ( .A(n9676), .ZN(n9677) );
  INV_X1 U11486 ( .A(n13029), .ZN(n10478) );
  AOI21_X1 U11487 ( .B1(n13088), .B2(n13207), .A(n13515), .ZN(n11878) );
  OAI22_X1 U11488 ( .A1(n14369), .A2(n19647), .B1(n19569), .B2(n11341), .ZN(
        n11342) );
  NAND2_X1 U11489 ( .A1(n13088), .A2(n13958), .ZN(n13293) );
  NOR2_X1 U11490 ( .A1(n14002), .A2(n21045), .ZN(n11932) );
  NAND3_X1 U11491 ( .A1(n10037), .A2(n10034), .A3(n10036), .ZN(n15593) );
  INV_X1 U11492 ( .A(n11655), .ZN(n10279) );
  NAND2_X1 U11493 ( .A1(n9881), .A2(n18315), .ZN(n9885) );
  NOR2_X1 U11494 ( .A1(n17717), .A2(n11103), .ZN(n11129) );
  INV_X2 U11495 ( .A(n11618), .ZN(n11667) );
  AOI21_X1 U11496 ( .B1(n9678), .B2(n10285), .A(n15654), .ZN(n9918) );
  CLKBUF_X1 U11497 ( .A(n11847), .Z(n12410) );
  AND2_X1 U11499 ( .A1(n11424), .A2(n11420), .ZN(n11418) );
  MUX2_X1 U11500 ( .A(n11003), .B(n13635), .S(n10495), .Z(n11417) );
  NAND2_X1 U11501 ( .A1(n10481), .A2(n10480), .ZN(n10482) );
  NAND2_X1 U11502 ( .A1(n11125), .A2(n17720), .ZN(n11103) );
  OAI21_X1 U11503 ( .B1(n11259), .B2(n19006), .A(n11258), .ZN(n11273) );
  INV_X1 U11504 ( .A(n14017), .ZN(n10240) );
  NAND2_X1 U11505 ( .A1(n10240), .A2(n14010), .ZN(n10239) );
  INV_X1 U11506 ( .A(n13614), .ZN(n12137) );
  OR2_X1 U11507 ( .A1(n13967), .A2(n21042), .ZN(n12260) );
  OR2_X1 U11508 ( .A1(n13875), .A2(n21042), .ZN(n12663) );
  NOR2_X1 U11509 ( .A1(n11713), .A2(n11712), .ZN(n11734) );
  INV_X1 U11510 ( .A(n12780), .ZN(n13344) );
  NAND2_X1 U11511 ( .A1(n12023), .A2(n12022), .ZN(n20581) );
  OR2_X1 U11512 ( .A1(n13514), .A2(n21045), .ZN(n12007) );
  INV_X1 U11513 ( .A(n12788), .ZN(n12796) );
  NOR2_X1 U11514 ( .A1(n10690), .A2(n19603), .ZN(n10458) );
  INV_X1 U11515 ( .A(n14139), .ZN(n9830) );
  NAND2_X1 U11516 ( .A1(n10474), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10532) );
  NOR2_X1 U11517 ( .A1(n15511), .A2(n15510), .ZN(n10977) );
  NOR2_X1 U11518 ( .A1(n15593), .A2(n10190), .ZN(n11609) );
  NOR2_X1 U11519 ( .A1(n10258), .A2(n15462), .ZN(n10257) );
  INV_X1 U11520 ( .A(n15385), .ZN(n10258) );
  INV_X1 U11521 ( .A(n13910), .ZN(n10102) );
  INV_X1 U11522 ( .A(n11430), .ZN(n9903) );
  NAND2_X1 U11523 ( .A1(n11380), .A2(n10493), .ZN(n11381) );
  NOR2_X1 U11524 ( .A1(n10719), .A2(n10718), .ZN(n10741) );
  NOR2_X1 U11525 ( .A1(n17976), .A2(n10002), .ZN(n10001) );
  NAND2_X1 U11526 ( .A1(n18029), .A2(n18398), .ZN(n18040) );
  NAND2_X1 U11527 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18127), .ZN(
        n11312) );
  AOI21_X1 U11528 ( .B1(n19014), .B2(n9716), .A(n16106), .ZN(n16201) );
  CLKBUF_X1 U11529 ( .A(n13088), .Z(n13423) );
  NOR2_X1 U11530 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  INV_X1 U11531 ( .A(n20276), .ZN(n13511) );
  AND2_X1 U11532 ( .A1(n21042), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12861) );
  AND2_X1 U11533 ( .A1(n10661), .A2(n10660), .ZN(n11690) );
  CLKBUF_X2 U11534 ( .A(n10737), .Z(n10989) );
  NAND2_X1 U11535 ( .A1(n10205), .A2(n10203), .ZN(n10202) );
  INV_X1 U11536 ( .A(n15438), .ZN(n10203) );
  NOR2_X1 U11537 ( .A1(n10691), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13056) );
  NAND2_X1 U11538 ( .A1(n10196), .A2(n15765), .ZN(n10195) );
  NAND2_X1 U11539 ( .A1(n9683), .A2(n11588), .ZN(n10031) );
  NOR2_X1 U11540 ( .A1(n10184), .A2(n15659), .ZN(n10185) );
  OAI21_X1 U11541 ( .B1(n16014), .B2(n10275), .A(n10272), .ZN(n16523) );
  INV_X1 U11542 ( .A(n10276), .ZN(n10275) );
  AOI21_X1 U11543 ( .B1(n10276), .B2(n10274), .A(n10273), .ZN(n10272) );
  NOR2_X1 U11544 ( .A1(n10189), .A2(n15998), .ZN(n10276) );
  INV_X1 U11545 ( .A(n12823), .ZN(n10253) );
  NAND2_X1 U11546 ( .A1(n15582), .A2(n9833), .ZN(n9835) );
  NOR2_X1 U11547 ( .A1(n15569), .A2(n9834), .ZN(n9833) );
  INV_X1 U11548 ( .A(n15580), .ZN(n9834) );
  OAI211_X1 U11549 ( .C1(n10028), .C2(n9912), .A(n9910), .B(n9720), .ZN(n11600) );
  OAI21_X1 U11550 ( .B1(n10265), .B2(n10271), .A(n10263), .ZN(n15672) );
  AND2_X1 U11551 ( .A1(n10266), .A2(n10264), .ZN(n10263) );
  NAND2_X1 U11552 ( .A1(n10270), .A2(n15657), .ZN(n10264) );
  AND2_X1 U11553 ( .A1(n15673), .A2(n10267), .ZN(n10266) );
  NAND2_X1 U11554 ( .A1(n10265), .A2(n15656), .ZN(n10269) );
  NAND2_X1 U11555 ( .A1(n16525), .A2(n9678), .ZN(n9917) );
  INV_X1 U11556 ( .A(n10288), .ZN(n10287) );
  OR2_X2 U11557 ( .A1(n15720), .A2(n15721), .ZN(n16014) );
  NAND2_X1 U11558 ( .A1(n11428), .A2(n10302), .ZN(n9900) );
  AND2_X1 U11559 ( .A1(n13128), .A2(n13332), .ZN(n13153) );
  INV_X1 U11560 ( .A(n19379), .ZN(n10362) );
  NAND2_X1 U11561 ( .A1(n10173), .A2(n10172), .ZN(n16174) );
  NAND2_X1 U11562 ( .A1(n11150), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10172) );
  NAND2_X1 U11563 ( .A1(n10175), .A2(n10174), .ZN(n10173) );
  AND2_X1 U11564 ( .A1(n9699), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10174) );
  NAND2_X1 U11565 ( .A1(n17971), .A2(n11144), .ZN(n17911) );
  NAND2_X1 U11566 ( .A1(n18011), .A2(n11141), .ZN(n11143) );
  AND2_X1 U11567 ( .A1(n18040), .A2(n18109), .ZN(n10168) );
  NAND2_X1 U11568 ( .A1(n11138), .A2(n10171), .ZN(n10170) );
  NAND2_X1 U11569 ( .A1(n18109), .A2(n11135), .ZN(n10171) );
  NAND2_X1 U11570 ( .A1(n9881), .A2(n9879), .ZN(n9882) );
  NOR2_X1 U11571 ( .A1(n9883), .A2(n9880), .ZN(n9879) );
  NAND2_X1 U11572 ( .A1(n15757), .A2(n16589), .ZN(n11703) );
  NAND2_X1 U11573 ( .A1(n11719), .A2(n13358), .ZN(n12603) );
  NAND2_X1 U11574 ( .A1(n13362), .A2(n13584), .ZN(n12608) );
  INV_X1 U11575 ( .A(n12802), .ZN(n12782) );
  NOR2_X1 U11576 ( .A1(n10192), .A2(n10191), .ZN(n11458) );
  NOR2_X1 U11577 ( .A1(n19895), .A2(n11439), .ZN(n10191) );
  NOR2_X1 U11578 ( .A1(n10512), .A2(n10459), .ZN(n10460) );
  OR2_X1 U11579 ( .A1(n11176), .A2(n11177), .ZN(n11169) );
  AOI22_X1 U11580 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11222) );
  AND3_X1 U11581 ( .A1(n13209), .A2(n11875), .A3(n14267), .ZN(n11876) );
  NAND2_X1 U11582 ( .A1(n10228), .A2(n10227), .ZN(n12149) );
  AND2_X1 U11583 ( .A1(n12129), .A2(n12139), .ZN(n10227) );
  NAND2_X1 U11584 ( .A1(n15224), .A2(n10155), .ZN(n9954) );
  NOR2_X1 U11585 ( .A1(n14322), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n10127) );
  AND2_X1 U11586 ( .A1(n13308), .A2(n14265), .ZN(n10147) );
  AOI22_X1 U11587 ( .A1(n11891), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11890), 
        .B2(n11889), .ZN(n11892) );
  OR2_X1 U11588 ( .A1(n12634), .A2(n11736), .ZN(n11737) );
  NOR2_X1 U11589 ( .A1(n12782), .A2(n13083), .ZN(n12793) );
  NAND2_X1 U11590 ( .A1(n13212), .A2(n12775), .ZN(n12792) );
  INV_X1 U11591 ( .A(n11464), .ZN(n10111) );
  NOR2_X1 U11592 ( .A1(n10100), .A2(n15904), .ZN(n10099) );
  INV_X1 U11593 ( .A(n12932), .ZN(n10100) );
  NOR2_X1 U11594 ( .A1(n20009), .A2(n11396), .ZN(n11399) );
  AOI21_X1 U11595 ( .B1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20229), .A(
        n10654), .ZN(n10669) );
  NOR2_X1 U11596 ( .A1(n11677), .A2(n11419), .ZN(n10654) );
  INV_X1 U11597 ( .A(n9850), .ZN(n9849) );
  OAI211_X1 U11598 ( .C1(n17557), .C2(n11051), .A(n9852), .B(n9851), .ZN(n9850) );
  NAND2_X1 U11599 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n9851) );
  NAND2_X1 U11600 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n9852) );
  NAND2_X1 U11601 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n9853) );
  AND2_X1 U11602 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  NAND2_X1 U11603 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n9858) );
  NAND2_X1 U11604 ( .A1(n17541), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n9859) );
  NAND2_X1 U11605 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n9855) );
  NOR2_X1 U11606 ( .A1(n17725), .A2(n11123), .ZN(n11125) );
  NOR2_X1 U11607 ( .A1(n17725), .A2(n11296), .ZN(n11285) );
  INV_X1 U11608 ( .A(n14771), .ZN(n12402) );
  NOR2_X1 U11609 ( .A1(n14888), .A2(n14800), .ZN(n10230) );
  INV_X1 U11610 ( .A(n12665), .ZN(n12627) );
  INV_X1 U11611 ( .A(n12260), .ZN(n12292) );
  NAND2_X1 U11612 ( .A1(n10132), .A2(n14325), .ZN(n10131) );
  NAND2_X1 U11613 ( .A1(n14814), .A2(n14826), .ZN(n10137) );
  INV_X1 U11614 ( .A(n12717), .ZN(n9930) );
  NAND2_X1 U11615 ( .A1(n9733), .A2(n12668), .ZN(n12727) );
  OR2_X1 U11616 ( .A1(n11951), .A2(n11950), .ZN(n12685) );
  NAND2_X1 U11617 ( .A1(n13523), .A2(n11907), .ZN(n11936) );
  AND2_X1 U11618 ( .A1(n11906), .A2(n11905), .ZN(n11907) );
  INV_X1 U11619 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13361) );
  NAND2_X1 U11620 ( .A1(n14002), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12008) );
  NAND2_X1 U11621 ( .A1(n10116), .A2(n10115), .ZN(n11544) );
  INV_X1 U11622 ( .A(n11542), .ZN(n10115) );
  INV_X1 U11623 ( .A(n15446), .ZN(n10218) );
  INV_X1 U11624 ( .A(n14031), .ZN(n10090) );
  NOR2_X1 U11625 ( .A1(n20258), .A2(n19603), .ZN(n14549) );
  NOR2_X1 U11626 ( .A1(n15629), .A2(n10062), .ZN(n10061) );
  INV_X1 U11627 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U11628 ( .A1(n16564), .A2(n10066), .ZN(n10065) );
  INV_X1 U11629 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10066) );
  INV_X1 U11630 ( .A(n13546), .ZN(n10252) );
  NOR2_X1 U11631 ( .A1(n16592), .A2(n10070), .ZN(n10069) );
  AND2_X1 U11632 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  INV_X1 U11633 ( .A(n15489), .ZN(n10107) );
  AND2_X1 U11634 ( .A1(n15595), .A2(n15783), .ZN(n10190) );
  INV_X1 U11635 ( .A(n15592), .ZN(n9908) );
  NOR2_X1 U11636 ( .A1(n12929), .A2(n11667), .ZN(n11576) );
  INV_X1 U11637 ( .A(n15452), .ZN(n10256) );
  AND2_X1 U11638 ( .A1(n13825), .A2(n13936), .ZN(n10249) );
  NOR2_X1 U11639 ( .A1(n16504), .A2(n10291), .ZN(n10290) );
  NOR2_X1 U11640 ( .A1(n10292), .A2(n15653), .ZN(n10291) );
  NAND2_X1 U11641 ( .A1(n10289), .A2(n16503), .ZN(n10288) );
  NAND2_X1 U11642 ( .A1(n10290), .A2(n15653), .ZN(n10289) );
  AND2_X1 U11643 ( .A1(n9723), .A2(n13485), .ZN(n10251) );
  INV_X1 U11644 ( .A(n10178), .ZN(n9902) );
  INV_X1 U11645 ( .A(n13288), .ZN(n10261) );
  OAI211_X1 U11646 ( .C1(n11416), .C2(n9962), .A(n9961), .B(n9773), .ZN(n11651) );
  NAND2_X1 U11647 ( .A1(n11415), .A2(n9963), .ZN(n9962) );
  NAND3_X1 U11648 ( .A1(n9960), .A2(n11416), .A3(n9963), .ZN(n9961) );
  INV_X1 U11649 ( .A(n14027), .ZN(n10555) );
  NAND2_X1 U11650 ( .A1(n9816), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9815) );
  NAND2_X1 U11651 ( .A1(n13278), .A2(n13277), .ZN(n13284) );
  AND2_X1 U11652 ( .A1(n14549), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13283) );
  INV_X1 U11653 ( .A(n13631), .ZN(n10092) );
  NAND2_X1 U11654 ( .A1(n10385), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9819) );
  NAND2_X1 U11655 ( .A1(n10386), .A2(n10680), .ZN(n9818) );
  NAND2_X1 U11656 ( .A1(n11688), .A2(n11687), .ZN(n13121) );
  OAI21_X1 U11657 ( .B1(n11686), .B2(n11685), .A(n11684), .ZN(n11688) );
  NAND2_X1 U11658 ( .A1(n9743), .A2(n9682), .ZN(n9973) );
  OR2_X1 U11659 ( .A1(n9710), .A2(n17527), .ZN(n10305) );
  INV_X1 U11660 ( .A(n10163), .ZN(n10162) );
  NAND2_X1 U11661 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9986) );
  NAND2_X1 U11662 ( .A1(n18318), .A2(n18011), .ZN(n17954) );
  NAND2_X1 U11663 ( .A1(n18136), .A2(n9681), .ZN(n10165) );
  NAND2_X1 U11664 ( .A1(n18148), .A2(n9681), .ZN(n10166) );
  NOR2_X1 U11665 ( .A1(n11249), .A2(n9989), .ZN(n12871) );
  XNOR2_X1 U11666 ( .A(n11302), .B(n11103), .ZN(n11128) );
  XNOR2_X1 U11667 ( .A(n11123), .B(n9886), .ZN(n11124) );
  INV_X1 U11668 ( .A(n17725), .ZN(n9886) );
  XNOR2_X1 U11669 ( .A(n11104), .B(n17735), .ZN(n11119) );
  INV_X1 U11670 ( .A(n11284), .ZN(n11104) );
  NOR3_X1 U11671 ( .A1(n11275), .A2(n11274), .A3(n11273), .ZN(n12872) );
  INV_X1 U11672 ( .A(n9863), .ZN(n16104) );
  NOR2_X1 U11673 ( .A1(n13954), .A2(n13308), .ZN(n13870) );
  AND2_X1 U11674 ( .A1(n10236), .A2(n14010), .ZN(n10232) );
  AND2_X1 U11675 ( .A1(n14108), .A2(n14075), .ZN(n10236) );
  NAND2_X1 U11676 ( .A1(n13299), .A2(n13298), .ZN(n13435) );
  OR2_X1 U11677 ( .A1(n16159), .A2(n13295), .ZN(n13299) );
  NAND2_X1 U11678 ( .A1(n13499), .A2(n13498), .ZN(n13246) );
  INV_X1 U11679 ( .A(n12663), .ZN(n12862) );
  AND2_X1 U11680 ( .A1(n12542), .A2(n10242), .ZN(n14679) );
  NOR2_X1 U11681 ( .A1(n10244), .A2(n14708), .ZN(n10242) );
  NAND2_X1 U11682 ( .A1(n10246), .A2(n10245), .ZN(n10244) );
  INV_X1 U11683 ( .A(n14681), .ZN(n10245) );
  NAND2_X1 U11684 ( .A1(n10040), .A2(n10039), .ZN(n10038) );
  NOR2_X1 U11685 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10039) );
  INV_X1 U11686 ( .A(n16184), .ZN(n10040) );
  NOR2_X1 U11687 ( .A1(n14016), .A2(n10239), .ZN(n10238) );
  NAND2_X1 U11688 ( .A1(n12151), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12150) );
  NOR2_X1 U11689 ( .A1(n14016), .A2(n14017), .ZN(n14105) );
  OAI21_X1 U11690 ( .B1(n15320), .B2(n12260), .A(n12127), .ZN(n13656) );
  INV_X1 U11691 ( .A(n15181), .ZN(n9926) );
  NOR2_X1 U11692 ( .A1(n15009), .A2(n15182), .ZN(n12755) );
  NAND2_X1 U11693 ( .A1(n15045), .A2(n15018), .ZN(n15036) );
  NAND2_X1 U11694 ( .A1(n15071), .A2(n15236), .ZN(n12747) );
  NAND2_X1 U11695 ( .A1(n15126), .A2(n12738), .ZN(n12740) );
  OAI211_X1 U11696 ( .C1(n10144), .C2(n10145), .A(n10143), .B(n13814), .ZN(
        n9932) );
  OR2_X1 U11697 ( .A1(n9708), .A2(n10146), .ZN(n10144) );
  OR2_X1 U11698 ( .A1(n13704), .A2(n9708), .ZN(n10143) );
  INV_X1 U11699 ( .A(n12699), .ZN(n10146) );
  NAND3_X1 U11700 ( .A1(n13871), .A2(n13870), .A3(n9933), .ZN(n13528) );
  NOR2_X1 U11701 ( .A1(n13499), .A2(n13958), .ZN(n9933) );
  NOR2_X1 U11702 ( .A1(n13528), .A2(n14267), .ZN(n13515) );
  AND4_X1 U11703 ( .A1(n11723), .A2(n11722), .A3(n11721), .A4(n11720), .ZN(
        n11732) );
  OR2_X1 U11704 ( .A1(n11998), .A2(n11997), .ZN(n11999) );
  INV_X1 U11705 ( .A(n20581), .ZN(n13942) );
  INV_X1 U11706 ( .A(n20464), .ZN(n15326) );
  AND2_X1 U11707 ( .A1(n11835), .A2(n13498), .ZN(n10149) );
  INV_X1 U11708 ( .A(n20521), .ZN(n20759) );
  NAND2_X1 U11709 ( .A1(n15321), .A2(n20582), .ZN(n21020) );
  OR2_X1 U11710 ( .A1(n20582), .A2(n13942), .ZN(n21022) );
  NOR2_X1 U11711 ( .A1(n20755), .A2(n15326), .ZN(n20849) );
  NAND2_X2 U11712 ( .A1(n12008), .A2(n12007), .ZN(n12802) );
  AND2_X1 U11713 ( .A1(n12801), .A2(n12800), .ZN(n12805) );
  OR2_X1 U11714 ( .A1(n12799), .A2(n12798), .ZN(n12801) );
  AOI21_X1 U11715 ( .B1(n12795), .B2(n13084), .A(n12794), .ZN(n10078) );
  NAND2_X1 U11716 ( .A1(n11604), .A2(n10119), .ZN(n11615) );
  INV_X1 U11717 ( .A(n15627), .ZN(n10054) );
  NAND2_X1 U11718 ( .A1(n11011), .A2(n11589), .ZN(n11594) );
  NAND2_X1 U11719 ( .A1(n9658), .A2(n10050), .ZN(n10049) );
  NAND2_X1 U11720 ( .A1(n19289), .A2(n15697), .ZN(n10050) );
  NOR2_X2 U11721 ( .A1(n11562), .A2(n11010), .ZN(n11552) );
  NAND2_X2 U11722 ( .A1(n11515), .A2(n10792), .ZN(n11602) );
  NOR2_X1 U11723 ( .A1(n11426), .A2(n11427), .ZN(n11465) );
  AND2_X1 U11724 ( .A1(n9697), .A2(n13605), .ZN(n10217) );
  OAI21_X1 U11725 ( .B1(n15396), .B2(n10208), .A(n10206), .ZN(n10211) );
  INV_X1 U11726 ( .A(n10213), .ZN(n10208) );
  AOI21_X1 U11727 ( .B1(n10213), .B2(n10207), .A(n14588), .ZN(n10206) );
  INV_X1 U11728 ( .A(n15409), .ZN(n10207) );
  NOR2_X1 U11729 ( .A1(n15392), .A2(n10214), .ZN(n10213) );
  INV_X1 U11730 ( .A(n15397), .ZN(n10214) );
  NAND2_X1 U11731 ( .A1(n14458), .A2(n9786), .ZN(n10201) );
  AND2_X1 U11732 ( .A1(n14458), .A2(n14483), .ZN(n10204) );
  XNOR2_X1 U11733 ( .A(n14457), .B(n14456), .ZN(n15439) );
  NOR2_X1 U11734 ( .A1(n15439), .A2(n15438), .ZN(n15437) );
  NOR2_X1 U11735 ( .A1(n16622), .A2(n16621), .ZN(n16007) );
  XNOR2_X1 U11736 ( .A(n10326), .B(n10325), .ZN(n11700) );
  NAND2_X1 U11737 ( .A1(n10328), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10331) );
  NAND2_X1 U11738 ( .A1(n11588), .A2(n9725), .ZN(n10033) );
  AND2_X1 U11739 ( .A1(n15982), .A2(n16522), .ZN(n10292) );
  NAND4_X1 U11740 ( .A1(n9941), .A2(n9829), .A3(n9828), .A4(n9827), .ZN(n16063) );
  NAND2_X1 U11741 ( .A1(n15582), .A2(n15580), .ZN(n15566) );
  NAND2_X1 U11742 ( .A1(n10194), .A2(n10196), .ZN(n15619) );
  INV_X1 U11743 ( .A(n15623), .ZN(n10035) );
  INV_X1 U11744 ( .A(n15634), .ZN(n9844) );
  NAND2_X1 U11745 ( .A1(n11600), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9845) );
  INV_X1 U11746 ( .A(n15871), .ZN(n10030) );
  INV_X1 U11747 ( .A(n15658), .ZN(n10267) );
  NAND2_X1 U11748 ( .A1(n9917), .A2(n9765), .ZN(n10265) );
  INV_X1 U11749 ( .A(n15703), .ZN(n9922) );
  AOI21_X1 U11750 ( .B1(n16525), .B2(n10290), .A(n10288), .ZN(n10280) );
  AND2_X1 U11751 ( .A1(n10582), .A2(n10581), .ZN(n13607) );
  AND3_X1 U11752 ( .A1(n10842), .A2(n10841), .A3(n10840), .ZN(n13910) );
  AND2_X1 U11753 ( .A1(n13619), .A2(n9762), .ZN(n16025) );
  NAND2_X1 U11754 ( .A1(n16047), .A2(n16048), .ZN(n9839) );
  AOI21_X1 U11755 ( .B1(n10022), .B2(n10024), .A(n10020), .ZN(n10019) );
  INV_X1 U11756 ( .A(n10027), .ZN(n10024) );
  AOI21_X1 U11757 ( .B1(n13637), .B2(n11618), .A(n15732), .ZN(n10027) );
  NAND2_X1 U11758 ( .A1(n13981), .A2(n13637), .ZN(n10021) );
  NOR2_X1 U11759 ( .A1(n10026), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10025) );
  CLKBUF_X1 U11760 ( .A(n10691), .Z(n16700) );
  NAND2_X1 U11761 ( .A1(n13284), .A2(n13283), .ZN(n13374) );
  NAND2_X1 U11762 ( .A1(n10087), .A2(n10091), .ZN(n13633) );
  NAND2_X1 U11763 ( .A1(n13050), .A2(n13270), .ZN(n13053) );
  AOI21_X1 U11764 ( .B1(n13174), .B2(n13270), .A(n13173), .ZN(n13175) );
  XNOR2_X1 U11765 ( .A(n13171), .B(n13181), .ZN(n13176) );
  INV_X1 U11766 ( .A(n11340), .ZN(n9842) );
  AND2_X1 U11767 ( .A1(n20204), .A2(n20234), .ZN(n19756) );
  AND2_X1 U11768 ( .A1(n20204), .A2(n19500), .ZN(n19788) );
  AND2_X1 U11769 ( .A1(n13903), .A2(n11354), .ZN(n11355) );
  NAND2_X1 U11770 ( .A1(n19854), .A2(n19500), .ZN(n19970) );
  OR2_X1 U11771 ( .A1(n20210), .A2(n20222), .ZN(n20049) );
  AND2_X1 U11772 ( .A1(n11694), .A2(n20256), .ZN(n20053) );
  OR2_X1 U11773 ( .A1(n20190), .A2(n11693), .ZN(n11694) );
  INV_X2 U11774 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20256) );
  NOR2_X1 U11775 ( .A1(n16909), .A2(n16910), .ZN(n16908) );
  INV_X1 U11776 ( .A(n18077), .ZN(n10006) );
  INV_X1 U11777 ( .A(n16885), .ZN(n17158) );
  INV_X1 U11778 ( .A(n18545), .ZN(n17195) );
  NAND2_X1 U11779 ( .A1(n9893), .A2(n9724), .ZN(n9889) );
  INV_X1 U11780 ( .A(n11045), .ZN(n9893) );
  AOI22_X1 U11781 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11046) );
  OAI21_X1 U11782 ( .B1(n16201), .B2(n16200), .A(n19206), .ZN(n16202) );
  NOR2_X1 U11783 ( .A1(n11276), .A2(n18202), .ZN(n16731) );
  NAND2_X1 U11784 ( .A1(n16731), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16719) );
  NOR2_X1 U11785 ( .A1(n17898), .A2(n17899), .ZN(n17882) );
  INV_X1 U11786 ( .A(n17945), .ZN(n10000) );
  NOR2_X1 U11787 ( .A1(n18014), .A2(n18015), .ZN(n17999) );
  AOI21_X1 U11788 ( .B1(n11313), .B2(n11312), .A(n11311), .ZN(n18118) );
  NOR2_X1 U11789 ( .A1(n18218), .A2(n11316), .ZN(n16724) );
  NAND2_X1 U11790 ( .A1(n10318), .A2(n11147), .ZN(n11148) );
  INV_X1 U11791 ( .A(n17881), .ZN(n9876) );
  NAND2_X1 U11792 ( .A1(n17956), .A2(n17961), .ZN(n17938) );
  INV_X1 U11793 ( .A(n10168), .ZN(n9971) );
  NOR2_X1 U11794 ( .A1(n18068), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18029) );
  NAND2_X1 U11795 ( .A1(n9977), .A2(n9794), .ZN(n9974) );
  XNOR2_X1 U11796 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n11128), .ZN(
        n18136) );
  INV_X1 U11797 ( .A(n18148), .ZN(n18151) );
  NAND2_X1 U11798 ( .A1(n18382), .A2(n19212), .ZN(n9866) );
  NAND2_X1 U11799 ( .A1(n12881), .A2(n12872), .ZN(n18987) );
  NAND2_X1 U11800 ( .A1(n19017), .A2(n16102), .ZN(n19014) );
  INV_X1 U11801 ( .A(n11259), .ZN(n18567) );
  NAND2_X1 U11802 ( .A1(n10077), .A2(n9766), .ZN(n13248) );
  INV_X1 U11803 ( .A(n16159), .ZN(n10077) );
  AND2_X1 U11804 ( .A1(n14099), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20348) );
  AND2_X1 U11805 ( .A1(n13683), .A2(n13679), .ZN(n20362) );
  AND2_X1 U11806 ( .A1(n13683), .A2(n13682), .ZN(n20360) );
  INV_X1 U11807 ( .A(n20360), .ZN(n20325) );
  OR2_X1 U11808 ( .A1(n16159), .A2(n13426), .ZN(n20416) );
  OR2_X2 U11809 ( .A1(n16159), .A2(n12810), .ZN(n20282) );
  NOR2_X1 U11810 ( .A1(n16159), .A2(n20760), .ZN(n15312) );
  INV_X1 U11811 ( .A(n20696), .ZN(n20717) );
  AND2_X1 U11812 ( .A1(n16672), .A2(n10991), .ZN(n12978) );
  NOR2_X1 U11813 ( .A1(n15363), .A2(n15588), .ZN(n15362) );
  NAND2_X1 U11814 ( .A1(n10059), .A2(n19411), .ZN(n10058) );
  OR2_X1 U11815 ( .A1(n20253), .A2(n10993), .ZN(n19416) );
  CLKBUF_X1 U11816 ( .A(n13828), .Z(n13604) );
  INV_X1 U11817 ( .A(n15479), .ZN(n15470) );
  OR2_X1 U11818 ( .A1(n15448), .A2(n10692), .ZN(n15479) );
  NAND2_X1 U11819 ( .A1(n15572), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11672) );
  OAI21_X1 U11820 ( .B1(n15575), .B2(n19564), .A(n15574), .ZN(n15576) );
  AND2_X1 U11821 ( .A1(n12824), .A2(n12825), .ZN(n15766) );
  OR2_X1 U11822 ( .A1(n19239), .A2(n10493), .ZN(n16586) );
  NAND3_X1 U11823 ( .A1(n20196), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20053), 
        .ZN(n19559) );
  XNOR2_X1 U11824 ( .A(n12825), .B(n10653), .ZN(n15757) );
  NAND2_X1 U11825 ( .A1(n9835), .A2(n9727), .ZN(n10017) );
  AOI211_X1 U11826 ( .C1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n15769), .A(
        n10104), .B(n15767), .ZN(n10103) );
  NOR2_X1 U11827 ( .A1(n15782), .A2(n15771), .ZN(n10104) );
  NAND2_X1 U11828 ( .A1(n12829), .A2(n12828), .ZN(n15768) );
  NOR2_X1 U11829 ( .A1(n15967), .A2(n9967), .ZN(n9966) );
  NAND2_X1 U11830 ( .A1(n9970), .A2(n9969), .ZN(n9968) );
  AND2_X1 U11831 ( .A1(n15945), .A2(n15977), .ZN(n9967) );
  NAND2_X1 U11832 ( .A1(n9919), .A2(n10281), .ZN(n15714) );
  NAND2_X1 U11833 ( .A1(n9921), .A2(n9920), .ZN(n9919) );
  AND2_X1 U11834 ( .A1(n13153), .A2(n13130), .ZN(n16645) );
  AND2_X1 U11835 ( .A1(n13153), .A2(n20241), .ZN(n16646) );
  INV_X1 U11836 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20209) );
  OR2_X1 U11837 ( .A1(n16906), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10012) );
  OR2_X1 U11838 ( .A1(n16904), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U11839 ( .A1(n10014), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10013) );
  OR2_X1 U11840 ( .A1(n16902), .A2(n17259), .ZN(n10014) );
  NAND2_X1 U11841 ( .A1(n17058), .A2(n10003), .ZN(n17001) );
  NAND2_X1 U11842 ( .A1(n16885), .A2(n17017), .ZN(n10003) );
  NAND4_X1 U11843 ( .A1(n16883), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n18551), 
        .A4(n16882), .ZN(n17249) );
  NOR2_X1 U11844 ( .A1(n17248), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9874) );
  INV_X1 U11845 ( .A(n17249), .ZN(n17258) );
  NAND2_X1 U11846 ( .A1(n17675), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n9994) );
  INV_X1 U11847 ( .A(n17738), .ZN(n17728) );
  INV_X1 U11848 ( .A(n17741), .ZN(n17736) );
  NAND2_X1 U11849 ( .A1(n17586), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17739) );
  NAND2_X1 U11850 ( .A1(n19006), .A2(n17586), .ZN(n17743) );
  INV_X1 U11851 ( .A(n16202), .ZN(n17586) );
  INV_X1 U11852 ( .A(n17743), .ZN(n17730) );
  NAND2_X1 U11853 ( .A1(n17870), .A2(n9883), .ZN(n9985) );
  INV_X1 U11854 ( .A(n17857), .ZN(n9982) );
  NAND2_X1 U11855 ( .A1(n17865), .A2(n9980), .ZN(n9979) );
  NAND2_X1 U11856 ( .A1(n17867), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9980) );
  AND2_X1 U11857 ( .A1(n18203), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n17970) );
  INV_X1 U11858 ( .A(n18199), .ZN(n18210) );
  AOI21_X1 U11859 ( .B1(n10175), .B2(n9699), .A(n11150), .ZN(n16175) );
  INV_X1 U11860 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19222) );
  INV_X1 U11861 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U11862 ( .A1(n13584), .A2(n11718), .ZN(n12492) );
  OAI21_X1 U11863 ( .B1(n11446), .B2(n11383), .A(n16700), .ZN(n11384) );
  OR2_X1 U11864 ( .A1(n12036), .A2(n12035), .ZN(n12710) );
  INV_X1 U11865 ( .A(n13308), .ZN(n11874) );
  OR2_X1 U11866 ( .A1(n11986), .A2(n11985), .ZN(n12684) );
  NAND2_X1 U11867 ( .A1(n15338), .A2(n14265), .ZN(n12780) );
  OAI21_X1 U11868 ( .B1(n21045), .B2(n14265), .A(n12782), .ZN(n12776) );
  NOR2_X1 U11869 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9909) );
  INV_X1 U11870 ( .A(n13982), .ZN(n9963) );
  NOR2_X1 U11871 ( .A1(n10642), .A2(n20136), .ZN(n10540) );
  OAI22_X1 U11872 ( .A1(n11368), .A2(n13719), .B1(n19758), .B2(n11367), .ZN(
        n11369) );
  AND2_X1 U11873 ( .A1(n11683), .A2(n11682), .ZN(n11686) );
  OAI21_X1 U11874 ( .B1(n9763), .B2(n11673), .A(n9905), .ZN(n11683) );
  AOI21_X1 U11875 ( .B1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n14248), .A(n9740), .ZN(n10163) );
  NAND2_X1 U11876 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10164) );
  NAND2_X1 U11877 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11067) );
  AOI22_X1 U11878 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9996) );
  AND2_X1 U11879 ( .A1(n11265), .A2(n11266), .ZN(n11168) );
  NOR2_X1 U11880 ( .A1(n11275), .A2(n18557), .ZN(n9987) );
  NAND2_X1 U11881 ( .A1(n9744), .A2(n9990), .ZN(n9988) );
  INV_X1 U11882 ( .A(n11122), .ZN(n10159) );
  AOI211_X1 U11883 ( .C1(n17497), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n11226), .B(n11225), .ZN(n11227) );
  NOR2_X1 U11884 ( .A1(n11017), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11266) );
  INV_X1 U11885 ( .A(n11848), .ZN(n10125) );
  NOR2_X1 U11886 ( .A1(n14695), .A2(n10247), .ZN(n10246) );
  INV_X1 U11887 ( .A(n14261), .ZN(n10247) );
  NOR2_X1 U11888 ( .A1(n14948), .A2(n14758), .ZN(n10241) );
  NAND2_X1 U11889 ( .A1(n10151), .A2(n12741), .ZN(n9938) );
  OAI21_X1 U11890 ( .B1(n15235), .B2(n10150), .A(n12748), .ZN(n9956) );
  NAND2_X1 U11891 ( .A1(n10153), .A2(n12741), .ZN(n10150) );
  AND2_X1 U11892 ( .A1(n13214), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12665) );
  INV_X1 U11893 ( .A(n12129), .ZN(n9939) );
  NOR2_X1 U11894 ( .A1(n14709), .A2(n10133), .ZN(n10132) );
  INV_X1 U11895 ( .A(n9953), .ZN(n9952) );
  OAI21_X1 U11896 ( .B1(n15062), .B2(n16163), .A(n9737), .ZN(n9953) );
  INV_X1 U11897 ( .A(n9951), .ZN(n9948) );
  BUF_X1 U11898 ( .A(n14093), .Z(n14291) );
  NAND2_X1 U11899 ( .A1(n14652), .A2(n10127), .ZN(n13535) );
  OR2_X1 U11900 ( .A1(n11965), .A2(n11964), .ZN(n12735) );
  NAND2_X1 U11901 ( .A1(n11792), .A2(n11791), .ZN(n11837) );
  NAND2_X1 U11902 ( .A1(n10147), .A2(n15338), .ZN(n11792) );
  NAND2_X1 U11903 ( .A1(n12006), .A2(n12005), .ZN(n20583) );
  OR2_X1 U11904 ( .A1(n11910), .A2(n11909), .ZN(n11917) );
  NOR2_X1 U11905 ( .A1(n12578), .A2(n11858), .ZN(n10085) );
  NAND2_X1 U11906 ( .A1(n11738), .A2(n11737), .ZN(n11739) );
  INV_X1 U11907 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20692) );
  NAND2_X1 U11908 ( .A1(n12796), .A2(n13081), .ZN(n10080) );
  OR2_X1 U11909 ( .A1(n11004), .A2(n10667), .ZN(n11685) );
  NAND2_X1 U11910 ( .A1(n10659), .A2(n10658), .ZN(n10663) );
  OR2_X1 U11911 ( .A1(n10666), .A2(n10664), .ZN(n10659) );
  INV_X1 U11912 ( .A(n11605), .ZN(n10120) );
  AND2_X1 U11913 ( .A1(n11604), .A2(n9700), .ZN(n11612) );
  AND2_X1 U11914 ( .A1(n10118), .A2(n10578), .ZN(n10117) );
  NAND2_X1 U11915 ( .A1(n11528), .A2(n11531), .ZN(n11556) );
  AND2_X1 U11916 ( .A1(n10570), .A2(n13489), .ZN(n10118) );
  OR2_X1 U11917 ( .A1(n11426), .A2(n9783), .ZN(n11505) );
  NAND2_X1 U11918 ( .A1(n15423), .A2(n14508), .ZN(n14526) );
  NAND2_X1 U11919 ( .A1(n10691), .A2(n20205), .ZN(n10856) );
  NAND2_X1 U11920 ( .A1(n10970), .A2(n10099), .ZN(n10098) );
  INV_X1 U11921 ( .A(n15428), .ZN(n10205) );
  INV_X1 U11922 ( .A(n15456), .ZN(n10219) );
  NAND2_X1 U11923 ( .A1(n10095), .A2(n14114), .ZN(n10094) );
  INV_X1 U11924 ( .A(n14043), .ZN(n10095) );
  NAND2_X1 U11925 ( .A1(n9679), .A2(n14159), .ZN(n10220) );
  INV_X1 U11926 ( .A(n15970), .ZN(n10096) );
  NAND2_X1 U11927 ( .A1(n9718), .A2(n10188), .ZN(n10187) );
  NOR2_X1 U11928 ( .A1(n10189), .A2(n11523), .ZN(n10188) );
  OR2_X1 U11929 ( .A1(n10346), .A2(n10322), .ZN(n10358) );
  INV_X1 U11930 ( .A(n11523), .ZN(n10274) );
  INV_X1 U11931 ( .A(n10349), .ZN(n10064) );
  AND2_X1 U11932 ( .A1(n14136), .A2(n11655), .ZN(n9958) );
  NAND2_X1 U11933 ( .A1(n11499), .A2(n11498), .ZN(n11656) );
  INV_X1 U11934 ( .A(n14136), .ZN(n9959) );
  INV_X1 U11935 ( .A(n10999), .ZN(n11642) );
  AND2_X1 U11936 ( .A1(n15400), .A2(n15354), .ZN(n10254) );
  NOR2_X1 U11937 ( .A1(n15840), .A2(n15821), .ZN(n10196) );
  AND2_X1 U11938 ( .A1(n10029), .A2(n15642), .ZN(n9911) );
  NOR2_X1 U11939 ( .A1(n10197), .A2(n9945), .ZN(n9944) );
  OR2_X1 U11940 ( .A1(n10198), .A2(n15855), .ZN(n10197) );
  NAND2_X1 U11941 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10198) );
  NAND2_X1 U11942 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9945) );
  INV_X1 U11943 ( .A(n10099), .ZN(n10097) );
  INV_X1 U11944 ( .A(n15963), .ZN(n10286) );
  NAND2_X1 U11945 ( .A1(n10545), .A2(n10544), .ZN(n10546) );
  INV_X1 U11946 ( .A(n14028), .ZN(n10262) );
  AOI21_X1 U11947 ( .B1(n10027), .B2(n10026), .A(n10023), .ZN(n10022) );
  INV_X1 U11948 ( .A(n13979), .ZN(n10023) );
  AND2_X1 U11949 ( .A1(n10025), .A2(n11618), .ZN(n10020) );
  NAND2_X1 U11950 ( .A1(n13189), .A2(n13184), .ZN(n10182) );
  NAND2_X1 U11951 ( .A1(n16662), .A2(n10086), .ZN(n10500) );
  AND2_X1 U11952 ( .A1(n10499), .A2(n10691), .ZN(n10086) );
  AND2_X1 U11953 ( .A1(n13163), .A2(n13164), .ZN(n10717) );
  OR2_X1 U11954 ( .A1(n13039), .A2(n13038), .ZN(n16665) );
  NAND2_X1 U11955 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20239), .ZN(
        n11419) );
  NAND2_X1 U11956 ( .A1(n19177), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11022) );
  NAND2_X1 U11957 ( .A1(n11017), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11023) );
  NAND2_X1 U11958 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n9892) );
  AOI21_X1 U11959 ( .B1(n17433), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(n9891), .ZN(n9890) );
  NOR2_X1 U11960 ( .A1(n9652), .A2(n11044), .ZN(n9891) );
  NAND2_X1 U11961 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11056) );
  AND2_X1 U11962 ( .A1(n12869), .A2(n11261), .ZN(n11258) );
  NOR2_X1 U11963 ( .A1(n17880), .A2(n11148), .ZN(n16744) );
  NOR2_X1 U11964 ( .A1(n9854), .A2(n9848), .ZN(n9847) );
  NAND2_X1 U11965 ( .A1(n9853), .A2(n9849), .ZN(n9848) );
  NAND2_X1 U11966 ( .A1(n11068), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n9856) );
  NOR2_X1 U11967 ( .A1(n11266), .A2(n9867), .ZN(n11264) );
  AND2_X1 U11968 ( .A1(n11017), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n9867) );
  AND2_X1 U11969 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11300), .ZN(
        n11301) );
  NOR2_X1 U11970 ( .A1(n11253), .A2(n11262), .ZN(n16102) );
  NOR2_X1 U11971 ( .A1(n10075), .A2(n10076), .ZN(n10072) );
  INV_X1 U11972 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n10075) );
  NOR2_X1 U11973 ( .A1(n20979), .A2(n10074), .ZN(n10073) );
  INV_X1 U11974 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20309) );
  INV_X1 U11975 ( .A(n14812), .ZN(n20307) );
  AND2_X1 U11976 ( .A1(n13683), .A2(n13681), .ZN(n20366) );
  AND2_X1 U11977 ( .A1(n12598), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12599) );
  NAND2_X1 U11978 ( .A1(n10243), .A2(n10246), .ZN(n14680) );
  AND2_X1 U11979 ( .A1(n12567), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12568) );
  NAND2_X1 U11980 ( .A1(n12568), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12597) );
  INV_X1 U11981 ( .A(n14722), .ZN(n12515) );
  NAND2_X1 U11982 ( .A1(n16167), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10155) );
  NOR2_X1 U11983 ( .A1(n12397), .A2(n16261), .ZN(n12398) );
  AND2_X1 U11984 ( .A1(n12377), .A2(n12376), .ZN(n14772) );
  CLKBUF_X1 U11985 ( .A(n14771), .Z(n14947) );
  NOR2_X1 U11986 ( .A1(n12339), .A2(n14802), .ZN(n12340) );
  NAND2_X1 U11987 ( .A1(n10230), .A2(n14781), .ZN(n10229) );
  NAND2_X1 U11988 ( .A1(n12320), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12339) );
  AND2_X1 U11989 ( .A1(n12300), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12320) );
  NOR2_X1 U11990 ( .A1(n12223), .A2(n12236), .ZN(n12300) );
  INV_X1 U11991 ( .A(n15236), .ZN(n15072) );
  NOR2_X1 U11992 ( .A1(n12263), .A2(n16216), .ZN(n12243) );
  NOR2_X1 U11993 ( .A1(n12207), .A2(n12206), .ZN(n12293) );
  NOR2_X1 U11994 ( .A1(n12172), .A2(n12171), .ZN(n12187) );
  NAND2_X1 U11995 ( .A1(n14009), .A2(n14075), .ZN(n10235) );
  NAND2_X1 U11996 ( .A1(n10234), .A2(n10233), .ZN(n10237) );
  INV_X1 U11997 ( .A(n10239), .ZN(n10233) );
  AOI21_X1 U11998 ( .B1(n12718), .B2(n12292), .A(n12154), .ZN(n14017) );
  INV_X1 U11999 ( .A(n13612), .ZN(n12147) );
  NOR2_X1 U12000 ( .A1(n12133), .A2(n13707), .ZN(n12142) );
  CLKBUF_X1 U12001 ( .A(n13612), .Z(n13838) );
  INV_X1 U12002 ( .A(n12100), .ZN(n12123) );
  NAND2_X1 U12003 ( .A1(n12123), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12133) );
  NAND2_X1 U12004 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12100) );
  OAI21_X1 U12005 ( .B1(n20582), .B2(n12260), .A(n12103), .ZN(n12104) );
  CLKBUF_X1 U12006 ( .A(n13647), .Z(n13657) );
  NAND2_X1 U12007 ( .A1(n12848), .A2(n15227), .ZN(n12849) );
  NAND2_X1 U12008 ( .A1(n10045), .A2(n10044), .ZN(n10043) );
  NOR2_X1 U12009 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10044) );
  INV_X1 U12010 ( .A(n14999), .ZN(n10045) );
  NOR2_X1 U12011 ( .A1(n9706), .A2(n10130), .ZN(n14698) );
  INV_X1 U12012 ( .A(n10132), .ZN(n10130) );
  NOR2_X1 U12013 ( .A1(n9706), .A2(n14709), .ZN(n14710) );
  OR3_X1 U12014 ( .A1(n16169), .A2(n16170), .A3(n14761), .ZN(n14762) );
  NAND2_X1 U12015 ( .A1(n14786), .A2(n14774), .ZN(n16169) );
  NAND2_X1 U12016 ( .A1(n10136), .A2(n10135), .ZN(n10134) );
  NOR2_X1 U12017 ( .A1(n14294), .A2(n10137), .ZN(n10136) );
  INV_X1 U12018 ( .A(n14840), .ZN(n10135) );
  NAND2_X1 U12019 ( .A1(n15018), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9949) );
  NOR3_X1 U12020 ( .A1(n10309), .A2(n14840), .A3(n10138), .ZN(n14828) );
  NOR2_X1 U12021 ( .A1(n10309), .A2(n14840), .ZN(n14839) );
  NOR2_X1 U12022 ( .A1(n14908), .A2(n14907), .ZN(n14910) );
  OR2_X1 U12023 ( .A1(n14170), .A2(n14169), .ZN(n14908) );
  NAND2_X1 U12024 ( .A1(n12740), .A2(n10152), .ZN(n15251) );
  OR2_X1 U12025 ( .A1(n15290), .A2(n14096), .ZN(n14170) );
  AND2_X1 U12026 ( .A1(n16403), .A2(n14085), .ZN(n16405) );
  AOI21_X1 U12027 ( .B1(n14015), .B2(n9930), .A(n9736), .ZN(n9929) );
  INV_X1 U12028 ( .A(n14015), .ZN(n9931) );
  OAI21_X1 U12029 ( .B1(n20518), .B2(n12697), .A(n12672), .ZN(n13491) );
  XNOR2_X1 U12030 ( .A(n11938), .B(n11937), .ZN(n12115) );
  XNOR2_X1 U12031 ( .A(n12107), .B(n12106), .ZN(n13595) );
  INV_X1 U12032 ( .A(n12105), .ZN(n12107) );
  INV_X1 U12033 ( .A(n12673), .ZN(n12106) );
  INV_X1 U12034 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10226) );
  AND3_X1 U12035 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13572) );
  OR2_X1 U12036 ( .A1(n21020), .A2(n20750), .ZN(n20756) );
  INV_X1 U12037 ( .A(n15339), .ZN(n13968) );
  INV_X1 U12038 ( .A(n20559), .ZN(n20661) );
  AND2_X1 U12039 ( .A1(n21021), .A2(n20518), .ZN(n20842) );
  INV_X1 U12040 ( .A(n21022), .ZN(n20884) );
  AOI21_X1 U12041 ( .B1(n20721), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n15326), 
        .ZN(n20888) );
  AND2_X1 U12042 ( .A1(n10498), .A2(n10468), .ZN(n9846) );
  NAND2_X1 U12043 ( .A1(n10691), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20258) );
  AOI22_X1 U12044 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n20229), .B2(n20194), .ZN(
        n11677) );
  NAND2_X1 U12045 ( .A1(n16434), .A2(n11602), .ZN(n11604) );
  AND2_X1 U12046 ( .A1(n9700), .A2(n11611), .ZN(n10119) );
  NAND2_X1 U12047 ( .A1(n10977), .A2(n10108), .ZN(n15501) );
  NAND2_X1 U12048 ( .A1(n16454), .A2(n11012), .ZN(n16434) );
  NAND2_X1 U12049 ( .A1(n10114), .A2(n10113), .ZN(n11539) );
  INV_X1 U12050 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10113) );
  NAND2_X1 U12051 ( .A1(n11602), .A2(n11549), .ZN(n11569) );
  NAND2_X1 U12052 ( .A1(n11552), .A2(n14071), .ZN(n11549) );
  AND2_X1 U12053 ( .A1(n11513), .A2(n10118), .ZN(n11527) );
  NOR2_X1 U12054 ( .A1(n10223), .A2(n13831), .ZN(n10222) );
  NAND2_X1 U12055 ( .A1(n15422), .A2(n15424), .ZN(n15423) );
  NOR2_X1 U12056 ( .A1(n15905), .A2(n15904), .ZN(n15907) );
  AND2_X1 U12057 ( .A1(n9762), .A2(n16026), .ZN(n10101) );
  AND2_X1 U12058 ( .A1(n10090), .A2(n14129), .ZN(n10089) );
  AND3_X1 U12059 ( .A1(n10778), .A2(n10777), .A3(n10776), .ZN(n14031) );
  NOR2_X1 U12060 ( .A1(n13323), .A2(n10088), .ZN(n14130) );
  NAND2_X1 U12061 ( .A1(n10091), .A2(n10090), .ZN(n10088) );
  INV_X1 U12062 ( .A(n12922), .ZN(n14116) );
  AND2_X1 U12063 ( .A1(n9693), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10060) );
  NAND2_X1 U12064 ( .A1(n13851), .A2(n10249), .ZN(n14069) );
  AND2_X1 U12065 ( .A1(n13851), .A2(n13825), .ZN(n13935) );
  NAND2_X1 U12066 ( .A1(n9687), .A2(n9775), .ZN(n10063) );
  AND2_X1 U12067 ( .A1(n13695), .A2(n9723), .ZN(n13547) );
  NOR2_X1 U12068 ( .A1(n15725), .A2(n10068), .ZN(n10067) );
  INV_X1 U12069 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15725) );
  NAND2_X1 U12070 ( .A1(n16063), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16062) );
  AND2_X1 U12071 ( .A1(n10564), .A2(n10563), .ZN(n13454) );
  INV_X1 U12072 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13983) );
  NAND2_X1 U12073 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10355) );
  AND2_X1 U12074 ( .A1(n10106), .A2(n15357), .ZN(n10105) );
  OR3_X1 U12075 ( .A1(n12838), .A2(n11667), .A3(n15764), .ZN(n15567) );
  NOR2_X1 U12076 ( .A1(n10190), .A2(n15597), .ZN(n9837) );
  NAND2_X1 U12077 ( .A1(n9944), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9943) );
  NOR2_X1 U12078 ( .A1(n15432), .A2(n15431), .ZN(n15433) );
  OR2_X1 U12079 ( .A1(n12959), .A2(n12958), .ZN(n15432) );
  INV_X1 U12080 ( .A(n9944), .ZN(n9942) );
  INV_X1 U12081 ( .A(n12931), .ZN(n10255) );
  INV_X1 U12082 ( .A(n10198), .ZN(n9823) );
  INV_X1 U12083 ( .A(n15667), .ZN(n9825) );
  OR2_X1 U12084 ( .A1(n9945), .A2(n10199), .ZN(n9822) );
  NAND2_X1 U12085 ( .A1(n11537), .A2(n10199), .ZN(n15651) );
  NAND2_X1 U12086 ( .A1(n15475), .A2(n10257), .ZN(n15464) );
  NAND2_X1 U12087 ( .A1(n15475), .A2(n9756), .ZN(n15454) );
  NAND2_X1 U12088 ( .A1(n13851), .A2(n9774), .ZN(n15474) );
  INV_X1 U12089 ( .A(n14070), .ZN(n10248) );
  NOR2_X2 U12090 ( .A1(n15474), .A2(n15473), .ZN(n15475) );
  INV_X1 U12091 ( .A(n15943), .ZN(n9970) );
  NAND2_X1 U12092 ( .A1(n16630), .A2(n15944), .ZN(n9969) );
  INV_X1 U12093 ( .A(n10282), .ZN(n10281) );
  OAI21_X1 U12094 ( .B1(n10288), .B2(n10283), .A(n15962), .ZN(n10282) );
  NAND2_X1 U12095 ( .A1(n10284), .A2(n10286), .ZN(n10283) );
  INV_X1 U12096 ( .A(n10290), .ZN(n10284) );
  INV_X1 U12097 ( .A(n16525), .ZN(n9921) );
  NOR2_X1 U12098 ( .A1(n15987), .A2(n14043), .ZN(n15969) );
  AND2_X1 U12099 ( .A1(n13695), .A2(n9750), .ZN(n13809) );
  INV_X1 U12100 ( .A(n13607), .ZN(n10250) );
  NAND2_X1 U12101 ( .A1(n13695), .A2(n10251), .ZN(n13606) );
  NAND2_X1 U12102 ( .A1(n13695), .A2(n13694), .ZN(n13696) );
  NOR2_X1 U12103 ( .A1(n14028), .A2(n10259), .ZN(n13457) );
  NAND2_X1 U12104 ( .A1(n9717), .A2(n10260), .ZN(n10259) );
  INV_X1 U12105 ( .A(n13454), .ZN(n10260) );
  AND2_X1 U12106 ( .A1(n13457), .A2(n13446), .ZN(n13695) );
  NAND2_X1 U12107 ( .A1(n14124), .A2(n9916), .ZN(n9840) );
  INV_X1 U12108 ( .A(n9898), .ZN(n9841) );
  XNOR2_X1 U12109 ( .A(n11508), .B(n16055), .ZN(n16048) );
  AND2_X2 U12110 ( .A1(n11653), .A2(n14024), .ZN(n14139) );
  AND2_X1 U12111 ( .A1(n10559), .A2(n10558), .ZN(n13288) );
  NAND2_X1 U12112 ( .A1(n10262), .A2(n9717), .ZN(n13455) );
  AND2_X1 U12113 ( .A1(n10554), .A2(n10553), .ZN(n14027) );
  NAND2_X1 U12114 ( .A1(n10262), .A2(n10555), .ZN(n14030) );
  INV_X1 U12115 ( .A(n16665), .ZN(n13136) );
  NAND2_X1 U12116 ( .A1(n10376), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9821) );
  NAND2_X1 U12117 ( .A1(n10375), .A2(n10680), .ZN(n9820) );
  NAND3_X1 U12118 ( .A1(n10315), .A2(n10424), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10431) );
  INV_X1 U12119 ( .A(n11365), .ZN(n9843) );
  INV_X1 U12120 ( .A(n20049), .ZN(n19795) );
  BUF_X1 U12121 ( .A(n10495), .Z(n19597) );
  NAND2_X1 U12122 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20053), .ZN(n19596) );
  NAND2_X1 U12123 ( .A1(n19854), .A2(n20234), .ZN(n20003) );
  INV_X1 U12124 ( .A(n19607), .ZN(n19609) );
  INV_X1 U12125 ( .A(n19608), .ZN(n19611) );
  INV_X1 U12126 ( .A(n19596), .ZN(n19613) );
  NAND2_X1 U12127 ( .A1(n13121), .A2(n11692), .ZN(n16668) );
  NOR2_X1 U12128 ( .A1(n16928), .A2(n17868), .ZN(n16927) );
  NOR2_X1 U12129 ( .A1(n16949), .A2(n16950), .ZN(n16948) );
  NOR2_X1 U12130 ( .A1(n17936), .A2(n16985), .ZN(n16984) );
  NOR2_X1 U12131 ( .A1(n16992), .A2(n16993), .ZN(n16991) );
  INV_X1 U12132 ( .A(n18153), .ZN(n10007) );
  INV_X1 U12133 ( .A(n16880), .ZN(n16883) );
  NAND2_X1 U12134 ( .A1(n9703), .A2(n9795), .ZN(n9995) );
  OAI211_X1 U12135 ( .C1(n11180), .C2(n18582), .A(n11034), .B(n11033), .ZN(
        n11302) );
  NOR2_X1 U12136 ( .A1(n9731), .A2(n9973), .ZN(n9972) );
  NOR2_X2 U12137 ( .A1(n18578), .A2(n11251), .ZN(n19006) );
  NOR2_X1 U12138 ( .A1(n17783), .A2(n17745), .ZN(n17763) );
  NOR2_X1 U12139 ( .A1(n17899), .A2(n16888), .ZN(n17853) );
  NOR2_X1 U12140 ( .A1(n9754), .A2(n9999), .ZN(n9998) );
  NAND2_X1 U12141 ( .A1(n17897), .A2(n18207), .ZN(n17964) );
  NOR2_X1 U12142 ( .A1(n18202), .A2(n11278), .ZN(n17975) );
  AOI21_X1 U12143 ( .B1(n11277), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18932), .ZN(n18052) );
  NAND2_X1 U12144 ( .A1(n10004), .A2(n10006), .ZN(n18051) );
  NOR2_X1 U12145 ( .A1(n18153), .A2(n10005), .ZN(n10004) );
  NAND2_X1 U12146 ( .A1(n9742), .A2(n10008), .ZN(n10005) );
  NAND2_X1 U12147 ( .A1(n10007), .A2(n10008), .ZN(n18112) );
  NOR2_X1 U12148 ( .A1(n11151), .A2(n10301), .ZN(n11153) );
  NAND2_X1 U12149 ( .A1(n17955), .A2(n11146), .ZN(n17920) );
  NOR2_X1 U12150 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11142), .ZN(
        n17956) );
  NOR2_X1 U12151 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n9883), .ZN(
        n17995) );
  OAI21_X1 U12152 ( .B1(n18040), .B2(n11135), .A(n18109), .ZN(n11140) );
  NAND2_X1 U12153 ( .A1(n9976), .A2(n9688), .ZN(n18068) );
  AND2_X1 U12154 ( .A1(n9794), .A2(n18375), .ZN(n9975) );
  NAND2_X1 U12155 ( .A1(n9863), .A2(n9860), .ZN(n19019) );
  NOR2_X1 U12156 ( .A1(n17785), .A2(n9686), .ZN(n9860) );
  AOI21_X1 U12157 ( .B1(n11263), .B2(n18551), .A(n11262), .ZN(n18996) );
  NOR2_X1 U12158 ( .A1(n11308), .A2(n11312), .ZN(n11314) );
  NAND2_X1 U12159 ( .A1(n9976), .A2(n9977), .ZN(n18096) );
  INV_X1 U12160 ( .A(n19023), .ZN(n18992) );
  NOR2_X1 U12161 ( .A1(n16102), .A2(n19019), .ZN(n19007) );
  AND2_X1 U12162 ( .A1(n9873), .A2(n9872), .ZN(n19187) );
  NAND2_X1 U12163 ( .A1(n19007), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9872) );
  NAND2_X1 U12164 ( .A1(n19009), .A2(n11017), .ZN(n9873) );
  INV_X1 U12165 ( .A(n19019), .ZN(n19017) );
  NOR2_X1 U12166 ( .A1(n19026), .A2(n11017), .ZN(n18995) );
  NAND2_X1 U12167 ( .A1(n19224), .A2(n16109), .ZN(n19023) );
  OAI211_X1 U12168 ( .C1(n17557), .C2(n18752), .A(n11220), .B(n11219), .ZN(
        n18545) );
  AOI211_X2 U12169 ( .C1(n16109), .C2(n16108), .A(n16201), .B(n16107), .ZN(
        n19029) );
  OAI21_X1 U12170 ( .B1(n9865), .B2(n9866), .A(n9772), .ZN(n18993) );
  NAND2_X1 U12171 ( .A1(n18400), .A2(n16108), .ZN(n9865) );
  NOR2_X1 U12172 ( .A1(n18551), .A2(n9862), .ZN(n19046) );
  INV_X1 U12173 ( .A(n13212), .ZN(n9934) );
  AND2_X1 U12174 ( .A1(n14717), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14705) );
  OR2_X1 U12175 ( .A1(n14753), .A2(n20995), .ZN(n14742) );
  NOR2_X1 U12176 ( .A1(n14773), .A2(n20990), .ZN(n16207) );
  AND2_X1 U12177 ( .A1(n16221), .A2(n10071), .ZN(n14804) );
  AND2_X1 U12178 ( .A1(n9704), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U12179 ( .A1(n16221), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n14844) );
  INV_X1 U12180 ( .A(n20348), .ZN(n20365) );
  NOR2_X1 U12181 ( .A1(n20343), .A2(n14077), .ZN(n16235) );
  INV_X1 U12182 ( .A(n20308), .ZN(n20346) );
  INV_X1 U12183 ( .A(n14864), .ZN(n20328) );
  NOR2_X1 U12184 ( .A1(n20960), .A2(n13805), .ZN(n20344) );
  NAND2_X1 U12185 ( .A1(n14099), .A2(n9935), .ZN(n13671) );
  OR2_X1 U12186 ( .A1(n20366), .A2(n13674), .ZN(n14812) );
  INV_X1 U12187 ( .A(n14914), .ZN(n20383) );
  INV_X1 U12188 ( .A(n14916), .ZN(n20382) );
  INV_X1 U12189 ( .A(n20387), .ZN(n14902) );
  OR2_X1 U12190 ( .A1(n13868), .A2(n20276), .ZN(n13874) );
  NAND2_X1 U12191 ( .A1(n20387), .A2(n14347), .ZN(n14916) );
  INV_X1 U12192 ( .A(n20383), .ZN(n14884) );
  INV_X1 U12193 ( .A(n14957), .ZN(n14969) );
  INV_X1 U12194 ( .A(n14987), .ZN(n14979) );
  INV_X1 U12195 ( .A(n20416), .ZN(n20388) );
  INV_X1 U12196 ( .A(n21049), .ZN(n20400) );
  XNOR2_X1 U12197 ( .A(n12865), .B(n12864), .ZN(n14651) );
  OAI21_X1 U12198 ( .B1(n15061), .B2(n10155), .A(n15224), .ZN(n15053) );
  AND2_X1 U12199 ( .A1(n16260), .A2(n13492), .ZN(n16285) );
  OAI22_X1 U12200 ( .A1(n9928), .A2(n9927), .B1(n12847), .B2(n12757), .ZN(
        n12758) );
  NAND2_X1 U12201 ( .A1(n16163), .A2(n12846), .ZN(n9927) );
  XNOR2_X1 U12202 ( .A(n10041), .B(n15001), .ZN(n15185) );
  OAI21_X1 U12203 ( .B1(n9722), .B2(n16163), .A(n10042), .ZN(n10041) );
  OAI21_X1 U12204 ( .B1(n15000), .B2(n10043), .A(n16163), .ZN(n10042) );
  AND2_X1 U12205 ( .A1(n16303), .A2(n15136), .ZN(n15191) );
  NAND2_X1 U12206 ( .A1(n15021), .A2(n15009), .ZN(n15008) );
  NOR2_X1 U12207 ( .A1(n16311), .A2(n16320), .ZN(n16303) );
  NAND2_X1 U12208 ( .A1(n12740), .A2(n12739), .ZN(n15117) );
  INV_X1 U12209 ( .A(n20446), .ZN(n16394) );
  NAND2_X1 U12210 ( .A1(n9932), .A2(n12717), .ZN(n14014) );
  NAND2_X1 U12211 ( .A1(n10142), .A2(n10141), .ZN(n13815) );
  OR2_X1 U12212 ( .A1(n13540), .A2(n13530), .ZN(n16407) );
  INV_X1 U12213 ( .A(n16407), .ZN(n20451) );
  OR2_X1 U12214 ( .A1(n13540), .A2(n13518), .ZN(n20446) );
  CLKBUF_X1 U12215 ( .A(n15296), .Z(n20693) );
  CLKBUF_X1 U12216 ( .A(n13569), .Z(n13570) );
  INV_X1 U12217 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21034) );
  INV_X1 U12218 ( .A(n10228), .ZN(n12130) );
  INV_X1 U12219 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20456) );
  CLKBUF_X1 U12220 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n15318) );
  INV_X1 U12221 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13370) );
  AND2_X1 U12222 ( .A1(n20552), .A2(n20842), .ZN(n20575) );
  OAI21_X1 U12223 ( .B1(n20603), .B2(n20588), .A(n20849), .ZN(n20606) );
  OAI211_X1 U12224 ( .C1(n20715), .C2(n20760), .A(n20759), .B(n20700), .ZN(
        n20718) );
  INV_X1 U12225 ( .A(n20751), .ZN(n20789) );
  NOR2_X1 U12226 ( .A1(n21022), .A2(n20457), .ZN(n20835) );
  OAI211_X1 U12227 ( .C1(n20867), .C2(n20850), .A(n20849), .B(n20848), .ZN(
        n20871) );
  INV_X1 U12228 ( .A(n20767), .ZN(n20880) );
  INV_X1 U12229 ( .A(n20770), .ZN(n20895) );
  INV_X1 U12230 ( .A(n20774), .ZN(n20901) );
  INV_X1 U12231 ( .A(n20777), .ZN(n20907) );
  INV_X1 U12232 ( .A(n20476), .ZN(n20908) );
  INV_X1 U12233 ( .A(n20781), .ZN(n20913) );
  INV_X1 U12234 ( .A(n20784), .ZN(n20919) );
  INV_X1 U12235 ( .A(n20481), .ZN(n20920) );
  INV_X1 U12236 ( .A(n20942), .ZN(n20928) );
  INV_X1 U12237 ( .A(n20787), .ZN(n20925) );
  INV_X1 U12238 ( .A(n20484), .ZN(n20926) );
  NAND2_X1 U12239 ( .A1(n20884), .A2(n20842), .ZN(n20942) );
  AND2_X1 U12240 ( .A1(n20464), .A2(n14939), .ZN(n20936) );
  OR2_X1 U12241 ( .A1(n12806), .A2(n13086), .ZN(n12807) );
  INV_X1 U12242 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16420) );
  AND2_X1 U12243 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16157), .ZN(n20945) );
  INV_X1 U12244 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21045) );
  NAND2_X1 U12246 ( .A1(n19393), .A2(n10054), .ZN(n10053) );
  NAND2_X1 U12247 ( .A1(n12954), .A2(n10337), .ZN(n10052) );
  NOR2_X1 U12248 ( .A1(n16472), .A2(n16473), .ZN(n16471) );
  NOR2_X1 U12249 ( .A1(n12954), .A2(n19393), .ZN(n16472) );
  INV_X1 U12250 ( .A(n19270), .ZN(n10048) );
  INV_X1 U12251 ( .A(n10049), .ZN(n19271) );
  OR2_X1 U12252 ( .A1(n19402), .A2(n20205), .ZN(n19386) );
  NAND2_X1 U12253 ( .A1(n12834), .A2(n12833), .ZN(n19406) );
  CLKBUF_X1 U12254 ( .A(n10363), .Z(n19411) );
  AND2_X1 U12255 ( .A1(n20253), .A2(n9796), .ZN(n19425) );
  INV_X1 U12256 ( .A(n12832), .ZN(n9904) );
  OR2_X1 U12257 ( .A1(n10887), .A2(n10886), .ZN(n13605) );
  OR2_X1 U12258 ( .A1(n10854), .A2(n10853), .ZN(n13545) );
  NAND2_X1 U12259 ( .A1(n10211), .A2(n10210), .ZN(n14610) );
  NAND2_X1 U12260 ( .A1(n10215), .A2(n10213), .ZN(n10212) );
  INV_X1 U12261 ( .A(n10216), .ZN(n10209) );
  NOR2_X1 U12262 ( .A1(n15410), .A2(n15409), .ZN(n15408) );
  NAND2_X1 U12263 ( .A1(n10201), .A2(n10200), .ZN(n15427) );
  OR2_X1 U12264 ( .A1(n13331), .A2(n13330), .ZN(n13333) );
  NOR2_X1 U12265 ( .A1(n19497), .A2(n19495), .ZN(n19473) );
  NOR2_X1 U12266 ( .A1(n13171), .A2(n13058), .ZN(n19500) );
  AND2_X1 U12267 ( .A1(n19466), .A2(n10692), .ZN(n19495) );
  INV_X1 U12268 ( .A(n19459), .ZN(n19503) );
  NAND2_X1 U12269 ( .A1(n15402), .A2(n15401), .ZN(n16423) );
  OAI21_X1 U12270 ( .B1(n15618), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15619), .ZN(n15818) );
  OR2_X1 U12271 ( .A1(n16014), .A2(n10033), .ZN(n10032) );
  AOI21_X1 U12272 ( .B1(n16525), .B2(n10292), .A(n15653), .ZN(n16507) );
  NAND2_X1 U12273 ( .A1(n19239), .A2(n11695), .ZN(n16593) );
  AND2_X1 U12274 ( .A1(n16593), .A2(n13067), .ZN(n16583) );
  INV_X1 U12275 ( .A(n16593), .ZN(n19551) );
  AOI21_X1 U12276 ( .B1(n15817), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15585) );
  XNOR2_X1 U12277 ( .A(n15817), .B(n15796), .ZN(n15801) );
  AND3_X1 U12278 ( .A1(n10037), .A2(n10036), .A3(n10035), .ZN(n15612) );
  NAND2_X1 U12279 ( .A1(n10037), .A2(n10036), .ZN(n15625) );
  INV_X1 U12280 ( .A(n11600), .ZN(n15636) );
  NAND2_X1 U12281 ( .A1(n9913), .A2(n10028), .ZN(n15643) );
  NAND2_X1 U12282 ( .A1(n16014), .A2(n10029), .ZN(n9913) );
  NAND2_X1 U12283 ( .A1(n10269), .A2(n10270), .ZN(n10268) );
  XNOR2_X1 U12284 ( .A(n9923), .B(n9759), .ZN(n15927) );
  INV_X1 U12285 ( .A(n10269), .ZN(n15692) );
  NAND2_X1 U12286 ( .A1(n9917), .A2(n9918), .ZN(n15704) );
  INV_X1 U12287 ( .A(n10280), .ZN(n15966) );
  NAND2_X1 U12288 ( .A1(n10186), .A2(n10277), .ZN(n16000) );
  NAND2_X1 U12289 ( .A1(n16014), .A2(n11523), .ZN(n10186) );
  INV_X1 U12290 ( .A(n15989), .ZN(n19364) );
  NAND2_X1 U12291 ( .A1(n9817), .A2(n11663), .ZN(n16570) );
  NAND2_X1 U12292 ( .A1(n13619), .A2(n13620), .ZN(n13909) );
  NAND2_X1 U12293 ( .A1(n9915), .A2(n9914), .ZN(n14125) );
  INV_X1 U12294 ( .A(n9916), .ZN(n9915) );
  OAI21_X1 U12295 ( .B1(n13981), .B2(n11618), .A(n10025), .ZN(n13978) );
  NAND2_X1 U12296 ( .A1(n10021), .A2(n10027), .ZN(n13977) );
  XNOR2_X1 U12297 ( .A(n13189), .B(n13184), .ZN(n11329) );
  INV_X1 U12298 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13155) );
  AND2_X1 U12299 ( .A1(n15944), .A2(n15940), .ZN(n16609) );
  INV_X1 U12300 ( .A(n13050), .ZN(n13162) );
  INV_X1 U12301 ( .A(n16645), .ZN(n16629) );
  INV_X1 U12302 ( .A(n19500), .ZN(n20234) );
  INV_X1 U12303 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20229) );
  INV_X1 U12304 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20219) );
  NAND2_X1 U12305 ( .A1(n13372), .A2(n13378), .ZN(n20204) );
  NAND2_X1 U12306 ( .A1(n13377), .A2(n13376), .ZN(n13378) );
  INV_X1 U12307 ( .A(n20196), .ZN(n20202) );
  NOR2_X1 U12308 ( .A1(n13323), .A2(n10742), .ZN(n13632) );
  OR2_X1 U12309 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  NAND2_X1 U12310 ( .A1(n13197), .A2(n13196), .ZN(n20210) );
  OR2_X1 U12311 ( .A1(n13282), .A2(n13281), .ZN(n13197) );
  INV_X1 U12312 ( .A(n20204), .ZN(n19854) );
  NOR2_X1 U12313 ( .A1(n10691), .A2(n10468), .ZN(n16659) );
  INV_X1 U12314 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16675) );
  OAI21_X1 U12315 ( .B1(n19568), .B2(n19615), .A(n20053), .ZN(n19618) );
  INV_X1 U12316 ( .A(n19636), .ZN(n19639) );
  INV_X1 U12317 ( .A(n19643), .ZN(n19669) );
  INV_X1 U12318 ( .A(n19698), .ZN(n19702) );
  INV_X1 U12319 ( .A(n19716), .ZN(n19734) );
  AND2_X1 U12320 ( .A1(n19788), .A2(n13723), .ZN(n19771) );
  OR2_X1 U12321 ( .A1(n20003), .A2(n19855), .ZN(n19886) );
  OAI21_X1 U12322 ( .B1(n19896), .B2(n19911), .A(n20053), .ZN(n19914) );
  INV_X1 U12323 ( .A(n19891), .ZN(n19913) );
  NOR2_X1 U12324 ( .A1(n20003), .A2(n20197), .ZN(n19939) );
  INV_X1 U12325 ( .A(n20067), .ZN(n19985) );
  INV_X1 U12326 ( .A(n20061), .ZN(n20018) );
  NOR2_X1 U12327 ( .A1(n19970), .A2(n19974), .ZN(n20026) );
  INV_X1 U12328 ( .A(n20026), .ZN(n20040) );
  OAI22_X1 U12329 ( .A1(n19586), .A2(n19611), .B1(n15503), .B2(n19609), .ZN(
        n20073) );
  AND2_X1 U12330 ( .A1(n10457), .A2(n19613), .ZN(n20071) );
  OAI22_X1 U12331 ( .A1(n16779), .A2(n19611), .B1(n18565), .B2(n19609), .ZN(
        n20079) );
  OAI22_X1 U12332 ( .A1(n19595), .A2(n19611), .B1(n19594), .B2(n19609), .ZN(
        n20085) );
  INV_X1 U12333 ( .A(n20106), .ZN(n20092) );
  OR2_X1 U12334 ( .A1(n19970), .A2(n20049), .ZN(n20106) );
  AND2_X1 U12335 ( .A1(n19614), .A2(n19613), .ZN(n20097) );
  INV_X1 U12336 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20205) );
  INV_X1 U12337 ( .A(n9861), .ZN(n16864) );
  AOI21_X1 U12338 ( .B1(n18984), .B2(n19014), .A(n17783), .ZN(n19226) );
  NAND2_X1 U12339 ( .A1(n18993), .A2(n19206), .ZN(n16865) );
  NOR2_X1 U12340 ( .A1(n16939), .A2(n16938), .ZN(n16937) );
  NOR2_X1 U12341 ( .A1(n17912), .A2(n16962), .ZN(n16961) );
  NOR2_X1 U12342 ( .A1(n16969), .A2(n17924), .ZN(n16968) );
  NOR2_X1 U12343 ( .A1(n17969), .A2(n17001), .ZN(n17000) );
  NAND2_X1 U12344 ( .A1(n16885), .A2(n10313), .ZN(n17058) );
  AND2_X1 U12345 ( .A1(n9801), .A2(n10006), .ZN(n17111) );
  INV_X1 U12346 ( .A(n17259), .ZN(n17244) );
  NOR2_X1 U12347 ( .A1(n17400), .A2(n17414), .ZN(n17385) );
  NAND2_X1 U12348 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17385), .ZN(n17384) );
  INV_X1 U12349 ( .A(n17711), .ZN(n18585) );
  NOR2_X1 U12350 ( .A1(n17811), .A2(n17610), .ZN(n17601) );
  NOR2_X1 U12351 ( .A1(n17807), .A2(n17619), .ZN(n17614) );
  NOR2_X1 U12352 ( .A1(n17623), .A2(n17803), .ZN(n17624) );
  NAND2_X1 U12353 ( .A1(n17624), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17619) );
  NAND2_X1 U12354 ( .A1(n17630), .A2(n17711), .ZN(n17623) );
  NOR2_X1 U12355 ( .A1(n17631), .A2(n17801), .ZN(n17630) );
  NOR2_X1 U12356 ( .A1(n17793), .A2(n17655), .ZN(n17650) );
  INV_X1 U12357 ( .A(n17660), .ZN(n17656) );
  NOR2_X1 U12358 ( .A1(n17787), .A2(n17672), .ZN(n17666) );
  INV_X1 U12359 ( .A(n17649), .ZN(n17664) );
  NAND2_X1 U12360 ( .A1(n9991), .A2(n9992), .ZN(n17672) );
  NOR2_X1 U12361 ( .A1(n9793), .A2(n9993), .ZN(n9992) );
  INV_X1 U12362 ( .A(n17739), .ZN(n9991) );
  NOR2_X1 U12363 ( .A1(n17739), .A2(n9793), .ZN(n17677) );
  INV_X1 U12364 ( .A(n11041), .ZN(n9887) );
  NOR2_X1 U12365 ( .A1(n11042), .A2(n9889), .ZN(n9888) );
  AND2_X1 U12366 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17724), .ZN(n17727) );
  AOI211_X1 U12367 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n11080), .B(n11079), .ZN(n11081) );
  OR2_X1 U12368 ( .A1(n17821), .A2(n17712), .ZN(n17732) );
  AOI211_X1 U12369 ( .C1(n9647), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n11050), .B(n11049), .ZN(n11061) );
  INV_X1 U12370 ( .A(n11284), .ZN(n17744) );
  NOR2_X1 U12371 ( .A1(n17739), .A2(n17819), .ZN(n17737) );
  NOR2_X1 U12372 ( .A1(n11115), .A2(n11114), .ZN(n11116) );
  INV_X1 U12373 ( .A(n11107), .ZN(n11117) );
  NOR2_X1 U12374 ( .A1(n17780), .A2(n17763), .ZN(n17760) );
  CLKBUF_X1 U12375 ( .A(n17760), .Z(n17779) );
  CLKBUF_X1 U12376 ( .A(n17845), .Z(n17848) );
  NOR2_X1 U12377 ( .A1(n17858), .A2(n17859), .ZN(n16735) );
  NAND2_X1 U12378 ( .A1(n17713), .A2(n18199), .ZN(n18058) );
  NOR2_X1 U12379 ( .A1(n11278), .A2(n9754), .ZN(n17926) );
  NOR2_X1 U12380 ( .A1(n11278), .A2(n17976), .ZN(n17965) );
  NOR2_X1 U12381 ( .A1(n18051), .A2(n18053), .ZN(n18037) );
  INV_X1 U12382 ( .A(n18776), .ZN(n18932) );
  OAI22_X1 U12383 ( .A1(n18404), .A2(n18211), .B1(n18058), .B2(n18081), .ZN(
        n18093) );
  INV_X1 U12384 ( .A(n18203), .ZN(n18099) );
  NOR2_X1 U12385 ( .A1(n18125), .A2(n18113), .ZN(n18110) );
  INV_X1 U12386 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18113) );
  INV_X1 U12387 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18125) );
  INV_X1 U12388 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18152) );
  NAND2_X1 U12389 ( .A1(n17199), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18153) );
  INV_X1 U12390 ( .A(n18207), .ZN(n18178) );
  INV_X1 U12391 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18177) );
  INV_X1 U12392 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18193) );
  INV_X1 U12393 ( .A(n17923), .ZN(n18190) );
  NOR2_X1 U12394 ( .A1(n18166), .A2(n18178), .ZN(n18203) );
  OR2_X1 U12395 ( .A1(n17970), .A2(n11277), .ZN(n17923) );
  NOR2_X2 U12396 ( .A1(n18551), .A2(n16865), .ZN(n18196) );
  OAI21_X1 U12397 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19205), .A(n16865), 
        .ZN(n18207) );
  NOR2_X1 U12398 ( .A1(n16753), .A2(n9895), .ZN(n9894) );
  AND2_X1 U12399 ( .A1(n18483), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n9895) );
  INV_X1 U12400 ( .A(n9983), .ZN(n17856) );
  NAND2_X1 U12401 ( .A1(n9876), .A2(n9800), .ZN(n9875) );
  NAND2_X1 U12402 ( .A1(n11148), .A2(n11149), .ZN(n9878) );
  INV_X1 U12403 ( .A(n18472), .ZN(n18493) );
  AND2_X1 U12404 ( .A1(n10169), .A2(n10167), .ZN(n18006) );
  NOR2_X1 U12405 ( .A1(n10168), .A2(n10170), .ZN(n10167) );
  OAI21_X1 U12406 ( .B1(n18997), .B2(n19019), .A(n18996), .ZN(n19015) );
  NOR2_X1 U12407 ( .A1(n18130), .A2(n9974), .ZN(n18074) );
  OAI221_X1 U12408 ( .B1(n12882), .B2(n18988), .C1(n12882), .C2(n12881), .A(
        n19206), .ZN(n18466) );
  NOR2_X1 U12409 ( .A1(n18149), .A2(n18151), .ZN(n18137) );
  NOR2_X1 U12410 ( .A1(n18165), .A2(n18164), .ZN(n18163) );
  NOR2_X1 U12411 ( .A1(n18171), .A2(n11122), .ZN(n18165) );
  NAND2_X1 U12412 ( .A1(n9864), .A2(n18400), .ZN(n18501) );
  INV_X1 U12413 ( .A(n9866), .ZN(n9864) );
  INV_X1 U12414 ( .A(n19007), .ZN(n19002) );
  INV_X1 U12415 ( .A(n18466), .ZN(n18521) );
  NOR2_X1 U12416 ( .A1(n18987), .A2(n18510), .ZN(n18525) );
  INV_X1 U12417 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19030) );
  NAND2_X1 U12418 ( .A1(n19187), .A2(n19223), .ZN(n9871) );
  INV_X1 U12419 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19079) );
  CLKBUF_X1 U12420 ( .A(n19144), .Z(n19137) );
  OR2_X1 U12422 ( .A1(n14921), .A2(n14864), .ZN(n10121) );
  INV_X1 U12423 ( .A(n14673), .ZN(n14692) );
  AND2_X1 U12424 ( .A1(n12841), .A2(n12840), .ZN(n12842) );
  NOR2_X1 U12425 ( .A1(n15364), .A2(n10056), .ZN(n10055) );
  OR2_X1 U12426 ( .A1(n10058), .A2(n15362), .ZN(n10057) );
  NOR2_X1 U12427 ( .A1(n15777), .A2(n19389), .ZN(n10056) );
  NOR2_X1 U12428 ( .A1(n11705), .A2(n11704), .ZN(n11706) );
  NOR2_X1 U12429 ( .A1(n15758), .A2(n16584), .ZN(n11705) );
  AOI21_X1 U12430 ( .B1(n15766), .B2(n16589), .A(n15576), .ZN(n15577) );
  OAI21_X1 U12431 ( .B1(n15768), .B2(n16624), .A(n9730), .ZN(n15772) );
  INV_X1 U12432 ( .A(n9964), .ZN(n15960) );
  OAI21_X1 U12433 ( .B1(n15956), .B2(n15958), .A(n9965), .ZN(n9964) );
  AOI21_X1 U12434 ( .B1(n15959), .B2(n15958), .A(n15957), .ZN(n9965) );
  OAI21_X1 U12435 ( .B1(n10015), .B2(n19061), .A(n10010), .ZN(P3_U2641) );
  AND2_X1 U12436 ( .A1(n10013), .A2(n9745), .ZN(n10010) );
  XNOR2_X1 U12437 ( .A(n9684), .B(n16901), .ZN(n10015) );
  AOI21_X1 U12438 ( .B1(n17256), .B2(P3_REIP_REG_0__SCAN_IN), .A(n9874), .ZN(
        n17262) );
  OR2_X1 U12439 ( .A1(n17739), .A2(n9994), .ZN(n17707) );
  AOI211_X1 U12440 ( .C1(n16723), .C2(n18104), .A(n16722), .B(n16721), .ZN(
        n16727) );
  OAI211_X1 U12441 ( .C1(n9981), .C2(n17855), .A(n9978), .B(n9735), .ZN(
        P3_U2802) );
  NOR2_X1 U12442 ( .A1(n17863), .A2(n9979), .ZN(n9978) );
  OAI21_X1 U12443 ( .B1(n9983), .B2(n9982), .A(n18104), .ZN(n9981) );
  AOI21_X1 U12444 ( .B1(n19190), .B2(n11017), .A(n9868), .ZN(P3_U3290) );
  NOR2_X1 U12445 ( .A1(n19190), .A2(n9869), .ZN(n9868) );
  NAND2_X1 U12446 ( .A1(n9871), .A2(n9870), .ZN(n9869) );
  AOI22_X1 U12447 ( .A1(n19186), .A2(n11017), .B1(P3_STATE2_REG_1__SCAN_IN), 
        .B2(n19188), .ZN(n9870) );
  INV_X1 U12448 ( .A(n12605), .ZN(n12649) );
  AND2_X1 U12449 ( .A1(n11718), .A2(n13358), .ZN(n11768) );
  AND2_X1 U12450 ( .A1(n10281), .A2(n11574), .ZN(n9678) );
  NAND2_X1 U12451 ( .A1(n10361), .A2(n9695), .ZN(n10342) );
  AND2_X1 U12452 ( .A1(n10222), .A2(n14066), .ZN(n9679) );
  NAND2_X1 U12453 ( .A1(n15460), .A2(n9698), .ZN(n9680) );
  INV_X2 U12454 ( .A(n10691), .ZN(n10493) );
  OR2_X2 U12455 ( .A1(n11022), .A2(n19020), .ZN(n17500) );
  NAND2_X1 U12456 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11128), .ZN(
        n9681) );
  OR2_X1 U12457 ( .A1(n11600), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10036) );
  NAND2_X1 U12458 ( .A1(n10231), .A2(n12319), .ZN(n14799) );
  NAND2_X1 U12459 ( .A1(n10356), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10353) );
  NAND2_X1 U12460 ( .A1(n10064), .A2(n10065), .ZN(n10348) );
  AND2_X1 U12461 ( .A1(n12402), .A2(n10241), .ZN(n14746) );
  NAND2_X1 U12462 ( .A1(n11654), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14137) );
  AND2_X1 U12463 ( .A1(n11072), .A2(n11063), .ZN(n9682) );
  NAND2_X1 U12464 ( .A1(n10185), .A2(n15651), .ZN(n9683) );
  AOI21_X1 U12465 ( .B1(n11523), .B2(n16565), .A(n9739), .ZN(n10277) );
  INV_X1 U12466 ( .A(n10277), .ZN(n10189) );
  OR2_X1 U12467 ( .A1(n16908), .A2(n17158), .ZN(n9684) );
  OR3_X1 U12468 ( .A1(n15987), .A2(n10094), .A3(n10096), .ZN(n9685) );
  AND3_X1 U12469 ( .A1(n11256), .A2(n19212), .A3(n11255), .ZN(n9686) );
  AND2_X1 U12470 ( .A1(n10065), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9687) );
  AND2_X1 U12471 ( .A1(n9977), .A2(n9975), .ZN(n9688) );
  NAND2_X1 U12472 ( .A1(n12516), .A2(n12515), .ZN(n14721) );
  AND2_X1 U12473 ( .A1(n10091), .A2(n10089), .ZN(n9689) );
  AND2_X1 U12474 ( .A1(n11913), .A2(n11912), .ZN(n9690) );
  AND2_X1 U12475 ( .A1(n12402), .A2(n9757), .ZN(n14734) );
  NOR2_X1 U12476 ( .A1(n10170), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9691) );
  AND2_X1 U12477 ( .A1(n10268), .A2(n10267), .ZN(n9692) );
  NOR2_X1 U12478 ( .A1(n11132), .A2(n9734), .ZN(n9977) );
  NAND2_X1 U12479 ( .A1(n10336), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10335) );
  NAND2_X1 U12480 ( .A1(n10221), .A2(n10222), .ZN(n14065) );
  AND2_X1 U12481 ( .A1(n15475), .A2(n9781), .ZN(n12930) );
  AND2_X1 U12482 ( .A1(n10061), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9693) );
  AND2_X1 U12483 ( .A1(n19376), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9694) );
  AND2_X1 U12484 ( .A1(n9758), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9695) );
  AND2_X1 U12485 ( .A1(n12104), .A2(n13658), .ZN(n9696) );
  AND2_X1 U12486 ( .A1(n13478), .A2(n13483), .ZN(n9697) );
  INV_X1 U12487 ( .A(n13637), .ZN(n10026) );
  NAND2_X1 U12488 ( .A1(n10336), .A2(n9693), .ZN(n10332) );
  AND2_X1 U12489 ( .A1(n10219), .A2(n15461), .ZN(n9698) );
  INV_X1 U12490 ( .A(n9637), .ZN(n11676) );
  AND2_X1 U12491 ( .A1(n9784), .A2(n18109), .ZN(n9699) );
  AND2_X1 U12492 ( .A1(n16437), .A2(n10120), .ZN(n9700) );
  AND2_X1 U12493 ( .A1(n9698), .A2(n10218), .ZN(n9701) );
  AND2_X1 U12494 ( .A1(n11676), .A2(n9797), .ZN(n9702) );
  AND4_X1 U12495 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n9703) );
  AND2_X1 U12496 ( .A1(n10073), .A2(n10072), .ZN(n9704) );
  AND2_X1 U12497 ( .A1(n9802), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n9705) );
  NOR2_X1 U12498 ( .A1(n9653), .A2(n14322), .ZN(n10128) );
  OR2_X1 U12499 ( .A1(n14739), .A2(n14723), .ZN(n9706) );
  NAND2_X2 U12500 ( .A1(n13335), .A2(n13056), .ZN(n10860) );
  INV_X1 U12501 ( .A(n12586), .ZN(n12639) );
  AND2_X2 U12502 ( .A1(n14594), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10779) );
  OR2_X1 U12503 ( .A1(n10309), .A2(n10134), .ZN(n9707) );
  NAND2_X1 U12504 ( .A1(n13358), .A2(n10047), .ZN(n11842) );
  BUF_X1 U12505 ( .A(n10477), .Z(n10792) );
  AND2_X1 U12506 ( .A1(n12707), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9708) );
  NAND2_X1 U12507 ( .A1(n9845), .A2(n9844), .ZN(n10037) );
  NAND2_X1 U12508 ( .A1(n17971), .A2(n17954), .ZN(n17955) );
  AND2_X2 U12509 ( .A1(n9660), .A2(n10680), .ZN(n10766) );
  NOR2_X1 U12510 ( .A1(n15694), .A2(n15899), .ZN(n15677) );
  AND2_X1 U12511 ( .A1(n10231), .A2(n10230), .ZN(n9711) );
  NAND2_X1 U12512 ( .A1(n11602), .A2(n11008), .ZN(n11513) );
  NAND2_X1 U12513 ( .A1(n12754), .A2(n15224), .ZN(n15019) );
  NOR2_X1 U12514 ( .A1(n10349), .A2(n16564), .ZN(n10350) );
  AND2_X1 U12515 ( .A1(n10356), .A2(n10069), .ZN(n9712) );
  OR2_X1 U12516 ( .A1(n11539), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n9713) );
  NOR2_X2 U12517 ( .A1(n17713), .A2(n18210), .ZN(n18104) );
  AND4_X1 U12518 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n9714) );
  OR2_X1 U12519 ( .A1(n10209), .A2(n10212), .ZN(n9715) );
  OR2_X1 U12520 ( .A1(n9862), .A2(n19212), .ZN(n9716) );
  AND2_X1 U12521 ( .A1(n10555), .A2(n10261), .ZN(n9717) );
  NOR2_X1 U12522 ( .A1(n17247), .A2(n11018), .ZN(n11068) );
  INV_X1 U12523 ( .A(n11068), .ZN(n14198) );
  NOR2_X1 U12524 ( .A1(n15998), .A2(n11535), .ZN(n9718) );
  NAND2_X1 U12525 ( .A1(n10352), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10349) );
  OR2_X1 U12526 ( .A1(n15224), .A2(n15275), .ZN(n9719) );
  AOI21_X1 U12527 ( .B1(n10530), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10531), .ZN(n13184) );
  INV_X1 U12528 ( .A(n13184), .ZN(n10183) );
  NAND2_X1 U12529 ( .A1(n15251), .A2(n12741), .ZN(n15069) );
  OR3_X1 U12530 ( .A1(n12957), .A2(n11667), .A3(n15855), .ZN(n9720) );
  INV_X1 U12531 ( .A(n17785), .ZN(n9862) );
  NAND2_X1 U12532 ( .A1(n10032), .A2(n10031), .ZN(n15870) );
  AND2_X1 U12533 ( .A1(n16525), .A2(n16522), .ZN(n9721) );
  NOR2_X1 U12534 ( .A1(n15905), .A2(n10097), .ZN(n12933) );
  AND3_X1 U12535 ( .A1(n15000), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9722) );
  XNOR2_X1 U12536 ( .A(n11998), .B(n11996), .ZN(n12105) );
  NAND2_X1 U12537 ( .A1(n13053), .A2(n13052), .ZN(n13171) );
  AND2_X1 U12538 ( .A1(n10252), .A2(n13694), .ZN(n9723) );
  AND3_X1 U12539 ( .A1(n11837), .A2(n11835), .A3(n11836), .ZN(n11887) );
  INV_X1 U12540 ( .A(n11352), .ZN(n13903) );
  NAND2_X1 U12541 ( .A1(n10175), .A2(n17857), .ZN(n16114) );
  NAND2_X1 U12542 ( .A1(n13498), .A2(n14002), .ZN(n13212) );
  AND3_X1 U12543 ( .A1(n9892), .A2(n11043), .A3(n9890), .ZN(n9724) );
  AND2_X1 U12544 ( .A1(n9718), .A2(n10277), .ZN(n9725) );
  NOR2_X1 U12545 ( .A1(n19212), .A2(n18545), .ZN(n11275) );
  AND4_X1 U12546 ( .A1(n11841), .A2(n11840), .A3(n11839), .A4(n11838), .ZN(
        n9726) );
  NAND2_X1 U12547 ( .A1(n9878), .A2(n9875), .ZN(n17869) );
  INV_X1 U12548 ( .A(n17869), .ZN(n9984) );
  INV_X1 U12549 ( .A(n14809), .ZN(n10231) );
  OR2_X1 U12550 ( .A1(n15694), .A2(n9942), .ZN(n9946) );
  AND2_X1 U12551 ( .A1(n15567), .A2(n15581), .ZN(n9727) );
  INV_X1 U12552 ( .A(n10129), .ZN(n14683) );
  NOR2_X1 U12553 ( .A1(n9706), .A2(n10131), .ZN(n10129) );
  AND2_X1 U12554 ( .A1(n11873), .A2(n11872), .ZN(n9728) );
  NOR2_X1 U12555 ( .A1(n15658), .A2(n11575), .ZN(n9729) );
  AND2_X1 U12556 ( .A1(n15770), .A2(n10103), .ZN(n9730) );
  OR2_X1 U12557 ( .A1(n10162), .A2(n10161), .ZN(n9731) );
  NOR2_X1 U12558 ( .A1(n15597), .A2(n9909), .ZN(n9732) );
  AND2_X1 U12559 ( .A1(n16744), .A2(n10317), .ZN(n16745) );
  AND2_X1 U12560 ( .A1(n12718), .A2(n13303), .ZN(n9733) );
  NAND2_X1 U12561 ( .A1(n18109), .A2(n18442), .ZN(n9734) );
  OR2_X1 U12562 ( .A1(n17874), .A2(n17866), .ZN(n9735) );
  AND2_X1 U12563 ( .A1(n12728), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9736) );
  AND2_X1 U12564 ( .A1(n9954), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9737) );
  NAND2_X1 U12565 ( .A1(n10499), .A2(n10481), .ZN(n10472) );
  AND2_X1 U12566 ( .A1(n12796), .A2(n13084), .ZN(n9738) );
  INV_X1 U12567 ( .A(n14707), .ZN(n10243) );
  NAND2_X1 U12568 ( .A1(n16550), .A2(n16548), .ZN(n9739) );
  NAND2_X1 U12569 ( .A1(n12402), .A2(n12401), .ZN(n14757) );
  AND2_X1 U12570 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17539), .ZN(n9740) );
  AND2_X1 U12571 ( .A1(n11069), .A2(n9986), .ZN(n9741) );
  AND2_X1 U12572 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n9742) );
  INV_X1 U12573 ( .A(n10153), .ZN(n10152) );
  NAND2_X1 U12574 ( .A1(n9719), .A2(n12739), .ZN(n10153) );
  AND3_X1 U12575 ( .A1(n11066), .A2(n10305), .A3(n11065), .ZN(n9743) );
  AND2_X1 U12576 ( .A1(n11259), .A2(n18573), .ZN(n9744) );
  AND3_X1 U12577 ( .A1(n10012), .A2(n16903), .A3(n10011), .ZN(n9745) );
  OR2_X1 U12578 ( .A1(n11119), .A2(n18508), .ZN(n9746) );
  AND3_X1 U12579 ( .A1(n19177), .A2(n19185), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9747) );
  OR2_X1 U12580 ( .A1(n11241), .A2(n18560), .ZN(n9748) );
  NAND2_X2 U12581 ( .A1(n10431), .A2(n10430), .ZN(n10481) );
  AND2_X1 U12582 ( .A1(n11513), .A2(n10570), .ZN(n9749) );
  AND2_X1 U12583 ( .A1(n10251), .A2(n10250), .ZN(n9750) );
  AND2_X1 U12584 ( .A1(n13143), .A2(n10494), .ZN(n10518) );
  INV_X1 U12585 ( .A(n9644), .ZN(n13178) );
  NAND2_X1 U12586 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11124), .ZN(
        n9751) );
  INV_X2 U12587 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19177) );
  OR2_X1 U12588 ( .A1(n11062), .A2(n17532), .ZN(n9752) );
  INV_X1 U12589 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13923) );
  INV_X1 U12590 ( .A(n11860), .ZN(n11798) );
  AND2_X1 U12591 ( .A1(n13572), .A2(n13370), .ZN(n11860) );
  INV_X1 U12592 ( .A(n12429), .ZN(n12546) );
  INV_X1 U12593 ( .A(n18109), .ZN(n9883) );
  INV_X1 U12594 ( .A(n15690), .ZN(n9924) );
  AND2_X1 U12595 ( .A1(n10361), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10344) );
  NOR2_X1 U12596 ( .A1(n18108), .A2(n11137), .ZN(n18028) );
  NAND2_X1 U12597 ( .A1(n15475), .A2(n15385), .ZN(n15384) );
  NAND2_X1 U12598 ( .A1(n15460), .A2(n15461), .ZN(n15455) );
  NOR2_X1 U12599 ( .A1(n16006), .A2(n13890), .ZN(n13889) );
  NOR2_X1 U12600 ( .A1(n10349), .A2(n10063), .ZN(n10347) );
  OR3_X1 U12601 ( .A1(n10309), .A2(n14840), .A3(n10137), .ZN(n9753) );
  NAND2_X1 U12602 ( .A1(n10001), .A2(n10000), .ZN(n9754) );
  AND2_X1 U12603 ( .A1(n16221), .A2(n10073), .ZN(n9755) );
  AND2_X1 U12604 ( .A1(n11887), .A2(n11853), .ZN(n13080) );
  AND2_X1 U12605 ( .A1(n10257), .A2(n10256), .ZN(n9756) );
  AND2_X1 U12606 ( .A1(n10238), .A2(n14009), .ZN(n14008) );
  NOR2_X1 U12607 ( .A1(n10235), .A2(n10237), .ZN(n14074) );
  NAND2_X1 U12608 ( .A1(n9841), .A2(n9840), .ZN(n16047) );
  NAND2_X1 U12609 ( .A1(n9839), .A2(n11509), .ZN(n15720) );
  AND2_X1 U12610 ( .A1(n14748), .A2(n10241), .ZN(n9757) );
  NAND2_X1 U12611 ( .A1(n12080), .A2(n12079), .ZN(n14009) );
  AND2_X1 U12612 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n9758) );
  AND2_X1 U12613 ( .A1(n15682), .A2(n15681), .ZN(n9759) );
  OR2_X1 U12614 ( .A1(n10792), .A2(n10590), .ZN(n9760) );
  NOR3_X1 U12615 ( .A1(n12946), .A2(n11667), .A3(n15882), .ZN(n9761) );
  INV_X1 U12616 ( .A(n10148), .ZN(n13300) );
  XNOR2_X1 U12617 ( .A(n14505), .B(n14506), .ZN(n15422) );
  NOR3_X1 U12618 ( .A1(n15987), .A2(n10096), .A3(n14043), .ZN(n14113) );
  NAND2_X1 U12619 ( .A1(n13183), .A2(n13182), .ZN(n13282) );
  AND2_X1 U12620 ( .A1(n10361), .A2(n9758), .ZN(n10343) );
  AND2_X1 U12621 ( .A1(n15460), .A2(n9701), .ZN(n15442) );
  AND2_X1 U12622 ( .A1(n10102), .A2(n13620), .ZN(n9762) );
  AND2_X1 U12623 ( .A1(n16700), .A2(n20263), .ZN(n9763) );
  XOR2_X1 U12624 ( .A(n15724), .B(n16040), .Z(n9764) );
  AND2_X1 U12625 ( .A1(n9918), .A2(n9922), .ZN(n9765) );
  NAND2_X1 U12626 ( .A1(n13176), .A2(n13175), .ZN(n13183) );
  AND2_X1 U12627 ( .A1(n13423), .A2(n13511), .ZN(n9766) );
  AND2_X1 U12628 ( .A1(n11531), .A2(n9760), .ZN(n9767) );
  NOR2_X1 U12629 ( .A1(n15437), .A2(n10204), .ZN(n9768) );
  INV_X1 U12630 ( .A(n19212), .ZN(n18551) );
  AND2_X1 U12631 ( .A1(n16221), .A2(n9704), .ZN(n9769) );
  NAND2_X1 U12632 ( .A1(n12004), .A2(n15325), .ZN(n9770) );
  OR2_X1 U12633 ( .A1(n10713), .A2(n10712), .ZN(n11001) );
  INV_X1 U12634 ( .A(n10285), .ZN(n9920) );
  NAND2_X1 U12635 ( .A1(n10287), .A2(n10286), .ZN(n10285) );
  AND2_X1 U12636 ( .A1(n10052), .A2(n9658), .ZN(n9771) );
  INV_X1 U12637 ( .A(n14826), .ZN(n10138) );
  OR2_X1 U12638 ( .A1(n18987), .A2(n12880), .ZN(n9772) );
  OR2_X1 U12639 ( .A1(n11648), .A2(n15732), .ZN(n9773) );
  AND2_X1 U12640 ( .A1(n10249), .A2(n10248), .ZN(n9774) );
  OR2_X1 U12641 ( .A1(n10873), .A2(n10872), .ZN(n13483) );
  AND2_X1 U12642 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9775) );
  INV_X1 U12643 ( .A(n14708), .ZN(n12541) );
  NAND2_X1 U12644 ( .A1(n9949), .A2(n15081), .ZN(n9950) );
  AND2_X1 U12645 ( .A1(n9901), .A2(n9694), .ZN(n9776) );
  INV_X1 U12646 ( .A(n10271), .ZN(n10270) );
  NAND2_X1 U12647 ( .A1(n9924), .A2(n15681), .ZN(n10271) );
  CLKBUF_X3 U12648 ( .A(n10362), .Z(n19393) );
  OR2_X1 U12649 ( .A1(n15905), .A2(n10098), .ZN(n9777) );
  AND2_X1 U12650 ( .A1(n9757), .A2(n14736), .ZN(n9778) );
  AND2_X1 U12651 ( .A1(n10064), .A2(n9687), .ZN(n9779) );
  OR2_X1 U12652 ( .A1(n10022), .A2(n10025), .ZN(n9780) );
  AND2_X1 U12653 ( .A1(n9756), .A2(n10255), .ZN(n9781) );
  AND2_X1 U12654 ( .A1(n9695), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9782) );
  OR2_X1 U12655 ( .A1(n11427), .A2(n10111), .ZN(n9783) );
  INV_X1 U12656 ( .A(n12538), .ZN(n12630) );
  INV_X1 U12657 ( .A(n12630), .ZN(n13667) );
  NAND2_X2 U12658 ( .A1(n11725), .A2(n13362), .ZN(n11822) );
  NOR2_X1 U12659 ( .A1(n10742), .A2(n10092), .ZN(n10091) );
  INV_X1 U12660 ( .A(n18315), .ZN(n9880) );
  INV_X1 U12661 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U12662 ( .A1(n13372), .A2(n13286), .ZN(n13479) );
  NAND2_X1 U12663 ( .A1(n13479), .A2(n13478), .ZN(n13481) );
  AND2_X1 U12664 ( .A1(n10340), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10338) );
  NOR2_X1 U12665 ( .A1(n13832), .A2(n13831), .ZN(n13933) );
  AND2_X1 U12666 ( .A1(n13479), .A2(n9697), .ZN(n13603) );
  NOR2_X1 U12667 ( .A1(n13832), .A2(n10220), .ZN(n14363) );
  AND2_X1 U12668 ( .A1(n10361), .A2(n9782), .ZN(n10340) );
  INV_X1 U12669 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10070) );
  AND2_X1 U12670 ( .A1(n17857), .A2(n16121), .ZN(n9784) );
  AND2_X1 U12671 ( .A1(n10336), .A2(n10061), .ZN(n9785) );
  AND2_X1 U12672 ( .A1(n14483), .A2(n10205), .ZN(n9786) );
  AND2_X1 U12673 ( .A1(n10338), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10336) );
  INV_X1 U12674 ( .A(n15997), .ZN(n10273) );
  NAND2_X1 U12675 ( .A1(n10221), .A2(n9679), .ZN(n10224) );
  NAND2_X1 U12676 ( .A1(n11876), .A2(n13521), .ZN(n10148) );
  NOR2_X1 U12677 ( .A1(n18137), .A2(n18136), .ZN(n9787) );
  NAND2_X1 U12678 ( .A1(n11993), .A2(n11992), .ZN(n13944) );
  INV_X1 U12679 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10068) );
  INV_X1 U12680 ( .A(n13832), .ZN(n10221) );
  OR2_X1 U12681 ( .A1(n10947), .A2(n10946), .ZN(n13934) );
  INV_X1 U12682 ( .A(n13934), .ZN(n10223) );
  NAND2_X1 U12683 ( .A1(n14483), .A2(n14482), .ZN(n9788) );
  OR2_X1 U12684 ( .A1(n18109), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9789) );
  AND2_X1 U12685 ( .A1(n9701), .A2(n15443), .ZN(n9790) );
  AND2_X1 U12686 ( .A1(n10054), .A2(n10337), .ZN(n9791) );
  AND2_X1 U12687 ( .A1(n10254), .A2(n10253), .ZN(n9792) );
  OR2_X1 U12688 ( .A1(n10775), .A2(n10774), .ZN(n11650) );
  NOR2_X1 U12689 ( .A1(n18152), .A2(n10009), .ZN(n10008) );
  NOR2_X1 U12690 ( .A1(n10331), .A2(n15586), .ZN(n10324) );
  AND2_X2 U12691 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13381) );
  AND2_X1 U12692 ( .A1(n10336), .A2(n10060), .ZN(n10328) );
  OR2_X1 U12693 ( .A1(n9994), .A2(n9995), .ZN(n9793) );
  AND2_X1 U12694 ( .A1(n11134), .A2(n11133), .ZN(n9794) );
  AND3_X1 U12695 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .ZN(n9795) );
  AND2_X1 U12696 ( .A1(n11676), .A2(n9904), .ZN(n9796) );
  AND2_X1 U12697 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12832), .ZN(n9797) );
  AND2_X1 U12698 ( .A1(n10119), .A2(n11613), .ZN(n9798) );
  NAND2_X1 U12699 ( .A1(n9997), .A2(n10001), .ZN(n17933) );
  NOR2_X1 U12700 ( .A1(n18153), .A2(n18152), .ZN(n17171) );
  AND2_X1 U12701 ( .A1(n10008), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9799) );
  NAND2_X1 U12702 ( .A1(n17999), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11278) );
  AND2_X1 U12703 ( .A1(n18228), .A2(n11149), .ZN(n9800) );
  AND2_X1 U12704 ( .A1(n10007), .A2(n9799), .ZN(n9801) );
  INV_X1 U12705 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n10076) );
  INV_X1 U12706 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n10074) );
  AND2_X1 U12707 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17199) );
  INV_X1 U12708 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n9993) );
  INV_X1 U12709 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9999) );
  INV_X1 U12710 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16176) );
  AND2_X1 U12711 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n9802) );
  AND2_X1 U12712 ( .A1(n9705), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n9803) );
  INV_X1 U12713 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U12714 ( .A1(n20239), .A2(n19710), .ZN(n9804) );
  INV_X1 U12715 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20239) );
  OAI22_X1 U12716 ( .A1(n21061), .A2(n15340), .B1(n16774), .B2(n15341), .ZN(
        n9805) );
  NAND2_X1 U12717 ( .A1(n16286), .A2(n14923), .ZN(n15341) );
  NAND3_X2 U12718 ( .A1(n19223), .A2(n19052), .A3(n19222), .ZN(n18522) );
  OAI22_X2 U12719 ( .A1(n16763), .A2(n15341), .B1(n21160), .B2(n15340), .ZN(
        n20921) );
  INV_X1 U12720 ( .A(n20891), .ZN(n9806) );
  INV_X1 U12721 ( .A(n9806), .ZN(n9807) );
  INV_X1 U12722 ( .A(n20927), .ZN(n9808) );
  INV_X1 U12723 ( .A(n9808), .ZN(n9809) );
  INV_X1 U12724 ( .A(n20897), .ZN(n9810) );
  INV_X1 U12725 ( .A(n9810), .ZN(n9811) );
  INV_X1 U12726 ( .A(n20903), .ZN(n9812) );
  INV_X1 U12727 ( .A(n9812), .ZN(n9813) );
  OAI22_X2 U12728 ( .A1(n16765), .A2(n15341), .B1(n21068), .B2(n15340), .ZN(
        n20915) );
  AOI22_X2 U12729 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19608), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19607), .ZN(n20107) );
  NOR3_X2 U12730 ( .A1(n18900), .A2(n18856), .A3(n18831), .ZN(n18825) );
  OAI22_X2 U12731 ( .A1(n21222), .A2(n15340), .B1(n19612), .B2(n15341), .ZN(
        n20869) );
  NAND2_X1 U12732 ( .A1(n9814), .A2(n10518), .ZN(n9816) );
  NAND2_X1 U12733 ( .A1(n10516), .A2(n11676), .ZN(n9814) );
  XNOR2_X1 U12734 ( .A(n10476), .B(n10477), .ZN(n13029) );
  OR2_X2 U12735 ( .A1(n15694), .A2(n9945), .ZN(n15667) );
  NAND2_X1 U12737 ( .A1(n9825), .A2(n9823), .ZN(n15868) );
  NAND2_X1 U12738 ( .A1(n15869), .A2(n15882), .ZN(n9824) );
  NAND2_X2 U12739 ( .A1(n9826), .A2(n9842), .ZN(n19569) );
  NAND2_X2 U12740 ( .A1(n9826), .A2(n11354), .ZN(n13760) );
  NAND2_X2 U12741 ( .A1(n9843), .A2(n9826), .ZN(n19647) );
  AND2_X2 U12742 ( .A1(n11339), .A2(n9675), .ZN(n9826) );
  NAND2_X1 U12743 ( .A1(n10278), .A2(n11656), .ZN(n9827) );
  NAND2_X1 U12744 ( .A1(n9831), .A2(n9959), .ZN(n9828) );
  NAND2_X1 U12745 ( .A1(n9831), .A2(n9830), .ZN(n9829) );
  NOR2_X2 U12746 ( .A1(n10278), .A2(n11655), .ZN(n9831) );
  XNOR2_X2 U12747 ( .A(n11327), .B(n11326), .ZN(n13271) );
  NAND2_X1 U12748 ( .A1(n10180), .A2(n11328), .ZN(n9832) );
  NAND2_X2 U12749 ( .A1(n10529), .A2(n10528), .ZN(n11328) );
  INV_X1 U12750 ( .A(n15593), .ZN(n9838) );
  NAND2_X2 U12751 ( .A1(n9846), .A2(n10458), .ZN(n10672) );
  INV_X1 U12752 ( .A(n13117), .ZN(n10501) );
  NAND2_X1 U12753 ( .A1(n10515), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10539) );
  OR2_X2 U12754 ( .A1(n11652), .A2(n11651), .ZN(n14024) );
  INV_X1 U12755 ( .A(n15235), .ZN(n10151) );
  NOR2_X1 U12756 ( .A1(n9938), .A2(n12740), .ZN(n9957) );
  INV_X1 U12757 ( .A(n16745), .ZN(n10177) );
  NAND2_X1 U12758 ( .A1(n11143), .A2(n10311), .ZN(n11144) );
  NOR2_X2 U12759 ( .A1(n18150), .A2(n18467), .ZN(n18149) );
  INV_X1 U12760 ( .A(n11544), .ZN(n10114) );
  INV_X1 U12761 ( .A(n11426), .ZN(n10110) );
  INV_X1 U12762 ( .A(n15642), .ZN(n9912) );
  OAI21_X1 U12763 ( .B1(n9957), .B2(n9956), .A(n12749), .ZN(n12752) );
  INV_X1 U12764 ( .A(n12098), .ZN(n9940) );
  NOR2_X2 U12765 ( .A1(n14809), .A2(n10229), .ZN(n14770) );
  NAND2_X1 U12766 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17415), .ZN(n17414) );
  OR2_X1 U12767 ( .A1(n19272), .A2(n11667), .ZN(n11545) );
  INV_X1 U12768 ( .A(n11650), .ZN(n11431) );
  NAND2_X1 U12769 ( .A1(n9911), .A2(n16014), .ZN(n9910) );
  INV_X1 U12770 ( .A(n10116), .ZN(n11548) );
  NAND2_X2 U12771 ( .A1(n14680), .A2(n14262), .ZN(n15003) );
  OR2_X2 U12772 ( .A1(n12097), .A2(n12098), .ZN(n12121) );
  NAND2_X1 U12773 ( .A1(n11910), .A2(n11892), .ZN(n11911) );
  NOR2_X1 U12774 ( .A1(n14707), .A2(n14695), .ZN(n14694) );
  OAI21_X1 U12775 ( .B1(n15185), .B2(n20282), .A(n15007), .ZN(P1_U2971) );
  NAND3_X1 U12776 ( .A1(n11242), .A2(n9847), .A3(n11243), .ZN(n11244) );
  NAND4_X1 U12777 ( .A1(n9857), .A2(n9856), .A3(n9748), .A4(n9855), .ZN(n9854)
         );
  AND2_X1 U12778 ( .A1(n18400), .A2(n18382), .ZN(n18440) );
  INV_X1 U12779 ( .A(n11137), .ZN(n9881) );
  NOR2_X1 U12780 ( .A1(n18432), .A2(n18109), .ZN(n18108) );
  INV_X1 U12781 ( .A(n18432), .ZN(n9884) );
  NOR2_X2 U12782 ( .A1(n18131), .A2(n18132), .ZN(n18130) );
  XNOR2_X1 U12783 ( .A(n11131), .B(n11130), .ZN(n18131) );
  OAI21_X1 U12784 ( .B1(n18149), .B2(n10166), .A(n10165), .ZN(n11131) );
  NAND3_X1 U12785 ( .A1(n9897), .A2(n18522), .A3(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9896) );
  OAI21_X1 U12786 ( .B1(n9899), .B2(n9902), .A(n11467), .ZN(n9898) );
  OAI21_X1 U12787 ( .B1(n11428), .B2(n9903), .A(n9776), .ZN(n9899) );
  NAND2_X1 U12788 ( .A1(n10178), .A2(n9694), .ZN(n9914) );
  NAND2_X1 U12789 ( .A1(n9900), .A2(n11430), .ZN(n14124) );
  OR2_X1 U12790 ( .A1(n10302), .A2(n9903), .ZN(n9901) );
  NAND2_X1 U12791 ( .A1(n10467), .A2(n9906), .ZN(n12972) );
  NAND2_X1 U12792 ( .A1(n11685), .A2(n9637), .ZN(n11684) );
  NOR2_X1 U12793 ( .A1(n16662), .A2(n9637), .ZN(n20245) );
  NAND2_X1 U12794 ( .A1(n9637), .A2(n11673), .ZN(n9905) );
  MUX2_X1 U12795 ( .A(n10999), .B(n11673), .S(n9637), .Z(n11622) );
  MUX2_X1 U12796 ( .A(n11002), .B(n11380), .S(n11676), .Z(n11003) );
  MUX2_X1 U12797 ( .A(n11431), .B(n11004), .S(n9637), .Z(n11005) );
  NAND2_X1 U12798 ( .A1(n10178), .A2(n19376), .ZN(n11466) );
  INV_X1 U12799 ( .A(n10265), .ZN(n15702) );
  INV_X1 U12800 ( .A(n9928), .ZN(n12845) );
  OAI21_X2 U12801 ( .B1(n9932), .B2(n9931), .A(n9929), .ZN(n16295) );
  NAND3_X1 U12802 ( .A1(n13498), .A2(n13870), .A3(n14002), .ZN(n13354) );
  NOR2_X1 U12803 ( .A1(n14322), .A2(n9934), .ZN(n13203) );
  NAND2_X1 U12804 ( .A1(n11899), .A2(n9934), .ZN(n13351) );
  NOR2_X1 U12805 ( .A1(n13212), .A2(n21042), .ZN(n9935) );
  XNOR2_X2 U12806 ( .A(n12001), .B(n20583), .ZN(n13342) );
  NAND2_X2 U12807 ( .A1(n9937), .A2(n9936), .ZN(n12001) );
  XNOR2_X1 U12808 ( .A(n10228), .B(n9939), .ZN(n12701) );
  AND3_X2 U12809 ( .A1(n10046), .A2(n9940), .A3(n20581), .ZN(n10228) );
  OAI21_X2 U12810 ( .B1(n15063), .B2(n10038), .A(n15018), .ZN(n15052) );
  OAI21_X2 U12811 ( .B1(n15063), .B2(n16163), .A(n9952), .ZN(n12754) );
  NAND2_X2 U12812 ( .A1(n12752), .A2(n12751), .ZN(n15063) );
  NAND2_X1 U12813 ( .A1(n9958), .A2(n14139), .ZN(n9941) );
  AND3_X2 U12814 ( .A1(n11416), .A2(n11650), .A3(n11415), .ZN(n11469) );
  NOR2_X2 U12815 ( .A1(n15619), .A2(n15783), .ZN(n15817) );
  OR2_X2 U12816 ( .A1(n15694), .A2(n9943), .ZN(n15630) );
  INV_X1 U12817 ( .A(n9946), .ZN(n15644) );
  NAND2_X2 U12818 ( .A1(n12668), .A2(n12670), .ZN(n12742) );
  NOR2_X1 U12819 ( .A1(n9950), .A2(n9947), .ZN(n15236) );
  INV_X1 U12820 ( .A(n16276), .ZN(n9947) );
  OAI21_X1 U12821 ( .B1(n15018), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15102), .ZN(n9951) );
  AND2_X2 U12822 ( .A1(n11718), .A2(n11725), .ZN(n11847) );
  AND2_X2 U12823 ( .A1(n9955), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11725) );
  INV_X2 U12824 ( .A(n13499), .ZN(n14002) );
  NAND2_X2 U12825 ( .A1(n10123), .A2(n11852), .ZN(n13499) );
  NAND3_X1 U12826 ( .A1(n13178), .A2(n13903), .A3(n11371), .ZN(n13858) );
  AND2_X2 U12827 ( .A1(n13271), .A2(n13162), .ZN(n11371) );
  NAND2_X1 U12828 ( .A1(n14139), .A2(n14136), .ZN(n11657) );
  NAND2_X1 U12829 ( .A1(n11416), .A2(n11415), .ZN(n11649) );
  INV_X1 U12830 ( .A(n11415), .ZN(n9960) );
  OAI21_X2 U12831 ( .B1(n11416), .B2(n11415), .A(n11649), .ZN(n13981) );
  NAND2_X2 U12832 ( .A1(n16572), .A2(n11670), .ZN(n16024) );
  NAND3_X1 U12833 ( .A1(n9971), .A2(n10169), .A3(n9691), .ZN(n18004) );
  NAND3_X1 U12834 ( .A1(n10160), .A2(n10158), .A3(n9751), .ZN(n11127) );
  INV_X1 U12835 ( .A(n18130), .ZN(n9976) );
  AND2_X2 U12836 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n9747), .ZN(
        n17547) );
  OAI211_X1 U12837 ( .C1(n9987), .C2(n12868), .A(n9988), .B(n11248), .ZN(n9989) );
  INV_X1 U12838 ( .A(n12868), .ZN(n9990) );
  NAND3_X1 U12839 ( .A1(n11161), .A2(n11160), .A3(n9996), .ZN(n11162) );
  INV_X1 U12840 ( .A(n11278), .ZN(n9997) );
  NAND2_X1 U12841 ( .A1(n9997), .A2(n9998), .ZN(n17898) );
  XNOR2_X2 U12842 ( .A(n16719), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16885) );
  INV_X1 U12843 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10009) );
  OAI21_X1 U12844 ( .B1(n15762), .B2(n16651), .A(n10016), .ZN(P2_U3015) );
  XNOR2_X1 U12845 ( .A(n10017), .B(n11621), .ZN(n15762) );
  NAND2_X1 U12846 ( .A1(n13981), .A2(n9780), .ZN(n10018) );
  NAND2_X1 U12847 ( .A1(n10018), .A2(n10019), .ZN(n14026) );
  INV_X1 U12848 ( .A(n12097), .ZN(n10046) );
  INV_X2 U12849 ( .A(n11842), .ZN(n11744) );
  NAND2_X2 U12850 ( .A1(n10126), .A2(n9728), .ZN(n13958) );
  NAND2_X1 U12851 ( .A1(n10051), .A2(n10053), .ZN(n15365) );
  NAND2_X1 U12852 ( .A1(n12954), .A2(n9791), .ZN(n10051) );
  NAND2_X1 U12853 ( .A1(n10057), .A2(n10055), .ZN(P2_U2826) );
  NAND2_X1 U12854 ( .A1(n15363), .A2(n15588), .ZN(n10059) );
  NAND3_X1 U12855 ( .A1(n10356), .A2(n10069), .A3(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10351) );
  NAND2_X1 U12856 ( .A1(n14717), .A2(n9705), .ZN(n14673) );
  AOI21_X1 U12857 ( .B1(n14717), .B2(n9803), .A(P1_REIP_REG_30__SCAN_IN), .ZN(
        n14675) );
  NAND2_X2 U12858 ( .A1(n21047), .A2(n13669), .ZN(n14099) );
  AND2_X2 U12859 ( .A1(n12808), .A2(n12807), .ZN(n16159) );
  AOI21_X1 U12860 ( .B1(n10079), .B2(n10078), .A(n9738), .ZN(n12797) );
  NAND2_X1 U12861 ( .A1(n10081), .A2(n10080), .ZN(n10079) );
  NAND2_X1 U12862 ( .A1(n10083), .A2(n10082), .ZN(n10081) );
  NAND2_X1 U12863 ( .A1(n12792), .A2(n12793), .ZN(n10082) );
  NAND2_X1 U12864 ( .A1(n12791), .A2(n12790), .ZN(n10083) );
  INV_X2 U12865 ( .A(n13958), .ZN(n13498) );
  INV_X1 U12866 ( .A(n13323), .ZN(n10087) );
  NAND2_X1 U12867 ( .A1(n10087), .A2(n9689), .ZN(n16052) );
  AND2_X1 U12868 ( .A1(n10977), .A2(n10106), .ZN(n15488) );
  NAND2_X1 U12869 ( .A1(n10977), .A2(n10105), .ZN(n12826) );
  INV_X1 U12870 ( .A(n10977), .ZN(n15513) );
  INV_X1 U12871 ( .A(n15499), .ZN(n10108) );
  NAND2_X1 U12872 ( .A1(n10110), .A2(n10109), .ZN(n11512) );
  NOR2_X2 U12873 ( .A1(n11512), .A2(n11510), .ZN(n11515) );
  MUX2_X1 U12874 ( .A(n11601), .B(P2_EBX_REG_25__SCAN_IN), .S(n10112), .Z(
        n11603) );
  NOR2_X2 U12875 ( .A1(n11571), .A2(n11546), .ZN(n10116) );
  NAND2_X1 U12876 ( .A1(n11513), .A2(n10117), .ZN(n11532) );
  NAND2_X1 U12877 ( .A1(n11604), .A2(n9798), .ZN(n11014) );
  NAND2_X1 U12878 ( .A1(n11604), .A2(n16437), .ZN(n16435) );
  NAND2_X1 U12879 ( .A1(n14678), .A2(n10121), .ZN(P1_U2810) );
  NAND3_X1 U12880 ( .A1(n11849), .A2(n11850), .A3(n11851), .ZN(n10124) );
  NAND2_X1 U12881 ( .A1(n10128), .A2(n14285), .ZN(n14288) );
  NAND2_X1 U12882 ( .A1(n10128), .A2(n14877), .ZN(n14300) );
  NAND2_X1 U12883 ( .A1(n10128), .A2(n13745), .ZN(n13748) );
  NAND2_X1 U12884 ( .A1(n10128), .A2(n20386), .ZN(n14083) );
  NAND2_X1 U12885 ( .A1(n10128), .A2(n20379), .ZN(n14090) );
  NAND2_X1 U12886 ( .A1(n10128), .A2(n14871), .ZN(n14317) );
  MUX2_X1 U12887 ( .A(n10128), .B(n14322), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13558) );
  MUX2_X1 U12888 ( .A(n10128), .B(n14322), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n14167) );
  MUX2_X1 U12889 ( .A(n10128), .B(n14322), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n14274) );
  MUX2_X1 U12890 ( .A(n10128), .B(n14322), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n14278) );
  MUX2_X1 U12891 ( .A(n10128), .B(n14322), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n14290) );
  MUX2_X1 U12892 ( .A(n10128), .B(n14322), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14305) );
  MUX2_X1 U12893 ( .A(n10128), .B(n14322), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14310) );
  MUX2_X1 U12894 ( .A(n10128), .B(n14322), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14324) );
  NOR3_X4 U12895 ( .A1(n9706), .A2(n10131), .A3(n14682), .ZN(n14685) );
  INV_X1 U12896 ( .A(n14696), .ZN(n10133) );
  NAND2_X1 U12897 ( .A1(n13552), .A2(n10139), .ZN(n12695) );
  XNOR2_X1 U12898 ( .A(n13552), .B(n10139), .ZN(n13653) );
  NAND2_X1 U12899 ( .A1(n12692), .A2(n12691), .ZN(n10139) );
  NAND2_X1 U12900 ( .A1(n16295), .A2(n16293), .ZN(n10140) );
  NAND2_X1 U12901 ( .A1(n10145), .A2(n13704), .ZN(n10141) );
  AOI21_X1 U12902 ( .B1(n13704), .B2(n10146), .A(n9708), .ZN(n10142) );
  INV_X1 U12903 ( .A(n12700), .ZN(n10145) );
  NAND2_X1 U12904 ( .A1(n12700), .A2(n12699), .ZN(n13705) );
  AND3_X2 U12905 ( .A1(n11876), .A2(n13521), .A3(n13499), .ZN(n13088) );
  NAND4_X1 U12906 ( .A1(n11853), .A2(n11837), .A3(n11836), .A4(n10149), .ZN(
        n13296) );
  INV_X1 U12907 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10154) );
  INV_X1 U12908 ( .A(n10156), .ZN(n18184) );
  NOR2_X1 U12909 ( .A1(n18197), .A2(n11118), .ZN(n18186) );
  NAND2_X1 U12910 ( .A1(n10157), .A2(n18171), .ZN(n10160) );
  INV_X1 U12911 ( .A(n18164), .ZN(n10157) );
  NAND3_X1 U12912 ( .A1(n9752), .A2(n11067), .A3(n10164), .ZN(n10161) );
  NAND2_X1 U12913 ( .A1(n17869), .A2(n17852), .ZN(n10176) );
  NAND2_X1 U12914 ( .A1(n10181), .A2(n10183), .ZN(n10180) );
  INV_X1 U12915 ( .A(n13189), .ZN(n10181) );
  NAND2_X1 U12916 ( .A1(n9729), .A2(n10187), .ZN(n10184) );
  NOR2_X1 U12917 ( .A1(n20009), .A2(n11438), .ZN(n10192) );
  OR2_X2 U12918 ( .A1(n11372), .A2(n9675), .ZN(n20009) );
  INV_X1 U12919 ( .A(n10193), .ZN(n11662) );
  NAND2_X1 U12920 ( .A1(n10193), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11661) );
  XNOR2_X1 U12921 ( .A(n11662), .B(n9764), .ZN(n16035) );
  NOR2_X1 U12922 ( .A1(n15630), .A2(n15840), .ZN(n15618) );
  INV_X1 U12923 ( .A(n15630), .ZN(n10194) );
  NOR2_X2 U12924 ( .A1(n15630), .A2(n10195), .ZN(n15572) );
  INV_X1 U12925 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U12926 ( .A1(n15396), .A2(n15409), .ZN(n10215) );
  NAND2_X1 U12927 ( .A1(n15396), .A2(n15410), .ZN(n10216) );
  NAND3_X1 U12928 ( .A1(n10216), .A2(n10215), .A3(n15397), .ZN(n15391) );
  NAND3_X1 U12929 ( .A1(n15396), .A2(n15410), .A3(n14587), .ZN(n10210) );
  NAND2_X1 U12930 ( .A1(n13479), .A2(n10217), .ZN(n13828) );
  INV_X1 U12931 ( .A(n10224), .ZN(n14158) );
  INV_X1 U12932 ( .A(n10225), .ZN(n11817) );
  NAND2_X2 U12933 ( .A1(n10225), .A2(n13875), .ZN(n11880) );
  NOR2_X4 U12934 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U12935 ( .A1(n10228), .A2(n12129), .ZN(n12140) );
  NAND2_X1 U12936 ( .A1(n12402), .A2(n9778), .ZN(n14720) );
  NAND2_X1 U12937 ( .A1(n15406), .A2(n10254), .ZN(n15356) );
  NAND2_X1 U12938 ( .A1(n15406), .A2(n9792), .ZN(n12825) );
  NAND3_X1 U12939 ( .A1(n11660), .A2(n11503), .A3(n11667), .ZN(n11507) );
  INV_X1 U12940 ( .A(n14137), .ZN(n10278) );
  NAND2_X1 U12941 ( .A1(n11658), .A2(n10279), .ZN(n11659) );
  AND2_X2 U12942 ( .A1(n11414), .A2(n11413), .ZN(n11415) );
  NAND2_X2 U12943 ( .A1(n11382), .A2(n11381), .ZN(n11416) );
  INV_X1 U12944 ( .A(n13828), .ZN(n13830) );
  CLKBUF_X1 U12945 ( .A(n14809), .Z(n14887) );
  INV_X1 U12946 ( .A(n13935), .ZN(n13826) );
  NAND2_X1 U12947 ( .A1(n12130), .A2(n12122), .ZN(n15320) );
  NAND2_X1 U12948 ( .A1(n14552), .A2(n14551), .ZN(n14553) );
  NAND2_X1 U12949 ( .A1(n12930), .A2(n12947), .ZN(n12959) );
  NAND2_X1 U12950 ( .A1(n15396), .A2(n14553), .ZN(n15410) );
  CLKBUF_X1 U12951 ( .A(n13613), .Z(n13661) );
  INV_X1 U12952 ( .A(n13613), .ZN(n12138) );
  NAND2_X1 U12953 ( .A1(n15433), .A2(n15367), .ZN(n15415) );
  OAI21_X1 U12954 ( .B1(n10495), .B2(n13054), .A(n10499), .ZN(n10485) );
  OAI22_X1 U12955 ( .A1(n11345), .A2(n13858), .B1(n19823), .B2(n11344), .ZN(
        n11360) );
  AOI21_X1 U12956 ( .B1(n13054), .B2(n10486), .A(n10692), .ZN(n10487) );
  INV_X1 U12957 ( .A(n19895), .ZN(n11374) );
  AOI21_X1 U12959 ( .B1(n14681), .B2(n14680), .A(n14679), .ZN(n14996) );
  AND2_X2 U12960 ( .A1(n16072), .A2(n13923), .ZN(n10444) );
  NAND2_X1 U12961 ( .A1(n10478), .A2(n10486), .ZN(n13034) );
  OR2_X1 U12962 ( .A1(n14694), .A2(n14261), .ZN(n14262) );
  AND2_X1 U12963 ( .A1(n14987), .A2(n14347), .ZN(n10293) );
  NOR2_X1 U12964 ( .A1(n20753), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10294) );
  OR2_X1 U12965 ( .A1(n11619), .A2(n19423), .ZN(n10295) );
  OR2_X1 U12966 ( .A1(n11667), .A2(n10951), .ZN(n10296) );
  INV_X1 U12967 ( .A(n10328), .ZN(n10333) );
  NAND2_X2 U12968 ( .A1(n13874), .A2(n13873), .ZN(n20387) );
  AND2_X1 U12969 ( .A1(n14525), .A2(n14549), .ZN(n10297) );
  OR2_X1 U12970 ( .A1(n13280), .A2(n13279), .ZN(n10298) );
  OR2_X1 U12971 ( .A1(n10461), .A2(n10460), .ZN(n10299) );
  OR2_X1 U12972 ( .A1(n15797), .A2(n15796), .ZN(n10300) );
  AND2_X1 U12973 ( .A1(n16176), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10301) );
  XOR2_X1 U12974 ( .A(n19387), .B(n14127), .Z(n10302) );
  INV_X1 U12975 ( .A(n17964), .ZN(n11277) );
  NAND4_X1 U12976 ( .A1(n10495), .A2(n19603), .A3(n10692), .A4(n10486), .ZN(
        n10480) );
  AND2_X1 U12977 ( .A1(n9669), .A2(n18585), .ZN(n17583) );
  AND3_X1 U12978 ( .A1(n19185), .A2(n19167), .A3(n19177), .ZN(n10303) );
  OR2_X1 U12979 ( .A1(n14198), .A2(n17419), .ZN(n10304) );
  NAND2_X1 U12980 ( .A1(n13830), .A2(n13829), .ZN(n13832) );
  OR2_X1 U12981 ( .A1(n14198), .A2(n14238), .ZN(n10306) );
  INV_X1 U12982 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13532) );
  AND3_X1 U12983 ( .A1(n10680), .A2(n13923), .A3(n20194), .ZN(n10307) );
  AND2_X1 U12984 ( .A1(n11060), .A2(n11059), .ZN(n10308) );
  OR2_X2 U12985 ( .A1(n14900), .A2(n14899), .ZN(n10309) );
  AND2_X1 U12986 ( .A1(n12669), .A2(n12684), .ZN(n10310) );
  INV_X1 U12987 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11133) );
  OR3_X1 U12988 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17938), .ZN(n10311) );
  AND2_X1 U12989 ( .A1(n10415), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10312) );
  OR2_X1 U12990 ( .A1(n17061), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10313) );
  OR3_X2 U12991 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19167), .A3(
        n19026), .ZN(n10314) );
  AND3_X1 U12992 ( .A1(n10423), .A2(n10422), .A3(n10421), .ZN(n10315) );
  INV_X1 U12993 ( .A(n10486), .ZN(n10479) );
  INV_X1 U12994 ( .A(n10697), .ZN(n10692) );
  NOR2_X1 U12995 ( .A1(n11149), .A2(n18109), .ZN(n10317) );
  OR2_X1 U12996 ( .A1(n17904), .A2(n18109), .ZN(n10318) );
  AND3_X1 U12997 ( .A1(n11743), .A2(n11742), .A3(n11741), .ZN(n10319) );
  NAND3_X1 U12998 ( .A1(n11863), .A2(n11862), .A3(n11861), .ZN(n10320) );
  NAND2_X1 U12999 ( .A1(n14437), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10767) );
  OR2_X1 U13000 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n12762), .ZN(
        n12761) );
  NAND2_X1 U13001 ( .A1(n11385), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11386) );
  AND2_X1 U13002 ( .A1(n11990), .A2(n11989), .ZN(n11996) );
  INV_X1 U13003 ( .A(n11656), .ZN(n11500) );
  AOI22_X1 U13004 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10423) );
  OR2_X1 U13005 ( .A1(n12772), .A2(n12778), .ZN(n12774) );
  INV_X1 U13006 ( .A(n12148), .ZN(n12069) );
  NAND2_X1 U13007 ( .A1(n11790), .A2(n13941), .ZN(n11791) );
  NAND2_X1 U13008 ( .A1(n10657), .A2(n10656), .ZN(n10666) );
  INV_X1 U13009 ( .A(n14506), .ZN(n14507) );
  AND4_X1 U13010 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10402) );
  AND2_X1 U13011 ( .A1(n13351), .A2(n11901), .ZN(n13523) );
  INV_X1 U13012 ( .A(n12685), .ZN(n12674) );
  AND2_X1 U13013 ( .A1(n13581), .A2(n13580), .ZN(n16125) );
  NAND2_X1 U13014 ( .A1(n14505), .A2(n14507), .ZN(n14508) );
  OAI22_X1 U13015 ( .A1(n10530), .A2(n10507), .B1(n10647), .B2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13016 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10384) );
  NOR3_X1 U13017 ( .A1(n16750), .A2(n18510), .A3(n16749), .ZN(n16751) );
  NOR2_X1 U13018 ( .A1(n12509), .A2(n15038), .ZN(n12510) );
  INV_X1 U13019 ( .A(n14888), .ZN(n12319) );
  INV_X1 U13020 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12846) );
  OR2_X1 U13021 ( .A1(n12021), .A2(n12020), .ZN(n12702) );
  AND2_X1 U13022 ( .A1(n13958), .A2(n14265), .ZN(n13303) );
  NOR2_X1 U13023 ( .A1(n13845), .A2(n13846), .ZN(n13829) );
  INV_X1 U13024 ( .A(n10860), .ZN(n10736) );
  AND2_X1 U13025 ( .A1(n10595), .A2(n10594), .ZN(n13848) );
  NAND2_X1 U13026 ( .A1(n11666), .A2(n11665), .ZN(n11670) );
  AND2_X1 U13027 ( .A1(n11690), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11687) );
  NOR2_X1 U13028 ( .A1(n17711), .A2(n18545), .ZN(n11256) );
  INV_X1 U13029 ( .A(n17450), .ZN(n17420) );
  NAND2_X1 U13030 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11112) );
  NAND2_X1 U13031 ( .A1(n9883), .A2(n11319), .ZN(n11147) );
  NAND2_X1 U13032 ( .A1(n9883), .A2(n18334), .ZN(n11138) );
  NOR2_X1 U13033 ( .A1(n11306), .A2(n18140), .ZN(n11309) );
  NAND2_X1 U13034 ( .A1(n11120), .A2(n17729), .ZN(n11123) );
  INV_X1 U13035 ( .A(n11936), .ZN(n11937) );
  NAND2_X1 U13036 ( .A1(n14322), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n13533) );
  INV_X1 U13037 ( .A(n13646), .ZN(n12120) );
  OR2_X1 U13038 ( .A1(n12855), .A2(n12854), .ZN(n12857) );
  NAND2_X1 U13039 ( .A1(n12599), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12855) );
  AND2_X1 U13040 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n12459), .ZN(
        n12460) );
  INV_X1 U13041 ( .A(n13837), .ZN(n12146) );
  INV_X1 U13042 ( .A(n15010), .ZN(n12756) );
  INV_X1 U13043 ( .A(n12805), .ZN(n13086) );
  AND2_X1 U13044 ( .A1(n12962), .A2(n12961), .ZN(n10970) );
  INV_X1 U13045 ( .A(n13483), .ZN(n13480) );
  INV_X1 U13046 ( .A(n10652), .ZN(n10646) );
  AND2_X1 U13047 ( .A1(n10574), .A2(n10573), .ZN(n13546) );
  INV_X1 U13048 ( .A(n16569), .ZN(n11669) );
  INV_X1 U13049 ( .A(n11001), .ZN(n11640) );
  AOI21_X1 U13050 ( .B1(n19012), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11168), .ZN(n11177) );
  NAND3_X1 U13051 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n19185), .ZN(n11026) );
  NAND2_X1 U13052 ( .A1(n18110), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18077) );
  NOR2_X1 U13053 ( .A1(n9883), .A2(n16115), .ZN(n11154) );
  OAI21_X1 U13054 ( .B1(n11129), .B2(n16746), .A(n18109), .ZN(n11130) );
  NOR2_X1 U13055 ( .A1(n11295), .A2(n18174), .ZN(n11297) );
  NAND2_X1 U13056 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n20366), .ZN(n13805) );
  AND4_X1 U13057 ( .A1(n11808), .A2(n11807), .A3(n11806), .A4(n11805), .ZN(
        n11814) );
  INV_X1 U13058 ( .A(n12863), .ZN(n12864) );
  NAND2_X1 U13059 ( .A1(n16285), .A2(n14671), .ZN(n12816) );
  NAND2_X1 U13060 ( .A1(n12460), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12509) );
  OR2_X1 U13061 ( .A1(n14107), .A2(n12205), .ZN(n14852) );
  NOR2_X1 U13062 ( .A1(n12150), .A2(n20309), .ZN(n12167) );
  INV_X1 U13063 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13707) );
  INV_X1 U13064 ( .A(n15145), .ZN(n15261) );
  INV_X1 U13065 ( .A(n20842), .ZN(n20750) );
  OR2_X1 U13066 ( .A1(n20582), .A2(n20581), .ZN(n21024) );
  OR2_X1 U13067 ( .A1(n21020), .A2(n20728), .ZN(n20751) );
  AOI21_X1 U13068 ( .B1(n21044), .B2(n16421), .A(n15312), .ZN(n13940) );
  OR2_X1 U13069 ( .A1(n21021), .A2(n15322), .ZN(n20457) );
  OR2_X1 U13070 ( .A1(n21021), .A2(n20518), .ZN(n20728) );
  INV_X1 U13071 ( .A(n13308), .ZN(n13941) );
  OR3_X1 U13072 ( .A1(n20760), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13940), 
        .ZN(n15339) );
  INV_X1 U13073 ( .A(n19423), .ZN(n12839) );
  NOR2_X1 U13074 ( .A1(n19393), .A2(n16443), .ZN(n16425) );
  NOR2_X1 U13075 ( .A1(n19393), .A2(n15365), .ZN(n16451) );
  OAI211_X1 U13076 ( .C1(n11328), .C2(n13195), .A(n13194), .B(n13193), .ZN(
        n13281) );
  OR2_X1 U13077 ( .A1(n19239), .A2(n16700), .ZN(n16584) );
  AND2_X1 U13078 ( .A1(n11592), .A2(n15882), .ZN(n15871) );
  AND2_X1 U13079 ( .A1(n11566), .A2(n16510), .ZN(n16504) );
  AND2_X1 U13080 ( .A1(n15737), .A2(n15736), .ZN(n16608) );
  INV_X1 U13081 ( .A(n19974), .ZN(n13723) );
  NAND2_X1 U13082 ( .A1(n20210), .A2(n20224), .ZN(n20197) );
  OR2_X1 U13083 ( .A1(n20210), .A2(n20224), .ZN(n19974) );
  INV_X1 U13084 ( .A(n16862), .ZN(n18986) );
  INV_X1 U13085 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17126) );
  NOR3_X1 U13086 ( .A1(n18567), .A2(n18585), .A3(n14173), .ZN(n14174) );
  INV_X1 U13087 ( .A(n9648), .ZN(n17522) );
  INV_X1 U13088 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17478) );
  AOI211_X1 U13089 ( .C1(n9641), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n11032), .B(n11031), .ZN(n11033) );
  NOR3_X1 U13090 ( .A1(n18578), .A2(n18567), .A3(n11252), .ZN(n17785) );
  NOR2_X1 U13091 ( .A1(n16990), .A2(n16886), .ZN(n17895) );
  NOR2_X1 U13092 ( .A1(n10002), .A2(n17017), .ZN(n16887) );
  INV_X1 U13093 ( .A(n17970), .ZN(n18063) );
  NAND2_X1 U13094 ( .A1(n17902), .A2(n18215), .ZN(n18218) );
  NOR2_X1 U13095 ( .A1(n18314), .A2(n18238), .ZN(n18293) );
  INV_X1 U13096 ( .A(n18272), .ZN(n18401) );
  NOR2_X1 U13097 ( .A1(n18118), .A2(n18442), .ZN(n18117) );
  NOR2_X1 U13098 ( .A1(n18141), .A2(n18457), .ZN(n18140) );
  NOR2_X1 U13099 ( .A1(n18480), .A2(n18160), .ZN(n18159) );
  XNOR2_X1 U13100 ( .A(n11119), .B(n18508), .ZN(n18185) );
  AOI211_X1 U13101 ( .C1(n9641), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n11218), .B(n11217), .ZN(n11219) );
  INV_X1 U13102 ( .A(n12141), .ZN(n12151) );
  NAND2_X1 U13103 ( .A1(n13435), .A2(n13511), .ZN(n13437) );
  INV_X1 U13104 ( .A(n13252), .ZN(n20426) );
  NAND2_X1 U13105 ( .A1(n12398), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12458) );
  NAND2_X1 U13106 ( .A1(n12340), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12397) );
  INV_X1 U13107 ( .A(n15129), .ZN(n20377) );
  INV_X1 U13108 ( .A(n16260), .ZN(n16291) );
  INV_X1 U13109 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12852) );
  NOR2_X1 U13110 ( .A1(n16374), .A2(n13562), .ZN(n16370) );
  INV_X1 U13111 ( .A(n16371), .ZN(n15147) );
  INV_X1 U13112 ( .A(n20453), .ZN(n16353) );
  AND2_X1 U13113 ( .A1(n15132), .A2(n16370), .ZN(n15281) );
  AND2_X1 U13114 ( .A1(n15320), .A2(n20582), .ZN(n20552) );
  AND2_X1 U13115 ( .A1(n20552), .A2(n20497), .ZN(n20541) );
  INV_X1 U13116 ( .A(n20558), .ZN(n20577) );
  NOR2_X2 U13117 ( .A1(n20560), .A2(n20559), .ZN(n20605) );
  NOR2_X2 U13118 ( .A1(n21024), .A2(n20728), .ZN(n20656) );
  NOR2_X2 U13119 ( .A1(n21024), .A2(n20750), .ZN(n20686) );
  INV_X1 U13120 ( .A(n21024), .ZN(n20665) );
  INV_X1 U13121 ( .A(n20457), .ZN(n20690) );
  INV_X1 U13122 ( .A(n20764), .ZN(n20790) );
  INV_X1 U13123 ( .A(n20756), .ZN(n20819) );
  NOR2_X1 U13124 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13940), .ZN(n20464) );
  NAND2_X1 U13125 ( .A1(n21021), .A2(n15322), .ZN(n20559) );
  INV_X1 U13126 ( .A(n20471), .ZN(n20896) );
  INV_X1 U13127 ( .A(n20931), .ZN(n20938) );
  AND2_X1 U13128 ( .A1(n11690), .A2(n10671), .ZN(n16672) );
  AND2_X1 U13129 ( .A1(n16672), .A2(n16664), .ZN(n16654) );
  NOR2_X1 U13130 ( .A1(n19393), .A2(n12926), .ZN(n12942) );
  AND2_X1 U13131 ( .A1(n19545), .A2(n10994), .ZN(n19420) );
  INV_X1 U13132 ( .A(n19416), .ZN(n19402) );
  INV_X1 U13133 ( .A(n19490), .ZN(n19497) );
  INV_X1 U13134 ( .A(n13020), .ZN(n13113) );
  NAND2_X1 U13135 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  INV_X1 U13136 ( .A(n10338), .ZN(n10341) );
  AND2_X1 U13137 ( .A1(n13549), .A2(n13548), .ZN(n19360) );
  INV_X1 U13138 ( .A(n16584), .ZN(n19554) );
  AND2_X1 U13139 ( .A1(n16531), .A2(n16530), .ZN(n16615) );
  NOR2_X1 U13140 ( .A1(n16638), .A2(n16636), .ZN(n16597) );
  INV_X1 U13141 ( .A(n16624), .ZN(n16643) );
  INV_X1 U13142 ( .A(n20053), .ZN(n19764) );
  NAND2_X1 U13143 ( .A1(n13183), .A2(n13177), .ZN(n20224) );
  AND2_X1 U13144 ( .A1(n16668), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20190) );
  OAI21_X1 U13145 ( .B1(n19573), .B2(n19572), .A(n19571), .ZN(n19617) );
  AND2_X1 U13146 ( .A1(n20210), .A2(n20222), .ZN(n19819) );
  INV_X1 U13147 ( .A(n20197), .ZN(n19674) );
  AND2_X1 U13148 ( .A1(n19788), .A2(n19674), .ZN(n19733) );
  AND2_X1 U13149 ( .A1(n19756), .A2(n13723), .ZN(n19751) );
  OR3_X1 U13150 ( .A1(n19766), .A2(n19765), .A3(n19764), .ZN(n19784) );
  INV_X1 U13151 ( .A(n19813), .ZN(n19815) );
  OAI21_X1 U13152 ( .B1(n19847), .B2(n19826), .A(n20053), .ZN(n19850) );
  INV_X1 U13153 ( .A(n19819), .ZN(n19855) );
  AND2_X1 U13154 ( .A1(n19924), .A2(n19922), .ZN(n19944) );
  INV_X1 U13155 ( .A(n20070), .ZN(n19982) );
  OAI21_X1 U13156 ( .B1(n20012), .B2(n20011), .A(n20010), .ZN(n20036) );
  AND2_X1 U13157 ( .A1(n10468), .A2(n19613), .ZN(n20046) );
  INV_X1 U13158 ( .A(n20095), .ZN(n20102) );
  NAND2_X1 U13159 ( .A1(n19045), .A2(n16883), .ZN(n17245) );
  INV_X1 U13160 ( .A(n17245), .ZN(n17237) );
  INV_X1 U13161 ( .A(n17646), .ZN(n17642) );
  NAND2_X1 U13162 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17656), .ZN(n17655) );
  NOR2_X1 U13163 ( .A1(n17837), .A2(n17699), .ZN(n17694) );
  NOR2_X1 U13164 ( .A1(n19006), .A2(n17728), .ZN(n17741) );
  INV_X1 U13165 ( .A(n18010), .ZN(n18021) );
  NAND2_X1 U13166 ( .A1(n18039), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18273) );
  NOR2_X1 U13167 ( .A1(n11314), .A2(n18117), .ZN(n18404) );
  NOR2_X1 U13168 ( .A1(n11319), .A2(n17894), .ZN(n18220) );
  NOR2_X1 U13169 ( .A1(n18273), .A2(n12884), .ZN(n17902) );
  NOR2_X1 U13170 ( .A1(n18987), .A2(n17713), .ZN(n18354) );
  XNOR2_X1 U13171 ( .A(n11284), .B(n19173), .ZN(n18198) );
  NOR2_X2 U13172 ( .A1(n18483), .A2(n18521), .ZN(n18520) );
  INV_X1 U13173 ( .A(n20362), .ZN(n20320) );
  NAND2_X1 U13174 ( .A1(n14099), .A2(n13670), .ZN(n14864) );
  INV_X1 U13175 ( .A(n20349), .ZN(n20375) );
  NAND2_X1 U13176 ( .A1(n20387), .A2(n13875), .ZN(n14914) );
  OAI21_X1 U13177 ( .B1(n14837), .B2(n14825), .A(n14824), .ZN(n16279) );
  NAND2_X1 U13178 ( .A1(n13437), .A2(n13436), .ZN(n14987) );
  NOR2_X1 U13179 ( .A1(n13248), .A2(n13247), .ZN(n13251) );
  INV_X1 U13180 ( .A(n12859), .ZN(n12867) );
  NAND2_X1 U13181 ( .A1(n20282), .A2(n12811), .ZN(n16260) );
  INV_X1 U13182 ( .A(n16285), .ZN(n16299) );
  INV_X1 U13183 ( .A(n16286), .ZN(n16263) );
  INV_X1 U13184 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20721) );
  NAND2_X1 U13185 ( .A1(n20552), .A2(n20690), .ZN(n20517) );
  AOI22_X1 U13186 ( .A1(n20520), .A2(n20524), .B1(n10294), .B2(n20755), .ZN(
        n20545) );
  NAND2_X1 U13187 ( .A1(n20665), .A2(n20690), .ZN(n20632) );
  NAND2_X1 U13188 ( .A1(n20665), .A2(n20661), .ZN(n20696) );
  NAND2_X1 U13189 ( .A1(n20691), .A2(n20690), .ZN(n20749) );
  INV_X1 U13190 ( .A(n20936), .ZN(n20793) );
  OR2_X1 U13191 ( .A1(n21020), .A2(n20559), .ZN(n20841) );
  NAND2_X1 U13192 ( .A1(n20884), .A2(n20661), .ZN(n20931) );
  INV_X1 U13193 ( .A(n21019), .ZN(n21015) );
  AND2_X1 U13194 ( .A1(n16654), .A2(n13332), .ZN(n20253) );
  INV_X1 U13195 ( .A(n12822), .ZN(n12843) );
  INV_X1 U13196 ( .A(n19406), .ZN(n19418) );
  INV_X1 U13197 ( .A(n19425), .ZN(n19389) );
  INV_X1 U13198 ( .A(n19420), .ZN(n19408) );
  AND2_X1 U13199 ( .A1(n13061), .A2(n13332), .ZN(n15449) );
  INV_X1 U13200 ( .A(n20224), .ZN(n20222) );
  AND2_X2 U13201 ( .A1(n13333), .A2(n13332), .ZN(n19466) );
  NAND2_X1 U13202 ( .A1(n19466), .A2(n13334), .ZN(n19490) );
  NAND2_X1 U13203 ( .A1(n13226), .A2(n20262), .ZN(n19542) );
  INV_X1 U13204 ( .A(n19545), .ZN(n13223) );
  INV_X1 U13205 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16592) );
  INV_X1 U13206 ( .A(n16583), .ZN(n19564) );
  AOI21_X1 U13207 ( .B1(n15801), .B2(n16646), .A(n15800), .ZN(n15802) );
  INV_X1 U13208 ( .A(n16646), .ZN(n16630) );
  INV_X1 U13209 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20194) );
  NAND2_X1 U13210 ( .A1(n19819), .A2(n19756), .ZN(n19636) );
  NAND2_X1 U13211 ( .A1(n19756), .A2(n19674), .ZN(n19698) );
  INV_X1 U13212 ( .A(n19733), .ZN(n19707) );
  INV_X1 U13213 ( .A(n19751), .ZN(n19748) );
  INV_X1 U13214 ( .A(n19771), .ZN(n19787) );
  NAND2_X1 U13215 ( .A1(n19795), .A2(n19756), .ZN(n19813) );
  NAND2_X1 U13216 ( .A1(n19788), .A2(n19795), .ZN(n19844) );
  OR2_X1 U13217 ( .A1(n19970), .A2(n19855), .ZN(n19891) );
  INV_X1 U13218 ( .A(n19939), .ZN(n19948) );
  AOI21_X1 U13219 ( .B1(n13860), .B2(n13861), .A(n13859), .ZN(n19969) );
  INV_X1 U13220 ( .A(n20085), .ZN(n19993) );
  INV_X1 U13221 ( .A(n20073), .ZN(n20024) );
  OR2_X1 U13222 ( .A1(n20003), .A2(n20049), .ZN(n20095) );
  INV_X1 U13223 ( .A(n17242), .ZN(n17205) );
  INV_X1 U13224 ( .A(n11302), .ZN(n17717) );
  INV_X1 U13225 ( .A(n17763), .ZN(n17782) );
  NAND2_X1 U13226 ( .A1(n12883), .A2(n18104), .ZN(n11325) );
  NAND2_X1 U13227 ( .A1(n18315), .A2(n18093), .ZN(n18010) );
  INV_X1 U13228 ( .A(n18104), .ZN(n18122) );
  INV_X1 U13230 ( .A(n18520), .ZN(n18511) );
  INV_X1 U13231 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19012) );
  INV_X1 U13232 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18560) );
  INV_X1 U13233 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18582) );
  INV_X1 U13234 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19160) );
  OAI21_X1 U13235 ( .B1(n14921), .B2(n16263), .A(n12820), .ZN(P1_U2969) );
  NAND2_X1 U13236 ( .A1(n11325), .A2(n11324), .ZN(P3_U2799) );
  INV_X1 U13237 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16564) );
  INV_X1 U13238 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16544) );
  NAND2_X1 U13239 ( .A1(n10347), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10346) );
  INV_X1 U13240 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10321) );
  INV_X1 U13241 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16502) );
  OR2_X1 U13242 ( .A1(n10321), .A2(n16502), .ZN(n10322) );
  INV_X1 U13243 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15705) );
  INV_X1 U13244 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15666) );
  INV_X1 U13245 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15629) );
  INV_X1 U13246 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15606) );
  INV_X1 U13247 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10329) );
  INV_X1 U13248 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15586) );
  INV_X1 U13249 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10323) );
  XNOR2_X1 U13250 ( .A(n10324), .B(n10323), .ZN(n15573) );
  NAND2_X1 U13251 ( .A1(n10324), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10326) );
  INV_X1 U13252 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10325) );
  INV_X1 U13253 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10651) );
  AND2_X1 U13254 ( .A1(n10331), .A2(n15586), .ZN(n10327) );
  NOR2_X1 U13255 ( .A1(n10324), .A2(n10327), .ZN(n15588) );
  NAND2_X1 U13256 ( .A1(n10333), .A2(n10329), .ZN(n10330) );
  NAND2_X1 U13257 ( .A1(n10331), .A2(n10330), .ZN(n15600) );
  INV_X1 U13258 ( .A(n15600), .ZN(n16426) );
  AOI21_X1 U13259 ( .B1(n15606), .B2(n10332), .A(n10328), .ZN(n16445) );
  OR2_X1 U13260 ( .A1(n9785), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10334) );
  NAND2_X1 U13261 ( .A1(n10332), .A2(n10334), .ZN(n15617) );
  INV_X1 U13262 ( .A(n15617), .ZN(n16452) );
  AOI21_X1 U13263 ( .B1(n15629), .B2(n10335), .A(n9785), .ZN(n15627) );
  OAI21_X1 U13264 ( .B1(n10336), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n10335), .ZN(n10337) );
  INV_X1 U13265 ( .A(n10337), .ZN(n16473) );
  NOR2_X1 U13266 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n10338), .ZN(
        n10339) );
  NOR2_X1 U13267 ( .A1(n10336), .A2(n10339), .ZN(n15647) );
  OAI21_X1 U13268 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10340), .A(
        n10341), .ZN(n16496) );
  INV_X1 U13269 ( .A(n16496), .ZN(n12943) );
  AOI21_X1 U13270 ( .B1(n15666), .B2(n10342), .A(n10340), .ZN(n15664) );
  OAI21_X1 U13271 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10343), .A(
        n10342), .ZN(n15676) );
  INV_X1 U13272 ( .A(n15676), .ZN(n19262) );
  NOR2_X1 U13273 ( .A1(n10344), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10345) );
  NOR2_X1 U13274 ( .A1(n10343), .A2(n10345), .ZN(n19270) );
  AOI21_X1 U13275 ( .B1(n15705), .B2(n10358), .A(n10361), .ZN(n19291) );
  NOR2_X1 U13276 ( .A1(n16502), .A2(n10346), .ZN(n10359) );
  AOI21_X1 U13277 ( .B1(n16502), .B2(n10346), .A(n10359), .ZN(n19313) );
  INV_X1 U13278 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16520) );
  NAND2_X1 U13279 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n9779), .ZN(
        n10357) );
  AOI21_X1 U13280 ( .B1(n16520), .B2(n10357), .A(n10347), .ZN(n19327) );
  AOI21_X1 U13281 ( .B1(n16544), .B2(n10348), .A(n9779), .ZN(n19339) );
  AOI21_X1 U13282 ( .B1(n16564), .B2(n10349), .A(n10350), .ZN(n19359) );
  AOI21_X1 U13283 ( .B1(n15725), .B2(n10351), .A(n10352), .ZN(n15726) );
  AOI21_X1 U13284 ( .B1(n16592), .B2(n10353), .A(n9712), .ZN(n19381) );
  AOI21_X1 U13285 ( .B1(n13983), .B2(n10355), .A(n10356), .ZN(n13985) );
  OAI22_X1 U13286 ( .A1(n20256), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n10354) );
  INV_X1 U13287 ( .A(n10354), .ZN(n19426) );
  AOI22_X1 U13288 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13155), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20256), .ZN(n16069) );
  NOR2_X1 U13289 ( .A1(n19426), .A2(n16069), .ZN(n16068) );
  OAI21_X1 U13290 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n10355), .ZN(n14644) );
  NAND2_X1 U13291 ( .A1(n16068), .A2(n14644), .ZN(n13629) );
  NOR2_X1 U13292 ( .A1(n13985), .A2(n13629), .ZN(n19392) );
  OAI21_X1 U13293 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10356), .A(
        n10353), .ZN(n19563) );
  NAND2_X1 U13294 ( .A1(n19392), .A2(n19563), .ZN(n19378) );
  NOR2_X1 U13295 ( .A1(n19381), .A2(n19378), .ZN(n19368) );
  OAI21_X1 U13296 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9712), .A(
        n10351), .ZN(n19369) );
  NAND2_X1 U13297 ( .A1(n19368), .A2(n19369), .ZN(n13617) );
  NOR2_X1 U13298 ( .A1(n15726), .A2(n13617), .ZN(n13906) );
  OAI21_X1 U13299 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10352), .A(
        n10349), .ZN(n16576) );
  NAND2_X1 U13300 ( .A1(n13906), .A2(n16576), .ZN(n19357) );
  NOR2_X1 U13301 ( .A1(n19359), .A2(n19357), .ZN(n19347) );
  OAI21_X1 U13302 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10350), .A(
        n10348), .ZN(n19348) );
  NAND2_X1 U13303 ( .A1(n19347), .A2(n19348), .ZN(n19337) );
  NOR2_X1 U13304 ( .A1(n19339), .A2(n19337), .ZN(n13883) );
  OAI21_X1 U13305 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9779), .A(
        n10357), .ZN(n16538) );
  NAND2_X1 U13306 ( .A1(n13883), .A2(n16538), .ZN(n19320) );
  NOR2_X1 U13307 ( .A1(n19327), .A2(n19320), .ZN(n19319) );
  OAI21_X1 U13308 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10347), .A(
        n10346), .ZN(n16513) );
  NAND2_X1 U13309 ( .A1(n19319), .A2(n16513), .ZN(n19311) );
  NOR2_X1 U13310 ( .A1(n19313), .A2(n19311), .ZN(n19298) );
  OAI21_X1 U13311 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10359), .A(
        n10358), .ZN(n19300) );
  NAND2_X1 U13312 ( .A1(n19298), .A2(n19300), .ZN(n19290) );
  NOR2_X1 U13313 ( .A1(n19291), .A2(n19290), .ZN(n19289) );
  INV_X1 U13314 ( .A(n10344), .ZN(n10360) );
  OAI21_X1 U13315 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n10361), .A(
        n10360), .ZN(n15697) );
  NOR2_X1 U13316 ( .A1(n19262), .A2(n19261), .ZN(n19260) );
  NOR2_X1 U13317 ( .A1(n19393), .A2(n19260), .ZN(n12927) );
  NOR2_X1 U13318 ( .A1(n15664), .A2(n12927), .ZN(n12926) );
  NOR2_X1 U13319 ( .A1(n12943), .A2(n12942), .ZN(n12941) );
  NOR2_X1 U13320 ( .A1(n19393), .A2(n12941), .ZN(n12955) );
  NOR2_X1 U13321 ( .A1(n15647), .A2(n12955), .ZN(n12954) );
  NOR2_X1 U13322 ( .A1(n16452), .A2(n16451), .ZN(n16450) );
  NOR2_X1 U13323 ( .A1(n19393), .A2(n16450), .ZN(n16444) );
  NOR2_X1 U13324 ( .A1(n16445), .A2(n16444), .ZN(n16443) );
  NOR2_X1 U13325 ( .A1(n16426), .A2(n16425), .ZN(n16424) );
  NOR2_X1 U13326 ( .A1(n19393), .A2(n16424), .ZN(n15363) );
  NOR2_X1 U13327 ( .A1(n19393), .A2(n15362), .ZN(n12821) );
  NOR2_X1 U13328 ( .A1(n15573), .A2(n12821), .ZN(n12844) );
  NOR4_X1 U13329 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n10598), .ZN(n10363) );
  INV_X1 U13330 ( .A(n19411), .ZN(n19394) );
  NOR2_X1 U13331 ( .A1(n19393), .A2(n19394), .ZN(n19427) );
  NAND2_X1 U13332 ( .A1(n12844), .A2(n19427), .ZN(n11016) );
  INV_X1 U13333 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10364) );
  AND2_X2 U13334 ( .A1(n10364), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10366) );
  NOR2_X2 U13335 ( .A1(n10364), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10365) );
  INV_X2 U13336 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16653) );
  AND2_X4 U13337 ( .A1(n10365), .A2(n16653), .ZN(n14595) );
  AOI22_X1 U13338 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10370) );
  AND2_X4 U13339 ( .A1(n16072), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14594) );
  AOI22_X1 U13340 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10369) );
  AND2_X4 U13341 ( .A1(n13380), .A2(n16653), .ZN(n14600) );
  AOI22_X1 U13342 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13343 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10367) );
  NAND4_X1 U13344 ( .A1(n10370), .A2(n10369), .A3(n10368), .A4(n10367), .ZN(
        n10376) );
  AOI22_X1 U13345 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13346 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13347 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13348 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10371) );
  NAND4_X1 U13349 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10375) );
  INV_X2 U13350 ( .A(n10477), .ZN(n10495) );
  AOI22_X1 U13351 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13352 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13353 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13354 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10377) );
  NAND4_X1 U13355 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10386) );
  AOI22_X1 U13356 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13357 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13358 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10381) );
  NAND4_X1 U13359 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10385) );
  AOI22_X1 U13360 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14577), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13361 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13362 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13363 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10387) );
  NAND4_X1 U13364 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10396) );
  AOI22_X1 U13365 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13366 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13367 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U13368 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10391) );
  NAND4_X1 U13369 ( .A1(n10394), .A2(n10393), .A3(n10392), .A4(n10391), .ZN(
        n10395) );
  AOI22_X1 U13370 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14577), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U13371 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U13372 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13373 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U13374 ( .A1(n10402), .A2(n10680), .ZN(n10409) );
  AOI22_X1 U13375 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14577), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13376 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13377 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U13378 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10403) );
  NAND4_X1 U13379 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        n10408) );
  AOI22_X1 U13380 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13381 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13382 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13383 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10412) );
  NAND3_X1 U13384 ( .A1(n10414), .A2(n10413), .A3(n10412), .ZN(n10420) );
  AOI22_X1 U13385 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U13386 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13387 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13388 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10416) );
  NAND4_X1 U13389 ( .A1(n10418), .A2(n10417), .A3(n10312), .A4(n10416), .ZN(
        n10419) );
  AOI22_X1 U13390 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U13391 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U13392 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U13393 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13394 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13395 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13396 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13397 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13398 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13399 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13400 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10432) );
  NAND4_X1 U13401 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        n10436) );
  NAND2_X1 U13402 ( .A1(n10436), .A2(n10680), .ZN(n10443) );
  AOI22_X1 U13403 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13404 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13405 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13406 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10437) );
  NAND4_X1 U13407 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10441) );
  NAND2_X1 U13408 ( .A1(n10441), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10442) );
  AOI22_X1 U13409 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13410 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13411 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9674), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13412 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10445) );
  NAND4_X1 U13413 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10454) );
  AOI22_X1 U13414 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13415 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13416 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9673), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U13417 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10449) );
  NAND4_X1 U13418 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10453) );
  MUX2_X2 U13419 ( .A(n10454), .B(n10453), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10468) );
  NAND2_X1 U13420 ( .A1(n13329), .A2(n11676), .ZN(n13059) );
  INV_X1 U13421 ( .A(n13059), .ZN(n10455) );
  NAND2_X2 U13422 ( .A1(n10455), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10533) );
  INV_X1 U13423 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10456) );
  INV_X1 U13424 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13076) );
  OAI22_X1 U13425 ( .A1(n10533), .A2(n10456), .B1(n10598), .B2(n13076), .ZN(
        n10461) );
  NAND2_X1 U13426 ( .A1(n10495), .A2(n10697), .ZN(n10690) );
  INV_X1 U13427 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U13428 ( .A1(n13116), .A2(n10481), .A3(n10486), .A4(n10477), .ZN(
        n10462) );
  NAND2_X1 U13429 ( .A1(n10697), .A2(n10476), .ZN(n10496) );
  NOR2_X2 U13430 ( .A1(n10462), .A2(n10496), .ZN(n10484) );
  INV_X1 U13431 ( .A(n10472), .ZN(n10463) );
  INV_X1 U13432 ( .A(n10496), .ZN(n13336) );
  NAND4_X1 U13433 ( .A1(n10463), .A2(n16659), .A3(n10495), .A4(n13336), .ZN(
        n10464) );
  NAND2_X1 U13434 ( .A1(n10673), .A2(n10464), .ZN(n10466) );
  INV_X1 U13435 ( .A(n10466), .ZN(n10465) );
  NAND2_X1 U13436 ( .A1(n10465), .A2(n10672), .ZN(n10502) );
  OAI21_X1 U13437 ( .B1(n10493), .B2(n10466), .A(n10502), .ZN(n10473) );
  OR2_X1 U13438 ( .A1(n10691), .A2(n10468), .ZN(n10467) );
  INV_X1 U13439 ( .A(n10692), .ZN(n19614) );
  NAND3_X1 U13440 ( .A1(n12972), .A2(n19614), .A3(n10479), .ZN(n10471) );
  NAND2_X2 U13441 ( .A1(n13054), .A2(n10477), .ZN(n10492) );
  NAND3_X1 U13442 ( .A1(n13054), .A2(n16663), .A3(n10495), .ZN(n10469) );
  MUX2_X2 U13443 ( .A(n10492), .B(n10469), .S(n10481), .Z(n10470) );
  NAND2_X1 U13444 ( .A1(n10473), .A2(n10508), .ZN(n10474) );
  NOR2_X1 U13445 ( .A1(n10532), .A2(n13155), .ZN(n10475) );
  NOR2_X1 U13446 ( .A1(n10299), .A2(n10475), .ZN(n10525) );
  NAND2_X1 U13447 ( .A1(n10492), .A2(n10479), .ZN(n13027) );
  NAND3_X1 U13448 ( .A1(n13034), .A2(n13027), .A3(n19614), .ZN(n13138) );
  NAND2_X1 U13449 ( .A1(n13138), .A2(n10457), .ZN(n10483) );
  NAND2_X1 U13450 ( .A1(n10483), .A2(n10482), .ZN(n10516) );
  INV_X1 U13451 ( .A(n10484), .ZN(n10491) );
  INV_X1 U13452 ( .A(n10485), .ZN(n10489) );
  NAND2_X1 U13453 ( .A1(n10492), .A2(n10457), .ZN(n10488) );
  NAND3_X1 U13454 ( .A1(n10489), .A2(n10488), .A3(n10487), .ZN(n10490) );
  NAND3_X1 U13455 ( .A1(n10491), .A2(n10490), .A3(n16663), .ZN(n13143) );
  NAND2_X1 U13456 ( .A1(n10493), .A2(n10492), .ZN(n10517) );
  NAND2_X1 U13457 ( .A1(n10517), .A2(n16663), .ZN(n10494) );
  NOR2_X1 U13458 ( .A1(n10496), .A2(n10495), .ZN(n10497) );
  NAND2_X1 U13459 ( .A1(n10501), .A2(n10500), .ZN(n13024) );
  NAND2_X1 U13460 ( .A1(n10468), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20263) );
  NAND2_X1 U13461 ( .A1(n10530), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10506) );
  NAND2_X1 U13463 ( .A1(n10598), .A2(n20256), .ZN(n20252) );
  NOR2_X1 U13464 ( .A1(n20252), .A2(n20229), .ZN(n10504) );
  AOI21_X1 U13465 ( .B1(n10503), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10504), 
        .ZN(n10505) );
  NAND2_X1 U13466 ( .A1(n10506), .A2(n10505), .ZN(n10524) );
  XNOR2_X1 U13467 ( .A(n10525), .B(n10524), .ZN(n11333) );
  AND3_X1 U13468 ( .A1(n10463), .A2(n11676), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10507) );
  INV_X4 U13469 ( .A(n10533), .ZN(n10647) );
  OAI22_X1 U13470 ( .A1(n10508), .A2(n20256), .B1(n20252), .B2(n20239), .ZN(
        n10509) );
  INV_X1 U13471 ( .A(n10509), .ZN(n10510) );
  NAND2_X1 U13472 ( .A1(n10511), .A2(n10510), .ZN(n11330) );
  AOI22_X1 U13473 ( .A1(n10647), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n10648), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n10523) );
  NAND2_X1 U13474 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10513) );
  AND3_X1 U13475 ( .A1(n10514), .A2(n20252), .A3(n10513), .ZN(n10522) );
  INV_X1 U13476 ( .A(n10532), .ZN(n10515) );
  NAND2_X1 U13477 ( .A1(n10515), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10521) );
  NAND2_X1 U13478 ( .A1(n10516), .A2(n10517), .ZN(n13137) );
  NAND2_X1 U13479 ( .A1(n13137), .A2(n10518), .ZN(n10519) );
  NAND2_X1 U13480 ( .A1(n10519), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10520) );
  NAND4_X1 U13481 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n11331) );
  NAND2_X1 U13482 ( .A1(n11330), .A2(n11331), .ZN(n11334) );
  NAND2_X1 U13483 ( .A1(n11333), .A2(n11334), .ZN(n10529) );
  INV_X1 U13484 ( .A(n10524), .ZN(n10527) );
  NAND2_X1 U13485 ( .A1(n10527), .A2(n10526), .ZN(n10528) );
  OAI21_X1 U13486 ( .B1(n20219), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10598), 
        .ZN(n10531) );
  INV_X1 U13487 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13198) );
  INV_X1 U13488 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n10598) );
  INV_X1 U13489 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10534) );
  OAI22_X1 U13490 ( .A1(n10606), .A2(n13198), .B1(n10598), .B2(n10534), .ZN(
        n10537) );
  INV_X1 U13491 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10535) );
  NOR2_X1 U13492 ( .A1(n10537), .A2(n10536), .ZN(n10538) );
  INV_X1 U13493 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13635) );
  OAI22_X1 U13494 ( .A1(n10606), .A2(n13635), .B1(n10598), .B2(n13983), .ZN(
        n10541) );
  NOR2_X1 U13495 ( .A1(n10541), .A2(n10540), .ZN(n10542) );
  NAND2_X1 U13496 ( .A1(n10530), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10545) );
  OR2_X1 U13497 ( .A1(n20252), .A2(n20209), .ZN(n10544) );
  XNOR2_X2 U13498 ( .A(n10547), .B(n10546), .ZN(n11326) );
  NAND2_X1 U13499 ( .A1(n11327), .A2(n11326), .ZN(n10550) );
  INV_X1 U13500 ( .A(n10546), .ZN(n10548) );
  NAND2_X1 U13501 ( .A1(n10548), .A2(n10547), .ZN(n10549) );
  NAND2_X1 U13502 ( .A1(n10550), .A2(n10549), .ZN(n14028) );
  INV_X1 U13503 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14127) );
  OR2_X1 U13504 ( .A1(n10652), .A2(n14127), .ZN(n10554) );
  INV_X1 U13505 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14343) );
  OAI22_X1 U13506 ( .A1(n10606), .A2(n14343), .B1(n10598), .B2(n10070), .ZN(
        n10552) );
  INV_X1 U13507 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10760) );
  NOR2_X1 U13508 ( .A1(n10642), .A2(n10760), .ZN(n10551) );
  NOR2_X1 U13509 ( .A1(n10552), .A2(n10551), .ZN(n10553) );
  INV_X1 U13510 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14128) );
  OR2_X1 U13511 ( .A1(n10652), .A2(n14128), .ZN(n10559) );
  INV_X1 U13512 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13289) );
  OAI22_X1 U13513 ( .A1(n10606), .A2(n13289), .B1(n10598), .B2(n16592), .ZN(
        n10557) );
  INV_X1 U13514 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10794) );
  NOR2_X1 U13515 ( .A1(n10642), .A2(n10794), .ZN(n10556) );
  NOR2_X1 U13516 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  INV_X1 U13517 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16055) );
  OR2_X1 U13518 ( .A1(n10652), .A2(n16055), .ZN(n10564) );
  INV_X1 U13519 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10560) );
  OAI22_X1 U13520 ( .A1(n10606), .A2(n10560), .B1(n10598), .B2(n10068), .ZN(
        n10562) );
  INV_X1 U13521 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n16058) );
  NOR2_X1 U13522 ( .A1(n10642), .A2(n16058), .ZN(n10561) );
  NOR2_X1 U13523 ( .A1(n10562), .A2(n10561), .ZN(n10563) );
  INV_X1 U13524 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10567) );
  INV_X1 U13525 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16040) );
  OR2_X1 U13526 ( .A1(n10652), .A2(n16040), .ZN(n10566) );
  AOI22_X1 U13527 ( .A1(n10647), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10565) );
  OAI211_X1 U13528 ( .C1(n10642), .C2(n10567), .A(n10566), .B(n10565), .ZN(
        n13446) );
  INV_X1 U13529 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13912) );
  INV_X1 U13530 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16639) );
  OR2_X1 U13531 ( .A1(n10652), .A2(n16639), .ZN(n10569) );
  AOI22_X1 U13532 ( .A1(n10647), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10568) );
  OAI211_X1 U13533 ( .C1(n10642), .C2(n13912), .A(n10569), .B(n10568), .ZN(
        n13694) );
  INV_X1 U13534 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16032) );
  OR2_X1 U13535 ( .A1(n10652), .A2(n16032), .ZN(n10574) );
  INV_X1 U13536 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10570) );
  OAI22_X1 U13537 ( .A1(n10606), .A2(n10570), .B1(n10598), .B2(n16564), .ZN(
        n10572) );
  INV_X1 U13538 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n10855) );
  NOR2_X1 U13539 ( .A1(n10642), .A2(n10855), .ZN(n10571) );
  NOR2_X1 U13540 ( .A1(n10572), .A2(n10571), .ZN(n10573) );
  INV_X1 U13541 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10577) );
  INV_X1 U13542 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11519) );
  OR2_X1 U13543 ( .A1(n10652), .A2(n11519), .ZN(n10576) );
  AOI22_X1 U13544 ( .A1(n10647), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10575) );
  OAI211_X1 U13545 ( .C1(n10642), .C2(n10577), .A(n10576), .B(n10575), .ZN(
        n13485) );
  INV_X1 U13546 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16003) );
  OR2_X1 U13547 ( .A1(n10652), .A2(n16003), .ZN(n10582) );
  INV_X1 U13548 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10578) );
  OAI22_X1 U13549 ( .A1(n10606), .A2(n10578), .B1(n10598), .B2(n16544), .ZN(
        n10580) );
  INV_X1 U13550 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10888) );
  NOR2_X1 U13551 ( .A1(n10642), .A2(n10888), .ZN(n10579) );
  NOR2_X1 U13552 ( .A1(n10580), .A2(n10579), .ZN(n10581) );
  INV_X1 U13553 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16528) );
  OR2_X1 U13554 ( .A1(n10652), .A2(n16528), .ZN(n10589) );
  INV_X1 U13555 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10584) );
  INV_X1 U13556 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10583) );
  OAI22_X1 U13557 ( .A1(n10606), .A2(n10584), .B1(n10598), .B2(n10583), .ZN(
        n10587) );
  INV_X1 U13558 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10585) );
  NOR2_X1 U13559 ( .A1(n10642), .A2(n10585), .ZN(n10586) );
  NOR2_X1 U13560 ( .A1(n10587), .A2(n10586), .ZN(n10588) );
  NAND2_X1 U13561 ( .A1(n10589), .A2(n10588), .ZN(n13810) );
  NAND2_X1 U13562 ( .A1(n13809), .A2(n13810), .ZN(n13849) );
  INV_X1 U13563 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11557) );
  OR2_X1 U13564 ( .A1(n10652), .A2(n11557), .ZN(n10595) );
  INV_X1 U13565 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10590) );
  OAI22_X1 U13566 ( .A1(n10606), .A2(n10590), .B1(n10598), .B2(n16520), .ZN(
        n10593) );
  INV_X1 U13567 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n10591) );
  NOR2_X1 U13568 ( .A1(n10642), .A2(n10591), .ZN(n10592) );
  NOR2_X1 U13569 ( .A1(n10593), .A2(n10592), .ZN(n10594) );
  INV_X1 U13570 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n14045) );
  INV_X1 U13571 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16510) );
  OR2_X1 U13572 ( .A1(n10652), .A2(n16510), .ZN(n10597) );
  AOI22_X1 U13573 ( .A1(n10647), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10596) );
  OAI211_X1 U13574 ( .C1(n10642), .C2(n14045), .A(n10597), .B(n10596), .ZN(
        n13825) );
  INV_X1 U13575 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15977) );
  OR2_X1 U13576 ( .A1(n10652), .A2(n15977), .ZN(n10603) );
  INV_X1 U13577 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10599) );
  OAI22_X1 U13578 ( .A1(n10606), .A2(n10599), .B1(n10598), .B2(n16502), .ZN(
        n10601) );
  INV_X1 U13579 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n10948) );
  NOR2_X1 U13580 ( .A1(n10642), .A2(n10948), .ZN(n10600) );
  NOR2_X1 U13581 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  NAND2_X1 U13582 ( .A1(n10603), .A2(n10602), .ZN(n13936) );
  INV_X1 U13583 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14071) );
  NAND2_X1 U13584 ( .A1(n10648), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10605) );
  NAND2_X1 U13585 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10604) );
  OAI211_X1 U13586 ( .C1(n14071), .C2(n10606), .A(n10605), .B(n10604), .ZN(
        n10607) );
  AOI21_X1 U13587 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10607), .ZN(n14070) );
  NAND2_X1 U13588 ( .A1(n10647), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U13589 ( .A1(n10648), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10608) );
  OAI211_X1 U13590 ( .C1(n10598), .C2(n15705), .A(n10609), .B(n10608), .ZN(
        n10610) );
  AOI21_X1 U13591 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10610), .ZN(n15473) );
  INV_X1 U13592 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15696) );
  INV_X1 U13593 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15934) );
  OR2_X1 U13594 ( .A1(n10652), .A2(n15934), .ZN(n10612) );
  AOI22_X1 U13595 ( .A1(n10647), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10611) );
  OAI211_X1 U13596 ( .C1(n10642), .C2(n15696), .A(n10612), .B(n10611), .ZN(
        n15385) );
  INV_X1 U13597 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20154) );
  NAND2_X1 U13598 ( .A1(n10647), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U13599 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10613) );
  OAI211_X1 U13600 ( .C1(n20154), .C2(n10642), .A(n10614), .B(n10613), .ZN(
        n10615) );
  AOI21_X1 U13601 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10615), .ZN(n15462) );
  INV_X1 U13602 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15674) );
  NAND2_X1 U13603 ( .A1(n10647), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U13604 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10616) );
  OAI211_X1 U13605 ( .C1(n15674), .C2(n10642), .A(n10617), .B(n10616), .ZN(
        n10618) );
  AOI21_X1 U13606 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10618), .ZN(n15452) );
  INV_X1 U13607 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20157) );
  NAND2_X1 U13608 ( .A1(n10647), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10620) );
  NAND2_X1 U13609 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10619) );
  OAI211_X1 U13610 ( .C1(n20157), .C2(n10642), .A(n10620), .B(n10619), .ZN(
        n10621) );
  AOI21_X1 U13611 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10621), .ZN(n12931) );
  INV_X1 U13612 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n10965) );
  INV_X1 U13613 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15882) );
  OR2_X1 U13614 ( .A1(n10652), .A2(n15882), .ZN(n10623) );
  AOI22_X1 U13615 ( .A1(n10647), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10622) );
  OAI211_X1 U13616 ( .C1(n10642), .C2(n10965), .A(n10623), .B(n10622), .ZN(
        n12947) );
  INV_X1 U13617 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15645) );
  NAND2_X1 U13618 ( .A1(n10647), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10625) );
  NAND2_X1 U13619 ( .A1(n10648), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10624) );
  OAI211_X1 U13620 ( .C1(n10598), .C2(n15645), .A(n10625), .B(n10624), .ZN(
        n10626) );
  AOI21_X1 U13621 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10626), .ZN(n12958) );
  INV_X1 U13622 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20162) );
  NAND2_X1 U13623 ( .A1(n10647), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10628) );
  NAND2_X1 U13624 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10627) );
  OAI211_X1 U13625 ( .C1(n20162), .C2(n10642), .A(n10628), .B(n10627), .ZN(
        n10629) );
  AOI21_X1 U13626 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10629), .ZN(n15431) );
  INV_X1 U13627 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20164) );
  INV_X1 U13628 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15840) );
  OR2_X1 U13629 ( .A1(n10652), .A2(n15840), .ZN(n10631) );
  AOI22_X1 U13630 ( .A1(n10647), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10630) );
  OAI211_X1 U13631 ( .C1(n10642), .C2(n20164), .A(n10631), .B(n10630), .ZN(
        n15367) );
  INV_X1 U13632 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15615) );
  NAND2_X1 U13633 ( .A1(n10647), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10633) );
  NAND2_X1 U13634 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10632) );
  OAI211_X1 U13635 ( .C1(n15615), .C2(n10642), .A(n10633), .B(n10632), .ZN(
        n10634) );
  AOI21_X1 U13636 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10634), .ZN(n15416) );
  INV_X1 U13637 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20168) );
  NAND2_X1 U13638 ( .A1(n10647), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10636) );
  NAND2_X1 U13639 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10635) );
  OAI211_X1 U13640 ( .C1(n20168), .C2(n10642), .A(n10636), .B(n10635), .ZN(
        n10637) );
  AOI21_X1 U13641 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10637), .ZN(n15405) );
  INV_X1 U13642 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20169) );
  INV_X1 U13643 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15796) );
  OR2_X1 U13644 ( .A1(n10652), .A2(n15796), .ZN(n10639) );
  AOI22_X1 U13645 ( .A1(n10647), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10638) );
  OAI211_X1 U13646 ( .C1(n10642), .C2(n20169), .A(n10639), .B(n10638), .ZN(
        n15400) );
  INV_X1 U13647 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20171) );
  INV_X1 U13648 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15787) );
  OR2_X1 U13649 ( .A1(n10652), .A2(n15787), .ZN(n10641) );
  AOI22_X1 U13650 ( .A1(n10647), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10640) );
  OAI211_X1 U13651 ( .C1(n10642), .C2(n20171), .A(n10641), .B(n10640), .ZN(
        n15354) );
  INV_X1 U13652 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20174) );
  NAND2_X1 U13653 ( .A1(n10647), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10644) );
  NAND2_X1 U13654 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10643) );
  OAI211_X1 U13655 ( .C1(n20174), .C2(n10642), .A(n10644), .B(n10643), .ZN(
        n10645) );
  AOI21_X1 U13656 ( .B1(n10646), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10645), .ZN(n12823) );
  AOI22_X1 U13657 ( .A1(n10647), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n10650) );
  NAND2_X1 U13658 ( .A1(n10648), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n10649) );
  OAI211_X1 U13659 ( .C1(n10652), .C2(n10651), .A(n10650), .B(n10649), .ZN(
        n10653) );
  NAND2_X1 U13660 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20219), .ZN(
        n10655) );
  NAND2_X1 U13661 ( .A1(n10669), .A2(n10655), .ZN(n10657) );
  NAND2_X1 U13662 ( .A1(n16653), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10656) );
  XNOR2_X1 U13663 ( .A(n10680), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10664) );
  NAND2_X1 U13664 ( .A1(n20209), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10658) );
  NAND2_X1 U13665 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16675), .ZN(
        n10662) );
  NAND2_X1 U13666 ( .A1(n10663), .A2(n10662), .ZN(n10661) );
  INV_X1 U13667 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16198) );
  NAND2_X1 U13668 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16198), .ZN(
        n10660) );
  XOR2_X1 U13669 ( .A(n11677), .B(n11419), .Z(n11674) );
  NOR2_X1 U13670 ( .A1(n10663), .A2(n10662), .ZN(n11004) );
  INV_X1 U13671 ( .A(n10664), .ZN(n10665) );
  XNOR2_X1 U13672 ( .A(n10666), .B(n10665), .ZN(n11002) );
  INV_X1 U13673 ( .A(n11002), .ZN(n10667) );
  INV_X1 U13674 ( .A(n11685), .ZN(n11626) );
  XNOR2_X1 U13675 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10668) );
  XNOR2_X1 U13676 ( .A(n10669), .B(n10668), .ZN(n11673) );
  NAND2_X1 U13677 ( .A1(n11626), .A2(n11673), .ZN(n11629) );
  INV_X1 U13678 ( .A(n11629), .ZN(n10670) );
  NAND2_X1 U13679 ( .A1(n11674), .A2(n10670), .ZN(n10671) );
  NAND2_X1 U13680 ( .A1(n10672), .A2(n10673), .ZN(n16664) );
  NAND2_X1 U13681 ( .A1(n10598), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20113) );
  INV_X1 U13682 ( .A(n20113), .ZN(n10674) );
  NAND2_X1 U13683 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10674), .ZN(n19237) );
  INV_X1 U13684 ( .A(n19237), .ZN(n13332) );
  NAND2_X1 U13685 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20257) );
  INV_X1 U13686 ( .A(n20257), .ZN(n20128) );
  OR2_X1 U13687 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20128), .ZN(n12832) );
  AND2_X2 U13688 ( .A1(n14602), .A2(n10680), .ZN(n14448) );
  AND2_X2 U13689 ( .A1(n14600), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10700) );
  AOI22_X1 U13690 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n14448), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13691 ( .A1(n14406), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13693 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10676) );
  AND2_X2 U13694 ( .A1(n14601), .A2(n10680), .ZN(n10701) );
  AOI22_X1 U13695 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10701), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10675) );
  NAND4_X1 U13696 ( .A1(n10678), .A2(n10677), .A3(n10676), .A4(n10675), .ZN(
        n10686) );
  AND2_X2 U13697 ( .A1(n14600), .A2(n10680), .ZN(n10720) );
  AND2_X2 U13698 ( .A1(n10307), .A2(n16653), .ZN(n14437) );
  AOI22_X1 U13699 ( .A1(n10720), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__0__SCAN_IN), .B2(n14437), .ZN(n10684) );
  AND2_X2 U13700 ( .A1(n14595), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14446) );
  NAND3_X1 U13701 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11631) );
  INV_X1 U13702 ( .A(n11631), .ZN(n10679) );
  INV_X1 U13703 ( .A(n14440), .ZN(n14407) );
  AOI22_X1 U13704 ( .A1(n14446), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__0__SCAN_IN), .B2(n14407), .ZN(n10683) );
  AOI22_X1 U13705 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10682) );
  AND2_X2 U13706 ( .A1(n14577), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10744) );
  AOI22_X1 U13707 ( .A1(n10744), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14398), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10681) );
  NAND4_X1 U13708 ( .A1(n10684), .A2(n10683), .A3(n10682), .A4(n10681), .ZN(
        n10685) );
  NOR2_X1 U13709 ( .A1(n10686), .A2(n10685), .ZN(n13065) );
  OR2_X1 U13710 ( .A1(n10856), .A2(n10492), .ZN(n10734) );
  MUX2_X1 U13711 ( .A(n10697), .B(n20239), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10687) );
  AND2_X1 U13712 ( .A1(n10734), .A2(n10687), .ZN(n10688) );
  NAND2_X1 U13713 ( .A1(n10689), .A2(n10688), .ZN(n13163) );
  INV_X1 U13714 ( .A(n10690), .ZN(n13335) );
  INV_X1 U13715 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19251) );
  OR2_X1 U13716 ( .A1(n10860), .A2(n19251), .ZN(n10696) );
  INV_X1 U13717 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U13718 ( .A1(n10692), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10693) );
  OAI211_X1 U13719 ( .C1(n10493), .C2(n13149), .A(n10693), .B(n20205), .ZN(
        n10694) );
  INV_X1 U13720 ( .A(n10694), .ZN(n10695) );
  NAND2_X1 U13721 ( .A1(n10696), .A2(n10695), .ZN(n13164) );
  OR2_X1 U13722 ( .A1(n10860), .A2(n10459), .ZN(n10699) );
  NOR2_X1 U13723 ( .A1(n10697), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10737) );
  INV_X2 U13724 ( .A(n10856), .ZN(n10984) );
  AOI22_X1 U13725 ( .A1(n10737), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10984), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10698) );
  NAND2_X1 U13726 ( .A1(n10699), .A2(n10698), .ZN(n10716) );
  XNOR2_X1 U13727 ( .A(n10717), .B(n10716), .ZN(n13135) );
  AOI22_X1 U13728 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13729 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13730 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13731 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10702) );
  NAND4_X1 U13732 ( .A1(n10705), .A2(n10704), .A3(n10703), .A4(n10702), .ZN(
        n10713) );
  AOI22_X1 U13733 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13734 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10710) );
  INV_X1 U13735 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11388) );
  NAND2_X1 U13736 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n14437), .ZN(
        n10706) );
  OAI21_X1 U13737 ( .B1(n14440), .B2(n11388), .A(n10706), .ZN(n10707) );
  AOI21_X1 U13738 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n10707), .ZN(n10709) );
  NAND2_X1 U13739 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10708) );
  NAND4_X1 U13740 ( .A1(n10711), .A2(n10710), .A3(n10709), .A4(n10708), .ZN(
        n10712) );
  NAND2_X1 U13741 ( .A1(n10492), .A2(n19614), .ZN(n10714) );
  MUX2_X1 U13742 ( .A(n10714), .B(n20229), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10715) );
  OAI21_X1 U13743 ( .B1(n11640), .B2(n10951), .A(n10715), .ZN(n13134) );
  NOR2_X1 U13744 ( .A1(n13135), .A2(n13134), .ZN(n10719) );
  NOR2_X1 U13745 ( .A1(n10717), .A2(n10716), .ZN(n10718) );
  AOI22_X1 U13746 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13747 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13748 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13749 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10701), .B1(
        n14398), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10721) );
  NAND4_X1 U13750 ( .A1(n10724), .A2(n10723), .A3(n10722), .A4(n10721), .ZN(
        n10733) );
  AOI22_X1 U13751 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10765), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13752 ( .A1(n14406), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10730) );
  INV_X1 U13753 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10726) );
  NAND2_X1 U13754 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n14437), .ZN(
        n10725) );
  OAI21_X1 U13755 ( .B1(n14440), .B2(n10726), .A(n10725), .ZN(n10727) );
  AOI21_X1 U13756 ( .B1(n9642), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n10727), .ZN(n10729) );
  NAND2_X1 U13757 ( .A1(n14448), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10728) );
  NAND4_X1 U13758 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10732) );
  NAND2_X1 U13759 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10735) );
  OAI211_X1 U13760 ( .C1(n10951), .C2(n11642), .A(n10735), .B(n10734), .ZN(
        n10740) );
  XNOR2_X1 U13761 ( .A(n10741), .B(n10740), .ZN(n13322) );
  OR2_X1 U13762 ( .A1(n10860), .A2(n10535), .ZN(n10739) );
  AOI22_X1 U13763 ( .A1(n10989), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10984), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10738) );
  NAND2_X1 U13764 ( .A1(n10739), .A2(n10738), .ZN(n13321) );
  NOR2_X1 U13765 ( .A1(n13322), .A2(n13321), .ZN(n13323) );
  NOR2_X1 U13766 ( .A1(n10741), .A2(n10740), .ZN(n10742) );
  AOI22_X1 U13767 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n14406), .B1(
        n9642), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13768 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n14407), .ZN(n10747) );
  AOI22_X1 U13769 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10743), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13770 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10745) );
  NAND4_X1 U13771 ( .A1(n10748), .A2(n10747), .A3(n10746), .A4(n10745), .ZN(
        n10754) );
  AOI22_X1 U13772 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U13773 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10701), .B1(
        n14398), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13774 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14448), .B1(
        n10720), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U13775 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14437), .ZN(n10749) );
  NAND4_X1 U13776 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        n10753) );
  INV_X1 U13777 ( .A(n11380), .ZN(n10759) );
  OR2_X1 U13778 ( .A1(n10860), .A2(n20136), .ZN(n10758) );
  AOI22_X1 U13779 ( .A1(n10984), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10756) );
  NAND2_X1 U13780 ( .A1(n10989), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10755) );
  AND2_X1 U13781 ( .A1(n10756), .A2(n10755), .ZN(n10757) );
  OAI211_X1 U13782 ( .C1(n10951), .C2(n10759), .A(n10758), .B(n10757), .ZN(
        n13631) );
  OR2_X1 U13783 ( .A1(n10860), .A2(n10760), .ZN(n10778) );
  AOI22_X1 U13784 ( .A1(n10989), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10984), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U13785 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10779), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13786 ( .A1(n14390), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13787 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13788 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10701), .B1(
        n14398), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10761) );
  NAND4_X1 U13789 ( .A1(n10764), .A2(n10763), .A3(n10762), .A4(n10761), .ZN(
        n10775) );
  AOI22_X1 U13790 ( .A1(n14436), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13791 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10772) );
  INV_X1 U13792 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10768) );
  OAI21_X1 U13793 ( .B1(n14440), .B2(n10768), .A(n10767), .ZN(n10769) );
  AOI21_X1 U13794 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n10769), .ZN(n10771) );
  NAND2_X1 U13795 ( .A1(n14448), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10770) );
  NAND4_X1 U13796 ( .A1(n10773), .A2(n10772), .A3(n10771), .A4(n10770), .ZN(
        n10774) );
  OR2_X1 U13797 ( .A1(n10951), .A2(n11431), .ZN(n10776) );
  AOI22_X1 U13798 ( .A1(n10989), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10984), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10797) );
  INV_X1 U13799 ( .A(n13056), .ZN(n10793) );
  AOI22_X1 U13800 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13801 ( .A1(n10744), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U13802 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10781) );
  AOI22_X1 U13803 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10780) );
  NAND4_X1 U13804 ( .A1(n10783), .A2(n10782), .A3(n10781), .A4(n10780), .ZN(
        n10791) );
  AOI22_X1 U13805 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13806 ( .A1(n14406), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10788) );
  INV_X1 U13807 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13451) );
  NAND2_X1 U13808 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n14437), .ZN(
        n10784) );
  OAI21_X1 U13809 ( .B1(n14440), .B2(n13451), .A(n10784), .ZN(n10785) );
  AOI21_X1 U13810 ( .B1(n9642), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n10785), .ZN(n10787) );
  NAND2_X1 U13811 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10786) );
  NAND4_X1 U13812 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        n10790) );
  NAND2_X1 U13813 ( .A1(n11460), .A2(n10792), .ZN(n11006) );
  OAI22_X1 U13814 ( .A1(n10860), .A2(n10794), .B1(n10793), .B2(n11006), .ZN(
        n10795) );
  INV_X1 U13815 ( .A(n10795), .ZN(n10796) );
  NAND2_X1 U13816 ( .A1(n10797), .A2(n10796), .ZN(n14129) );
  AOI22_X1 U13817 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n9639), .B1(
        n14406), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10803) );
  INV_X1 U13818 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U13819 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n14437), .ZN(
        n10798) );
  OAI21_X1 U13820 ( .B1(n14440), .B2(n11481), .A(n10798), .ZN(n10799) );
  AOI21_X1 U13821 ( .B1(n10743), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n10799), .ZN(n10802) );
  AOI22_X1 U13822 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10765), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10801) );
  NAND2_X1 U13823 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10800) );
  NAND4_X1 U13824 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(
        n10809) );
  AOI22_X1 U13825 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10766), .B1(
        n9642), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13826 ( .A1(n10744), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13827 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13828 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10804) );
  NAND4_X1 U13829 ( .A1(n10807), .A2(n10806), .A3(n10805), .A4(n10804), .ZN(
        n10808) );
  NOR2_X1 U13830 ( .A1(n10809), .A2(n10808), .ZN(n11497) );
  OR2_X1 U13831 ( .A1(n10951), .A2(n11497), .ZN(n16050) );
  NAND2_X1 U13832 ( .A1(n16052), .A2(n16050), .ZN(n10812) );
  OR2_X1 U13833 ( .A1(n10860), .A2(n16058), .ZN(n10811) );
  AOI22_X1 U13834 ( .A1(n10989), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10984), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10810) );
  NAND2_X1 U13835 ( .A1(n10811), .A2(n10810), .ZN(n16049) );
  NAND2_X1 U13836 ( .A1(n10812), .A2(n16049), .ZN(n16054) );
  AOI22_X1 U13837 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U13838 ( .A1(n10779), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13839 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13840 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10813) );
  NAND4_X1 U13841 ( .A1(n10816), .A2(n10815), .A3(n10814), .A4(n10813), .ZN(
        n10825) );
  AOI22_X1 U13842 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13843 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10822) );
  INV_X1 U13844 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10818) );
  NAND2_X1 U13845 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14437), .ZN(
        n10817) );
  OAI21_X1 U13846 ( .B1(n14440), .B2(n10818), .A(n10817), .ZN(n10819) );
  AOI21_X1 U13847 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n10819), .ZN(n10821) );
  NAND2_X1 U13848 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10820) );
  NAND4_X1 U13849 ( .A1(n10823), .A2(n10822), .A3(n10821), .A4(n10820), .ZN(
        n10824) );
  OR2_X1 U13850 ( .A1(n10860), .A2(n10567), .ZN(n10827) );
  AOI22_X1 U13851 ( .A1(n10989), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10984), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13852 ( .A1(n10827), .A2(n10826), .ZN(n13620) );
  OR2_X1 U13853 ( .A1(n10860), .A2(n13912), .ZN(n10842) );
  AOI22_X1 U13854 ( .A1(n10989), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10984), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13855 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13856 ( .A1(n14406), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13857 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13858 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n14398), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10828) );
  NAND4_X1 U13859 ( .A1(n10831), .A2(n10830), .A3(n10829), .A4(n10828), .ZN(
        n10839) );
  AOI22_X1 U13860 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U13861 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10836) );
  INV_X1 U13862 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n19624) );
  NAND2_X1 U13863 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n14437), .ZN(
        n10832) );
  OAI21_X1 U13864 ( .B1(n14440), .B2(n19624), .A(n10832), .ZN(n10833) );
  AOI21_X1 U13865 ( .B1(n10765), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n10833), .ZN(n10835) );
  NAND2_X1 U13866 ( .A1(n10701), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10834) );
  NAND4_X1 U13867 ( .A1(n10837), .A2(n10836), .A3(n10835), .A4(n10834), .ZN(
        n10838) );
  OR2_X1 U13868 ( .A1(n10839), .A2(n10838), .ZN(n13475) );
  INV_X1 U13869 ( .A(n13475), .ZN(n13700) );
  OR2_X1 U13870 ( .A1(n10951), .A2(n13700), .ZN(n10840) );
  AOI22_X1 U13871 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13872 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13873 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13874 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n14448), .B1(
        n10701), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10843) );
  NAND4_X1 U13875 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10854) );
  AOI22_X1 U13876 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U13877 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10851) );
  INV_X1 U13878 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11391) );
  NAND2_X1 U13879 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14437), .ZN(
        n10847) );
  OAI21_X1 U13880 ( .B1(n14440), .B2(n11391), .A(n10847), .ZN(n10848) );
  AOI21_X1 U13881 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n10848), .ZN(n10850) );
  NAND2_X1 U13882 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10849) );
  NAND4_X1 U13883 ( .A1(n10852), .A2(n10851), .A3(n10850), .A4(n10849), .ZN(
        n10853) );
  INV_X1 U13884 ( .A(n13545), .ZN(n10859) );
  OR2_X1 U13885 ( .A1(n10860), .A2(n10855), .ZN(n10858) );
  AOI22_X1 U13886 ( .A1(n10989), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10984), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10857) );
  OAI211_X1 U13887 ( .C1(n10951), .C2(n10859), .A(n10858), .B(n10857), .ZN(
        n16026) );
  AOI22_X1 U13888 ( .A1(n14406), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U13889 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U13890 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13891 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n14448), .B1(
        n10701), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10861) );
  NAND4_X1 U13892 ( .A1(n10864), .A2(n10863), .A3(n10862), .A4(n10861), .ZN(
        n10873) );
  AOI22_X1 U13893 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13894 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10870) );
  INV_X1 U13895 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10866) );
  NAND2_X1 U13896 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14437), .ZN(
        n10865) );
  OAI21_X1 U13897 ( .B1(n14440), .B2(n10866), .A(n10865), .ZN(n10867) );
  AOI21_X1 U13898 ( .B1(n10766), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n10867), .ZN(n10869) );
  NAND2_X1 U13899 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10868) );
  NAND4_X1 U13900 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .ZN(
        n10872) );
  AOI22_X1 U13901 ( .A1(n10989), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10874) );
  OAI21_X1 U13902 ( .B1(n10951), .B2(n13480), .A(n10874), .ZN(n10875) );
  AOI21_X1 U13903 ( .B1(n10736), .B2(P2_REIP_REG_10__SCAN_IN), .A(n10875), 
        .ZN(n16621) );
  AOI22_X1 U13904 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13905 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13906 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13907 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n14448), .B1(
        n10701), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10876) );
  NAND4_X1 U13908 ( .A1(n10879), .A2(n10878), .A3(n10877), .A4(n10876), .ZN(
        n10887) );
  AOI22_X1 U13909 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U13910 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10884) );
  INV_X1 U13911 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11363) );
  NAND2_X1 U13912 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14437), .ZN(
        n10880) );
  OAI21_X1 U13913 ( .B1(n14440), .B2(n11363), .A(n10880), .ZN(n10881) );
  AOI21_X1 U13914 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n10881), .ZN(n10883) );
  NAND2_X1 U13915 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10882) );
  NAND4_X1 U13916 ( .A1(n10885), .A2(n10884), .A3(n10883), .A4(n10882), .ZN(
        n10886) );
  INV_X1 U13917 ( .A(n13605), .ZN(n10891) );
  OR2_X1 U13918 ( .A1(n10860), .A2(n10888), .ZN(n10890) );
  AOI22_X1 U13919 ( .A1(n10989), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10889) );
  OAI211_X1 U13920 ( .C1(n10951), .C2(n10891), .A(n10890), .B(n10889), .ZN(
        n16008) );
  NAND2_X1 U13921 ( .A1(n16007), .A2(n16008), .ZN(n16006) );
  AOI22_X1 U13922 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13923 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13924 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13925 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10892) );
  NAND4_X1 U13926 ( .A1(n10895), .A2(n10894), .A3(n10893), .A4(n10892), .ZN(
        n10903) );
  AOI22_X1 U13927 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U13928 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10900) );
  INV_X1 U13929 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13767) );
  NAND2_X1 U13930 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14437), .ZN(
        n10896) );
  OAI21_X1 U13931 ( .B1(n14440), .B2(n13767), .A(n10896), .ZN(n10897) );
  AOI21_X1 U13932 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n10897), .ZN(n10899) );
  NAND2_X1 U13933 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10898) );
  NAND4_X1 U13934 ( .A1(n10901), .A2(n10900), .A3(n10899), .A4(n10898), .ZN(
        n10902) );
  NOR2_X1 U13935 ( .A1(n10903), .A2(n10902), .ZN(n13846) );
  AOI22_X1 U13936 ( .A1(n10989), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10904) );
  OAI21_X1 U13937 ( .B1(n10951), .B2(n13846), .A(n10904), .ZN(n10905) );
  AOI21_X1 U13938 ( .B1(n10736), .B2(P2_REIP_REG_12__SCAN_IN), .A(n10905), 
        .ZN(n13890) );
  AOI22_X1 U13939 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13940 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U13941 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U13942 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n14448), .B1(
        n10701), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10906) );
  NAND4_X1 U13943 ( .A1(n10909), .A2(n10908), .A3(n10907), .A4(n10906), .ZN(
        n10917) );
  AOI22_X1 U13944 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13945 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10914) );
  INV_X1 U13946 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14401) );
  NAND2_X1 U13947 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n14437), .ZN(
        n10910) );
  OAI21_X1 U13948 ( .B1(n14440), .B2(n14401), .A(n10910), .ZN(n10911) );
  AOI21_X1 U13949 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n10911), .ZN(n10913) );
  NAND2_X1 U13950 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10912) );
  NAND4_X1 U13951 ( .A1(n10915), .A2(n10914), .A3(n10913), .A4(n10912), .ZN(
        n10916) );
  NOR2_X1 U13952 ( .A1(n10917), .A2(n10916), .ZN(n13845) );
  NAND2_X1 U13953 ( .A1(n10736), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U13954 ( .A1(n10989), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10918) );
  OAI211_X1 U13955 ( .C1(n13845), .C2(n10951), .A(n10919), .B(n10918), .ZN(
        n15988) );
  NAND2_X1 U13956 ( .A1(n13889), .A2(n15988), .ZN(n15987) );
  INV_X1 U13957 ( .A(n10951), .ZN(n10934) );
  AOI22_X1 U13958 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n9639), .B1(
        n14406), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10925) );
  INV_X1 U13959 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11473) );
  NAND2_X1 U13960 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14437), .ZN(
        n10920) );
  OAI21_X1 U13961 ( .B1(n14440), .B2(n11473), .A(n10920), .ZN(n10921) );
  AOI21_X1 U13962 ( .B1(n10765), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n10921), .ZN(n10924) );
  AOI22_X1 U13963 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U13964 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10922) );
  NAND4_X1 U13965 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n10931) );
  AOI22_X1 U13966 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13967 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13968 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13969 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n14448), .B1(
        n10701), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10926) );
  NAND4_X1 U13970 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n10930) );
  NOR2_X1 U13971 ( .A1(n10931), .A2(n10930), .ZN(n13831) );
  INV_X1 U13972 ( .A(n13831), .ZN(n13834) );
  AOI22_X1 U13973 ( .A1(n10989), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10932) );
  OAI21_X1 U13974 ( .B1(n10860), .B2(n14045), .A(n10932), .ZN(n10933) );
  AOI21_X1 U13975 ( .B1(n10934), .B2(n13834), .A(n10933), .ZN(n14043) );
  AOI22_X1 U13976 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13977 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13978 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13979 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n14448), .B1(
        n10701), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10935) );
  NAND4_X1 U13980 ( .A1(n10938), .A2(n10937), .A3(n10936), .A4(n10935), .ZN(
        n10947) );
  AOI22_X1 U13981 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U13982 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10944) );
  INV_X1 U13983 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10940) );
  NAND2_X1 U13984 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14437), .ZN(
        n10939) );
  OAI21_X1 U13985 ( .B1(n14440), .B2(n10940), .A(n10939), .ZN(n10941) );
  AOI21_X1 U13986 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n10941), .ZN(n10943) );
  NAND2_X1 U13987 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10942) );
  NAND4_X1 U13988 ( .A1(n10945), .A2(n10944), .A3(n10943), .A4(n10942), .ZN(
        n10946) );
  OR2_X1 U13989 ( .A1(n10860), .A2(n10948), .ZN(n10950) );
  AOI22_X1 U13990 ( .A1(n10989), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10949) );
  OAI211_X1 U13991 ( .C1(n10951), .C2(n10223), .A(n10950), .B(n10949), .ZN(
        n15970) );
  INV_X1 U13992 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n10952) );
  OR2_X1 U13993 ( .A1(n10860), .A2(n10952), .ZN(n10954) );
  AOI22_X1 U13994 ( .A1(n10989), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10953) );
  NAND2_X1 U13995 ( .A1(n10954), .A2(n10953), .ZN(n14114) );
  INV_X1 U13996 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20151) );
  OR2_X1 U13997 ( .A1(n10860), .A2(n20151), .ZN(n10956) );
  AOI22_X1 U13998 ( .A1(n10989), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10955) );
  AND2_X1 U13999 ( .A1(n10956), .A2(n10955), .ZN(n14160) );
  OR2_X1 U14000 ( .A1(n10860), .A2(n15696), .ZN(n10958) );
  AOI22_X1 U14001 ( .A1(n10989), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10957) );
  NAND2_X1 U14002 ( .A1(n10958), .A2(n10957), .ZN(n15380) );
  NAND2_X1 U14003 ( .A1(n15381), .A2(n15380), .ZN(n15379) );
  OR2_X1 U14004 ( .A1(n10860), .A2(n20154), .ZN(n10960) );
  AOI22_X1 U14005 ( .A1(n10989), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10959) );
  AND2_X1 U14006 ( .A1(n10960), .A2(n10959), .ZN(n15555) );
  OR2_X1 U14007 ( .A1(n10860), .A2(n15674), .ZN(n10962) );
  AOI22_X1 U14008 ( .A1(n10989), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10961) );
  AND2_X1 U14009 ( .A1(n10962), .A2(n10961), .ZN(n15904) );
  OR2_X1 U14010 ( .A1(n10860), .A2(n20157), .ZN(n10964) );
  AOI22_X1 U14011 ( .A1(n10989), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10963) );
  NAND2_X1 U14012 ( .A1(n10964), .A2(n10963), .ZN(n12932) );
  OR2_X1 U14013 ( .A1(n10860), .A2(n10965), .ZN(n10967) );
  AOI22_X1 U14014 ( .A1(n10989), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10966) );
  NAND2_X1 U14015 ( .A1(n10967), .A2(n10966), .ZN(n12962) );
  INV_X1 U14016 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20160) );
  OR2_X1 U14017 ( .A1(n10860), .A2(n20160), .ZN(n10969) );
  AOI22_X1 U14018 ( .A1(n10989), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U14019 ( .A1(n10969), .A2(n10968), .ZN(n12961) );
  OR2_X1 U14020 ( .A1(n10860), .A2(n20162), .ZN(n10972) );
  AOI22_X1 U14021 ( .A1(n10989), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10971) );
  AND2_X1 U14022 ( .A1(n10972), .A2(n10971), .ZN(n15525) );
  OR2_X1 U14023 ( .A1(n10860), .A2(n20164), .ZN(n10974) );
  AOI22_X1 U14024 ( .A1(n10989), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10973) );
  NAND2_X1 U14025 ( .A1(n10974), .A2(n10973), .ZN(n15369) );
  NAND2_X1 U14026 ( .A1(n15527), .A2(n15369), .ZN(n15511) );
  OR2_X1 U14027 ( .A1(n10860), .A2(n15615), .ZN(n10976) );
  AOI22_X1 U14028 ( .A1(n10989), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10975) );
  AND2_X1 U14029 ( .A1(n10976), .A2(n10975), .ZN(n15510) );
  OR2_X1 U14030 ( .A1(n10860), .A2(n20168), .ZN(n10979) );
  AOI22_X1 U14031 ( .A1(n10989), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10978) );
  AND2_X1 U14032 ( .A1(n10979), .A2(n10978), .ZN(n15499) );
  OR2_X1 U14033 ( .A1(n10860), .A2(n20169), .ZN(n10981) );
  AOI22_X1 U14034 ( .A1(n10989), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10980) );
  AND2_X1 U14035 ( .A1(n10981), .A2(n10980), .ZN(n15489) );
  OR2_X1 U14036 ( .A1(n10860), .A2(n20171), .ZN(n10983) );
  AOI22_X1 U14037 ( .A1(n10989), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U14038 ( .A1(n10983), .A2(n10982), .ZN(n15357) );
  INV_X1 U14039 ( .A(n12826), .ZN(n10988) );
  OR2_X1 U14040 ( .A1(n10860), .A2(n20174), .ZN(n10986) );
  AOI22_X1 U14041 ( .A1(n10989), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10985) );
  AND2_X1 U14042 ( .A1(n10986), .A2(n10985), .ZN(n12827) );
  INV_X1 U14043 ( .A(n12827), .ZN(n10987) );
  NAND2_X1 U14044 ( .A1(n10988), .A2(n10987), .ZN(n12829) );
  AOI222_X1 U14045 ( .A1(n10736), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n10984), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n10989), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n10990) );
  NOR2_X1 U14046 ( .A1(n10672), .A2(n19237), .ZN(n10991) );
  AND2_X2 U14047 ( .A1(n12978), .A2(n10493), .ZN(n19545) );
  NOR2_X1 U14048 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20124) );
  AOI211_X1 U14049 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n20124), .ZN(n20262) );
  NAND2_X1 U14050 ( .A1(n20262), .A2(n20257), .ZN(n13043) );
  NOR2_X1 U14051 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13043), .ZN(n10994) );
  NOR2_X1 U14052 ( .A1(n19435), .A2(n19408), .ZN(n10998) );
  NOR2_X1 U14053 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20198) );
  INV_X1 U14054 ( .A(n20198), .ZN(n19233) );
  NOR2_X1 U14055 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19233), .ZN(n12974) );
  NAND2_X1 U14056 ( .A1(n12974), .A2(n20256), .ZN(n19333) );
  NOR3_X1 U14057 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20113), .A3(n20205), 
        .ZN(n16698) );
  NOR2_X1 U14058 ( .A1(n16698), .A2(n19411), .ZN(n10992) );
  NAND2_X1 U14059 ( .A1(n19364), .A2(n10992), .ZN(n10993) );
  INV_X1 U14060 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n11698) );
  INV_X2 U14061 ( .A(n19386), .ZN(n19431) );
  NAND2_X1 U14062 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19431), .ZN(
        n10996) );
  INV_X1 U14063 ( .A(n10994), .ZN(n16701) );
  NAND3_X1 U14064 ( .A1(n19545), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n16701), 
        .ZN(n10995) );
  OAI211_X1 U14065 ( .C1(n19416), .C2(n11698), .A(n10996), .B(n10995), .ZN(
        n10997) );
  AOI211_X1 U14066 ( .C1(n15757), .C2(n19425), .A(n10998), .B(n10997), .ZN(
        n11015) );
  MUX2_X1 U14067 ( .A(n13198), .B(n11622), .S(n10792), .Z(n11424) );
  NOR2_X1 U14068 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11000) );
  MUX2_X1 U14069 ( .A(n11001), .B(n11000), .S(n10495), .Z(n11420) );
  OAI21_X1 U14070 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n10792), .A(n11006), .ZN(
        n11464) );
  MUX2_X1 U14071 ( .A(n11497), .B(P2_EBX_REG_6__SCAN_IN), .S(n10495), .Z(
        n11504) );
  MUX2_X1 U14072 ( .A(n11667), .B(P2_EBX_REG_7__SCAN_IN), .S(n10495), .Z(
        n11510) );
  INV_X1 U14073 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U14074 ( .A1(n11515), .A2(n11007), .ZN(n11008) );
  INV_X1 U14075 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13489) );
  NAND2_X1 U14076 ( .A1(n19597), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11531) );
  NOR2_X1 U14077 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(P2_EBX_REG_15__SCAN_IN), 
        .ZN(n11009) );
  NOR2_X1 U14078 ( .A1(n10792), .A2(n11009), .ZN(n11010) );
  NAND2_X1 U14079 ( .A1(n19597), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11568) );
  AND2_X1 U14080 ( .A1(n19597), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11546) );
  AND2_X1 U14081 ( .A1(n19597), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U14082 ( .A1(n11602), .A2(n9713), .ZN(n11011) );
  NAND2_X1 U14083 ( .A1(n19597), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11589) );
  AND2_X1 U14084 ( .A1(n19597), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11593) );
  INV_X1 U14085 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11012) );
  NAND2_X1 U14086 ( .A1(n19597), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16437) );
  INV_X1 U14087 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11013) );
  NOR2_X1 U14088 ( .A1(n10792), .A2(n11013), .ZN(n11605) );
  NAND2_X1 U14089 ( .A1(n19597), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11611) );
  MUX2_X1 U14090 ( .A(n11014), .B(n11604), .S(n10792), .Z(n11619) );
  NAND2_X1 U14091 ( .A1(n20253), .A2(n9702), .ZN(n19423) );
  NAND3_X1 U14092 ( .A1(n11016), .A2(n11015), .A3(n10295), .ZN(P2_U2824) );
  OR3_X2 U14093 ( .A1(n19177), .A2(n19167), .A3(n19020), .ZN(n11180) );
  INV_X2 U14094 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19185) );
  OR2_X2 U14095 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11026), .ZN(
        n17274) );
  AOI22_X1 U14096 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11034) );
  INV_X1 U14097 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U14098 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11020) );
  INV_X2 U14099 ( .A(n10316), .ZN(n14248) );
  AOI22_X1 U14100 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11019) );
  OAI211_X1 U14101 ( .C1(n17526), .C2(n17330), .A(n11020), .B(n11019), .ZN(
        n11032) );
  AOI22_X1 U14102 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U14103 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14104 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U14105 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11027) );
  NAND4_X1 U14106 ( .A1(n11030), .A2(n11029), .A3(n11028), .A4(n11027), .ZN(
        n11031) );
  INV_X1 U14107 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17361) );
  AOI22_X1 U14108 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11035) );
  OAI21_X1 U14109 ( .B1(n11241), .B2(n17361), .A(n11035), .ZN(n11045) );
  INV_X1 U14110 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U14111 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11043) );
  AOI22_X1 U14112 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11037) );
  OAI21_X1 U14113 ( .B1(n17500), .B2(n17478), .A(n11037), .ZN(n11042) );
  INV_X1 U14114 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U14115 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U14116 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11038) );
  OAI211_X1 U14117 ( .C1(n17526), .C2(n11040), .A(n11039), .B(n11038), .ZN(
        n11041) );
  OAI21_X1 U14118 ( .B1(n11180), .B2(n18560), .A(n11046), .ZN(n11050) );
  INV_X1 U14119 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U14120 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11047) );
  OAI21_X1 U14121 ( .B1(n9710), .B2(n11048), .A(n11047), .ZN(n11049) );
  INV_X1 U14122 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U14123 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11055) );
  INV_X1 U14124 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11052) );
  INV_X1 U14125 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11051) );
  OAI22_X1 U14126 ( .A1(n10316), .A2(n11052), .B1(n17388), .B2(n11051), .ZN(
        n11053) );
  INV_X1 U14127 ( .A(n11053), .ZN(n11054) );
  OAI211_X1 U14128 ( .C1(n17526), .C2(n17507), .A(n11055), .B(n11054), .ZN(
        n11058) );
  INV_X1 U14129 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14238) );
  NAND2_X1 U14130 ( .A1(n11056), .A2(n10306), .ZN(n11057) );
  NOR2_X1 U14131 ( .A1(n11058), .A2(n11057), .ZN(n11060) );
  AOI22_X1 U14132 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14133 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17501), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17433), .ZN(n11063) );
  INV_X1 U14134 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17532) );
  INV_X4 U14135 ( .A(n17274), .ZN(n17538) );
  AOI22_X1 U14136 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17541), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11066) );
  INV_X1 U14137 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17527) );
  NAND2_X1 U14138 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11065) );
  INV_X1 U14139 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14202) );
  NAND2_X1 U14140 ( .A1(n11068), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11069) );
  INV_X1 U14141 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14206) );
  INV_X2 U14142 ( .A(n17500), .ZN(n17520) );
  AOI22_X1 U14143 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17520), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11070) );
  OAI21_X1 U14144 ( .B1(n9709), .B2(n14206), .A(n11070), .ZN(n11071) );
  INV_X1 U14145 ( .A(n11071), .ZN(n11072) );
  INV_X1 U14146 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U14147 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17545), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11082) );
  INV_X1 U14148 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17486) );
  AOI22_X1 U14149 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14150 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11073) );
  OAI211_X1 U14151 ( .C1(n10314), .C2(n17486), .A(n11074), .B(n11073), .ZN(
        n11080) );
  AOI22_X1 U14152 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U14153 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14154 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U14155 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11075) );
  NAND4_X1 U14156 ( .A1(n11078), .A2(n11077), .A3(n11076), .A4(n11075), .ZN(
        n11079) );
  INV_X1 U14157 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18796) );
  AOI22_X1 U14158 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11092) );
  INV_X1 U14159 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14179) );
  AOI22_X1 U14160 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14161 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11083) );
  OAI211_X1 U14162 ( .C1(n17526), .C2(n14179), .A(n11084), .B(n11083), .ZN(
        n11090) );
  AOI22_X1 U14163 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14164 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U14165 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11086) );
  NAND2_X1 U14166 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11085) );
  NAND4_X1 U14167 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n11089) );
  OAI211_X1 U14168 ( .C1(n17557), .C2(n18796), .A(n11092), .B(n11091), .ZN(
        n17720) );
  INV_X1 U14169 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14234) );
  AOI22_X1 U14170 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11102) );
  INV_X1 U14171 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U14172 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U14173 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11093) );
  OAI211_X1 U14174 ( .C1(n17526), .C2(n17282), .A(n11094), .B(n11093), .ZN(
        n11100) );
  AOI22_X1 U14175 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14176 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14177 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11096) );
  NAND2_X1 U14178 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11095) );
  NAND4_X1 U14179 ( .A1(n11098), .A2(n11097), .A3(n11096), .A4(n11095), .ZN(
        n11099) );
  AOI211_X1 U14180 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11100), .B(n11099), .ZN(n11101) );
  OAI211_X1 U14181 ( .C1(n17274), .C2(n14234), .A(n11102), .B(n11101), .ZN(
        n16746) );
  INV_X1 U14182 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17905) );
  INV_X1 U14183 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18490) );
  INV_X1 U14184 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18508) );
  INV_X1 U14185 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19173) );
  NOR2_X1 U14186 ( .A1(n11284), .A2(n19173), .ZN(n11118) );
  INV_X1 U14187 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U14188 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14189 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11105) );
  OAI211_X1 U14190 ( .C1(n17526), .C2(n17556), .A(n11106), .B(n11105), .ZN(
        n11107) );
  AOI22_X1 U14191 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U14192 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U14193 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11109) );
  NAND2_X1 U14194 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11108) );
  NAND4_X1 U14195 ( .A1(n11111), .A2(n11110), .A3(n11109), .A4(n11108), .ZN(
        n11115) );
  AOI22_X1 U14196 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11113) );
  INV_X1 U14197 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17419) );
  NAND3_X1 U14198 ( .A1(n11113), .A2(n11112), .A3(n10304), .ZN(n11114) );
  NAND2_X1 U14199 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18205), .ZN(
        n18204) );
  NOR2_X1 U14200 ( .A1(n18198), .A2(n18204), .ZN(n18197) );
  XNOR2_X1 U14201 ( .A(n17729), .B(n11120), .ZN(n18172) );
  NOR2_X1 U14202 ( .A1(n11121), .A2(n18490), .ZN(n11122) );
  XNOR2_X1 U14203 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11124), .ZN(
        n18164) );
  XOR2_X1 U14204 ( .A(n17720), .B(n11125), .Z(n11126) );
  NOR2_X1 U14205 ( .A1(n11127), .A2(n11126), .ZN(n18150) );
  INV_X1 U14206 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18467) );
  INV_X1 U14207 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18132) );
  NOR2_X1 U14208 ( .A1(n11131), .A2(n11130), .ZN(n11132) );
  INV_X1 U14209 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18442) );
  INV_X1 U14210 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11134) );
  INV_X1 U14211 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18375) );
  INV_X1 U14212 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18398) );
  INV_X1 U14213 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18361) );
  INV_X1 U14214 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18345) );
  NAND2_X1 U14215 ( .A1(n18361), .A2(n18345), .ZN(n11135) );
  NAND2_X1 U14216 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18418) );
  NOR2_X1 U14217 ( .A1(n18418), .A2(n18375), .ZN(n18378) );
  NAND3_X1 U14218 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18378), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18347) );
  NOR2_X1 U14219 ( .A1(n18347), .A2(n18361), .ZN(n18335) );
  INV_X1 U14220 ( .A(n18335), .ZN(n11315) );
  NOR2_X1 U14221 ( .A1(n11315), .A2(n18345), .ZN(n18315) );
  INV_X1 U14222 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18334) );
  INV_X1 U14223 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18005) );
  NAND2_X1 U14224 ( .A1(n11139), .A2(n11140), .ZN(n18011) );
  NOR2_X1 U14225 ( .A1(n18334), .A2(n18005), .ZN(n18318) );
  INV_X1 U14226 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17988) );
  INV_X1 U14227 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17961) );
  NAND2_X1 U14228 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17958) );
  NOR3_X1 U14229 ( .A1(n17988), .A2(n17961), .A3(n17958), .ZN(n11145) );
  NAND2_X1 U14230 ( .A1(n18318), .A2(n11145), .ZN(n18276) );
  INV_X1 U14231 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17940) );
  NOR2_X1 U14232 ( .A1(n18276), .A2(n17940), .ZN(n18213) );
  NAND2_X1 U14233 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18213), .ZN(
        n18252) );
  INV_X1 U14234 ( .A(n18252), .ZN(n11141) );
  INV_X1 U14235 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17986) );
  NAND2_X1 U14236 ( .A1(n17995), .A2(n17986), .ZN(n11142) );
  NOR2_X2 U14237 ( .A1(n17911), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17910) );
  AND2_X1 U14238 ( .A1(n11145), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11146) );
  INV_X1 U14239 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18254) );
  NOR3_X2 U14240 ( .A1(n17910), .A2(n17920), .A3(n18254), .ZN(n17904) );
  NAND2_X1 U14241 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11319) );
  INV_X1 U14242 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11149) );
  INV_X1 U14243 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17852) );
  NOR2_X1 U14244 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18109), .ZN(
        n16754) );
  AOI21_X1 U14245 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18109), .A(
        n16754), .ZN(n17857) );
  NAND2_X1 U14246 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16729) );
  INV_X1 U14247 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16121) );
  NOR2_X1 U14248 ( .A1(n16729), .A2(n16121), .ZN(n16173) );
  INV_X1 U14249 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19172) );
  AOI22_X1 U14250 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n9883), .B1(
        n18109), .B2(n19172), .ZN(n11152) );
  OAI21_X1 U14251 ( .B1(n11154), .B2(n16174), .A(n11152), .ZN(n11158) );
  INV_X1 U14252 ( .A(n11150), .ZN(n11151) );
  NOR2_X1 U14253 ( .A1(n16176), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12887) );
  INV_X1 U14254 ( .A(n11154), .ZN(n11155) );
  NAND2_X1 U14255 ( .A1(n11156), .A2(n11155), .ZN(n11157) );
  NAND2_X1 U14256 ( .A1(n11158), .A2(n11157), .ZN(n12883) );
  INV_X1 U14257 ( .A(n16746), .ZN(n17713) );
  INV_X1 U14258 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U14259 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17544), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11159) );
  OAI21_X1 U14260 ( .B1(n9709), .B2(n17411), .A(n11159), .ZN(n11167) );
  INV_X1 U14261 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U14262 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11165) );
  INV_X1 U14263 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14211) );
  OAI22_X1 U14264 ( .A1(n9652), .A2(n14206), .B1(n10316), .B2(n14211), .ZN(
        n11163) );
  AOI22_X1 U14265 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11161) );
  AOI22_X1 U14266 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11160) );
  AOI211_X1 U14267 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n11163), .B(n11162), .ZN(n11164) );
  OAI211_X1 U14268 ( .C1(n17274), .C2(n17519), .A(n11165), .B(n11164), .ZN(
        n11166) );
  AOI211_X4 U14269 ( .C1(n9647), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n11167), .B(n11166), .ZN(n19212) );
  INV_X1 U14270 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19171) );
  NAND2_X1 U14271 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19171), .ZN(n19055) );
  NOR2_X1 U14272 ( .A1(n19055), .A2(n19222), .ZN(n19206) );
  INV_X1 U14273 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18540) );
  OAI22_X1 U14274 ( .A1(n19177), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19030), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14275 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19012), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19185), .ZN(n11265) );
  OAI21_X1 U14276 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19177), .A(
        n11169), .ZN(n11170) );
  NAND2_X1 U14277 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11170), .ZN(
        n11172) );
  OAI22_X1 U14278 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18540), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11170), .ZN(n11174) );
  AOI21_X1 U14279 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11172), .A(
        n11174), .ZN(n11171) );
  AOI21_X1 U14280 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18540), .A(
        n11171), .ZN(n11267) );
  NOR2_X1 U14281 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18540), .ZN(
        n11173) );
  AOI22_X1 U14282 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11174), .B1(
        n11173), .B2(n11172), .ZN(n11178) );
  NAND2_X1 U14283 ( .A1(n11177), .A2(n11176), .ZN(n11175) );
  OAI211_X1 U14284 ( .C1(n11177), .C2(n11176), .A(n11178), .B(n11175), .ZN(
        n11270) );
  NAND3_X1 U14285 ( .A1(n11265), .A2(n11178), .A3(n11264), .ZN(n11179) );
  NAND3_X1 U14286 ( .A1(n11267), .A2(n11270), .A3(n11179), .ZN(n18991) );
  INV_X1 U14287 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17469) );
  OAI22_X1 U14288 ( .A1(n9709), .A2(n17478), .B1(n11021), .B2(n17469), .ZN(
        n11190) );
  INV_X1 U14289 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U14290 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11188) );
  INV_X1 U14291 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18571) );
  AOI22_X1 U14292 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11181) );
  OAI21_X1 U14293 ( .B1(n17522), .B2(n18571), .A(n11181), .ZN(n11186) );
  AOI22_X1 U14294 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14295 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14296 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11182) );
  NAND3_X1 U14297 ( .A1(n11184), .A2(n11183), .A3(n11182), .ZN(n11185) );
  AOI211_X1 U14298 ( .C1(n17545), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n11186), .B(n11185), .ZN(n11187) );
  OAI211_X1 U14299 ( .C1(n14198), .C2(n17467), .A(n11188), .B(n11187), .ZN(
        n11189) );
  INV_X1 U14300 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18790) );
  AOI22_X1 U14301 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U14302 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11191) );
  OAI211_X1 U14303 ( .C1(n17526), .C2(n18790), .A(n11192), .B(n11191), .ZN(
        n11200) );
  INV_X1 U14304 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18760) );
  AOI22_X1 U14305 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11198) );
  INV_X1 U14306 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18564) );
  AOI22_X1 U14307 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11193) );
  OAI21_X1 U14308 ( .B1(n17522), .B2(n18564), .A(n11193), .ZN(n11196) );
  INV_X1 U14309 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U14310 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11194) );
  OAI21_X1 U14311 ( .B1(n11036), .B2(n17484), .A(n11194), .ZN(n11195) );
  OAI211_X1 U14312 ( .C1(n17557), .C2(n18760), .A(n11198), .B(n11197), .ZN(
        n11199) );
  AOI211_X2 U14313 ( .C1(n9641), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n11200), .B(n11199), .ZN(n11254) );
  INV_X1 U14314 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18806) );
  AOI22_X1 U14315 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14316 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11201) );
  OAI211_X1 U14317 ( .C1(n17526), .C2(n18806), .A(n11202), .B(n11201), .ZN(
        n11210) );
  INV_X1 U14318 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U14319 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11208) );
  INV_X1 U14320 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18590) );
  AOI22_X1 U14321 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11203) );
  OAI21_X1 U14322 ( .B1(n17522), .B2(n18590), .A(n11203), .ZN(n11206) );
  INV_X1 U14323 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U14324 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11204) );
  OAI21_X1 U14325 ( .B1(n17388), .B2(n17273), .A(n11204), .ZN(n11205) );
  AOI211_X1 U14326 ( .C1(n17545), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n11206), .B(n11205), .ZN(n11207) );
  OAI211_X1 U14327 ( .C1(n9709), .C2(n17442), .A(n11208), .B(n11207), .ZN(
        n11209) );
  AOI211_X4 U14328 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n11210), .B(n11209), .ZN(n17711) );
  INV_X1 U14329 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18752) );
  AOI22_X1 U14330 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11220) );
  INV_X1 U14331 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18782) );
  AOI22_X1 U14332 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14333 ( .A1(n14248), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11211) );
  OAI211_X1 U14334 ( .C1(n17526), .C2(n18782), .A(n11212), .B(n11211), .ZN(
        n11218) );
  AOI22_X1 U14335 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14336 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14337 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U14338 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11213) );
  NAND4_X1 U14339 ( .A1(n11216), .A2(n11215), .A3(n11214), .A4(n11213), .ZN(
        n11217) );
  INV_X1 U14340 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17459) );
  AOI22_X1 U14341 ( .A1(n14248), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11221) );
  OAI21_X1 U14342 ( .B1(n11180), .B2(n17459), .A(n11221), .ZN(n11230) );
  INV_X1 U14343 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U14344 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11228) );
  INV_X1 U14345 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17329) );
  OAI22_X1 U14346 ( .A1(n11062), .A2(n17329), .B1(n11241), .B2(n18582), .ZN(
        n11226) );
  AOI22_X1 U14347 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9655), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14348 ( .A1(n11068), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11223) );
  NAND3_X1 U14349 ( .A1(n11224), .A2(n11223), .A3(n11222), .ZN(n11225) );
  OAI211_X1 U14350 ( .C1(n17500), .C2(n17449), .A(n11228), .B(n11227), .ZN(
        n11229) );
  AOI22_X1 U14351 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11232) );
  AOI22_X1 U14352 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11231) );
  OAI211_X1 U14353 ( .C1(n17526), .C2(n18796), .A(n11232), .B(n11231), .ZN(
        n11240) );
  AOI22_X1 U14354 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17545), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11238) );
  AOI22_X1 U14355 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11237) );
  INV_X1 U14356 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18576) );
  INV_X1 U14357 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16085) );
  OAI22_X1 U14358 ( .A1(n11241), .A2(n18576), .B1(n11180), .B2(n16085), .ZN(
        n11235) );
  INV_X1 U14359 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17347) );
  AOI22_X1 U14360 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11233) );
  OAI21_X1 U14361 ( .B1(n11036), .B2(n17347), .A(n11233), .ZN(n11234) );
  AOI211_X1 U14362 ( .C1(n9651), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n11235), .B(n11234), .ZN(n11236) );
  NAND3_X1 U14363 ( .A1(n11238), .A2(n11237), .A3(n11236), .ZN(n11239) );
  AOI211_X2 U14364 ( .C1(n9641), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n11240), .B(n11239), .ZN(n11251) );
  NOR2_X1 U14365 ( .A1(n9663), .A2(n11251), .ZN(n12868) );
  NAND4_X1 U14366 ( .A1(n11259), .A2(n11254), .A3(n11256), .A4(n12868), .ZN(
        n11253) );
  INV_X1 U14367 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17499) );
  INV_X1 U14368 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17498) );
  OAI22_X1 U14369 ( .A1(n9652), .A2(n17499), .B1(n11180), .B2(n17498), .ZN(
        n11245) );
  AOI22_X1 U14370 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14371 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11242) );
  NAND2_X1 U14372 ( .A1(n9663), .A2(n18567), .ZN(n18998) );
  NAND2_X1 U14373 ( .A1(n11251), .A2(n18578), .ZN(n11272) );
  NAND3_X1 U14374 ( .A1(n12869), .A2(n18998), .A3(n11272), .ZN(n11247) );
  INV_X1 U14375 ( .A(n11251), .ZN(n18573) );
  NAND2_X1 U14376 ( .A1(n12869), .A2(n18573), .ZN(n12877) );
  NOR2_X1 U14377 ( .A1(n18551), .A2(n17195), .ZN(n11257) );
  OAI21_X1 U14378 ( .B1(n17711), .B2(n19006), .A(n11257), .ZN(n11246) );
  INV_X1 U14379 ( .A(n11246), .ZN(n12874) );
  AOI21_X1 U14380 ( .B1(n11247), .B2(n12877), .A(n12874), .ZN(n11250) );
  INV_X1 U14381 ( .A(n11254), .ZN(n18561) );
  OAI22_X1 U14382 ( .A1(n11256), .A2(n18561), .B1(n18545), .B2(n11247), .ZN(
        n11249) );
  INV_X1 U14383 ( .A(n12869), .ZN(n18557) );
  OAI21_X1 U14384 ( .B1(n12868), .B2(n17711), .A(n18567), .ZN(n11248) );
  NOR2_X1 U14385 ( .A1(n17711), .A2(n11254), .ZN(n11261) );
  NAND3_X1 U14386 ( .A1(n11258), .A2(n11251), .A3(n18545), .ZN(n11252) );
  NOR2_X1 U14387 ( .A1(n12869), .A2(n11253), .ZN(n12870) );
  NAND2_X1 U14388 ( .A1(n12869), .A2(n11254), .ZN(n18997) );
  INV_X1 U14389 ( .A(n14173), .ZN(n11255) );
  NOR2_X1 U14390 ( .A1(n11275), .A2(n11257), .ZN(n19224) );
  INV_X1 U14391 ( .A(n18984), .ZN(n11260) );
  NOR2_X1 U14392 ( .A1(n11261), .A2(n11260), .ZN(n11263) );
  INV_X1 U14393 ( .A(n11264), .ZN(n11269) );
  XNOR2_X1 U14394 ( .A(n11266), .B(n11265), .ZN(n11268) );
  OAI21_X1 U14395 ( .B1(n11268), .B2(n11270), .A(n11267), .ZN(n16862) );
  OAI21_X1 U14396 ( .B1(n11270), .B2(n11269), .A(n18986), .ZN(n12880) );
  NAND2_X1 U14397 ( .A1(n12869), .A2(n18551), .ZN(n12875) );
  NOR2_X1 U14398 ( .A1(n9663), .A2(n12875), .ZN(n12881) );
  INV_X1 U14399 ( .A(n11272), .ZN(n11274) );
  INV_X1 U14400 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19211) );
  NOR2_X1 U14401 ( .A1(n19171), .A2(n19211), .ZN(n18166) );
  NOR2_X1 U14402 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19223) );
  INV_X1 U14403 ( .A(n19223), .ZN(n19162) );
  NAND2_X1 U14404 ( .A1(n19222), .A2(n19160), .ZN(n16859) );
  NAND2_X1 U14405 ( .A1(n19162), .A2(n16859), .ZN(n18533) );
  INV_X1 U14406 ( .A(n18533), .ZN(n19205) );
  NAND2_X1 U14407 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18053) );
  NAND2_X1 U14408 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18037), .ZN(
        n18014) );
  NAND2_X1 U14409 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18015) );
  NAND2_X1 U14410 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17976) );
  NAND2_X1 U14411 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17945) );
  NAND2_X1 U14412 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17899) );
  NAND2_X1 U14413 ( .A1(n17882), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17858) );
  NAND2_X1 U14414 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17859) );
  NAND2_X1 U14415 ( .A1(n16735), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11276) );
  INV_X1 U14416 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18202) );
  INV_X1 U14417 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19141) );
  INV_X1 U14418 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19052) );
  NOR2_X1 U14419 ( .A1(n19141), .A2(n18522), .ZN(n12893) );
  INV_X1 U14420 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16718) );
  NOR2_X1 U14421 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19222), .ZN(n17897) );
  NOR2_X1 U14422 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19160), .ZN(
        n19186) );
  AOI221_X1 U14423 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19171), .C1(n19222), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n19186), .ZN(n18544) );
  NOR3_X1 U14424 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19211), .ZN(n18853) );
  OR2_X1 U14425 ( .A1(n11276), .A2(n18052), .ZN(n16717) );
  NOR2_X1 U14426 ( .A1(n16718), .A2(n16717), .ZN(n11282) );
  NOR2_X1 U14427 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17964), .ZN(
        n16733) );
  NOR2_X1 U14428 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16717), .ZN(
        n11280) );
  INV_X1 U14429 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17872) );
  INV_X1 U14430 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16990) );
  NAND3_X1 U14431 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n17975), .ZN(n17017) );
  NAND2_X1 U14432 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16887), .ZN(
        n16886) );
  NAND2_X1 U14433 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17895), .ZN(
        n16888) );
  NAND2_X1 U14434 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17853), .ZN(
        n16893) );
  NOR2_X1 U14435 ( .A1(n17872), .A2(n16893), .ZN(n16892) );
  NAND2_X1 U14436 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16892), .ZN(
        n16884) );
  AOI22_X1 U14437 ( .A1(n17897), .A2(n16884), .B1(n18932), .B2(n11276), .ZN(
        n11279) );
  NAND2_X1 U14438 ( .A1(n11279), .A2(n18207), .ZN(n16734) );
  NOR3_X1 U14439 ( .A1(n16733), .A2(n11280), .A3(n16734), .ZN(n16716) );
  INV_X1 U14440 ( .A(n16716), .ZN(n11281) );
  MUX2_X1 U14441 ( .A(n11282), .B(n11281), .S(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n11283) );
  AOI211_X1 U14442 ( .C1(n17970), .C2(n16885), .A(n12893), .B(n11283), .ZN(
        n11323) );
  NAND2_X1 U14443 ( .A1(n18205), .A2(n11284), .ZN(n11287) );
  NAND2_X1 U14444 ( .A1(n17735), .A2(n11287), .ZN(n11286) );
  NAND2_X1 U14445 ( .A1(n11286), .A2(n17729), .ZN(n11296) );
  NAND2_X1 U14446 ( .A1(n11285), .A2(n17720), .ZN(n11303) );
  NOR2_X1 U14447 ( .A1(n17717), .A2(n11303), .ZN(n11307) );
  NAND2_X1 U14448 ( .A1(n11307), .A2(n16746), .ZN(n11308) );
  XOR2_X1 U14449 ( .A(n11285), .B(n17720), .Z(n11300) );
  XOR2_X1 U14450 ( .A(n11286), .B(n17729), .Z(n11294) );
  AND2_X1 U14451 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11294), .ZN(
        n11295) );
  XOR2_X1 U14452 ( .A(n17735), .B(n11287), .Z(n11288) );
  NOR2_X1 U14453 ( .A1(n11288), .A2(n18508), .ZN(n11293) );
  XNOR2_X1 U14454 ( .A(n18508), .B(n11288), .ZN(n18188) );
  INV_X1 U14455 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19188) );
  NOR2_X1 U14456 ( .A1(n17744), .A2(n19188), .ZN(n11291) );
  INV_X1 U14457 ( .A(n18205), .ZN(n11290) );
  NAND3_X1 U14458 ( .A1(n11290), .A2(n17744), .A3(n19188), .ZN(n11289) );
  OAI221_X1 U14459 ( .B1(n11291), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n11290), .C2(n17744), .A(n11289), .ZN(n18187) );
  NOR2_X1 U14460 ( .A1(n18188), .A2(n18187), .ZN(n11292) );
  NOR2_X1 U14461 ( .A1(n11293), .A2(n11292), .ZN(n18176) );
  XNOR2_X1 U14462 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11294), .ZN(
        n18175) );
  NOR2_X1 U14463 ( .A1(n18176), .A2(n18175), .ZN(n18174) );
  XNOR2_X1 U14464 ( .A(n11296), .B(n17725), .ZN(n11298) );
  NOR2_X1 U14465 ( .A1(n11297), .A2(n11298), .ZN(n11299) );
  INV_X1 U14466 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18480) );
  XNOR2_X1 U14467 ( .A(n11298), .B(n11297), .ZN(n18160) );
  XNOR2_X1 U14468 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11300), .ZN(
        n18146) );
  XOR2_X1 U14469 ( .A(n11303), .B(n11302), .Z(n11305) );
  NOR2_X1 U14470 ( .A1(n11304), .A2(n11305), .ZN(n11306) );
  XNOR2_X1 U14471 ( .A(n11305), .B(n11304), .ZN(n18141) );
  INV_X1 U14472 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18457) );
  XOR2_X1 U14473 ( .A(n11307), .B(n17713), .Z(n11310) );
  NAND2_X1 U14474 ( .A1(n11309), .A2(n11310), .ZN(n18127) );
  INV_X1 U14475 ( .A(n11308), .ZN(n11313) );
  OR2_X1 U14476 ( .A1(n11310), .A2(n11309), .ZN(n18128) );
  OAI21_X1 U14477 ( .B1(n11313), .B2(n11312), .A(n18128), .ZN(n11311) );
  NOR2_X2 U14478 ( .A1(n18404), .A2(n11315), .ZN(n18039) );
  INV_X1 U14479 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18256) );
  NOR2_X1 U14480 ( .A1(n18252), .A2(n18256), .ZN(n18239) );
  INV_X1 U14481 ( .A(n18239), .ZN(n12884) );
  INV_X1 U14482 ( .A(n11319), .ZN(n18215) );
  INV_X1 U14483 ( .A(n16173), .ZN(n11316) );
  NAND2_X1 U14484 ( .A1(n16724), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11317) );
  XNOR2_X1 U14485 ( .A(n11317), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12894) );
  NAND2_X1 U14486 ( .A1(n18335), .A2(n11318), .ZN(n18344) );
  NAND2_X1 U14487 ( .A1(n18239), .A2(n18343), .ZN(n17894) );
  NAND3_X1 U14488 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18220), .A3(
        n16173), .ZN(n11320) );
  XOR2_X1 U14489 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11320), .Z(
        n12897) );
  NOR2_X1 U14490 ( .A1(n12897), .A2(n18058), .ZN(n11321) );
  AOI21_X1 U14491 ( .B1(n12894), .B2(n18196), .A(n11321), .ZN(n11322) );
  AND2_X1 U14492 ( .A1(n11323), .A2(n11322), .ZN(n11324) );
  INV_X1 U14493 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15783) );
  NAND2_X1 U14494 ( .A1(n16435), .A2(n11618), .ZN(n15595) );
  INV_X1 U14495 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11338) );
  OR2_X1 U14496 ( .A1(n11331), .A2(n11330), .ZN(n11332) );
  INV_X1 U14498 ( .A(n11336), .ZN(n11351) );
  INV_X1 U14499 ( .A(n11334), .ZN(n11335) );
  OR2_X1 U14500 ( .A1(n13050), .A2(n9644), .ZN(n11340) );
  NAND2_X1 U14501 ( .A1(n13050), .A2(n11336), .ZN(n11361) );
  INV_X1 U14502 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11337) );
  OAI22_X1 U14503 ( .A1(n11338), .A2(n19709), .B1(n19789), .B2(n11337), .ZN(
        n11343) );
  INV_X1 U14504 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14369) );
  INV_X1 U14505 ( .A(n13271), .ZN(n11339) );
  NAND2_X1 U14506 ( .A1(n9644), .A2(n13162), .ZN(n11365) );
  INV_X1 U14507 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11341) );
  NOR2_X1 U14508 ( .A1(n11343), .A2(n11342), .ZN(n11378) );
  INV_X1 U14509 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11345) );
  NAND3_X1 U14510 ( .A1(n11371), .A2(n13178), .A3(n9675), .ZN(n19823) );
  INV_X1 U14511 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11344) );
  INV_X1 U14512 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11350) );
  BUF_X2 U14513 ( .A(n13271), .Z(n13379) );
  INV_X1 U14514 ( .A(n11361), .ZN(n11347) );
  AND2_X1 U14515 ( .A1(n9675), .A2(n11347), .ZN(n11346) );
  INV_X1 U14516 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11349) );
  OAI22_X1 U14517 ( .A1(n11350), .A2(n19920), .B1(n11447), .B2(n11349), .ZN(
        n11359) );
  INV_X1 U14518 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11357) );
  NAND2_X1 U14519 ( .A1(n11351), .A2(n13050), .ZN(n11364) );
  INV_X1 U14520 ( .A(n11364), .ZN(n11354) );
  AND2_X1 U14521 ( .A1(n9675), .A2(n11354), .ZN(n11353) );
  INV_X1 U14522 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11356) );
  OAI22_X1 U14523 ( .A1(n11357), .A2(n11446), .B1(n11450), .B2(n11356), .ZN(
        n11358) );
  NOR3_X1 U14524 ( .A1(n11360), .A2(n11359), .A3(n11358), .ZN(n11377) );
  INV_X1 U14525 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11362) );
  INV_X1 U14526 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11368) );
  OR2_X2 U14527 ( .A1(n11366), .A2(n11364), .ZN(n13719) );
  OR2_X2 U14528 ( .A1(n11366), .A2(n11365), .ZN(n19758) );
  INV_X1 U14529 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11367) );
  NOR2_X1 U14530 ( .A1(n11370), .A2(n11369), .ZN(n11376) );
  NAND2_X1 U14531 ( .A1(n11371), .A2(n9644), .ZN(n11372) );
  INV_X1 U14532 ( .A(n20009), .ZN(n11373) );
  AOI22_X1 U14533 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n11374), .B1(
        n11373), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11375) );
  NAND4_X1 U14534 ( .A1(n11378), .A2(n11377), .A3(n11376), .A4(n11375), .ZN(
        n11379) );
  NAND2_X1 U14535 ( .A1(n11379), .A2(n16700), .ZN(n11382) );
  INV_X1 U14536 ( .A(n19895), .ZN(n19888) );
  INV_X1 U14537 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11383) );
  INV_X1 U14538 ( .A(n11384), .ZN(n11387) );
  INV_X1 U14539 ( .A(n19920), .ZN(n11385) );
  OAI211_X1 U14540 ( .C1(n19569), .C2(n11388), .A(n11387), .B(n11386), .ZN(
        n11389) );
  AOI21_X1 U14541 ( .B1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n19888), .A(
        n11389), .ZN(n11411) );
  INV_X1 U14542 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11390) );
  OAI22_X1 U14543 ( .A1(n11391), .A2(n13760), .B1(n19758), .B2(n11390), .ZN(
        n11395) );
  INV_X1 U14544 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11393) );
  INV_X1 U14545 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11392) );
  OAI22_X1 U14546 ( .A1(n11393), .A2(n19709), .B1(n19676), .B2(n11392), .ZN(
        n11394) );
  NOR2_X1 U14547 ( .A1(n11395), .A2(n11394), .ZN(n11410) );
  INV_X1 U14548 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11396) );
  INV_X1 U14549 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14150) );
  INV_X1 U14550 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11397) );
  OAI22_X1 U14551 ( .A1(n14150), .A2(n19647), .B1(n19789), .B2(n11397), .ZN(
        n11398) );
  NOR2_X1 U14552 ( .A1(n11399), .A2(n11398), .ZN(n11409) );
  INV_X1 U14553 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11401) );
  INV_X1 U14554 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11400) );
  OAI22_X1 U14555 ( .A1(n11401), .A2(n13719), .B1(n19823), .B2(n11400), .ZN(
        n11407) );
  INV_X1 U14556 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11402) );
  NOR2_X1 U14557 ( .A1(n13858), .A2(n11402), .ZN(n11406) );
  INV_X1 U14558 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11404) );
  INV_X1 U14559 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11403) );
  OAI22_X1 U14560 ( .A1(n11404), .A2(n11450), .B1(n11447), .B2(n11403), .ZN(
        n11405) );
  NOR3_X1 U14561 ( .A1(n11407), .A2(n11406), .A3(n11405), .ZN(n11408) );
  NAND4_X1 U14562 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(
        n11414) );
  NOR2_X1 U14563 ( .A1(n13065), .A2(n11640), .ZN(n11412) );
  NAND2_X1 U14564 ( .A1(n10493), .A2(n11412), .ZN(n11643) );
  NAND2_X1 U14565 ( .A1(n11643), .A2(n11642), .ZN(n11413) );
  OAI21_X1 U14566 ( .B1(n11418), .B2(n11417), .A(n11426), .ZN(n13637) );
  OAI21_X1 U14567 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20239), .A(
        n11419), .ZN(n11678) );
  MUX2_X1 U14568 ( .A(n11678), .B(n13065), .S(n11676), .Z(n11624) );
  INV_X1 U14569 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n19417) );
  MUX2_X1 U14570 ( .A(n11624), .B(n19417), .S(n19597), .Z(n19422) );
  NOR2_X1 U14571 ( .A1(n19422), .A2(n13149), .ZN(n13063) );
  INV_X1 U14572 ( .A(n13063), .ZN(n13071) );
  INV_X1 U14573 ( .A(n11420), .ZN(n11423) );
  NAND3_X1 U14574 ( .A1(n19597), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11421) );
  NAND2_X1 U14575 ( .A1(n11423), .A2(n11421), .ZN(n19404) );
  NOR2_X1 U14576 ( .A1(n13071), .A2(n19404), .ZN(n11422) );
  NAND2_X1 U14577 ( .A1(n13071), .A2(n19404), .ZN(n13070) );
  OAI21_X1 U14578 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11422), .A(
        n13070), .ZN(n14637) );
  XNOR2_X1 U14579 ( .A(n11424), .B(n11423), .ZN(n13898) );
  XNOR2_X1 U14580 ( .A(n13898), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14636) );
  OR2_X1 U14581 ( .A1(n14637), .A2(n14636), .ZN(n14648) );
  NAND2_X1 U14582 ( .A1(n13898), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11425) );
  AND2_X1 U14583 ( .A1(n14648), .A2(n11425), .ZN(n13979) );
  INV_X1 U14584 ( .A(n14026), .ZN(n11428) );
  XNOR2_X1 U14585 ( .A(n11427), .B(n11426), .ZN(n19387) );
  INV_X1 U14586 ( .A(n19387), .ZN(n11429) );
  NAND2_X1 U14587 ( .A1(n11429), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11430) );
  INV_X1 U14588 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11433) );
  INV_X1 U14589 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11432) );
  OAI22_X1 U14590 ( .A1(n11433), .A2(n19676), .B1(n19758), .B2(n11432), .ZN(
        n11437) );
  INV_X1 U14591 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11435) );
  INV_X1 U14592 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11434) );
  OAI22_X1 U14593 ( .A1(n11435), .A2(n13719), .B1(n19789), .B2(n11434), .ZN(
        n11436) );
  NOR2_X1 U14594 ( .A1(n11437), .A2(n11436), .ZN(n11459) );
  INV_X1 U14595 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11439) );
  INV_X1 U14596 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11438) );
  INV_X1 U14597 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11441) );
  INV_X1 U14598 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11440) );
  OAI22_X1 U14599 ( .A1(n11441), .A2(n19709), .B1(n19647), .B2(n11440), .ZN(
        n11443) );
  OAI22_X1 U14600 ( .A1(n14401), .A2(n13760), .B1(n19569), .B2(n13451), .ZN(
        n11442) );
  NOR2_X1 U14601 ( .A1(n11443), .A2(n11442), .ZN(n11457) );
  INV_X1 U14602 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11445) );
  INV_X1 U14603 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11444) );
  OAI22_X1 U14604 ( .A1(n11445), .A2(n13858), .B1(n19823), .B2(n11444), .ZN(
        n11455) );
  INV_X1 U14605 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11449) );
  INV_X1 U14606 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11448) );
  OAI22_X1 U14607 ( .A1(n11449), .A2(n11446), .B1(n11447), .B2(n11448), .ZN(
        n11454) );
  INV_X1 U14608 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11452) );
  INV_X1 U14609 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11451) );
  OAI22_X1 U14610 ( .A1(n11452), .A2(n11450), .B1(n19920), .B2(n11451), .ZN(
        n11453) );
  NOR3_X1 U14611 ( .A1(n11455), .A2(n11454), .A3(n11453), .ZN(n11456) );
  NAND4_X1 U14612 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11463) );
  INV_X1 U14613 ( .A(n11460), .ZN(n11461) );
  NAND2_X1 U14614 ( .A1(n11461), .A2(n10493), .ZN(n11462) );
  OAI21_X1 U14615 ( .B1(n11465), .B2(n11464), .A(n11505), .ZN(n19376) );
  NAND2_X1 U14616 ( .A1(n11466), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11467) );
  INV_X1 U14617 ( .A(n11502), .ZN(n11501) );
  INV_X1 U14618 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11471) );
  INV_X1 U14619 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11470) );
  OAI22_X1 U14620 ( .A1(n11471), .A2(n19676), .B1(n19758), .B2(n11470), .ZN(
        n11475) );
  INV_X1 U14621 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11472) );
  OAI22_X1 U14622 ( .A1(n11473), .A2(n13760), .B1(n13719), .B2(n11472), .ZN(
        n11474) );
  NOR2_X1 U14623 ( .A1(n11475), .A2(n11474), .ZN(n11496) );
  INV_X1 U14624 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11477) );
  INV_X1 U14625 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11476) );
  OAI22_X1 U14626 ( .A1(n11477), .A2(n19895), .B1(n20009), .B2(n11476), .ZN(
        n11478) );
  INV_X1 U14627 ( .A(n11478), .ZN(n11495) );
  INV_X1 U14628 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11480) );
  INV_X1 U14629 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11479) );
  OAI22_X1 U14630 ( .A1(n11480), .A2(n19709), .B1(n19789), .B2(n11479), .ZN(
        n11484) );
  INV_X1 U14631 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11482) );
  OAI22_X1 U14632 ( .A1(n11482), .A2(n19647), .B1(n19569), .B2(n11481), .ZN(
        n11483) );
  NOR2_X1 U14633 ( .A1(n11484), .A2(n11483), .ZN(n11494) );
  INV_X1 U14634 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11486) );
  INV_X1 U14635 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11485) );
  OAI22_X1 U14636 ( .A1(n11486), .A2(n13858), .B1(n19823), .B2(n11485), .ZN(
        n11492) );
  INV_X1 U14637 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11488) );
  INV_X1 U14638 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11487) );
  OAI22_X1 U14639 ( .A1(n11488), .A2(n11450), .B1(n19920), .B2(n11487), .ZN(
        n11491) );
  INV_X1 U14640 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11489) );
  INV_X1 U14641 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14409) );
  OAI22_X1 U14642 ( .A1(n11489), .A2(n11446), .B1(n11447), .B2(n14409), .ZN(
        n11490) );
  NOR3_X1 U14643 ( .A1(n11492), .A2(n11491), .A3(n11490), .ZN(n11493) );
  NAND4_X1 U14644 ( .A1(n11496), .A2(n11495), .A3(n11494), .A4(n11493), .ZN(
        n11499) );
  NAND2_X1 U14645 ( .A1(n11497), .A2(n10493), .ZN(n11498) );
  NAND2_X1 U14646 ( .A1(n11502), .A2(n11656), .ZN(n11503) );
  NAND2_X1 U14647 ( .A1(n11505), .A2(n11504), .ZN(n11506) );
  NAND2_X1 U14648 ( .A1(n11512), .A2(n11506), .ZN(n19365) );
  NAND2_X1 U14649 ( .A1(n11507), .A2(n19365), .ZN(n11508) );
  NAND2_X1 U14650 ( .A1(n11508), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11509) );
  INV_X1 U14651 ( .A(n11510), .ZN(n11511) );
  XNOR2_X1 U14652 ( .A(n11512), .B(n11511), .ZN(n13621) );
  AND2_X1 U14653 ( .A1(n13621), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15721) );
  NAND2_X1 U14654 ( .A1(n19597), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11514) );
  NOR2_X1 U14655 ( .A1(n11515), .A2(n11514), .ZN(n11516) );
  OR2_X1 U14656 ( .A1(n11513), .A2(n11516), .ZN(n13913) );
  NAND2_X1 U14657 ( .A1(n11618), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11664) );
  NOR2_X1 U14658 ( .A1(n13913), .A2(n11664), .ZN(n16565) );
  NAND2_X1 U14659 ( .A1(n19597), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11517) );
  OAI21_X1 U14660 ( .B1(n9749), .B2(n11517), .A(n11602), .ZN(n11518) );
  OR2_X1 U14661 ( .A1(n11527), .A2(n11518), .ZN(n19345) );
  OAI21_X1 U14662 ( .B1(n19345), .B2(n11667), .A(n11519), .ZN(n16551) );
  AND2_X1 U14663 ( .A1(n19597), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11520) );
  XNOR2_X1 U14664 ( .A(n11513), .B(n11520), .ZN(n11525) );
  NAND2_X1 U14665 ( .A1(n11525), .A2(n11618), .ZN(n11521) );
  NAND2_X1 U14666 ( .A1(n11521), .A2(n16032), .ZN(n16019) );
  INV_X1 U14667 ( .A(n13621), .ZN(n11522) );
  NAND2_X1 U14668 ( .A1(n11522), .A2(n16040), .ZN(n16015) );
  OAI21_X1 U14669 ( .B1(n13913), .B2(n11667), .A(n16639), .ZN(n16016) );
  AND4_X1 U14670 ( .A1(n16551), .A2(n16019), .A3(n16015), .A4(n16016), .ZN(
        n11523) );
  NAND2_X1 U14671 ( .A1(n11618), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11524) );
  OR2_X1 U14672 ( .A1(n19345), .A2(n11524), .ZN(n16550) );
  INV_X1 U14673 ( .A(n11525), .ZN(n19354) );
  OR3_X1 U14674 ( .A1(n19354), .A2(n11667), .A3(n16032), .ZN(n16548) );
  NAND2_X1 U14675 ( .A1(n19597), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11526) );
  OR2_X1 U14676 ( .A1(n11527), .A2(n11526), .ZN(n11530) );
  INV_X1 U14677 ( .A(n11528), .ZN(n11529) );
  NAND2_X1 U14678 ( .A1(n11530), .A2(n11529), .ZN(n19334) );
  NOR2_X1 U14679 ( .A1(n19334), .A2(n11667), .ZN(n11560) );
  AND2_X1 U14680 ( .A1(n11560), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15998) );
  INV_X1 U14681 ( .A(n11531), .ZN(n11533) );
  NAND2_X1 U14682 ( .A1(n11533), .A2(n11532), .ZN(n11534) );
  NAND2_X1 U14683 ( .A1(n11556), .A2(n11534), .ZN(n13885) );
  OR3_X1 U14684 ( .A1(n13885), .A2(n11667), .A3(n16528), .ZN(n16521) );
  INV_X1 U14685 ( .A(n16521), .ZN(n11535) );
  NAND3_X1 U14686 ( .A1(n11539), .A2(n19597), .A3(P2_EBX_REG_21__SCAN_IN), 
        .ZN(n11536) );
  OAI211_X1 U14687 ( .C1(n11539), .C2(P2_EBX_REG_21__SCAN_IN), .A(n11536), .B(
        n11602), .ZN(n12929) );
  INV_X1 U14688 ( .A(n11576), .ZN(n11537) );
  NAND2_X1 U14689 ( .A1(n19597), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11538) );
  MUX2_X1 U14690 ( .A(n19597), .B(n11538), .S(n11544), .Z(n11540) );
  NAND2_X1 U14691 ( .A1(n11540), .A2(n11539), .ZN(n19264) );
  NOR2_X1 U14692 ( .A1(n19264), .A2(n11667), .ZN(n11586) );
  INV_X1 U14693 ( .A(n11586), .ZN(n11541) );
  INV_X1 U14694 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15902) );
  AND2_X1 U14695 ( .A1(n11541), .A2(n15902), .ZN(n15659) );
  NAND2_X1 U14696 ( .A1(n11548), .A2(n11542), .ZN(n11543) );
  NAND2_X1 U14697 ( .A1(n11544), .A2(n11543), .ZN(n19272) );
  INV_X1 U14698 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15899) );
  NAND2_X1 U14699 ( .A1(n11545), .A2(n15899), .ZN(n15682) );
  NAND2_X1 U14700 ( .A1(n11571), .A2(n11546), .ZN(n11547) );
  NAND2_X1 U14701 ( .A1(n11548), .A2(n11547), .ZN(n15390) );
  OR2_X1 U14702 ( .A1(n15390), .A2(n11667), .ZN(n11577) );
  NAND2_X1 U14703 ( .A1(n11577), .A2(n15934), .ZN(n15683) );
  NAND2_X1 U14704 ( .A1(n15682), .A2(n15683), .ZN(n15658) );
  NAND2_X1 U14705 ( .A1(n19597), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11550) );
  OAI211_X1 U14706 ( .C1(n11552), .C2(n11550), .A(n11602), .B(n11549), .ZN(
        n19296) );
  OR2_X1 U14707 ( .A1(n19296), .A2(n11667), .ZN(n11551) );
  INV_X1 U14708 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15958) );
  XNOR2_X1 U14709 ( .A(n11551), .B(n15958), .ZN(n15713) );
  INV_X1 U14710 ( .A(n15713), .ZN(n11574) );
  INV_X1 U14711 ( .A(n11552), .ZN(n11554) );
  OR2_X1 U14712 ( .A1(n11562), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11564) );
  NAND3_X1 U14713 ( .A1(n11564), .A2(n19597), .A3(P2_EBX_REG_15__SCAN_IN), 
        .ZN(n11553) );
  AND2_X1 U14714 ( .A1(n11554), .A2(n11553), .ZN(n11578) );
  NAND2_X1 U14715 ( .A1(n11578), .A2(n11618), .ZN(n11555) );
  NAND2_X1 U14716 ( .A1(n11555), .A2(n15977), .ZN(n15962) );
  XNOR2_X1 U14717 ( .A(n11556), .B(n9760), .ZN(n19321) );
  AND2_X1 U14718 ( .A1(n19321), .A2(n11618), .ZN(n11581) );
  INV_X1 U14719 ( .A(n11581), .ZN(n11558) );
  NAND2_X1 U14720 ( .A1(n11558), .A2(n11557), .ZN(n15982) );
  OR2_X1 U14721 ( .A1(n13885), .A2(n11667), .ZN(n11559) );
  NAND2_X1 U14722 ( .A1(n11559), .A2(n16528), .ZN(n16522) );
  INV_X1 U14723 ( .A(n11560), .ZN(n11561) );
  NAND2_X1 U14724 ( .A1(n11561), .A2(n16003), .ZN(n15997) );
  NAND4_X1 U14725 ( .A1(n15962), .A2(n15982), .A3(n16522), .A4(n15997), .ZN(
        n11567) );
  NAND2_X1 U14726 ( .A1(n19597), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11563) );
  MUX2_X1 U14727 ( .A(n19597), .B(n11563), .S(n11562), .Z(n11565) );
  AND2_X1 U14728 ( .A1(n11565), .A2(n11564), .ZN(n14040) );
  AND2_X1 U14729 ( .A1(n14040), .A2(n11618), .ZN(n11580) );
  INV_X1 U14730 ( .A(n11580), .ZN(n11566) );
  NOR2_X1 U14731 ( .A1(n11567), .A2(n16504), .ZN(n11573) );
  OR2_X1 U14732 ( .A1(n11569), .A2(n11568), .ZN(n11570) );
  NAND2_X1 U14733 ( .A1(n11571), .A2(n11570), .ZN(n19281) );
  OR2_X1 U14734 ( .A1(n19281), .A2(n11667), .ZN(n11572) );
  INV_X1 U14735 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15947) );
  NAND2_X1 U14736 ( .A1(n11572), .A2(n15947), .ZN(n15656) );
  NAND3_X1 U14737 ( .A1(n11574), .A2(n11573), .A3(n15656), .ZN(n11575) );
  NAND2_X1 U14738 ( .A1(n11576), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15652) );
  NOR2_X1 U14739 ( .A1(n11577), .A2(n15934), .ZN(n15690) );
  INV_X1 U14740 ( .A(n11578), .ZN(n19308) );
  NAND2_X1 U14741 ( .A1(n11618), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11579) );
  NOR2_X1 U14742 ( .A1(n19308), .A2(n11579), .ZN(n15963) );
  NOR2_X1 U14743 ( .A1(n15654), .A2(n15963), .ZN(n11582) );
  OR3_X1 U14744 ( .A1(n19281), .A2(n11667), .A3(n15947), .ZN(n15655) );
  NAND2_X1 U14745 ( .A1(n11580), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16503) );
  AND2_X1 U14746 ( .A1(n11581), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15653) );
  INV_X1 U14747 ( .A(n15653), .ZN(n15983) );
  NAND4_X1 U14748 ( .A1(n11582), .A2(n15655), .A3(n16503), .A4(n15983), .ZN(
        n11583) );
  NOR2_X1 U14749 ( .A1(n15690), .A2(n11583), .ZN(n11585) );
  NAND2_X1 U14750 ( .A1(n11618), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11584) );
  OR2_X1 U14751 ( .A1(n19272), .A2(n11584), .ZN(n15681) );
  NAND3_X1 U14752 ( .A1(n15652), .A2(n11585), .A3(n15681), .ZN(n11587) );
  AND2_X1 U14753 ( .A1(n11586), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15660) );
  NOR2_X1 U14754 ( .A1(n11587), .A2(n15660), .ZN(n11588) );
  INV_X1 U14755 ( .A(n11589), .ZN(n11590) );
  NAND2_X1 U14756 ( .A1(n11590), .A2(n9713), .ZN(n11591) );
  NAND2_X1 U14757 ( .A1(n11594), .A2(n11591), .ZN(n12946) );
  OR2_X1 U14758 ( .A1(n12946), .A2(n11667), .ZN(n11592) );
  NAND2_X1 U14759 ( .A1(n11594), .A2(n11593), .ZN(n11595) );
  OR2_X1 U14760 ( .A1(n12957), .A2(n11667), .ZN(n11596) );
  XNOR2_X1 U14761 ( .A(n11596), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15642) );
  INV_X1 U14762 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15855) );
  INV_X1 U14763 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15819) );
  NAND2_X1 U14764 ( .A1(n19597), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11598) );
  MUX2_X1 U14765 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n11598), .S(n11597), .Z(
        n11599) );
  NAND2_X1 U14766 ( .A1(n11599), .A2(n11602), .ZN(n16465) );
  NOR2_X1 U14767 ( .A1(n16465), .A2(n11667), .ZN(n15634) );
  NAND2_X1 U14768 ( .A1(n19597), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11601) );
  AND2_X1 U14769 ( .A1(n11603), .A2(n11602), .ZN(n11607) );
  AOI21_X1 U14770 ( .B1(n11607), .B2(n11618), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15623) );
  INV_X1 U14771 ( .A(n11604), .ZN(n16453) );
  AOI21_X1 U14772 ( .B1(n11605), .B2(n16435), .A(n11612), .ZN(n16427) );
  NAND2_X1 U14773 ( .A1(n16427), .A2(n11618), .ZN(n15597) );
  INV_X1 U14774 ( .A(n11606), .ZN(n11608) );
  NOR3_X1 U14775 ( .A1(n15376), .A2(n11667), .A3(n15840), .ZN(n15624) );
  AOI21_X1 U14776 ( .B1(n11608), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15624), .ZN(n15592) );
  NAND2_X1 U14777 ( .A1(n11609), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11610) );
  XNOR2_X1 U14778 ( .A(n11612), .B(n11611), .ZN(n11617) );
  OAI21_X1 U14779 ( .B1(n11617), .B2(n11667), .A(n15787), .ZN(n15580) );
  INV_X1 U14780 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11613) );
  NOR2_X1 U14781 ( .A1(n10792), .A2(n11613), .ZN(n11614) );
  XNOR2_X1 U14782 ( .A(n11615), .B(n11614), .ZN(n12838) );
  INV_X1 U14783 ( .A(n12838), .ZN(n11616) );
  AOI21_X1 U14784 ( .B1(n11616), .B2(n11618), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15569) );
  INV_X1 U14785 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15764) );
  INV_X1 U14786 ( .A(n11617), .ZN(n15359) );
  NAND3_X1 U14787 ( .A1(n15359), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11618), .ZN(n15581) );
  NOR2_X1 U14788 ( .A1(n11619), .A2(n11667), .ZN(n11620) );
  XOR2_X1 U14789 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11620), .Z(
        n11621) );
  INV_X1 U14790 ( .A(n11622), .ZN(n11623) );
  OAI21_X1 U14791 ( .B1(n11624), .B2(n11677), .A(n11623), .ZN(n11627) );
  INV_X1 U14792 ( .A(n11690), .ZN(n11625) );
  AOI21_X1 U14793 ( .B1(n11627), .B2(n11626), .A(n11625), .ZN(n20249) );
  AND2_X1 U14794 ( .A1(n10493), .A2(n10468), .ZN(n13030) );
  INV_X1 U14795 ( .A(n13030), .ZN(n11628) );
  NOR2_X1 U14796 ( .A1(n16662), .A2(n11628), .ZN(n20241) );
  NAND2_X1 U14797 ( .A1(n20249), .A2(n20241), .ZN(n11636) );
  INV_X1 U14798 ( .A(n16662), .ZN(n11634) );
  OAI21_X1 U14799 ( .B1(n11678), .B2(n11629), .A(n16672), .ZN(n11630) );
  INV_X1 U14800 ( .A(n11630), .ZN(n11633) );
  NAND2_X1 U14801 ( .A1(n16675), .A2(n11631), .ZN(n16658) );
  INV_X1 U14802 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11632) );
  OAI21_X1 U14803 ( .B1(n9643), .B2(n16658), .A(n11632), .ZN(n20230) );
  MUX2_X1 U14804 ( .A(n11633), .B(n20230), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20243) );
  NAND3_X1 U14805 ( .A1(n11634), .A2(n16700), .A3(n20243), .ZN(n11635) );
  NAND2_X1 U14806 ( .A1(n11636), .A2(n11635), .ZN(n13127) );
  AND2_X1 U14807 ( .A1(n10468), .A2(n13332), .ZN(n11637) );
  NAND2_X1 U14808 ( .A1(n13127), .A2(n11637), .ZN(n19239) );
  NAND2_X1 U14809 ( .A1(n13065), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13064) );
  INV_X1 U14810 ( .A(n13064), .ZN(n11638) );
  NAND2_X1 U14811 ( .A1(n11638), .A2(n11001), .ZN(n11641) );
  AND2_X1 U14812 ( .A1(n13149), .A2(n13065), .ZN(n11639) );
  XOR2_X1 U14813 ( .A(n11640), .B(n11639), .Z(n13074) );
  NAND2_X1 U14814 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13074), .ZN(
        n13073) );
  NAND2_X1 U14815 ( .A1(n11641), .A2(n13073), .ZN(n11644) );
  XOR2_X1 U14816 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11644), .Z(
        n14633) );
  XNOR2_X1 U14817 ( .A(n11643), .B(n11642), .ZN(n14631) );
  NAND2_X1 U14818 ( .A1(n14633), .A2(n14631), .ZN(n11646) );
  NAND2_X1 U14819 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11644), .ZN(
        n11645) );
  NAND2_X1 U14820 ( .A1(n11646), .A2(n11645), .ZN(n11647) );
  XNOR2_X1 U14821 ( .A(n11647), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13982) );
  INV_X1 U14822 ( .A(n11647), .ZN(n11648) );
  XNOR2_X1 U14823 ( .A(n11650), .B(n11649), .ZN(n11652) );
  NAND2_X1 U14824 ( .A1(n11651), .A2(n11652), .ZN(n14023) );
  NAND2_X1 U14825 ( .A1(n14023), .A2(n14127), .ZN(n11653) );
  NAND2_X1 U14826 ( .A1(n11657), .A2(n14137), .ZN(n11658) );
  XNOR2_X1 U14827 ( .A(n11660), .B(n11667), .ZN(n15724) );
  INV_X1 U14828 ( .A(n11660), .ZN(n11666) );
  INV_X1 U14829 ( .A(n11664), .ZN(n11665) );
  OAI21_X1 U14830 ( .B1(n11660), .B2(n11667), .A(n16639), .ZN(n11668) );
  NAND2_X1 U14831 ( .A1(n11670), .A2(n11668), .ZN(n16569) );
  NAND2_X1 U14832 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16001) );
  NOR2_X1 U14833 ( .A1(n16032), .A2(n16001), .ZN(n16610) );
  AND3_X1 U14834 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n16610), .ZN(n16594) );
  NAND2_X1 U14835 ( .A1(n16594), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15709) );
  AND2_X1 U14836 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15928) );
  NAND2_X1 U14837 ( .A1(n15928), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11671) );
  NOR2_X1 U14838 ( .A1(n15709), .A2(n11671), .ZN(n15693) );
  AND2_X1 U14839 ( .A1(n15693), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15903) );
  NAND2_X2 U14840 ( .A1(n16024), .A2(n15903), .ZN(n15694) );
  NAND3_X1 U14841 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15763) );
  XOR2_X1 U14842 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11672), .Z(
        n15758) );
  NOR2_X2 U14843 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20196) );
  NAND2_X1 U14844 ( .A1(n11673), .A2(n16659), .ZN(n11681) );
  NAND2_X1 U14845 ( .A1(n10493), .A2(n11678), .ZN(n11675) );
  NAND3_X1 U14846 ( .A1(n11675), .A2(n16663), .A3(n11674), .ZN(n11680) );
  OAI21_X1 U14847 ( .B1(n11678), .B2(n11677), .A(n11676), .ZN(n11679) );
  NAND3_X1 U14848 ( .A1(n11681), .A2(n11680), .A3(n11679), .ZN(n11682) );
  NAND2_X1 U14849 ( .A1(n20256), .A2(n16675), .ZN(n11689) );
  OAI21_X1 U14850 ( .B1(n11690), .B2(n20263), .A(n11689), .ZN(n11691) );
  INV_X1 U14851 ( .A(n11691), .ZN(n11692) );
  NAND2_X1 U14852 ( .A1(n10598), .A2(n19761), .ZN(n16196) );
  NAND2_X1 U14853 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n20231) );
  AND2_X1 U14854 ( .A1(n16196), .A2(n20231), .ZN(n11693) );
  INV_X1 U14855 ( .A(n19559), .ZN(n16589) );
  OR2_X1 U14856 ( .A1(n20196), .A2(n20198), .ZN(n20220) );
  NAND2_X1 U14857 ( .A1(n20220), .A2(n20256), .ZN(n11695) );
  AND2_X1 U14858 ( .A1(n20256), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13270) );
  INV_X1 U14859 ( .A(n13270), .ZN(n11697) );
  INV_X1 U14860 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19820) );
  NAND2_X1 U14861 ( .A1(n19820), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U14862 ( .A1(n11697), .A2(n11696), .ZN(n13067) );
  NOR2_X1 U14863 ( .A1(n19364), .A2(n11698), .ZN(n15748) );
  AOI21_X1 U14864 ( .B1(n19551), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15748), .ZN(n11699) );
  OAI21_X1 U14865 ( .B1(n19564), .B2(n11700), .A(n11699), .ZN(n11701) );
  INV_X1 U14866 ( .A(n11701), .ZN(n11702) );
  OAI21_X1 U14867 ( .B1(n15762), .B2(n16586), .A(n11706), .ZN(P2_U2983) );
  NAND2_X1 U14868 ( .A1(n11768), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11710) );
  NAND2_X1 U14869 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11709) );
  NAND2_X1 U14870 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11708) );
  NAND2_X1 U14871 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11707) );
  NAND4_X1 U14872 ( .A1(n11710), .A2(n11709), .A3(n11708), .A4(n11707), .ZN(
        n11713) );
  INV_X1 U14873 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11711) );
  NOR2_X1 U14874 ( .A1(n11798), .A2(n11711), .ZN(n11712) );
  NAND2_X1 U14875 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11717) );
  NAND2_X1 U14876 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11716) );
  NAND2_X1 U14877 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11715) );
  AND2_X2 U14878 ( .A1(n13584), .A2(n11719), .ZN(n12429) );
  NAND2_X1 U14879 ( .A1(n12429), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11714) );
  NAND2_X1 U14880 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11723) );
  NAND2_X1 U14881 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11722) );
  NAND2_X1 U14882 ( .A1(n12648), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U14883 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11720) );
  INV_X1 U14884 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U14885 ( .A1(n12586), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11728) );
  INV_X2 U14886 ( .A(n12637), .ZN(n12585) );
  NAND2_X1 U14887 ( .A1(n12615), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11727) );
  OAI211_X1 U14888 ( .C1(n12578), .C2(n11729), .A(n11728), .B(n11727), .ZN(
        n11730) );
  INV_X1 U14889 ( .A(n11730), .ZN(n11731) );
  NAND2_X1 U14890 ( .A1(n12648), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11743) );
  NAND2_X1 U14891 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11742) );
  INV_X1 U14892 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11735) );
  NOR2_X1 U14893 ( .A1(n11798), .A2(n11735), .ZN(n11740) );
  NAND2_X1 U14894 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11738) );
  INV_X1 U14895 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11736) );
  NOR2_X1 U14896 ( .A1(n11740), .A2(n11739), .ZN(n11741) );
  INV_X1 U14897 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U14898 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11746) );
  NAND2_X1 U14899 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11745) );
  OAI211_X1 U14900 ( .C1(n12647), .C2(n11747), .A(n11746), .B(n11745), .ZN(
        n11758) );
  NAND2_X1 U14901 ( .A1(n11768), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11751) );
  NAND2_X1 U14902 ( .A1(n12616), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11750) );
  NAND2_X1 U14903 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U14904 ( .A1(n12429), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U14905 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11755) );
  NAND2_X1 U14906 ( .A1(n12615), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11754) );
  NAND2_X1 U14907 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11753) );
  NAND2_X1 U14908 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11752) );
  INV_X1 U14909 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U14910 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11761) );
  NAND2_X1 U14911 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11760) );
  OAI211_X1 U14912 ( .C1(n12578), .C2(n11762), .A(n11761), .B(n11760), .ZN(
        n11763) );
  INV_X1 U14913 ( .A(n11763), .ZN(n11767) );
  INV_X2 U14914 ( .A(n11822), .ZN(n12614) );
  AOI22_X1 U14915 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14916 ( .A1(n12648), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11765) );
  NAND2_X1 U14917 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11764) );
  NAND4_X1 U14918 ( .A1(n11767), .A2(n11766), .A3(n11765), .A4(n11764), .ZN(
        n11775) );
  INV_X1 U14919 ( .A(n11768), .ZN(n12605) );
  AOI22_X1 U14920 ( .A1(n11768), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11773) );
  INV_X2 U14921 ( .A(n12639), .ZN(n12411) );
  AOI22_X1 U14922 ( .A1(n12586), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11772) );
  INV_X2 U14923 ( .A(n12603), .ZN(n12642) );
  AOI22_X1 U14924 ( .A1(n9657), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14925 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11770) );
  NAND4_X1 U14926 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n11774) );
  INV_X1 U14927 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12604) );
  NAND2_X1 U14928 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U14929 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11777) );
  OAI211_X1 U14930 ( .C1(n12647), .C2(n12604), .A(n11778), .B(n11777), .ZN(
        n11779) );
  INV_X1 U14931 ( .A(n11779), .ZN(n11783) );
  AOI22_X1 U14932 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14933 ( .A1(n12648), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11781) );
  NAND2_X1 U14934 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11780) );
  NAND4_X1 U14935 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11789) );
  AOI22_X1 U14936 ( .A1(n12586), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14937 ( .A1(n11768), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14938 ( .A1(n9657), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14939 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U14940 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11788) );
  NAND2_X1 U14941 ( .A1(n14265), .A2(n13967), .ZN(n11790) );
  INV_X1 U14942 ( .A(n11834), .ZN(n11900) );
  NAND2_X1 U14943 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11796) );
  NAND2_X1 U14944 ( .A1(n12615), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11795) );
  NAND2_X1 U14945 ( .A1(n9657), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11794) );
  NAND2_X1 U14946 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11793) );
  NAND4_X1 U14947 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11800) );
  INV_X1 U14948 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11797) );
  NOR2_X1 U14949 ( .A1(n11798), .A2(n11797), .ZN(n11799) );
  NOR2_X1 U14950 ( .A1(n11800), .A2(n11799), .ZN(n11816) );
  NAND2_X1 U14951 ( .A1(n11768), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11804) );
  NAND2_X1 U14952 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11803) );
  NAND2_X1 U14953 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11802) );
  NAND2_X1 U14954 ( .A1(n12429), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11801) );
  NAND2_X1 U14955 ( .A1(n12648), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U14956 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11807) );
  NAND2_X1 U14957 ( .A1(n12586), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11806) );
  NAND2_X1 U14958 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11805) );
  INV_X1 U14959 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U14960 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U14961 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11809) );
  OAI211_X1 U14962 ( .C1(n12647), .C2(n11811), .A(n11810), .B(n11809), .ZN(
        n11812) );
  INV_X1 U14963 ( .A(n11812), .ZN(n11813) );
  NAND2_X1 U14964 ( .A1(n11817), .A2(n11833), .ZN(n11882) );
  INV_X1 U14965 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11820) );
  NAND2_X1 U14966 ( .A1(n11768), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U14967 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11818) );
  OAI211_X1 U14968 ( .C1(n12647), .C2(n11820), .A(n11819), .B(n11818), .ZN(
        n11821) );
  INV_X1 U14969 ( .A(n11821), .ZN(n11826) );
  AOI22_X1 U14970 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12648), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14971 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U14972 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11823) );
  NAND4_X1 U14973 ( .A1(n11826), .A2(n11825), .A3(n11824), .A4(n11823), .ZN(
        n11832) );
  AOI22_X1 U14974 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11776), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14975 ( .A1(n12586), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14976 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14977 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11827) );
  NAND4_X1 U14978 ( .A1(n11830), .A2(n11829), .A3(n11828), .A4(n11827), .ZN(
        n11831) );
  NAND2_X1 U14979 ( .A1(n11882), .A2(n13954), .ZN(n11836) );
  NAND2_X1 U14980 ( .A1(n11875), .A2(n14267), .ZN(n11835) );
  NAND2_X1 U14981 ( .A1(n12648), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11841) );
  NAND2_X1 U14982 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11840) );
  NAND2_X1 U14983 ( .A1(n12615), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11839) );
  NAND2_X1 U14984 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11838) );
  AOI22_X1 U14985 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11845) );
  NAND2_X1 U14986 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11844) );
  NAND2_X1 U14987 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11843) );
  AOI22_X1 U14988 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11768), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U14989 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11776), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14990 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14991 ( .A1(n12586), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11848) );
  NOR2_X1 U14992 ( .A1(n12780), .A2(n13499), .ZN(n11853) );
  NAND2_X1 U14993 ( .A1(n12648), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11857) );
  NAND2_X1 U14994 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U14995 ( .A1(n12615), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U14996 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11854) );
  NAND4_X1 U14997 ( .A1(n11857), .A2(n11856), .A3(n11855), .A4(n11854), .ZN(
        n11859) );
  INV_X1 U14998 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11858) );
  NAND2_X1 U14999 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11863) );
  NAND2_X1 U15000 ( .A1(n12429), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11862) );
  NAND2_X1 U15001 ( .A1(n11768), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11861) );
  NAND2_X1 U15002 ( .A1(n11769), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11867) );
  NAND2_X1 U15003 ( .A1(n12616), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11866) );
  NAND2_X1 U15004 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11865) );
  NAND2_X1 U15005 ( .A1(n11776), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U15006 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11871) );
  NAND2_X1 U15007 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11870) );
  NAND2_X1 U15008 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11869) );
  NAND2_X1 U15009 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11868) );
  NAND2_X2 U15010 ( .A1(n11880), .A2(n11875), .ZN(n13521) );
  INV_X1 U15011 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n11877) );
  XNOR2_X1 U15012 ( .A(n11877), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n13207) );
  INV_X1 U15013 ( .A(n14265), .ZN(n13871) );
  NAND2_X2 U15014 ( .A1(n11879), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11910) );
  INV_X1 U15015 ( .A(n11880), .ZN(n13438) );
  AOI21_X1 U15016 ( .B1(n13871), .B2(n13967), .A(n13514), .ZN(n11881) );
  NAND2_X1 U15017 ( .A1(n13438), .A2(n11881), .ZN(n13305) );
  NAND2_X1 U15018 ( .A1(n13305), .A2(n15302), .ZN(n11886) );
  INV_X1 U15019 ( .A(n13954), .ZN(n11883) );
  NAND2_X4 U15020 ( .A1(n11883), .A2(n13499), .ZN(n14318) );
  INV_X1 U15021 ( .A(n13209), .ZN(n13211) );
  NAND2_X1 U15022 ( .A1(n14656), .A2(n13211), .ZN(n13348) );
  INV_X4 U15023 ( .A(n14093), .ZN(n14322) );
  NAND2_X1 U15024 ( .A1(n13344), .A2(n14322), .ZN(n11884) );
  NAND2_X1 U15025 ( .A1(n13499), .A2(n13308), .ZN(n13520) );
  NAND2_X1 U15026 ( .A1(n21043), .A2(n13514), .ZN(n11885) );
  NAND4_X1 U15027 ( .A1(n11886), .A2(n13348), .A3(n13349), .A4(n11885), .ZN(
        n11891) );
  INV_X1 U15028 ( .A(n12008), .ZN(n11890) );
  INV_X1 U15029 ( .A(n13870), .ZN(n11888) );
  NAND3_X1 U15030 ( .A1(n11887), .A2(n13498), .A3(n11888), .ZN(n11889) );
  NAND2_X1 U15031 ( .A1(n11911), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11895) );
  NOR2_X1 U15032 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13367) );
  NAND2_X1 U15033 ( .A1(n13367), .A2(n21045), .ZN(n12812) );
  NAND2_X1 U15034 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11915) );
  OAI21_X1 U15035 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11915), .ZN(n20753) );
  NAND2_X1 U15036 ( .A1(n16420), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20944) );
  NAND2_X1 U15037 ( .A1(n20944), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11908) );
  OAI21_X1 U15038 ( .B1(n12812), .B2(n20753), .A(n11908), .ZN(n11893) );
  INV_X1 U15039 ( .A(n11893), .ZN(n11894) );
  NAND2_X1 U15040 ( .A1(n11895), .A2(n11894), .ZN(n11896) );
  XNOR2_X2 U15041 ( .A(n11896), .B(n11910), .ZN(n20547) );
  NAND2_X1 U15042 ( .A1(n11911), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11898) );
  INV_X1 U15043 ( .A(n20944), .ZN(n16149) );
  MUX2_X1 U15044 ( .A(n16149), .B(n12812), .S(n20721), .Z(n11897) );
  INV_X1 U15045 ( .A(n11887), .ZN(n11899) );
  NAND2_X1 U15046 ( .A1(n13870), .A2(n11900), .ZN(n11901) );
  INV_X1 U15047 ( .A(n15302), .ZN(n13214) );
  NAND2_X1 U15048 ( .A1(n13214), .A2(n13958), .ZN(n13506) );
  NAND3_X1 U15049 ( .A1(n13506), .A2(n13212), .A3(n13305), .ZN(n11906) );
  INV_X1 U15050 ( .A(n13349), .ZN(n11904) );
  NAND2_X1 U15051 ( .A1(n13367), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20279) );
  INV_X1 U15052 ( .A(n20279), .ZN(n11902) );
  NAND2_X1 U15053 ( .A1(n14002), .A2(n13958), .ZN(n13676) );
  NAND3_X1 U15054 ( .A1(n14318), .A2(n11902), .A3(n13676), .ZN(n11903) );
  NOR2_X1 U15055 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  AND2_X1 U15056 ( .A1(n11908), .A2(n13361), .ZN(n11909) );
  NAND2_X1 U15057 ( .A1(n12002), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11913) );
  NAND2_X1 U15058 ( .A1(n20944), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11912) );
  INV_X1 U15059 ( .A(n12812), .ZN(n12004) );
  INV_X1 U15060 ( .A(n11915), .ZN(n11914) );
  INV_X1 U15061 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12762) );
  NAND2_X1 U15062 ( .A1(n11914), .A2(n12762), .ZN(n20795) );
  NAND2_X1 U15063 ( .A1(n11915), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11916) );
  NAND2_X1 U15064 ( .A1(n20795), .A2(n11916), .ZN(n15325) );
  NAND4_X1 U15065 ( .A1(n11994), .A2(n9690), .A3(n11917), .A4(n9770), .ZN(
        n11918) );
  NAND2_X1 U15066 ( .A1(n12001), .A2(n11918), .ZN(n13569) );
  INV_X1 U15067 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12490) );
  NAND2_X1 U15068 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U15069 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11919) );
  OAI211_X1 U15070 ( .C1(n12578), .C2(n12490), .A(n11920), .B(n11919), .ZN(
        n11921) );
  INV_X1 U15071 ( .A(n11921), .ZN(n11925) );
  AOI22_X1 U15072 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15073 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11923) );
  NAND2_X1 U15074 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11922) );
  NAND4_X1 U15075 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11931) );
  AOI22_X1 U15076 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15077 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U15078 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U15079 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11926) );
  NAND4_X1 U15080 ( .A1(n11929), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n11930) );
  NOR2_X1 U15081 ( .A1(n11931), .A2(n11930), .ZN(n12687) );
  NAND2_X1 U15082 ( .A1(n12788), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11933) );
  OAI21_X1 U15083 ( .B1(n12687), .B2(n12008), .A(n11933), .ZN(n11934) );
  NAND2_X1 U15084 ( .A1(n12115), .A2(n21045), .ZN(n11967) );
  INV_X1 U15085 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12438) );
  NAND2_X1 U15086 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11940) );
  NAND2_X1 U15087 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11939) );
  OAI211_X1 U15088 ( .C1(n12647), .C2(n12438), .A(n11940), .B(n11939), .ZN(
        n11941) );
  INV_X1 U15089 ( .A(n11941), .ZN(n11945) );
  AOI22_X1 U15090 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U15091 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11943) );
  NAND2_X1 U15092 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11942) );
  NAND4_X1 U15093 ( .A1(n11945), .A2(n11944), .A3(n11943), .A4(n11942), .ZN(
        n11951) );
  AOI22_X1 U15094 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12411), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15095 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15096 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U15097 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11946) );
  NAND4_X1 U15098 ( .A1(n11949), .A2(n11948), .A3(n11947), .A4(n11946), .ZN(
        n11950) );
  INV_X1 U15099 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11954) );
  NAND2_X1 U15100 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11953) );
  NAND2_X1 U15101 ( .A1(n12403), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11952) );
  OAI211_X1 U15102 ( .C1(n12647), .C2(n11954), .A(n11953), .B(n11952), .ZN(
        n11955) );
  INV_X1 U15103 ( .A(n11955), .ZN(n11959) );
  AOI22_X1 U15104 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U15105 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11957) );
  NAND2_X1 U15106 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11956) );
  NAND4_X1 U15107 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11965) );
  AOI22_X1 U15108 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12649), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15109 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15110 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15111 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11960) );
  NAND4_X1 U15112 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11964) );
  XNOR2_X1 U15113 ( .A(n12674), .B(n12735), .ZN(n11966) );
  INV_X1 U15114 ( .A(n12007), .ZN(n12669) );
  NAND2_X1 U15115 ( .A1(n11966), .A2(n12669), .ZN(n12114) );
  NAND2_X1 U15116 ( .A1(n11967), .A2(n12114), .ZN(n12113) );
  NAND2_X1 U15117 ( .A1(n13514), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11968) );
  MUX2_X1 U15118 ( .A(n11968), .B(n12674), .S(n14002), .Z(n11970) );
  AOI21_X1 U15119 ( .B1(n15338), .B2(n12735), .A(n21045), .ZN(n11969) );
  NAND2_X1 U15120 ( .A1(n11970), .A2(n11969), .ZN(n12112) );
  NAND2_X1 U15121 ( .A1(n12113), .A2(n12112), .ZN(n11972) );
  NAND2_X1 U15122 ( .A1(n12669), .A2(n12735), .ZN(n11971) );
  NAND2_X1 U15123 ( .A1(n12788), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11990) );
  INV_X1 U15124 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11975) );
  NAND2_X1 U15125 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11974) );
  NAND2_X1 U15126 ( .A1(n12403), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11973) );
  OAI211_X1 U15127 ( .C1(n12578), .C2(n11975), .A(n11974), .B(n11973), .ZN(
        n11976) );
  INV_X1 U15128 ( .A(n11976), .ZN(n11980) );
  AOI22_X1 U15129 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15130 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U15131 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11977) );
  NAND4_X1 U15132 ( .A1(n11980), .A2(n11979), .A3(n11978), .A4(n11977), .ZN(
        n11986) );
  AOI22_X1 U15133 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12651), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15134 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12411), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15135 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15136 ( .A1(n12616), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11981) );
  NAND4_X1 U15137 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n11985) );
  INV_X1 U15138 ( .A(n12684), .ZN(n11987) );
  OAI22_X1 U15139 ( .A1(n12008), .A2(n11987), .B1(n12007), .B2(n12735), .ZN(
        n11988) );
  INV_X1 U15140 ( .A(n11988), .ZN(n11989) );
  INV_X1 U15141 ( .A(n20547), .ZN(n11993) );
  INV_X1 U15142 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U15143 ( .A1(n11994), .A2(n13944), .ZN(n15296) );
  NAND2_X1 U15144 ( .A1(n12105), .A2(n12673), .ZN(n12000) );
  INV_X1 U15145 ( .A(n11996), .ZN(n11997) );
  NAND2_X1 U15146 ( .A1(n12000), .A2(n11999), .ZN(n12097) );
  NAND2_X1 U15147 ( .A1(n12002), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12006) );
  NOR3_X1 U15148 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12762), .A3(
        n20692), .ZN(n20669) );
  NAND2_X1 U15149 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20669), .ZN(
        n20662) );
  NAND2_X1 U15150 ( .A1(n21034), .A2(n20662), .ZN(n12003) );
  NAND3_X1 U15151 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20879) );
  INV_X1 U15152 ( .A(n20879), .ZN(n20890) );
  NAND2_X1 U15153 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20890), .ZN(
        n20877) );
  AND2_X1 U15154 ( .A1(n12003), .A2(n20877), .ZN(n20461) );
  AOI22_X1 U15155 ( .A1(n12004), .A2(n20461), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20944), .ZN(n12005) );
  NAND2_X1 U15156 ( .A1(n13342), .A2(n21045), .ZN(n12023) );
  INV_X1 U15157 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U15158 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12010) );
  NAND2_X1 U15159 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12009) );
  OAI211_X1 U15160 ( .C1(n12647), .C2(n12527), .A(n12010), .B(n12009), .ZN(
        n12011) );
  INV_X1 U15161 ( .A(n12011), .ZN(n12015) );
  AOI22_X1 U15162 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12014) );
  INV_X1 U15163 ( .A(n12634), .ZN(n12447) );
  AOI22_X1 U15164 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12013) );
  NAND2_X1 U15165 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12012) );
  NAND4_X1 U15166 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12021) );
  AOI22_X1 U15167 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15168 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15169 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15170 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U15171 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12020) );
  AOI22_X1 U15172 ( .A1(n12788), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12802), .B2(n12702), .ZN(n12022) );
  NAND2_X1 U15173 ( .A1(n12788), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12038) );
  INV_X1 U15174 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12543) );
  NAND2_X1 U15175 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12025) );
  NAND2_X1 U15176 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12024) );
  OAI211_X1 U15177 ( .C1(n12578), .C2(n12543), .A(n12025), .B(n12024), .ZN(
        n12026) );
  INV_X1 U15178 ( .A(n12026), .ZN(n12030) );
  AOI22_X1 U15179 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15180 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12028) );
  INV_X2 U15181 ( .A(n11798), .ZN(n13359) );
  NAND2_X1 U15182 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12027) );
  NAND4_X1 U15183 ( .A1(n12030), .A2(n12029), .A3(n12028), .A4(n12027), .ZN(
        n12036) );
  AOI22_X1 U15184 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12585), .B1(
        n12411), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15185 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n9666), .B1(
        n12342), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15186 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9668), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15187 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12031) );
  NAND4_X1 U15188 ( .A1(n12034), .A2(n12033), .A3(n12032), .A4(n12031), .ZN(
        n12035) );
  NAND2_X1 U15189 ( .A1(n12802), .A2(n12710), .ZN(n12037) );
  NAND2_X1 U15190 ( .A1(n12038), .A2(n12037), .ZN(n12129) );
  NAND2_X1 U15191 ( .A1(n12788), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12054) );
  INV_X1 U15192 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12041) );
  NAND2_X1 U15193 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12040) );
  NAND2_X1 U15194 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12039) );
  OAI211_X1 U15195 ( .C1(n12578), .C2(n12041), .A(n12040), .B(n12039), .ZN(
        n12042) );
  INV_X1 U15196 ( .A(n12042), .ZN(n12046) );
  AOI22_X1 U15197 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15198 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12044) );
  NAND2_X1 U15199 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12043) );
  NAND4_X1 U15200 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12052) );
  AOI22_X1 U15201 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15202 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15203 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12048) );
  INV_X1 U15204 ( .A(n12546), .ZN(n12403) );
  AOI22_X1 U15205 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15206 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12051) );
  OR2_X1 U15207 ( .A1(n12052), .A2(n12051), .ZN(n12720) );
  NAND2_X1 U15208 ( .A1(n12802), .A2(n12720), .ZN(n12053) );
  NAND2_X1 U15209 ( .A1(n12054), .A2(n12053), .ZN(n12139) );
  INV_X1 U15210 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12057) );
  NAND2_X1 U15211 ( .A1(n12403), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12056) );
  NAND2_X1 U15212 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12055) );
  OAI211_X1 U15213 ( .C1(n12647), .C2(n12057), .A(n12056), .B(n12055), .ZN(
        n12058) );
  INV_X1 U15214 ( .A(n12058), .ZN(n12062) );
  AOI22_X1 U15215 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15216 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12060) );
  NAND2_X1 U15217 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12059) );
  NAND4_X1 U15218 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12068) );
  INV_X1 U15219 ( .A(n12605), .ZN(n12342) );
  AOI22_X1 U15220 ( .A1(n12649), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12616), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15221 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15222 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12411), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15223 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U15224 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12067) );
  OR2_X1 U15225 ( .A1(n12068), .A2(n12067), .ZN(n12724) );
  AOI22_X1 U15226 ( .A1(n12788), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12802), .B2(n12724), .ZN(n12148) );
  NAND2_X1 U15227 ( .A1(n12788), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12072) );
  NAND2_X1 U15228 ( .A1(n12802), .A2(n12735), .ZN(n12071) );
  NAND2_X1 U15229 ( .A1(n12072), .A2(n12071), .ZN(n12073) );
  XNOR2_X1 U15230 ( .A(n12668), .B(n12073), .ZN(n12729) );
  INV_X2 U15231 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21042) );
  NAND2_X1 U15232 ( .A1(n12729), .A2(n12292), .ZN(n12080) );
  INV_X1 U15233 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12077) );
  NOR2_X1 U15234 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12538) );
  NAND2_X1 U15235 ( .A1(n12142), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12141) );
  INV_X1 U15236 ( .A(n12150), .ZN(n12075) );
  INV_X1 U15237 ( .A(n12167), .ZN(n12074) );
  OAI21_X1 U15238 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12075), .A(
        n12074), .ZN(n20319) );
  AOI22_X1 U15239 ( .A1(n13667), .A2(n20319), .B1(n12861), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12076) );
  OAI21_X1 U15240 ( .B1(n12663), .B2(n12077), .A(n12076), .ZN(n12078) );
  INV_X1 U15241 ( .A(n12078), .ZN(n12079) );
  AOI22_X1 U15242 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12082) );
  NAND2_X1 U15243 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12081) );
  AND2_X1 U15244 ( .A1(n12082), .A2(n12081), .ZN(n12086) );
  AOI22_X1 U15245 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15246 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12084) );
  NAND2_X1 U15247 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12083) );
  NAND4_X1 U15248 ( .A1(n12086), .A2(n12085), .A3(n12084), .A4(n12083), .ZN(
        n12092) );
  AOI22_X1 U15249 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12649), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15250 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U15251 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15252 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12087) );
  NAND4_X1 U15253 ( .A1(n12090), .A2(n12089), .A3(n12088), .A4(n12087), .ZN(
        n12091) );
  NOR2_X1 U15254 ( .A1(n12092), .A2(n12091), .ZN(n12096) );
  NAND2_X1 U15255 ( .A1(n12862), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12095) );
  XOR2_X1 U15256 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12167), .Z(n20301) );
  INV_X1 U15257 ( .A(n20301), .ZN(n12093) );
  AOI22_X1 U15258 ( .A1(n12861), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13667), .B2(n12093), .ZN(n12094) );
  OAI211_X1 U15259 ( .C1(n12096), .C2(n12260), .A(n12095), .B(n12094), .ZN(
        n14010) );
  NAND2_X1 U15260 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  INV_X1 U15261 ( .A(n14267), .ZN(n13526) );
  AND2_X1 U15262 ( .A1(n13526), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12131) );
  INV_X1 U15263 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20412) );
  OAI21_X1 U15264 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n12100), .ZN(n13687) );
  OAI21_X1 U15265 ( .B1(n13687), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21042), 
        .ZN(n12101) );
  OAI21_X1 U15266 ( .B1(n12663), .B2(n20412), .A(n12101), .ZN(n12102) );
  AOI21_X1 U15267 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n12131), .A(
        n12102), .ZN(n12103) );
  NAND2_X1 U15268 ( .A1(n12861), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13658) );
  NAND2_X1 U15269 ( .A1(n13595), .A2(n12292), .ZN(n12111) );
  INV_X1 U15270 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12108) );
  INV_X1 U15271 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13462) );
  OAI22_X1 U15272 ( .A1(n12663), .A2(n12108), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13462), .ZN(n12109) );
  AOI21_X1 U15273 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12131), .A(
        n12109), .ZN(n12110) );
  NAND2_X1 U15274 ( .A1(n12111), .A2(n12110), .ZN(n13443) );
  MUX2_X1 U15275 ( .A(n12114), .B(n12113), .S(n12112), .Z(n20518) );
  AOI21_X1 U15276 ( .B1(n20518), .B2(n11900), .A(n21042), .ZN(n13440) );
  NAND2_X1 U15277 ( .A1(n20546), .A2(n12292), .ZN(n12119) );
  INV_X1 U15278 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n12116) );
  INV_X1 U15279 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13794) );
  OAI22_X1 U15280 ( .A1(n12663), .A2(n12116), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13794), .ZN(n12117) );
  AOI21_X1 U15281 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12131), .A(
        n12117), .ZN(n12118) );
  NAND2_X1 U15282 ( .A1(n12119), .A2(n12118), .ZN(n13439) );
  MUX2_X1 U15283 ( .A(n13667), .B(n13440), .S(n13439), .Z(n13442) );
  NAND2_X1 U15284 ( .A1(n13443), .A2(n13442), .ZN(n13646) );
  NAND2_X1 U15285 ( .A1(n9696), .A2(n12120), .ZN(n13647) );
  NAND2_X1 U15286 ( .A1(n13647), .A2(n13658), .ZN(n12128) );
  NAND2_X1 U15287 ( .A1(n12121), .A2(n13942), .ZN(n12122) );
  INV_X1 U15288 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n12125) );
  OAI21_X1 U15289 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12123), .A(
        n12133), .ZN(n13802) );
  AOI22_X1 U15290 ( .A1(n13667), .A2(n13802), .B1(n12861), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12124) );
  OAI21_X1 U15291 ( .B1(n12663), .B2(n12125), .A(n12124), .ZN(n12126) );
  AOI21_X1 U15292 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12131), .A(
        n12126), .ZN(n12127) );
  NAND2_X1 U15293 ( .A1(n12128), .A2(n13656), .ZN(n13613) );
  NAND2_X1 U15294 ( .A1(n12131), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12135) );
  AOI21_X1 U15295 ( .B1(n13707), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12132) );
  AOI21_X1 U15296 ( .B1(n12862), .B2(P1_EAX_REG_4__SCAN_IN), .A(n12132), .ZN(
        n12134) );
  AOI21_X1 U15297 ( .B1(n13707), .B2(n12133), .A(n12142), .ZN(n20350) );
  AOI22_X1 U15298 ( .A1(n12135), .A2(n12134), .B1(n13667), .B2(n20350), .ZN(
        n12136) );
  AOI21_X1 U15299 ( .B1(n12701), .B2(n12292), .A(n12136), .ZN(n13614) );
  NAND2_X1 U15300 ( .A1(n12138), .A2(n12137), .ZN(n13612) );
  XNOR2_X1 U15301 ( .A(n12140), .B(n12139), .ZN(n12708) );
  INV_X1 U15302 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12144) );
  OAI21_X1 U15303 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12142), .A(
        n12141), .ZN(n20332) );
  AOI22_X1 U15304 ( .A1(n13667), .A2(n20332), .B1(n12861), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12143) );
  OAI21_X1 U15305 ( .B1(n12663), .B2(n12144), .A(n12143), .ZN(n12145) );
  AOI21_X1 U15306 ( .B1(n12708), .B2(n12292), .A(n12145), .ZN(n13837) );
  NAND2_X2 U15307 ( .A1(n12147), .A2(n12146), .ZN(n14016) );
  NAND2_X1 U15308 ( .A1(n12149), .A2(n12148), .ZN(n12718) );
  INV_X1 U15309 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12153) );
  OAI21_X1 U15310 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12151), .A(
        n12150), .ZN(n20330) );
  AOI22_X1 U15311 ( .A1(n13667), .A2(n20330), .B1(n12861), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12152) );
  OAI21_X1 U15312 ( .B1(n12663), .B2(n12153), .A(n12152), .ZN(n12154) );
  INV_X1 U15313 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U15314 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15315 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15316 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15317 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12155) );
  AND4_X1 U15318 ( .A1(n12158), .A2(n12157), .A3(n12156), .A4(n12155), .ZN(
        n12165) );
  AOI22_X1 U15319 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12342), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15320 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15321 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12160) );
  NAND2_X1 U15322 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12159) );
  AND3_X1 U15323 ( .A1(n12161), .A2(n12160), .A3(n12159), .ZN(n12163) );
  NAND2_X1 U15324 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12162) );
  NAND4_X1 U15325 ( .A1(n12165), .A2(n12164), .A3(n12163), .A4(n12162), .ZN(
        n12166) );
  NAND2_X1 U15326 ( .A1(n12292), .A2(n12166), .ZN(n12170) );
  NAND2_X1 U15327 ( .A1(n12167), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12172) );
  INV_X1 U15328 ( .A(n12172), .ZN(n12168) );
  XNOR2_X1 U15329 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12168), .ZN(
        n15120) );
  AOI22_X1 U15330 ( .A1(n13667), .A2(n15120), .B1(n12861), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12169) );
  OAI211_X1 U15331 ( .C1(n12663), .C2(n14111), .A(n12170), .B(n12169), .ZN(
        n14075) );
  INV_X1 U15332 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16239) );
  INV_X1 U15333 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12171) );
  XNOR2_X1 U15334 ( .A(n16239), .B(n12187), .ZN(n16284) );
  AOI22_X1 U15335 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12342), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15336 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15337 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15338 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12173) );
  AND4_X1 U15339 ( .A1(n12176), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(
        n12183) );
  AOI22_X1 U15340 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15341 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12178) );
  NAND2_X1 U15342 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12177) );
  AND3_X1 U15343 ( .A1(n12179), .A2(n12178), .A3(n12177), .ZN(n12182) );
  AOI22_X1 U15344 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12181) );
  NAND2_X1 U15345 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12180) );
  NAND4_X1 U15346 ( .A1(n12183), .A2(n12182), .A3(n12181), .A4(n12180), .ZN(
        n12184) );
  AOI22_X1 U15347 ( .A1(n12292), .A2(n12184), .B1(n12861), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12186) );
  NAND2_X1 U15348 ( .A1(n12862), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12185) );
  OAI211_X1 U15349 ( .C1(n16284), .C2(n12630), .A(n12186), .B(n12185), .ZN(
        n14108) );
  NAND2_X1 U15350 ( .A1(n12187), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12207) );
  INV_X1 U15351 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12206) );
  XNOR2_X1 U15352 ( .A(n12207), .B(n12206), .ZN(n16229) );
  NAND2_X1 U15353 ( .A1(n16229), .A2(n13667), .ZN(n12190) );
  INV_X1 U15354 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20397) );
  INV_X1 U15355 ( .A(n12861), .ZN(n12237) );
  OAI22_X1 U15356 ( .A1(n12663), .A2(n20397), .B1(n12237), .B2(n12206), .ZN(
        n12188) );
  INV_X1 U15357 ( .A(n12188), .ZN(n12189) );
  NAND2_X1 U15358 ( .A1(n12190), .A2(n12189), .ZN(n12204) );
  AOI22_X1 U15359 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12192) );
  NAND2_X1 U15360 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12191) );
  AND2_X1 U15361 ( .A1(n12192), .A2(n12191), .ZN(n12196) );
  AOI22_X1 U15362 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15363 ( .A1(n12649), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12194) );
  NAND2_X1 U15364 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12193) );
  NAND4_X1 U15365 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12202) );
  AOI22_X1 U15366 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12366), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15367 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15368 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15369 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U15370 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12201) );
  NOR2_X1 U15371 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  NOR2_X1 U15372 ( .A1(n12260), .A2(n12203), .ZN(n14911) );
  INV_X1 U15373 ( .A(n12204), .ZN(n12205) );
  NAND2_X1 U15374 ( .A1(n14850), .A2(n14852), .ZN(n14807) );
  NAND2_X1 U15375 ( .A1(n12293), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12263) );
  INV_X1 U15376 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16216) );
  NAND2_X1 U15377 ( .A1(n12243), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12223) );
  XNOR2_X1 U15378 ( .A(n12300), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15076) );
  AOI22_X1 U15379 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15380 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12209) );
  NAND2_X1 U15381 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12208) );
  AND3_X1 U15382 ( .A1(n12210), .A2(n12209), .A3(n12208), .ZN(n12218) );
  AOI22_X1 U15383 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15384 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15385 ( .A1(n12649), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15386 ( .A1(n12616), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12211) );
  AND4_X1 U15387 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12217) );
  AOI22_X1 U15388 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12216) );
  NAND2_X1 U15389 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12215) );
  NAND4_X1 U15390 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12219) );
  NAND2_X1 U15391 ( .A1(n12665), .A2(n12219), .ZN(n12221) );
  AOI22_X1 U15392 ( .A1(n12862), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21042), .ZN(n12220) );
  AOI21_X1 U15393 ( .B1(n12221), .B2(n12220), .A(n13667), .ZN(n12222) );
  AOI21_X1 U15394 ( .B1(n15076), .B2(n13667), .A(n12222), .ZN(n14810) );
  INV_X1 U15395 ( .A(n14810), .ZN(n12298) );
  XNOR2_X1 U15396 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12223), .ZN(
        n16280) );
  AOI22_X1 U15397 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12225) );
  NAND2_X1 U15398 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12224) );
  AND2_X1 U15399 ( .A1(n12225), .A2(n12224), .ZN(n12229) );
  AOI22_X1 U15400 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15401 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12227) );
  NAND2_X1 U15402 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12226) );
  NAND4_X1 U15403 ( .A1(n12229), .A2(n12228), .A3(n12227), .A4(n12226), .ZN(
        n12235) );
  AOI22_X1 U15404 ( .A1(n12649), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15405 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15406 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15407 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12230) );
  NAND4_X1 U15408 ( .A1(n12233), .A2(n12232), .A3(n12231), .A4(n12230), .ZN(
        n12234) );
  NOR2_X1 U15409 ( .A1(n12235), .A2(n12234), .ZN(n12238) );
  INV_X1 U15410 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12236) );
  OAI22_X1 U15411 ( .A1(n12260), .A2(n12238), .B1(n12237), .B2(n12236), .ZN(
        n12241) );
  INV_X1 U15412 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n12239) );
  NOR2_X1 U15413 ( .A1(n12663), .A2(n12239), .ZN(n12240) );
  NOR2_X1 U15414 ( .A1(n12241), .A2(n12240), .ZN(n12242) );
  OAI21_X1 U15415 ( .B1(n16280), .B2(n12630), .A(n12242), .ZN(n14825) );
  XNOR2_X1 U15416 ( .A(n12243), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15086) );
  INV_X1 U15417 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12246) );
  NAND2_X1 U15418 ( .A1(n12403), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12245) );
  NAND2_X1 U15419 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12244) );
  OAI211_X1 U15420 ( .C1(n12578), .C2(n12246), .A(n12245), .B(n12244), .ZN(
        n12247) );
  INV_X1 U15421 ( .A(n12247), .ZN(n12251) );
  AOI22_X1 U15422 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15423 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12249) );
  NAND2_X1 U15424 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12248) );
  NAND4_X1 U15425 ( .A1(n12251), .A2(n12250), .A3(n12249), .A4(n12248), .ZN(
        n12257) );
  AOI22_X1 U15426 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15427 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15428 ( .A1(n12649), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15429 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12252) );
  NAND4_X1 U15430 ( .A1(n12255), .A2(n12254), .A3(n12253), .A4(n12252), .ZN(
        n12256) );
  NOR2_X1 U15431 ( .A1(n12257), .A2(n12256), .ZN(n12261) );
  NAND2_X1 U15432 ( .A1(n12862), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12259) );
  NAND2_X1 U15433 ( .A1(n12861), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12258) );
  OAI211_X1 U15434 ( .C1(n12261), .C2(n12260), .A(n12259), .B(n12258), .ZN(
        n12262) );
  AOI21_X1 U15435 ( .B1(n15086), .B2(n13667), .A(n12262), .ZN(n14838) );
  INV_X1 U15436 ( .A(n14838), .ZN(n12297) );
  XNOR2_X1 U15437 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12263), .ZN(
        n16220) );
  INV_X1 U15438 ( .A(n16220), .ZN(n15096) );
  AOI22_X1 U15439 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15440 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15441 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15442 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12264) );
  NAND4_X1 U15443 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12275) );
  AOI22_X1 U15444 ( .A1(n12649), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12269) );
  NAND2_X1 U15445 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12268) );
  AND2_X1 U15446 ( .A1(n12269), .A2(n12268), .ZN(n12273) );
  AOI22_X1 U15447 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15448 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12271) );
  NAND2_X1 U15449 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12270) );
  NAND4_X1 U15450 ( .A1(n12273), .A2(n12272), .A3(n12271), .A4(n12270), .ZN(
        n12274) );
  OAI21_X1 U15451 ( .B1(n12275), .B2(n12274), .A(n12292), .ZN(n12278) );
  NAND2_X1 U15452 ( .A1(n12862), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12277) );
  NAND2_X1 U15453 ( .A1(n12861), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12276) );
  NAND3_X1 U15454 ( .A1(n12278), .A2(n12277), .A3(n12276), .ZN(n12279) );
  AOI21_X1 U15455 ( .B1(n15096), .B2(n13667), .A(n12279), .ZN(n14898) );
  INV_X1 U15456 ( .A(n14898), .ZN(n12296) );
  INV_X1 U15457 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14984) );
  AOI22_X1 U15458 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12342), .B1(
        n12616), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15459 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15460 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15461 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12411), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12280) );
  AND4_X1 U15462 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12290) );
  AOI22_X1 U15463 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15464 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15465 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12285) );
  NAND2_X1 U15466 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12284) );
  AND3_X1 U15467 ( .A1(n12286), .A2(n12285), .A3(n12284), .ZN(n12288) );
  NAND2_X1 U15468 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12287) );
  NAND4_X1 U15469 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(
        n12291) );
  NAND2_X1 U15470 ( .A1(n12292), .A2(n12291), .ZN(n12295) );
  XNOR2_X1 U15471 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12293), .ZN(
        n15106) );
  AOI22_X1 U15472 ( .A1(n13667), .A2(n15106), .B1(n12861), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12294) );
  OAI211_X1 U15473 ( .C1(n12663), .C2(n14984), .A(n12295), .B(n12294), .ZN(
        n14851) );
  AND2_X1 U15474 ( .A1(n12296), .A2(n14851), .ZN(n14836) );
  AND2_X1 U15475 ( .A1(n12297), .A2(n14836), .ZN(n14823) );
  AND2_X1 U15476 ( .A1(n14825), .A2(n14823), .ZN(n14808) );
  AND2_X1 U15477 ( .A1(n12298), .A2(n14808), .ZN(n12299) );
  NAND2_X1 U15478 ( .A1(n14807), .A2(n12299), .ZN(n14809) );
  XOR2_X1 U15479 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12320), .Z(
        n16269) );
  INV_X1 U15480 ( .A(n16269), .ZN(n12318) );
  INV_X1 U15481 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U15482 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12302) );
  NAND2_X1 U15483 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12301) );
  OAI211_X1 U15484 ( .C1(n12578), .C2(n12303), .A(n12302), .B(n12301), .ZN(
        n12304) );
  INV_X1 U15485 ( .A(n12304), .ZN(n12308) );
  AOI22_X1 U15486 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15487 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12306) );
  NAND2_X1 U15488 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12305) );
  NAND4_X1 U15489 ( .A1(n12308), .A2(n12307), .A3(n12306), .A4(n12305), .ZN(
        n12314) );
  AOI22_X1 U15490 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12411), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15491 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15492 ( .A1(n12649), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15493 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12309) );
  NAND4_X1 U15494 ( .A1(n12312), .A2(n12311), .A3(n12310), .A4(n12309), .ZN(
        n12313) );
  NOR2_X1 U15495 ( .A1(n12314), .A2(n12313), .ZN(n12316) );
  AOI22_X1 U15496 ( .A1(n12862), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12861), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12315) );
  OAI21_X1 U15497 ( .B1(n12627), .B2(n12316), .A(n12315), .ZN(n12317) );
  AOI21_X1 U15498 ( .B1(n12318), .B2(n12538), .A(n12317), .ZN(n14888) );
  XNOR2_X1 U15499 ( .A(n12339), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15066) );
  NAND2_X1 U15500 ( .A1(n15066), .A2(n13667), .ZN(n12338) );
  INV_X1 U15501 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12493) );
  NAND2_X1 U15502 ( .A1(n12403), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12322) );
  NAND2_X1 U15503 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12321) );
  OAI211_X1 U15504 ( .C1(n12647), .C2(n12493), .A(n12322), .B(n12321), .ZN(
        n12323) );
  INV_X1 U15505 ( .A(n12323), .ZN(n12327) );
  AOI22_X1 U15506 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15507 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U15508 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12324) );
  NAND4_X1 U15509 ( .A1(n12327), .A2(n12326), .A3(n12325), .A4(n12324), .ZN(
        n12333) );
  AOI22_X1 U15510 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12411), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15511 ( .A1(n12649), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15512 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15513 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12328) );
  NAND4_X1 U15514 ( .A1(n12331), .A2(n12330), .A3(n12329), .A4(n12328), .ZN(
        n12332) );
  NOR2_X1 U15515 ( .A1(n12333), .A2(n12332), .ZN(n12336) );
  INV_X1 U15516 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14802) );
  AOI21_X1 U15517 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14802), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12334) );
  AOI21_X1 U15518 ( .B1(n12862), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12334), .ZN(
        n12335) );
  OAI21_X1 U15519 ( .B1(n12627), .B2(n12336), .A(n12335), .ZN(n12337) );
  NAND2_X1 U15520 ( .A1(n12338), .A2(n12337), .ZN(n14800) );
  OR2_X1 U15521 ( .A1(n12340), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12341) );
  NAND2_X1 U15522 ( .A1(n12341), .A2(n12397), .ZN(n16268) );
  INV_X1 U15523 ( .A(n16268), .ZN(n14788) );
  AOI22_X1 U15524 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12651), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15525 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12616), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15526 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15527 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12343) );
  AND4_X1 U15528 ( .A1(n12346), .A2(n12345), .A3(n12344), .A4(n12343), .ZN(
        n12353) );
  AOI22_X1 U15529 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15530 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12348) );
  NAND2_X1 U15531 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12347) );
  AND3_X1 U15532 ( .A1(n12349), .A2(n12348), .A3(n12347), .ZN(n12352) );
  AOI22_X1 U15533 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12351) );
  NAND2_X1 U15534 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12350) );
  NAND4_X1 U15535 ( .A1(n12353), .A2(n12352), .A3(n12351), .A4(n12350), .ZN(
        n12356) );
  INV_X1 U15536 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14956) );
  NAND2_X1 U15537 ( .A1(n21042), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12354) );
  OAI211_X1 U15538 ( .C1(n12663), .C2(n14956), .A(n12630), .B(n12354), .ZN(
        n12355) );
  AOI21_X1 U15539 ( .B1(n12665), .B2(n12356), .A(n12355), .ZN(n12357) );
  AOI21_X1 U15540 ( .B1(n14788), .B2(n12538), .A(n12357), .ZN(n14781) );
  INV_X1 U15541 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12548) );
  NAND2_X1 U15542 ( .A1(n12403), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12359) );
  NAND2_X1 U15543 ( .A1(n12649), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12358) );
  OAI211_X1 U15544 ( .C1(n12578), .C2(n12548), .A(n12359), .B(n12358), .ZN(
        n12360) );
  INV_X1 U15545 ( .A(n12360), .ZN(n12364) );
  AOI22_X1 U15546 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11847), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15547 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12362) );
  NAND2_X1 U15548 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12361) );
  NAND4_X1 U15549 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .ZN(
        n12372) );
  AOI22_X1 U15550 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15551 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12411), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15552 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15553 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9665), .B1(
        n12378), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12367) );
  NAND4_X1 U15554 ( .A1(n12370), .A2(n12369), .A3(n12368), .A4(n12367), .ZN(
        n12371) );
  NOR2_X1 U15555 ( .A1(n12372), .A2(n12371), .ZN(n12375) );
  INV_X1 U15556 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16261) );
  AOI21_X1 U15557 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n16261), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12373) );
  AOI21_X1 U15558 ( .B1(n12862), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12373), .ZN(
        n12374) );
  OAI21_X1 U15559 ( .B1(n12627), .B2(n12375), .A(n12374), .ZN(n12377) );
  XNOR2_X1 U15560 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12397), .ZN(
        n16257) );
  NAND2_X1 U15561 ( .A1(n16257), .A2(n12538), .ZN(n12376) );
  NAND2_X1 U15562 ( .A1(n14770), .A2(n14772), .ZN(n14771) );
  NAND2_X1 U15563 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12382) );
  NAND2_X1 U15564 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12381) );
  NAND2_X1 U15565 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12380) );
  NAND2_X1 U15566 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12379) );
  AND4_X1 U15567 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12386) );
  AOI22_X1 U15568 ( .A1(n12616), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12385) );
  NAND2_X1 U15569 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12384) );
  NAND2_X1 U15570 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12383) );
  NAND4_X1 U15571 ( .A1(n12386), .A2(n12385), .A3(n12384), .A4(n12383), .ZN(
        n12392) );
  AOI22_X1 U15572 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12649), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12390) );
  AOI22_X1 U15573 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15574 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15575 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12387) );
  NAND4_X1 U15576 ( .A1(n12390), .A2(n12389), .A3(n12388), .A4(n12387), .ZN(
        n12391) );
  NOR2_X1 U15577 ( .A1(n12392), .A2(n12391), .ZN(n12396) );
  NAND2_X1 U15578 ( .A1(n21042), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12393) );
  NAND2_X1 U15579 ( .A1(n12630), .A2(n12393), .ZN(n12394) );
  AOI21_X1 U15580 ( .B1(n12862), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12394), .ZN(
        n12395) );
  OAI21_X1 U15581 ( .B1(n12627), .B2(n12396), .A(n12395), .ZN(n12400) );
  OAI21_X1 U15582 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12398), .A(
        n12458), .ZN(n16253) );
  OR2_X1 U15583 ( .A1(n12630), .A2(n16253), .ZN(n12399) );
  NAND2_X1 U15584 ( .A1(n12400), .A2(n12399), .ZN(n14948) );
  INV_X1 U15585 ( .A(n14948), .ZN(n12401) );
  AOI22_X1 U15586 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12405) );
  NAND2_X1 U15587 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12404) );
  AND2_X1 U15588 ( .A1(n12405), .A2(n12404), .ZN(n12409) );
  AOI22_X1 U15589 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15590 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12407) );
  NAND2_X1 U15591 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12406) );
  NAND4_X1 U15592 ( .A1(n12409), .A2(n12408), .A3(n12407), .A4(n12406), .ZN(
        n12417) );
  AOI22_X1 U15593 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15594 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12651), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15595 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15596 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12412) );
  NAND4_X1 U15597 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12416) );
  NOR2_X1 U15598 ( .A1(n12417), .A2(n12416), .ZN(n12421) );
  NAND2_X1 U15599 ( .A1(n21042), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12418) );
  NAND2_X1 U15600 ( .A1(n12630), .A2(n12418), .ZN(n12419) );
  AOI21_X1 U15601 ( .B1(n12862), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12419), .ZN(
        n12420) );
  OAI21_X1 U15602 ( .B1(n12627), .B2(n12421), .A(n12420), .ZN(n12423) );
  XNOR2_X1 U15603 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12458), .ZN(
        n15055) );
  NAND2_X1 U15604 ( .A1(n12538), .A2(n15055), .ZN(n12422) );
  NAND2_X1 U15605 ( .A1(n12423), .A2(n12422), .ZN(n14758) );
  INV_X1 U15606 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12638) );
  INV_X1 U15607 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12636) );
  INV_X1 U15608 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12424) );
  OAI22_X1 U15609 ( .A1(n11822), .A2(n12636), .B1(n12634), .B2(n12424), .ZN(
        n12428) );
  INV_X1 U15610 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12426) );
  INV_X1 U15611 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12425) );
  OAI22_X1 U15612 ( .A1(n12639), .A2(n12426), .B1(n12637), .B2(n12425), .ZN(
        n12427) );
  AOI211_X1 U15613 ( .C1(n13359), .C2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n12428), .B(n12427), .ZN(n12431) );
  AOI22_X1 U15614 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12430) );
  OAI211_X1 U15615 ( .C1(n12578), .C2(n12638), .A(n12431), .B(n12430), .ZN(
        n12437) );
  AOI22_X1 U15616 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15617 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15618 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15619 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12432) );
  NAND4_X1 U15620 ( .A1(n12435), .A2(n12434), .A3(n12433), .A4(n12432), .ZN(
        n12436) );
  NOR2_X1 U15621 ( .A1(n12437), .A2(n12436), .ZN(n12465) );
  INV_X1 U15622 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12446) );
  INV_X1 U15623 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12439) );
  OAI22_X1 U15624 ( .A1(n12639), .A2(n12439), .B1(n9654), .B2(n12438), .ZN(
        n12443) );
  INV_X1 U15625 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12441) );
  INV_X1 U15626 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12440) );
  OAI22_X1 U15627 ( .A1(n11822), .A2(n12441), .B1(n12608), .B2(n12440), .ZN(
        n12442) );
  AOI211_X1 U15628 ( .C1(n11744), .C2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n12443), .B(n12442), .ZN(n12445) );
  AOI22_X1 U15629 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12444) );
  OAI211_X1 U15630 ( .C1(n11798), .C2(n12446), .A(n12445), .B(n12444), .ZN(
        n12453) );
  AOI22_X1 U15631 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15632 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15633 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15634 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12448) );
  NAND4_X1 U15635 ( .A1(n12451), .A2(n12450), .A3(n12449), .A4(n12448), .ZN(
        n12452) );
  NOR2_X1 U15636 ( .A1(n12453), .A2(n12452), .ZN(n12466) );
  XNOR2_X1 U15637 ( .A(n12465), .B(n12466), .ZN(n12457) );
  NAND2_X1 U15638 ( .A1(n21042), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12454) );
  NAND2_X1 U15639 ( .A1(n12630), .A2(n12454), .ZN(n12455) );
  AOI21_X1 U15640 ( .B1(n12862), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12455), .ZN(
        n12456) );
  OAI21_X1 U15641 ( .B1(n12457), .B2(n12627), .A(n12456), .ZN(n12464) );
  INV_X1 U15642 ( .A(n12458), .ZN(n12459) );
  INV_X1 U15643 ( .A(n12460), .ZN(n12461) );
  INV_X1 U15644 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15046) );
  NAND2_X1 U15645 ( .A1(n12461), .A2(n15046), .ZN(n12462) );
  AND2_X1 U15646 ( .A1(n12509), .A2(n12462), .ZN(n15050) );
  NAND2_X1 U15647 ( .A1(n15050), .A2(n12538), .ZN(n12463) );
  AND2_X1 U15648 ( .A1(n12464), .A2(n12463), .ZN(n14748) );
  NOR2_X1 U15649 ( .A1(n12466), .A2(n12465), .ZN(n12489) );
  INV_X1 U15650 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12469) );
  NAND2_X1 U15651 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12468) );
  NAND2_X1 U15652 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12467) );
  OAI211_X1 U15653 ( .C1(n12647), .C2(n12469), .A(n12468), .B(n12467), .ZN(
        n12470) );
  INV_X1 U15654 ( .A(n12470), .ZN(n12474) );
  AOI22_X1 U15655 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15656 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12472) );
  NAND2_X1 U15657 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12471) );
  NAND4_X1 U15658 ( .A1(n12474), .A2(n12473), .A3(n12472), .A4(n12471), .ZN(
        n12480) );
  AOI22_X1 U15659 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15660 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12616), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15661 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15662 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12475) );
  NAND4_X1 U15663 ( .A1(n12478), .A2(n12477), .A3(n12476), .A4(n12475), .ZN(
        n12479) );
  OR2_X1 U15664 ( .A1(n12480), .A2(n12479), .ZN(n12488) );
  INV_X1 U15665 ( .A(n12488), .ZN(n12481) );
  XNOR2_X1 U15666 ( .A(n12489), .B(n12481), .ZN(n12482) );
  NAND2_X1 U15667 ( .A1(n12482), .A2(n12665), .ZN(n12487) );
  NAND2_X1 U15668 ( .A1(n21042), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12483) );
  NAND2_X1 U15669 ( .A1(n12630), .A2(n12483), .ZN(n12484) );
  AOI21_X1 U15670 ( .B1(n12862), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12484), .ZN(
        n12486) );
  XNOR2_X1 U15671 ( .A(n12509), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15042) );
  AND2_X1 U15672 ( .A1(n15042), .A2(n12538), .ZN(n12485) );
  AOI21_X1 U15673 ( .B1(n12487), .B2(n12486), .A(n12485), .ZN(n14736) );
  INV_X1 U15674 ( .A(n14720), .ZN(n12516) );
  NAND2_X1 U15675 ( .A1(n12489), .A2(n12488), .ZN(n12517) );
  INV_X1 U15676 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12499) );
  INV_X1 U15677 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12491) );
  OAI22_X1 U15678 ( .A1(n12492), .A2(n12491), .B1(n9654), .B2(n12490), .ZN(
        n12496) );
  INV_X1 U15679 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12494) );
  OAI22_X1 U15680 ( .A1(n11822), .A2(n12494), .B1(n12639), .B2(n12493), .ZN(
        n12495) );
  AOI211_X1 U15681 ( .C1(n13359), .C2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n12496), .B(n12495), .ZN(n12498) );
  AOI22_X1 U15682 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12497) );
  OAI211_X1 U15683 ( .C1(n12647), .C2(n12499), .A(n12498), .B(n12497), .ZN(
        n12505) );
  AOI22_X1 U15684 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U15685 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12651), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15686 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15687 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12500) );
  NAND4_X1 U15688 ( .A1(n12503), .A2(n12502), .A3(n12501), .A4(n12500), .ZN(
        n12504) );
  NOR2_X1 U15689 ( .A1(n12505), .A2(n12504), .ZN(n12518) );
  XNOR2_X1 U15690 ( .A(n12517), .B(n12518), .ZN(n12508) );
  INV_X1 U15691 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14727) );
  AOI21_X1 U15692 ( .B1(n14727), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12506) );
  AOI21_X1 U15693 ( .B1(n12862), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12506), .ZN(
        n12507) );
  OAI21_X1 U15694 ( .B1(n12508), .B2(n12627), .A(n12507), .ZN(n12514) );
  INV_X1 U15695 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15038) );
  NAND2_X1 U15696 ( .A1(n12510), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12566) );
  INV_X1 U15697 ( .A(n12510), .ZN(n12511) );
  NAND2_X1 U15698 ( .A1(n12511), .A2(n14727), .ZN(n12512) );
  NAND2_X1 U15699 ( .A1(n12566), .A2(n12512), .ZN(n15032) );
  OR2_X1 U15700 ( .A1(n15032), .A2(n12630), .ZN(n12513) );
  NAND2_X1 U15701 ( .A1(n12514), .A2(n12513), .ZN(n14722) );
  NOR2_X1 U15702 ( .A1(n12518), .A2(n12517), .ZN(n12561) );
  INV_X1 U15703 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12521) );
  NAND2_X1 U15704 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12520) );
  NAND2_X1 U15705 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12519) );
  OAI211_X1 U15706 ( .C1(n12647), .C2(n12521), .A(n12520), .B(n12519), .ZN(
        n12522) );
  INV_X1 U15707 ( .A(n12522), .ZN(n12526) );
  AOI22_X1 U15708 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15709 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12524) );
  NAND2_X1 U15710 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12523) );
  NAND4_X1 U15711 ( .A1(n12526), .A2(n12525), .A3(n12524), .A4(n12523), .ZN(
        n12533) );
  AOI22_X1 U15712 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15713 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15714 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15715 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12528) );
  NAND4_X1 U15716 ( .A1(n12531), .A2(n12530), .A3(n12529), .A4(n12528), .ZN(
        n12532) );
  OR2_X1 U15717 ( .A1(n12533), .A2(n12532), .ZN(n12560) );
  XNOR2_X1 U15718 ( .A(n12561), .B(n12560), .ZN(n12537) );
  NAND2_X1 U15719 ( .A1(n21042), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12534) );
  NAND2_X1 U15720 ( .A1(n12630), .A2(n12534), .ZN(n12535) );
  AOI21_X1 U15721 ( .B1(n12862), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12535), .ZN(
        n12536) );
  OAI21_X1 U15722 ( .B1(n12537), .B2(n12627), .A(n12536), .ZN(n12540) );
  XNOR2_X1 U15723 ( .A(n12566), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15023) );
  NAND2_X1 U15724 ( .A1(n15023), .A2(n12538), .ZN(n12539) );
  NAND2_X1 U15725 ( .A1(n12540), .A2(n12539), .ZN(n14708) );
  INV_X1 U15726 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12553) );
  INV_X1 U15727 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12545) );
  OAI22_X1 U15728 ( .A1(n12546), .A2(n12545), .B1(n9654), .B2(n12543), .ZN(
        n12550) );
  INV_X1 U15729 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12547) );
  OAI22_X1 U15730 ( .A1(n12548), .A2(n12639), .B1(n12634), .B2(n12547), .ZN(
        n12549) );
  AOI211_X1 U15731 ( .C1(n13359), .C2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n12550), .B(n12549), .ZN(n12552) );
  AOI22_X1 U15732 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12651), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12551) );
  OAI211_X1 U15733 ( .C1(n12578), .C2(n12553), .A(n12552), .B(n12551), .ZN(
        n12559) );
  AOI22_X1 U15734 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15735 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12585), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15736 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12649), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15737 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12554) );
  NAND4_X1 U15738 ( .A1(n12557), .A2(n12556), .A3(n12555), .A4(n12554), .ZN(
        n12558) );
  NOR2_X1 U15739 ( .A1(n12559), .A2(n12558), .ZN(n12574) );
  NAND2_X1 U15740 ( .A1(n12561), .A2(n12560), .ZN(n12573) );
  XNOR2_X1 U15741 ( .A(n12574), .B(n12573), .ZN(n12565) );
  NAND2_X1 U15742 ( .A1(n21042), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12562) );
  NAND2_X1 U15743 ( .A1(n12630), .A2(n12562), .ZN(n12563) );
  AOI21_X1 U15744 ( .B1(n12862), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12563), .ZN(
        n12564) );
  OAI21_X1 U15745 ( .B1(n12565), .B2(n12627), .A(n12564), .ZN(n12572) );
  INV_X1 U15746 ( .A(n12566), .ZN(n12567) );
  INV_X1 U15747 ( .A(n12568), .ZN(n12569) );
  INV_X1 U15748 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14699) );
  NAND2_X1 U15749 ( .A1(n12569), .A2(n14699), .ZN(n12570) );
  NAND2_X1 U15750 ( .A1(n12597), .A2(n12570), .ZN(n15014) );
  OR2_X1 U15751 ( .A1(n15014), .A2(n12630), .ZN(n12571) );
  NAND2_X1 U15752 ( .A1(n12572), .A2(n12571), .ZN(n14695) );
  XNOR2_X1 U15753 ( .A(n12597), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15006) );
  INV_X1 U15754 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15002) );
  OAI21_X1 U15755 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15002), .A(n12630), 
        .ZN(n12595) );
  NOR2_X1 U15756 ( .A1(n12574), .A2(n12573), .ZN(n12624) );
  INV_X1 U15757 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12577) );
  NAND2_X1 U15758 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12576) );
  NAND2_X1 U15759 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12575) );
  OAI211_X1 U15760 ( .C1(n12578), .C2(n12577), .A(n12576), .B(n12575), .ZN(
        n12579) );
  INV_X1 U15761 ( .A(n12579), .ZN(n12584) );
  AOI22_X1 U15762 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12580), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15763 ( .A1(n9664), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12582) );
  NAND2_X1 U15764 ( .A1(n13359), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12581) );
  NAND4_X1 U15765 ( .A1(n12584), .A2(n12583), .A3(n12582), .A4(n12581), .ZN(
        n12592) );
  AOI22_X1 U15766 ( .A1(n12411), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12585), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15767 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15768 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U15769 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12587) );
  NAND4_X1 U15770 ( .A1(n12590), .A2(n12589), .A3(n12588), .A4(n12587), .ZN(
        n12591) );
  OR2_X1 U15771 ( .A1(n12592), .A2(n12591), .ZN(n12623) );
  XNOR2_X1 U15772 ( .A(n12624), .B(n12623), .ZN(n12593) );
  NOR2_X1 U15773 ( .A1(n12593), .A2(n12627), .ZN(n12594) );
  AOI211_X1 U15774 ( .C1(n12862), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12595), .B(
        n12594), .ZN(n12596) );
  AOI21_X1 U15775 ( .B1(n12538), .B2(n15006), .A(n12596), .ZN(n14261) );
  INV_X1 U15776 ( .A(n12597), .ZN(n12598) );
  INV_X1 U15777 ( .A(n12599), .ZN(n12600) );
  INV_X1 U15778 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14686) );
  NAND2_X1 U15779 ( .A1(n12600), .A2(n14686), .ZN(n12601) );
  NAND2_X1 U15780 ( .A1(n12855), .A2(n12601), .ZN(n14994) );
  INV_X1 U15781 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12613) );
  INV_X1 U15782 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12602) );
  OAI22_X1 U15783 ( .A1(n12605), .A2(n12604), .B1(n12603), .B2(n12602), .ZN(
        n12610) );
  INV_X1 U15784 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12607) );
  INV_X1 U15785 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12606) );
  OAI22_X1 U15786 ( .A1(n12608), .A2(n12607), .B1(n12639), .B2(n12606), .ZN(
        n12609) );
  AOI211_X1 U15787 ( .C1(n13359), .C2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12610), .B(n12609), .ZN(n12612) );
  AOI22_X1 U15788 ( .A1(n12650), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12611) );
  OAI211_X1 U15789 ( .C1(n12647), .C2(n12613), .A(n12612), .B(n12611), .ZN(
        n12622) );
  AOI22_X1 U15790 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12614), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15791 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12651), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U15792 ( .A1(n12585), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12447), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15793 ( .A1(n12616), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9668), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12617) );
  NAND4_X1 U15794 ( .A1(n12620), .A2(n12619), .A3(n12618), .A4(n12617), .ZN(
        n12621) );
  NOR2_X1 U15795 ( .A1(n12622), .A2(n12621), .ZN(n12632) );
  NAND2_X1 U15796 ( .A1(n12624), .A2(n12623), .ZN(n12631) );
  XNOR2_X1 U15797 ( .A(n12632), .B(n12631), .ZN(n12628) );
  AOI21_X1 U15798 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21042), .A(
        n13667), .ZN(n12626) );
  NAND2_X1 U15799 ( .A1(n12862), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12625) );
  OAI211_X1 U15800 ( .C1(n12628), .C2(n12627), .A(n12626), .B(n12625), .ZN(
        n12629) );
  OAI21_X1 U15801 ( .B1(n12630), .B2(n14994), .A(n12629), .ZN(n14681) );
  XNOR2_X1 U15802 ( .A(n12855), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14671) );
  NOR2_X1 U15803 ( .A1(n12632), .A2(n12631), .ZN(n12660) );
  INV_X1 U15804 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12646) );
  INV_X1 U15805 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12635) );
  INV_X1 U15806 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12633) );
  OAI22_X1 U15807 ( .A1(n11822), .A2(n12635), .B1(n12634), .B2(n12633), .ZN(
        n12641) );
  OAI22_X1 U15808 ( .A1(n12639), .A2(n12638), .B1(n12637), .B2(n12636), .ZN(
        n12640) );
  AOI211_X1 U15809 ( .C1(n13359), .C2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n12641), .B(n12640), .ZN(n12645) );
  AOI22_X1 U15810 ( .A1(n9668), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12644) );
  OAI211_X1 U15811 ( .C1(n12647), .C2(n12646), .A(n12645), .B(n12644), .ZN(
        n12658) );
  AOI22_X1 U15812 ( .A1(n12410), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9664), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U15813 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12616), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15814 ( .A1(n12651), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12650), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U15815 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12429), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12653) );
  NAND4_X1 U15816 ( .A1(n12656), .A2(n12655), .A3(n12654), .A4(n12653), .ZN(
        n12657) );
  NOR2_X1 U15817 ( .A1(n12658), .A2(n12657), .ZN(n12659) );
  XNOR2_X1 U15818 ( .A(n12660), .B(n12659), .ZN(n12666) );
  INV_X1 U15819 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12662) );
  INV_X1 U15820 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21172) );
  NOR2_X1 U15821 ( .A1(n21172), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12661) );
  OAI22_X1 U15822 ( .A1(n12663), .A2(n12662), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12661), .ZN(n12664) );
  AOI21_X1 U15823 ( .B1(n12666), .B2(n12665), .A(n12664), .ZN(n12667) );
  AOI21_X1 U15824 ( .B1(n12538), .B2(n14671), .A(n12667), .ZN(n12860) );
  XNOR2_X1 U15825 ( .A(n14679), .B(n12860), .ZN(n14921) );
  NOR2_X2 U15826 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20889) );
  AND2_X1 U15827 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20889), .ZN(n21030) );
  AND3_X2 U15828 ( .A1(n21030), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n21045), 
        .ZN(n16286) );
  AND3_X1 U15829 ( .A1(n12669), .A2(n13303), .A3(n12735), .ZN(n12670) );
  NAND2_X1 U15830 ( .A1(n15224), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12757) );
  INV_X1 U15831 ( .A(n13303), .ZN(n12697) );
  NAND2_X1 U15832 ( .A1(n14002), .A2(n13954), .ZN(n12688) );
  OAI21_X1 U15833 ( .B1(n13246), .B2(n12685), .A(n12688), .ZN(n12671) );
  INV_X1 U15834 ( .A(n12671), .ZN(n12672) );
  NAND2_X1 U15835 ( .A1(n13491), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13490) );
  NAND2_X1 U15836 ( .A1(n12673), .A2(n13958), .ZN(n12678) );
  XNOR2_X1 U15837 ( .A(n12674), .B(n12684), .ZN(n12676) );
  NAND2_X1 U15838 ( .A1(n13941), .A2(n14265), .ZN(n12675) );
  AOI21_X1 U15839 ( .B1(n21043), .B2(n12676), .A(n12675), .ZN(n12677) );
  NAND2_X1 U15840 ( .A1(n12678), .A2(n12677), .ZN(n12679) );
  XNOR2_X1 U15841 ( .A(n13490), .B(n12679), .ZN(n13460) );
  NAND2_X1 U15842 ( .A1(n13460), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12682) );
  INV_X1 U15843 ( .A(n13490), .ZN(n12680) );
  NAND2_X1 U15844 ( .A1(n12680), .A2(n12679), .ZN(n12681) );
  NAND2_X1 U15845 ( .A1(n12682), .A2(n12681), .ZN(n12693) );
  INV_X1 U15846 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12683) );
  XNOR2_X1 U15847 ( .A(n12693), .B(n12683), .ZN(n13552) );
  OR2_X1 U15848 ( .A1(n20582), .A2(n12697), .ZN(n12692) );
  NAND2_X1 U15849 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  NAND2_X1 U15850 ( .A1(n12686), .A2(n12687), .ZN(n12703) );
  OAI21_X1 U15851 ( .B1(n12687), .B2(n12686), .A(n12703), .ZN(n12690) );
  INV_X1 U15852 ( .A(n12688), .ZN(n12689) );
  AOI21_X1 U15853 ( .B1(n21043), .B2(n12690), .A(n12689), .ZN(n12691) );
  NAND2_X1 U15854 ( .A1(n12693), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12694) );
  NAND2_X1 U15855 ( .A1(n12695), .A2(n12694), .ZN(n13654) );
  XNOR2_X1 U15856 ( .A(n12703), .B(n12702), .ZN(n12696) );
  INV_X1 U15857 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13741) );
  XNOR2_X1 U15858 ( .A(n12698), .B(n13741), .ZN(n13655) );
  NAND2_X1 U15859 ( .A1(n13654), .A2(n13655), .ZN(n12700) );
  NAND2_X1 U15860 ( .A1(n12698), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12699) );
  NAND2_X1 U15861 ( .A1(n12701), .A2(n13303), .ZN(n12706) );
  NAND2_X1 U15862 ( .A1(n12703), .A2(n12702), .ZN(n12709) );
  XNOR2_X1 U15863 ( .A(n12709), .B(n12710), .ZN(n12704) );
  NAND2_X1 U15864 ( .A1(n12704), .A2(n21043), .ZN(n12705) );
  NAND2_X1 U15865 ( .A1(n12706), .A2(n12705), .ZN(n12707) );
  INV_X1 U15866 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13742) );
  XNOR2_X1 U15867 ( .A(n12707), .B(n13742), .ZN(n13704) );
  NAND2_X1 U15868 ( .A1(n12708), .A2(n13303), .ZN(n12714) );
  INV_X1 U15869 ( .A(n12709), .ZN(n12711) );
  NAND2_X1 U15870 ( .A1(n12711), .A2(n12710), .ZN(n12719) );
  XNOR2_X1 U15871 ( .A(n12719), .B(n12720), .ZN(n12712) );
  NAND2_X1 U15872 ( .A1(n12712), .A2(n21043), .ZN(n12713) );
  NAND2_X1 U15873 ( .A1(n12714), .A2(n12713), .ZN(n12716) );
  INV_X1 U15874 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12715) );
  XNOR2_X1 U15875 ( .A(n12716), .B(n12715), .ZN(n13814) );
  NAND2_X1 U15876 ( .A1(n12716), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12717) );
  INV_X1 U15877 ( .A(n12719), .ZN(n12721) );
  NAND2_X1 U15878 ( .A1(n12721), .A2(n12720), .ZN(n12723) );
  INV_X1 U15879 ( .A(n12723), .ZN(n12725) );
  INV_X1 U15880 ( .A(n12724), .ZN(n12722) );
  OR2_X1 U15881 ( .A1(n12723), .A2(n12722), .ZN(n12734) );
  OAI211_X1 U15882 ( .C1(n12725), .C2(n12724), .A(n12734), .B(n21043), .ZN(
        n12726) );
  NAND2_X1 U15883 ( .A1(n12727), .A2(n12726), .ZN(n12728) );
  INV_X1 U15884 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16414) );
  XNOR2_X1 U15885 ( .A(n12728), .B(n16414), .ZN(n14015) );
  NAND2_X1 U15886 ( .A1(n12729), .A2(n13303), .ZN(n12732) );
  XNOR2_X1 U15887 ( .A(n12734), .B(n12735), .ZN(n12730) );
  NAND2_X1 U15888 ( .A1(n12730), .A2(n21043), .ZN(n12731) );
  NAND2_X1 U15889 ( .A1(n12732), .A2(n12731), .ZN(n12733) );
  OR2_X1 U15890 ( .A1(n12733), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16293) );
  NAND2_X1 U15891 ( .A1(n12733), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16292) );
  INV_X1 U15892 ( .A(n12734), .ZN(n12736) );
  NAND3_X1 U15893 ( .A1(n12736), .A2(n21043), .A3(n12735), .ZN(n12737) );
  NAND2_X1 U15894 ( .A1(n12742), .A2(n12737), .ZN(n15124) );
  OR2_X1 U15895 ( .A1(n15124), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12738) );
  NAND2_X1 U15896 ( .A1(n15124), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12739) );
  INV_X1 U15897 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15275) );
  INV_X2 U15898 ( .A(n12742), .ZN(n16163) );
  INV_X2 U15899 ( .A(n16163), .ZN(n15227) );
  NAND2_X1 U15900 ( .A1(n15227), .A2(n15275), .ZN(n12741) );
  NAND2_X1 U15901 ( .A1(n16163), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15081) );
  INV_X1 U15902 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16357) );
  NAND2_X1 U15903 ( .A1(n15224), .A2(n16357), .ZN(n12743) );
  NAND2_X1 U15904 ( .A1(n15081), .A2(n12743), .ZN(n15093) );
  NAND2_X1 U15905 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12744) );
  INV_X1 U15906 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12745) );
  NAND2_X1 U15907 ( .A1(n15224), .A2(n12745), .ZN(n15102) );
  NAND2_X1 U15908 ( .A1(n15018), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16276) );
  XNOR2_X1 U15909 ( .A(n15224), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15074) );
  INV_X1 U15910 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14280) );
  NAND2_X1 U15911 ( .A1(n15224), .A2(n14280), .ZN(n16275) );
  AND2_X1 U15912 ( .A1(n15074), .A2(n16275), .ZN(n12746) );
  NAND2_X1 U15913 ( .A1(n12747), .A2(n12746), .ZN(n15235) );
  OAI21_X1 U15914 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(n15018), .ZN(n12748) );
  INV_X1 U15915 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15247) );
  NAND2_X1 U15916 ( .A1(n15227), .A2(n15247), .ZN(n12749) );
  INV_X1 U15917 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15266) );
  INV_X1 U15918 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16389) );
  NAND2_X1 U15919 ( .A1(n15266), .A2(n16389), .ZN(n12750) );
  NAND2_X1 U15920 ( .A1(n15018), .A2(n12750), .ZN(n15100) );
  NAND2_X1 U15921 ( .A1(n16163), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15103) );
  NAND2_X1 U15922 ( .A1(n15100), .A2(n15103), .ZN(n15092) );
  NOR2_X1 U15923 ( .A1(n15072), .A2(n15092), .ZN(n12751) );
  XNOR2_X1 U15924 ( .A(n15227), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15062) );
  AND2_X1 U15925 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16167) );
  INV_X1 U15926 ( .A(n16167), .ZN(n16185) );
  INV_X1 U15927 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14301) );
  INV_X1 U15928 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15220) );
  INV_X1 U15929 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U15930 ( .A1(n15220), .A2(n12753), .ZN(n16184) );
  AND2_X1 U15931 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15195) );
  NAND2_X1 U15932 ( .A1(n15195), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15151) );
  NAND2_X1 U15933 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15182) );
  NAND2_X1 U15934 ( .A1(n12756), .A2(n12755), .ZN(n12847) );
  INV_X1 U15935 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16302) );
  INV_X1 U15936 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16301) );
  INV_X1 U15937 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15205) );
  NAND3_X1 U15938 ( .A1(n16302), .A2(n16301), .A3(n15205), .ZN(n14999) );
  INV_X1 U15939 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15190) );
  INV_X1 U15940 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15001) );
  NAND2_X1 U15941 ( .A1(n15190), .A2(n15001), .ZN(n15181) );
  XNOR2_X1 U15942 ( .A(n12758), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15167) );
  NAND2_X1 U15943 ( .A1(n20692), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12760) );
  NAND2_X1 U15944 ( .A1(n13361), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12759) );
  NAND2_X1 U15945 ( .A1(n12760), .A2(n12759), .ZN(n12772) );
  NAND2_X1 U15946 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20721), .ZN(
        n12778) );
  NAND2_X1 U15947 ( .A1(n12774), .A2(n12760), .ZN(n12770) );
  NAND2_X1 U15948 ( .A1(n12770), .A2(n12761), .ZN(n12764) );
  NAND2_X1 U15949 ( .A1(n12762), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12763) );
  NAND2_X1 U15950 ( .A1(n12764), .A2(n12763), .ZN(n12768) );
  XNOR2_X1 U15951 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U15952 ( .A1(n12768), .A2(n12767), .ZN(n12766) );
  NAND2_X1 U15953 ( .A1(n21034), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12765) );
  NAND2_X1 U15954 ( .A1(n12766), .A2(n12765), .ZN(n12799) );
  NOR3_X1 U15955 ( .A1(n12799), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n20456), .ZN(n13084) );
  XNOR2_X1 U15956 ( .A(n12768), .B(n12767), .ZN(n13081) );
  INV_X1 U15957 ( .A(n13081), .ZN(n12769) );
  NOR2_X1 U15958 ( .A1(n12806), .A2(n12769), .ZN(n12794) );
  MUX2_X1 U15959 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n12762), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12771) );
  XOR2_X1 U15960 ( .A(n12771), .B(n12770), .Z(n13083) );
  NAND2_X1 U15961 ( .A1(n13498), .A2(n14265), .ZN(n12775) );
  NAND2_X1 U15962 ( .A1(n12772), .A2(n12778), .ZN(n12773) );
  NAND2_X1 U15963 ( .A1(n12774), .A2(n12773), .ZN(n13082) );
  AOI22_X1 U15964 ( .A1(n12776), .A2(n12775), .B1(n12788), .B2(n13082), .ZN(
        n12787) );
  INV_X1 U15965 ( .A(n13082), .ZN(n12777) );
  NOR2_X1 U15966 ( .A1(n12795), .A2(n12777), .ZN(n12786) );
  OAI21_X1 U15967 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20721), .A(
        n12778), .ZN(n12781) );
  INV_X1 U15968 ( .A(n12781), .ZN(n12779) );
  OAI21_X1 U15969 ( .B1(n12780), .B2(n14002), .A(n12779), .ZN(n12784) );
  OAI21_X1 U15970 ( .B1(n12782), .B2(n12781), .A(n12806), .ZN(n12783) );
  OAI21_X1 U15971 ( .B1(n12784), .B2(n12792), .A(n12783), .ZN(n12785) );
  AOI222_X1 U15972 ( .A1(n12787), .A2(n12786), .B1(n12787), .B2(n12785), .C1(
        n12786), .C2(n12785), .ZN(n12791) );
  AND2_X1 U15973 ( .A1(n12788), .A2(n13083), .ZN(n12789) );
  AOI21_X1 U15974 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21045), .A(
        n12797), .ZN(n12804) );
  INV_X1 U15975 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13319) );
  NOR2_X1 U15976 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13319), .ZN(
        n12798) );
  OR2_X1 U15977 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20456), .ZN(
        n12800) );
  NAND2_X1 U15978 ( .A1(n12805), .A2(n12802), .ZN(n12803) );
  NAND2_X1 U15979 ( .A1(n12804), .A2(n12803), .ZN(n12808) );
  NAND2_X1 U15980 ( .A1(n15302), .A2(n14002), .ZN(n12809) );
  AND3_X1 U15981 ( .A1(n12809), .A2(n13209), .A3(n13521), .ZN(n13306) );
  NAND2_X1 U15982 ( .A1(n13306), .A2(n13344), .ZN(n16140) );
  OR2_X1 U15983 ( .A1(n20944), .A2(n21045), .ZN(n20276) );
  OR2_X1 U15984 ( .A1(n16140), .A2(n20276), .ZN(n12810) );
  NOR2_X1 U15985 ( .A1(n15167), .A2(n20282), .ZN(n12819) );
  INV_X1 U15986 ( .A(n20889), .ZN(n20883) );
  AND2_X1 U15987 ( .A1(n12812), .A2(n20883), .ZN(n21048) );
  OR2_X1 U15988 ( .A1(n21048), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12811) );
  INV_X1 U15989 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12854) );
  OR2_X1 U15990 ( .A1(n12812), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16406) );
  INV_X2 U15991 ( .A(n16406), .ZN(n16391) );
  NAND2_X1 U15992 ( .A1(n16391), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15159) );
  OAI21_X1 U15993 ( .B1(n16260), .B2(n12854), .A(n15159), .ZN(n12813) );
  INV_X1 U15994 ( .A(n12813), .ZN(n12817) );
  NAND2_X1 U15995 ( .A1(n21045), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12815) );
  NAND2_X1 U15996 ( .A1(n21172), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U15997 ( .A1(n12815), .A2(n12814), .ZN(n13492) );
  NAND2_X1 U15998 ( .A1(n12817), .A2(n12816), .ZN(n12818) );
  AOI21_X1 U15999 ( .B1(n12821), .B2(n15573), .A(n19394), .ZN(n12822) );
  NAND2_X1 U16000 ( .A1(n15356), .A2(n12823), .ZN(n12824) );
  NAND2_X1 U16001 ( .A1(n12826), .A2(n12827), .ZN(n12828) );
  NAND2_X1 U16002 ( .A1(n19545), .A2(n16701), .ZN(n12834) );
  INV_X1 U16003 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12830) );
  AND2_X1 U16004 ( .A1(n12830), .A2(n12978), .ZN(n12831) );
  NAND2_X1 U16005 ( .A1(n12832), .A2(n12831), .ZN(n12833) );
  NAND2_X1 U16006 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19406), .ZN(n12836) );
  AOI22_X1 U16007 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19431), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19402), .ZN(n12835) );
  OAI211_X1 U16008 ( .C1(n15768), .C2(n19408), .A(n12836), .B(n12835), .ZN(
        n12837) );
  AOI21_X1 U16009 ( .B1(n15766), .B2(n19425), .A(n12837), .ZN(n12841) );
  NAND2_X1 U16010 ( .A1(n11616), .A2(n12839), .ZN(n12840) );
  OAI21_X1 U16011 ( .B1(n12844), .B2(n12843), .A(n12842), .ZN(P2_U2825) );
  INV_X1 U16012 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15137) );
  NAND2_X1 U16013 ( .A1(n15018), .A2(n12846), .ZN(n12850) );
  NOR2_X1 U16014 ( .A1(n12847), .A2(n15137), .ZN(n12848) );
  OAI21_X1 U16015 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15137), .A(
        n12851), .ZN(n12853) );
  XNOR2_X1 U16016 ( .A(n12853), .B(n12852), .ZN(n15158) );
  INV_X1 U16017 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12856) );
  XNOR2_X1 U16018 ( .A(n12857), .B(n12856), .ZN(n13685) );
  INV_X1 U16019 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21165) );
  NOR2_X1 U16020 ( .A1(n16406), .A2(n21165), .ZN(n15139) );
  AOI21_X1 U16021 ( .B1(n16291), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15139), .ZN(n12858) );
  OAI21_X1 U16022 ( .B1(n16299), .B2(n13685), .A(n12858), .ZN(n12859) );
  NAND2_X1 U16023 ( .A1(n14679), .A2(n12860), .ZN(n12865) );
  AOI22_X1 U16024 ( .A1(n12862), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12861), .ZN(n12863) );
  NAND2_X1 U16025 ( .A1(n14651), .A2(n16286), .ZN(n12866) );
  OAI211_X1 U16026 ( .C1(n15158), .C2(n20282), .A(n12867), .B(n12866), .ZN(
        P1_U2968) );
  AOI21_X1 U16027 ( .B1(n12869), .B2(n12868), .A(n18567), .ZN(n12879) );
  AOI21_X1 U16028 ( .B1(n12872), .B2(n12871), .A(n12870), .ZN(n12873) );
  NOR2_X1 U16029 ( .A1(n12874), .A2(n12873), .ZN(n16105) );
  NAND2_X1 U16030 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19079), .ZN(n19220) );
  NAND2_X1 U16031 ( .A1(n19151), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19144) );
  INV_X1 U16032 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19073) );
  INV_X1 U16033 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19081) );
  NAND2_X1 U16034 ( .A1(n19073), .A2(n19081), .ZN(n16861) );
  NAND3_X1 U16035 ( .A1(n19079), .A2(n19137), .A3(n16861), .ZN(n19210) );
  INV_X1 U16036 ( .A(n19210), .ZN(n16103) );
  AOI21_X1 U16037 ( .B1(n19212), .B2(n18557), .A(n16103), .ZN(n12876) );
  NAND2_X1 U16038 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19213) );
  INV_X1 U16039 ( .A(n19213), .ZN(n19208) );
  AOI21_X1 U16040 ( .B1(n12876), .B2(n12875), .A(n19208), .ZN(n16863) );
  NAND3_X1 U16041 ( .A1(n18986), .A2(n16863), .A3(n12877), .ZN(n12878) );
  OAI211_X1 U16042 ( .C1(n12879), .C2(n18991), .A(n16105), .B(n12878), .ZN(
        n12882) );
  INV_X1 U16043 ( .A(n12880), .ZN(n18988) );
  NAND2_X1 U16044 ( .A1(n12883), .A2(n9631), .ZN(n12900) );
  NAND2_X1 U16045 ( .A1(n17713), .A2(n18525), .ZN(n18431) );
  NOR2_X1 U16046 ( .A1(n18440), .A2(n18510), .ZN(n18515) );
  NAND2_X1 U16047 ( .A1(n19007), .A2(n18400), .ZN(n18472) );
  NOR3_X1 U16048 ( .A1(n18132), .A2(n18457), .A3(n18442), .ZN(n18313) );
  NAND3_X1 U16049 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18441) );
  NAND2_X1 U16050 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18471) );
  NOR2_X1 U16051 ( .A1(n18441), .A2(n18471), .ZN(n18437) );
  NAND2_X1 U16052 ( .A1(n18313), .A2(n18437), .ZN(n18414) );
  NOR2_X1 U16053 ( .A1(n9880), .A2(n18414), .ZN(n18212) );
  INV_X1 U16054 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18228) );
  NAND3_X1 U16055 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17887) );
  NOR2_X1 U16056 ( .A1(n18228), .A2(n17887), .ZN(n16715) );
  NAND3_X1 U16057 ( .A1(n18213), .A2(n18212), .A3(n16715), .ZN(n12888) );
  AOI21_X1 U16058 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18498) );
  NOR2_X1 U16059 ( .A1(n18498), .A2(n18441), .ZN(n18438) );
  NAND2_X1 U16060 ( .A1(n18438), .A2(n18313), .ZN(n18376) );
  NOR2_X1 U16061 ( .A1(n9880), .A2(n18376), .ZN(n18319) );
  INV_X1 U16062 ( .A(n18319), .ZN(n18253) );
  NOR2_X1 U16063 ( .A1(n12884), .A2(n18253), .ZN(n18236) );
  NAND2_X1 U16064 ( .A1(n18215), .A2(n18236), .ZN(n12889) );
  AND2_X1 U16065 ( .A1(n12889), .A2(n18992), .ZN(n18217) );
  AOI21_X1 U16066 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n18400), .ZN(n12885) );
  AOI211_X1 U16067 ( .C1(n18472), .C2(n12888), .A(n18217), .B(n12885), .ZN(
        n16117) );
  OAI21_X1 U16068 ( .B1(n18440), .B2(n16173), .A(n16117), .ZN(n12886) );
  INV_X2 U16069 ( .A(n18522), .ZN(n18483) );
  AOI21_X1 U16070 ( .B1(n18521), .B2(n12886), .A(n18520), .ZN(n16178) );
  NAND2_X1 U16071 ( .A1(n16173), .A2(n12887), .ZN(n12891) );
  AOI21_X1 U16072 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19015), .A(
        n19002), .ZN(n18491) );
  OAI22_X1 U16073 ( .A1(n19023), .A2(n12889), .B1(n12888), .B2(n18491), .ZN(
        n12890) );
  NAND2_X1 U16074 ( .A1(n18521), .A2(n12890), .ZN(n16119) );
  OAI22_X1 U16075 ( .A1(n16178), .A2(n19172), .B1(n12891), .B2(n16119), .ZN(
        n12892) );
  AOI211_X1 U16076 ( .C1(n10301), .C2(n18515), .A(n12893), .B(n12892), .ZN(
        n12896) );
  NOR2_X1 U16077 ( .A1(n18501), .A2(n18510), .ZN(n18527) );
  NAND2_X1 U16078 ( .A1(n12894), .A2(n18527), .ZN(n12895) );
  OAI211_X1 U16079 ( .C1(n12897), .C2(n18431), .A(n12896), .B(n12895), .ZN(
        n12898) );
  INV_X1 U16080 ( .A(n12898), .ZN(n12899) );
  NAND2_X1 U16081 ( .A1(n12900), .A2(n12899), .ZN(P3_U2831) );
  NOR4_X1 U16082 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12904) );
  NOR4_X1 U16083 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12903) );
  NOR4_X1 U16084 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12902) );
  NOR4_X1 U16085 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12901) );
  AND4_X1 U16086 ( .A1(n12904), .A2(n12903), .A3(n12902), .A4(n12901), .ZN(
        n12909) );
  NOR4_X1 U16087 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12907) );
  NOR4_X1 U16088 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12906) );
  NOR4_X1 U16089 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12905) );
  INV_X1 U16090 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20962) );
  AND4_X1 U16091 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n20962), .ZN(
        n12908) );
  NAND2_X1 U16092 ( .A1(n12909), .A2(n12908), .ZN(n12910) );
  AND2_X2 U16093 ( .A1(n12910), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14923)
         );
  INV_X1 U16094 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21093) );
  NOR3_X1 U16095 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21093), .ZN(n12912) );
  NOR4_X1 U16096 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12911)
         );
  NAND4_X1 U16097 ( .A1(n14923), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12912), .A4(
        n12911), .ZN(U214) );
  NOR4_X1 U16098 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12916) );
  NOR4_X1 U16099 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12915) );
  NOR4_X1 U16100 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12914) );
  NOR4_X1 U16101 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12913) );
  NAND4_X1 U16102 ( .A1(n12916), .A2(n12915), .A3(n12914), .A4(n12913), .ZN(
        n12921) );
  NOR4_X1 U16103 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12919) );
  NOR4_X1 U16104 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12918) );
  NOR4_X1 U16105 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12917) );
  INV_X1 U16106 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20137) );
  NAND4_X1 U16107 ( .A1(n12919), .A2(n12918), .A3(n12917), .A4(n20137), .ZN(
        n12920) );
  OAI21_X1 U16108 ( .B1(n12921), .B2(n12920), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12922) );
  NOR2_X1 U16109 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12924) );
  NOR4_X1 U16110 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12923) );
  NAND4_X1 U16111 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12924), .A4(n12923), .ZN(n12925) );
  NOR2_X1 U16112 ( .A1(n14611), .A2(n12925), .ZN(n16760) );
  NAND2_X1 U16113 ( .A1(n16760), .A2(U214), .ZN(U212) );
  NOR2_X1 U16114 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12925), .ZN(n16845)
         );
  AOI211_X1 U16115 ( .C1(n15664), .C2(n12927), .A(n12926), .B(n19394), .ZN(
        n12940) );
  OAI22_X1 U16116 ( .A1(n15666), .A2(n19386), .B1(n20157), .B2(n19416), .ZN(
        n12939) );
  INV_X1 U16117 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12928) );
  OAI22_X1 U16118 ( .A1(n12929), .A2(n19423), .B1(n19418), .B2(n12928), .ZN(
        n12938) );
  AOI21_X1 U16119 ( .B1(n12931), .B2(n15454), .A(n12930), .ZN(n15891) );
  INV_X1 U16120 ( .A(n15891), .ZN(n12936) );
  OR2_X1 U16121 ( .A1(n15907), .A2(n12932), .ZN(n12935) );
  INV_X1 U16122 ( .A(n12933), .ZN(n12934) );
  NAND2_X1 U16123 ( .A1(n12935), .A2(n12934), .ZN(n15886) );
  OAI22_X1 U16124 ( .A1(n12936), .A2(n19389), .B1(n15886), .B2(n19408), .ZN(
        n12937) );
  OR4_X1 U16125 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        P2_U2834) );
  AOI211_X1 U16126 ( .C1(n12943), .C2(n12942), .A(n12941), .B(n19394), .ZN(
        n12953) );
  INV_X1 U16127 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12944) );
  OAI22_X1 U16128 ( .A1(n12944), .A2(n19386), .B1(n10965), .B2(n19416), .ZN(
        n12952) );
  INV_X1 U16129 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12945) );
  OAI22_X1 U16130 ( .A1(n12946), .A2(n19423), .B1(n19418), .B2(n12945), .ZN(
        n12951) );
  OR2_X1 U16131 ( .A1(n12930), .A2(n12947), .ZN(n12948) );
  AND2_X1 U16132 ( .A1(n12948), .A2(n12959), .ZN(n16492) );
  INV_X1 U16133 ( .A(n16492), .ZN(n12949) );
  XNOR2_X1 U16134 ( .A(n12962), .B(n12933), .ZN(n15878) );
  OAI22_X1 U16135 ( .A1(n12949), .A2(n19389), .B1(n19408), .B2(n15878), .ZN(
        n12950) );
  OR4_X1 U16136 ( .A1(n12953), .A2(n12952), .A3(n12951), .A4(n12950), .ZN(
        P2_U2833) );
  AOI211_X1 U16137 ( .C1(n15647), .C2(n12955), .A(n12954), .B(n19394), .ZN(
        n12969) );
  OAI22_X1 U16138 ( .A1(n15645), .A2(n19386), .B1(n20160), .B2(n19416), .ZN(
        n12968) );
  INV_X1 U16139 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12956) );
  OAI22_X1 U16140 ( .A1(n12957), .A2(n19423), .B1(n19418), .B2(n12956), .ZN(
        n12967) );
  NAND2_X1 U16141 ( .A1(n12959), .A2(n12958), .ZN(n12960) );
  NAND2_X1 U16142 ( .A1(n15432), .A2(n12960), .ZN(n15862) );
  INV_X1 U16143 ( .A(n12961), .ZN(n12964) );
  NAND2_X1 U16144 ( .A1(n12962), .A2(n12933), .ZN(n12963) );
  NAND2_X1 U16145 ( .A1(n12964), .A2(n12963), .ZN(n12965) );
  NAND2_X1 U16146 ( .A1(n9777), .A2(n12965), .ZN(n15859) );
  OAI22_X1 U16147 ( .A1(n15862), .A2(n19389), .B1(n19408), .B2(n15859), .ZN(
        n12966) );
  OR4_X1 U16148 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        P2_U2832) );
  NOR2_X1 U16149 ( .A1(n10673), .A2(n19237), .ZN(n13222) );
  AND2_X1 U16150 ( .A1(n16672), .A2(n13222), .ZN(n19428) );
  INV_X1 U16151 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20273) );
  INV_X1 U16152 ( .A(n12978), .ZN(n12971) );
  INV_X1 U16153 ( .A(n12974), .ZN(n12970) );
  OAI211_X1 U16154 ( .C1(n19428), .C2(n20273), .A(n12971), .B(n12970), .ZN(
        P2_U2814) );
  INV_X1 U16155 ( .A(n12972), .ZN(n12977) );
  INV_X1 U16156 ( .A(n20253), .ZN(n12976) );
  OAI21_X1 U16157 ( .B1(n12974), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n12976), 
        .ZN(n12975) );
  OAI21_X1 U16158 ( .B1(n12977), .B2(n12976), .A(n12975), .ZN(P2_U3612) );
  OAI21_X1 U16159 ( .B1(n10493), .B2(n20257), .A(n12978), .ZN(n19544) );
  AOI22_X1 U16160 ( .A1(n19545), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n19544), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n12980) );
  NAND3_X1 U16161 ( .A1(n12978), .A2(n20257), .A3(n16700), .ZN(n13019) );
  INV_X1 U16162 ( .A(n13019), .ZN(n19547) );
  AOI22_X1 U16163 ( .A1(n14116), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14611), .ZN(n19616) );
  INV_X1 U16164 ( .A(n19616), .ZN(n12979) );
  NAND2_X1 U16165 ( .A1(n19547), .A2(n12979), .ZN(n13097) );
  NAND2_X1 U16166 ( .A1(n12980), .A2(n13097), .ZN(P2_U2974) );
  INV_X1 U16167 ( .A(n19544), .ZN(n13020) );
  AOI22_X1 U16168 ( .A1(n19545), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13113), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n12982) );
  AOI22_X1 U16169 ( .A1(n14116), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14611), .ZN(n19598) );
  INV_X1 U16170 ( .A(n19598), .ZN(n12981) );
  NAND2_X1 U16171 ( .A1(n19547), .A2(n12981), .ZN(n13103) );
  NAND2_X1 U16172 ( .A1(n12982), .A2(n13103), .ZN(P2_U2972) );
  AOI22_X1 U16173 ( .A1(P2_EAX_REG_18__SCAN_IN), .A2(n19545), .B1(n13113), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n12983) );
  INV_X1 U16174 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16811) );
  INV_X1 U16175 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18556) );
  AOI22_X1 U16176 ( .A1(n14116), .A2(n16811), .B1(n18556), .B2(n14611), .ZN(
        n16484) );
  INV_X1 U16177 ( .A(n16484), .ZN(n19583) );
  OR2_X1 U16178 ( .A1(n13019), .A2(n19583), .ZN(n13000) );
  NAND2_X1 U16179 ( .A1(n12983), .A2(n13000), .ZN(P2_U2954) );
  AOI22_X1 U16180 ( .A1(P2_EAX_REG_16__SCAN_IN), .A2(n19545), .B1(n13113), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16181 ( .A1(n14116), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14611), .ZN(n19504) );
  INV_X1 U16182 ( .A(n19504), .ZN(n12984) );
  NAND2_X1 U16183 ( .A1(n19547), .A2(n12984), .ZN(n13105) );
  NAND2_X1 U16184 ( .A1(n12985), .A2(n13105), .ZN(P2_U2952) );
  AOI22_X1 U16185 ( .A1(P2_EAX_REG_20__SCAN_IN), .A2(n19545), .B1(n13113), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n12986) );
  OAI22_X1 U16186 ( .A1(n14611), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14116), .ZN(n19480) );
  INV_X1 U16187 ( .A(n19480), .ZN(n16479) );
  NAND2_X1 U16188 ( .A1(n19547), .A2(n16479), .ZN(n13004) );
  NAND2_X1 U16189 ( .A1(n12986), .A2(n13004), .ZN(P2_U2956) );
  AOI22_X1 U16190 ( .A1(P2_EAX_REG_22__SCAN_IN), .A2(n19545), .B1(n13113), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16191 ( .A1(n14116), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14611), .ZN(n19604) );
  INV_X1 U16192 ( .A(n19604), .ZN(n12987) );
  NAND2_X1 U16193 ( .A1(n19547), .A2(n12987), .ZN(n12998) );
  NAND2_X1 U16194 ( .A1(n12988), .A2(n12998), .ZN(P2_U2958) );
  AOI22_X1 U16195 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n19545), .B1(n13113), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12992) );
  INV_X1 U16196 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16797) );
  OR2_X1 U16197 ( .A1(n14611), .A2(n16797), .ZN(n12990) );
  NAND2_X1 U16198 ( .A1(n14611), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12989) );
  AND2_X1 U16199 ( .A1(n12990), .A2(n12989), .ZN(n19456) );
  INV_X1 U16200 ( .A(n19456), .ZN(n12991) );
  NAND2_X1 U16201 ( .A1(n19547), .A2(n12991), .ZN(n13095) );
  NAND2_X1 U16202 ( .A1(n12992), .A2(n13095), .ZN(P2_U2961) );
  AOI22_X1 U16203 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(n19545), .B1(n13113), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12997) );
  INV_X1 U16204 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12993) );
  OR2_X1 U16205 ( .A1(n14611), .A2(n12993), .ZN(n12995) );
  NAND2_X1 U16206 ( .A1(n14611), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12994) );
  AND2_X1 U16207 ( .A1(n12995), .A2(n12994), .ZN(n19451) );
  INV_X1 U16208 ( .A(n19451), .ZN(n12996) );
  NAND2_X1 U16209 ( .A1(n19547), .A2(n12996), .ZN(n13109) );
  NAND2_X1 U16210 ( .A1(n12997), .A2(n13109), .ZN(P2_U2963) );
  AOI22_X1 U16211 ( .A1(n19545), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13113), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16212 ( .A1(n12999), .A2(n12998), .ZN(P2_U2973) );
  AOI22_X1 U16213 ( .A1(n19545), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13113), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13001) );
  NAND2_X1 U16214 ( .A1(n13001), .A2(n13000), .ZN(P2_U2969) );
  AOI22_X1 U16215 ( .A1(n19545), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13113), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U16216 ( .A1(n14116), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14611), .ZN(n19587) );
  INV_X1 U16217 ( .A(n19587), .ZN(n13002) );
  NAND2_X1 U16218 ( .A1(n19547), .A2(n13002), .ZN(n13091) );
  NAND2_X1 U16219 ( .A1(n13003), .A2(n13091), .ZN(P2_U2970) );
  AOI22_X1 U16220 ( .A1(n19545), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13113), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U16221 ( .A1(n13005), .A2(n13004), .ZN(P2_U2971) );
  AOI22_X1 U16222 ( .A1(n19545), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13113), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13008) );
  INV_X1 U16223 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16790) );
  NOR2_X1 U16224 ( .A1(n14611), .A2(n16790), .ZN(n13006) );
  AOI21_X1 U16225 ( .B1(n14611), .B2(BUF2_REG_13__SCAN_IN), .A(n13006), .ZN(
        n19446) );
  INV_X1 U16226 ( .A(n19446), .ZN(n13007) );
  NAND2_X1 U16227 ( .A1(n19547), .A2(n13007), .ZN(n13111) );
  NAND2_X1 U16228 ( .A1(n13008), .A2(n13111), .ZN(P2_U2980) );
  INV_X1 U16229 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13243) );
  NAND2_X1 U16230 ( .A1(n14611), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13010) );
  INV_X1 U16231 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16795) );
  OR2_X1 U16232 ( .A1(n14611), .A2(n16795), .ZN(n13009) );
  NAND2_X1 U16233 ( .A1(n13010), .A2(n13009), .ZN(n19453) );
  NAND2_X1 U16234 ( .A1(n19547), .A2(n19453), .ZN(n13013) );
  NAND2_X1 U16235 ( .A1(n19544), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13011) );
  OAI211_X1 U16236 ( .C1(n13223), .C2(n13243), .A(n13013), .B(n13011), .ZN(
        P2_U2962) );
  INV_X1 U16237 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19521) );
  NAND2_X1 U16238 ( .A1(n19544), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13012) );
  OAI211_X1 U16239 ( .C1(n13223), .C2(n19521), .A(n13013), .B(n13012), .ZN(
        P2_U2977) );
  INV_X1 U16240 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19525) );
  NAND2_X1 U16241 ( .A1(n14611), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13015) );
  INV_X1 U16242 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16799) );
  OR2_X1 U16243 ( .A1(n14611), .A2(n16799), .ZN(n13014) );
  NAND2_X1 U16244 ( .A1(n13015), .A2(n13014), .ZN(n19460) );
  NAND2_X1 U16245 ( .A1(n19547), .A2(n19460), .ZN(n13018) );
  NAND2_X1 U16246 ( .A1(n19544), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13016) );
  OAI211_X1 U16247 ( .C1(n13223), .C2(n19525), .A(n13018), .B(n13016), .ZN(
        P2_U2975) );
  INV_X1 U16248 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13245) );
  NAND2_X1 U16249 ( .A1(n19544), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13017) );
  OAI211_X1 U16250 ( .C1(n13223), .C2(n13245), .A(n13018), .B(n13017), .ZN(
        P2_U2960) );
  INV_X1 U16251 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13022) );
  INV_X1 U16252 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16253 ( .A1(n14116), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14611), .ZN(n19441) );
  OAI222_X1 U16254 ( .A1(n13022), .A2(n13223), .B1(n13021), .B2(n13020), .C1(
        n13019), .C2(n19441), .ZN(P2_U2982) );
  NAND2_X1 U16255 ( .A1(n13023), .A2(n13024), .ZN(n16666) );
  OR2_X1 U16256 ( .A1(n16668), .A2(n16666), .ZN(n13060) );
  INV_X1 U16257 ( .A(n13043), .ZN(n16656) );
  NAND3_X1 U16258 ( .A1(n16672), .A2(n13117), .A3(n16656), .ZN(n13036) );
  NAND2_X1 U16259 ( .A1(n10479), .A2(n10493), .ZN(n13038) );
  NAND2_X1 U16260 ( .A1(n13038), .A2(n16663), .ZN(n13025) );
  NAND2_X1 U16261 ( .A1(n13025), .A2(n19614), .ZN(n13026) );
  AOI21_X1 U16262 ( .B1(n13026), .B2(n10499), .A(n10463), .ZN(n13033) );
  NAND2_X1 U16263 ( .A1(n13027), .A2(n10499), .ZN(n13028) );
  NAND2_X1 U16264 ( .A1(n10673), .A2(n13028), .ZN(n13032) );
  NAND2_X1 U16265 ( .A1(n13029), .A2(n19614), .ZN(n13031) );
  NAND2_X1 U16266 ( .A1(n13031), .A2(n13030), .ZN(n13139) );
  NAND4_X1 U16267 ( .A1(n13034), .A2(n13033), .A3(n13032), .A4(n13139), .ZN(
        n13039) );
  INV_X1 U16268 ( .A(n13039), .ZN(n13035) );
  NAND2_X1 U16269 ( .A1(n13036), .A2(n13035), .ZN(n13120) );
  INV_X1 U16270 ( .A(n13120), .ZN(n13037) );
  NAND2_X1 U16271 ( .A1(n13060), .A2(n13037), .ZN(n13042) );
  NAND2_X1 U16272 ( .A1(n16668), .A2(n13136), .ZN(n13041) );
  AND2_X1 U16273 ( .A1(n12972), .A2(n20257), .ZN(n16655) );
  NAND2_X1 U16274 ( .A1(n16654), .A2(n16655), .ZN(n13040) );
  NAND2_X1 U16275 ( .A1(n13041), .A2(n13040), .ZN(n13331) );
  NOR2_X1 U16276 ( .A1(n13042), .A2(n13331), .ZN(n13045) );
  NAND2_X1 U16277 ( .A1(n16668), .A2(n16700), .ZN(n13225) );
  OR2_X1 U16278 ( .A1(n13225), .A2(n13043), .ZN(n13125) );
  OR2_X1 U16279 ( .A1(n13125), .A2(n10673), .ZN(n13044) );
  NAND2_X1 U16280 ( .A1(n13045), .A2(n13044), .ZN(n16685) );
  NAND2_X1 U16281 ( .A1(n16685), .A2(n13332), .ZN(n13047) );
  NOR2_X1 U16282 ( .A1(n20256), .A2(n20231), .ZN(n16699) );
  AOI22_X1 U16283 ( .A1(n20256), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(
        P2_FLUSH_REG_SCAN_IN), .B2(n16699), .ZN(n13046) );
  NAND2_X1 U16284 ( .A1(n13047), .A2(n13046), .ZN(n20192) );
  AND4_X1 U16285 ( .A1(n10484), .A2(n16659), .A3(n20198), .A4(n16658), .ZN(
        n13048) );
  NAND2_X1 U16286 ( .A1(n20192), .A2(n13048), .ZN(n13049) );
  OAI21_X1 U16287 ( .B1(n20192), .B2(n16675), .A(n13049), .ZN(P2_U3595) );
  NAND2_X1 U16288 ( .A1(n19603), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13051) );
  NAND2_X1 U16289 ( .A1(n13051), .A2(n20205), .ZN(n13276) );
  AOI22_X1 U16290 ( .A1(n13276), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20196), .B2(n20239), .ZN(n13052) );
  NOR2_X1 U16291 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13055) );
  OAI211_X1 U16292 ( .C1(n13056), .C2(n13055), .A(P2_STATE2_REG_0__SCAN_IN), 
        .B(n13054), .ZN(n13057) );
  INV_X1 U16293 ( .A(n13057), .ZN(n13058) );
  NAND2_X1 U16294 ( .A1(n13060), .A2(n13384), .ZN(n13061) );
  MUX2_X1 U16295 ( .A(n13162), .B(n19417), .S(n15448), .Z(n13062) );
  OAI21_X1 U16296 ( .B1(n20234), .B2(n15479), .A(n13062), .ZN(P2_U2887) );
  INV_X1 U16297 ( .A(n16586), .ZN(n19552) );
  AOI21_X1 U16298 ( .B1(n13149), .B2(n19422), .A(n13063), .ZN(n13168) );
  OAI21_X1 U16299 ( .B1(n13065), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13064), .ZN(n13165) );
  OR2_X1 U16300 ( .A1(n19333), .A2(n19251), .ZN(n13161) );
  OAI21_X1 U16301 ( .B1(n16584), .B2(n13165), .A(n13161), .ZN(n13066) );
  AOI21_X1 U16302 ( .B1(n19552), .B2(n13168), .A(n13066), .ZN(n13069) );
  OAI21_X1 U16303 ( .B1(n19551), .B2(n13067), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13068) );
  OAI211_X1 U16304 ( .C1(n19559), .C2(n13162), .A(n13069), .B(n13068), .ZN(
        P2_U3014) );
  OAI21_X1 U16305 ( .B1(n19404), .B2(n13071), .A(n13070), .ZN(n13072) );
  XNOR2_X1 U16306 ( .A(n13072), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13158) );
  OAI21_X1 U16307 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13074), .A(
        n13073), .ZN(n13131) );
  NOR2_X1 U16308 ( .A1(n19333), .A2(n10459), .ZN(n13157) );
  INV_X1 U16309 ( .A(n13157), .ZN(n13075) );
  OAI21_X1 U16310 ( .B1(n16584), .B2(n13131), .A(n13075), .ZN(n13078) );
  MUX2_X1 U16311 ( .A(n19551), .B(n16583), .S(n13076), .Z(n13077) );
  AOI211_X1 U16312 ( .C1(n19552), .C2(n13158), .A(n13078), .B(n13077), .ZN(
        n13079) );
  OAI21_X1 U16313 ( .B1(n13178), .B2(n19559), .A(n13079), .ZN(P2_U3013) );
  OR4_X1 U16314 ( .A1(n13084), .A2(n13083), .A3(n13082), .A4(n13081), .ZN(
        n13085) );
  NAND2_X1 U16315 ( .A1(n13086), .A2(n13085), .ZN(n13297) );
  NOR2_X1 U16316 ( .A1(n13297), .A2(n20276), .ZN(n13087) );
  NAND2_X1 U16317 ( .A1(n13080), .A2(n13087), .ZN(n13200) );
  INV_X1 U16318 ( .A(n13200), .ZN(n13090) );
  INV_X1 U16319 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21081) );
  NOR2_X1 U16320 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20883), .ZN(n13201) );
  INV_X1 U16321 ( .A(n13201), .ZN(n13089) );
  OAI211_X1 U16322 ( .C1(n13090), .C2(n21081), .A(n13248), .B(n13089), .ZN(
        P1_U2801) );
  AOI22_X1 U16323 ( .A1(n19545), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19544), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13092) );
  NAND2_X1 U16324 ( .A1(n13092), .A2(n13091), .ZN(P2_U2955) );
  AOI22_X1 U16325 ( .A1(n19545), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13113), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16326 ( .A1(n14116), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14611), .ZN(n19578) );
  INV_X1 U16327 ( .A(n19578), .ZN(n13093) );
  NAND2_X1 U16328 ( .A1(n19547), .A2(n13093), .ZN(n13107) );
  NAND2_X1 U16329 ( .A1(n13094), .A2(n13107), .ZN(P2_U2953) );
  AOI22_X1 U16330 ( .A1(n19545), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n19544), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13096) );
  NAND2_X1 U16331 ( .A1(n13096), .A2(n13095), .ZN(P2_U2976) );
  AOI22_X1 U16332 ( .A1(n19545), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13113), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13098) );
  NAND2_X1 U16333 ( .A1(n13098), .A2(n13097), .ZN(P2_U2959) );
  AOI22_X1 U16334 ( .A1(n19545), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n19544), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13102) );
  INV_X1 U16335 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16792) );
  OR2_X1 U16336 ( .A1(n14611), .A2(n16792), .ZN(n13100) );
  NAND2_X1 U16337 ( .A1(n14611), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13099) );
  AND2_X1 U16338 ( .A1(n13100), .A2(n13099), .ZN(n19449) );
  INV_X1 U16339 ( .A(n19449), .ZN(n13101) );
  NAND2_X1 U16340 ( .A1(n19547), .A2(n13101), .ZN(n13114) );
  NAND2_X1 U16341 ( .A1(n13102), .A2(n13114), .ZN(P2_U2979) );
  AOI22_X1 U16342 ( .A1(n19545), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13113), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13104) );
  NAND2_X1 U16343 ( .A1(n13104), .A2(n13103), .ZN(P2_U2957) );
  AOI22_X1 U16344 ( .A1(n19545), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n13113), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13106) );
  NAND2_X1 U16345 ( .A1(n13106), .A2(n13105), .ZN(P2_U2967) );
  AOI22_X1 U16346 ( .A1(n19545), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13113), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13108) );
  NAND2_X1 U16347 ( .A1(n13108), .A2(n13107), .ZN(P2_U2968) );
  AOI22_X1 U16348 ( .A1(n19545), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n19544), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13110) );
  NAND2_X1 U16349 ( .A1(n13110), .A2(n13109), .ZN(P2_U2978) );
  AOI22_X1 U16350 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n19545), .B1(n13113), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13112) );
  NAND2_X1 U16351 ( .A1(n13112), .A2(n13111), .ZN(P2_U2965) );
  AOI22_X1 U16352 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(n19545), .B1(n13113), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13115) );
  NAND2_X1 U16353 ( .A1(n13115), .A2(n13114), .ZN(P2_U2964) );
  MUX2_X1 U16354 ( .A(n13117), .B(n13116), .S(n10493), .Z(n13118) );
  AND3_X1 U16355 ( .A1(n16672), .A2(n13118), .A3(n20257), .ZN(n13119) );
  NOR2_X1 U16356 ( .A1(n13120), .A2(n13119), .ZN(n13124) );
  NAND2_X1 U16357 ( .A1(n16663), .A2(n13121), .ZN(n13122) );
  NAND3_X1 U16358 ( .A1(n13225), .A2(n10479), .A3(n13122), .ZN(n13123) );
  OAI211_X1 U16359 ( .C1(n13125), .C2(n10499), .A(n13124), .B(n13123), .ZN(
        n13126) );
  OR2_X1 U16360 ( .A1(n13127), .A2(n13126), .ZN(n13128) );
  NAND2_X1 U16361 ( .A1(n10503), .A2(n10493), .ZN(n13129) );
  NAND2_X1 U16362 ( .A1(n13129), .A2(n10508), .ZN(n13130) );
  INV_X1 U16363 ( .A(n13131), .ZN(n13152) );
  NAND2_X1 U16364 ( .A1(n16664), .A2(n16700), .ZN(n13132) );
  NAND2_X1 U16365 ( .A1(n16666), .A2(n13132), .ZN(n13133) );
  NAND2_X1 U16366 ( .A1(n13153), .A2(n13133), .ZN(n16624) );
  XNOR2_X1 U16367 ( .A(n13135), .B(n13134), .ZN(n20227) );
  INV_X1 U16368 ( .A(n20227), .ZN(n19409) );
  NOR2_X1 U16369 ( .A1(n16624), .A2(n19409), .ZN(n13151) );
  NOR2_X1 U16370 ( .A1(n13149), .A2(n13155), .ZN(n14625) );
  NAND2_X1 U16371 ( .A1(n13153), .A2(n13136), .ZN(n15944) );
  NAND2_X1 U16372 ( .A1(n13137), .A2(n12972), .ZN(n13147) );
  NAND2_X1 U16373 ( .A1(n13138), .A2(n16700), .ZN(n13921) );
  NAND2_X1 U16374 ( .A1(n13921), .A2(n13139), .ZN(n13140) );
  NAND2_X1 U16375 ( .A1(n13140), .A2(n10457), .ZN(n13145) );
  OAI22_X1 U16376 ( .A1(n12972), .A2(n10486), .B1(n10499), .B2(n16663), .ZN(
        n13141) );
  INV_X1 U16377 ( .A(n13141), .ZN(n13142) );
  AND2_X1 U16378 ( .A1(n13143), .A2(n13142), .ZN(n13144) );
  NAND2_X1 U16379 ( .A1(n13145), .A2(n13144), .ZN(n13146) );
  AOI21_X1 U16380 ( .B1(n13147), .B2(n10463), .A(n13146), .ZN(n16076) );
  NAND2_X1 U16381 ( .A1(n16076), .A2(n13384), .ZN(n13148) );
  NAND2_X1 U16382 ( .A1(n13153), .A2(n13148), .ZN(n15940) );
  AOI211_X1 U16383 ( .C1(n13155), .C2(n13149), .A(n14625), .B(n16609), .ZN(
        n13150) );
  AOI211_X1 U16384 ( .C1(n16646), .C2(n13152), .A(n13151), .B(n13150), .ZN(
        n13160) );
  NAND2_X2 U16385 ( .A1(n13153), .A2(n20245), .ZN(n16651) );
  INV_X1 U16386 ( .A(n16651), .ZN(n16600) );
  INV_X1 U16387 ( .A(n13153), .ZN(n13154) );
  NAND2_X1 U16388 ( .A1(n13154), .A2(n19333), .ZN(n14629) );
  NOR2_X1 U16389 ( .A1(n14629), .A2(n13155), .ZN(n13156) );
  AOI211_X1 U16390 ( .C1(n13158), .C2(n16600), .A(n13157), .B(n13156), .ZN(
        n13159) );
  OAI211_X1 U16391 ( .C1(n13178), .C2(n16629), .A(n13160), .B(n13159), .ZN(
        P2_U3045) );
  OAI21_X1 U16392 ( .B1(n16629), .B2(n13162), .A(n13161), .ZN(n13167) );
  XNOR2_X1 U16393 ( .A(n13163), .B(n13164), .ZN(n19415) );
  OAI22_X1 U16394 ( .A1(n16630), .A2(n13165), .B1(n16624), .B2(n19415), .ZN(
        n13166) );
  AOI211_X1 U16395 ( .C1(n16600), .C2(n13168), .A(n13167), .B(n13166), .ZN(
        n13170) );
  MUX2_X1 U16396 ( .A(n16609), .B(n14629), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13169) );
  NAND2_X1 U16397 ( .A1(n13170), .A2(n13169), .ZN(P2_U3046) );
  NAND2_X1 U16398 ( .A1(n14549), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13181) );
  NAND2_X1 U16399 ( .A1(n13276), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13172) );
  XNOR2_X1 U16400 ( .A(n20239), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13854) );
  NAND2_X1 U16401 ( .A1(n13854), .A2(n20196), .ZN(n19890) );
  NAND2_X1 U16402 ( .A1(n13172), .A2(n19890), .ZN(n13173) );
  NOR2_X1 U16403 ( .A1(n13178), .A2(n15448), .ZN(n13179) );
  AOI21_X1 U16404 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n15448), .A(n13179), .ZN(
        n13180) );
  OAI21_X1 U16405 ( .B1(n20222), .B2(n15479), .A(n13180), .ZN(P2_U2886) );
  INV_X1 U16406 ( .A(n13171), .ZN(n13925) );
  NAND2_X1 U16407 ( .A1(n13925), .A2(n13181), .ZN(n13182) );
  NAND2_X1 U16408 ( .A1(n14549), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13280) );
  NAND2_X1 U16409 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19917) );
  NAND2_X1 U16410 ( .A1(n19917), .A2(n20219), .ZN(n13185) );
  NAND2_X1 U16411 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20048) );
  INV_X1 U16412 ( .A(n20048), .ZN(n20042) );
  NAND2_X1 U16413 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20042), .ZN(
        n13272) );
  NAND2_X1 U16414 ( .A1(n13185), .A2(n13272), .ZN(n13855) );
  NOR2_X1 U16415 ( .A1(n20202), .A2(n13855), .ZN(n13186) );
  AOI21_X1 U16416 ( .B1(n13276), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13186), .ZN(n13279) );
  AND2_X1 U16417 ( .A1(n13280), .A2(n13279), .ZN(n13187) );
  NAND2_X1 U16418 ( .A1(n10183), .A2(n13187), .ZN(n13195) );
  INV_X1 U16419 ( .A(n13187), .ZN(n13188) );
  OAI22_X1 U16420 ( .A1(n13195), .A2(n13189), .B1(n10183), .B2(n13188), .ZN(
        n13190) );
  NAND2_X1 U16421 ( .A1(n11328), .A2(n13190), .ZN(n13194) );
  INV_X1 U16422 ( .A(n13279), .ZN(n13192) );
  OAI21_X1 U16423 ( .B1(n13192), .B2(n13270), .A(n13280), .ZN(n13191) );
  OAI21_X1 U16424 ( .B1(n13280), .B2(n13192), .A(n13191), .ZN(n13193) );
  NAND2_X1 U16425 ( .A1(n13282), .A2(n13281), .ZN(n13196) );
  MUX2_X1 U16426 ( .A(n13198), .B(n9675), .S(n15449), .Z(n13199) );
  OAI21_X1 U16427 ( .B1(n20210), .B2(n15479), .A(n13199), .ZN(P2_U2885) );
  OAI21_X1 U16428 ( .B1(n13201), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n21047), 
        .ZN(n13202) );
  OAI21_X1 U16429 ( .B1(n21047), .B2(n13203), .A(n13202), .ZN(P1_U3487) );
  INV_X1 U16430 ( .A(n13297), .ZN(n13204) );
  AOI21_X1 U16431 ( .B1(n13080), .B2(n13204), .A(n13423), .ZN(n13205) );
  AOI21_X1 U16432 ( .B1(n16159), .B2(n13212), .A(n13205), .ZN(n20275) );
  INV_X1 U16433 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U16434 ( .A1(n13207), .A2(n13206), .ZN(n16182) );
  NAND3_X1 U16435 ( .A1(n13212), .A2(n16182), .A3(n9653), .ZN(n13208) );
  NAND2_X1 U16436 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n16416) );
  NAND2_X1 U16437 ( .A1(n13208), .A2(n16416), .ZN(n21041) );
  AND2_X1 U16438 ( .A1(n20275), .A2(n21041), .ZN(n16138) );
  NOR2_X1 U16439 ( .A1(n16138), .A2(n20276), .ZN(n20284) );
  INV_X1 U16440 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21162) );
  INV_X1 U16441 ( .A(n13531), .ZN(n14652) );
  NAND2_X1 U16442 ( .A1(n14652), .A2(n13209), .ZN(n13210) );
  NOR2_X1 U16443 ( .A1(n13210), .A2(n15302), .ZN(n13302) );
  INV_X1 U16444 ( .A(n13302), .ZN(n13525) );
  OR2_X1 U16445 ( .A1(n16159), .A2(n13525), .ZN(n13219) );
  NAND2_X1 U16446 ( .A1(n13080), .A2(n13297), .ZN(n13218) );
  INV_X1 U16447 ( .A(n13423), .ZN(n13215) );
  NOR2_X1 U16448 ( .A1(n13212), .A2(n13211), .ZN(n13213) );
  AND2_X1 U16449 ( .A1(n13214), .A2(n13213), .ZN(n13513) );
  INV_X1 U16450 ( .A(n13513), .ZN(n13357) );
  NAND3_X1 U16451 ( .A1(n13215), .A2(n16140), .A3(n13357), .ZN(n13216) );
  NAND2_X1 U16452 ( .A1(n16159), .A2(n13216), .ZN(n13217) );
  AND3_X1 U16453 ( .A1(n13219), .A2(n13218), .A3(n13217), .ZN(n16141) );
  INV_X1 U16454 ( .A(n16141), .ZN(n13220) );
  NAND2_X1 U16455 ( .A1(n20284), .A2(n13220), .ZN(n13221) );
  OAI21_X1 U16456 ( .B1(n20284), .B2(n21162), .A(n13221), .ZN(P1_U3484) );
  INV_X1 U16457 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15534) );
  INV_X1 U16458 ( .A(n13222), .ZN(n13224) );
  OAI21_X1 U16459 ( .B1(n13225), .B2(n13224), .A(n13223), .ZN(n13226) );
  OR2_X1 U16460 ( .A1(n19542), .A2(n20263), .ZN(n19506) );
  OR2_X1 U16461 ( .A1(n20231), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13227) );
  INV_X2 U16462 ( .A(n13227), .ZN(n20255) );
  NAND2_X1 U16463 ( .A1(n19542), .A2(n13227), .ZN(n19509) );
  INV_X2 U16464 ( .A(n19509), .ZN(n19540) );
  AOI22_X1 U16465 ( .A1(n20255), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13228) );
  OAI21_X1 U16466 ( .B1(n15534), .B2(n19506), .A(n13228), .ZN(P2_U2928) );
  INV_X1 U16467 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15541) );
  AOI22_X1 U16468 ( .A1(n20255), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13229) );
  OAI21_X1 U16469 ( .B1(n15541), .B2(n19506), .A(n13229), .ZN(P2_U2929) );
  INV_X1 U16470 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15548) );
  AOI22_X1 U16471 ( .A1(n20255), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13230) );
  OAI21_X1 U16472 ( .B1(n15548), .B2(n19506), .A(n13230), .ZN(P2_U2930) );
  INV_X1 U16473 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13232) );
  AOI22_X1 U16474 ( .A1(n20255), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13231) );
  OAI21_X1 U16475 ( .B1(n13232), .B2(n19506), .A(n13231), .ZN(P2_U2931) );
  INV_X1 U16476 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15557) );
  AOI22_X1 U16477 ( .A1(n20255), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13233) );
  OAI21_X1 U16478 ( .B1(n15557), .B2(n19506), .A(n13233), .ZN(P2_U2932) );
  INV_X1 U16479 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U16480 ( .A1(n20255), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13234) );
  OAI21_X1 U16481 ( .B1(n13235), .B2(n19506), .A(n13234), .ZN(P2_U2933) );
  INV_X1 U16482 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U16483 ( .A1(n20255), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13236) );
  OAI21_X1 U16484 ( .B1(n14162), .B2(n19506), .A(n13236), .ZN(P2_U2934) );
  INV_X1 U16485 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14115) );
  AOI22_X1 U16486 ( .A1(n20255), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13237) );
  OAI21_X1 U16487 ( .B1(n14115), .B2(n19506), .A(n13237), .ZN(P2_U2935) );
  INV_X1 U16488 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U16489 ( .A1(n20255), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13238) );
  OAI21_X1 U16490 ( .B1(n15518), .B2(n19506), .A(n13238), .ZN(P2_U2926) );
  INV_X1 U16491 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15482) );
  AOI22_X1 U16492 ( .A1(n20255), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13239) );
  OAI21_X1 U16493 ( .B1(n15482), .B2(n19506), .A(n13239), .ZN(P2_U2922) );
  INV_X1 U16494 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15492) );
  AOI22_X1 U16495 ( .A1(n20255), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13240) );
  OAI21_X1 U16496 ( .B1(n15492), .B2(n19506), .A(n13240), .ZN(P2_U2923) );
  INV_X1 U16497 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15502) );
  AOI22_X1 U16498 ( .A1(n20255), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13241) );
  OAI21_X1 U16499 ( .B1(n15502), .B2(n19506), .A(n13241), .ZN(P2_U2924) );
  AOI22_X1 U16500 ( .A1(n20255), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13242) );
  OAI21_X1 U16501 ( .B1(n13243), .B2(n19506), .A(n13242), .ZN(P2_U2925) );
  AOI22_X1 U16502 ( .A1(n20255), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13244) );
  OAI21_X1 U16503 ( .B1(n13245), .B2(n19506), .A(n13244), .ZN(P2_U2927) );
  INV_X1 U16504 ( .A(n16416), .ZN(n21050) );
  AND2_X1 U16505 ( .A1(n13246), .A2(n21050), .ZN(n13247) );
  NAND2_X1 U16506 ( .A1(n13251), .A2(n13498), .ZN(n13393) );
  NAND2_X1 U16507 ( .A1(n13251), .A2(n13958), .ZN(n13252) );
  INV_X1 U16508 ( .A(DATAI_15_), .ZN(n13250) );
  INV_X1 U16509 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13249) );
  MUX2_X1 U16510 ( .A(n13250), .B(n13249), .S(n14923), .Z(n14976) );
  INV_X1 U16511 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20390) );
  OAI222_X1 U16512 ( .A1(n13393), .A2(n12239), .B1(n13252), .B2(n14976), .C1(
        n13251), .C2(n20390), .ZN(P1_U2967) );
  INV_X2 U16513 ( .A(n13251), .ZN(n20438) );
  AOI22_X1 U16514 ( .A1(n20439), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13255) );
  INV_X1 U16515 ( .A(DATAI_3_), .ZN(n13254) );
  NAND2_X1 U16516 ( .A1(n14923), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13253) );
  OAI21_X1 U16517 ( .B1(n14923), .B2(n13254), .A(n13253), .ZN(n14959) );
  NAND2_X1 U16518 ( .A1(n20426), .A2(n14959), .ZN(n13397) );
  NAND2_X1 U16519 ( .A1(n13255), .A2(n13397), .ZN(P1_U2955) );
  AOI22_X1 U16520 ( .A1(n20439), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13258) );
  INV_X1 U16521 ( .A(n14923), .ZN(n14263) );
  INV_X1 U16522 ( .A(DATAI_4_), .ZN(n21168) );
  NAND2_X1 U16523 ( .A1(n14263), .A2(n21168), .ZN(n13257) );
  INV_X1 U16524 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16807) );
  NAND2_X1 U16525 ( .A1(n14923), .A2(n16807), .ZN(n13256) );
  AND2_X1 U16526 ( .A1(n13257), .A2(n13256), .ZN(n15337) );
  NAND2_X1 U16527 ( .A1(n20426), .A2(n15337), .ZN(n13419) );
  NAND2_X1 U16528 ( .A1(n13258), .A2(n13419), .ZN(P1_U2956) );
  AOI22_X1 U16529 ( .A1(n20439), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13260) );
  INV_X1 U16530 ( .A(DATAI_7_), .ZN(n21221) );
  NAND2_X1 U16531 ( .A1(n14923), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13259) );
  OAI21_X1 U16532 ( .B1(n14923), .B2(n21221), .A(n13259), .ZN(n14939) );
  NAND2_X1 U16533 ( .A1(n20426), .A2(n14939), .ZN(n13421) );
  NAND2_X1 U16534 ( .A1(n13260), .A2(n13421), .ZN(P1_U2959) );
  AOI22_X1 U16535 ( .A1(n20439), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13263) );
  INV_X1 U16536 ( .A(DATAI_5_), .ZN(n21157) );
  NAND2_X1 U16537 ( .A1(n14263), .A2(n21157), .ZN(n13262) );
  INV_X1 U16538 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16805) );
  NAND2_X1 U16539 ( .A1(n14923), .A2(n16805), .ZN(n13261) );
  AND2_X1 U16540 ( .A1(n13262), .A2(n13261), .ZN(n14950) );
  NAND2_X1 U16541 ( .A1(n20426), .A2(n14950), .ZN(n13401) );
  NAND2_X1 U16542 ( .A1(n13263), .A2(n13401), .ZN(P1_U2957) );
  AOI22_X1 U16543 ( .A1(n20439), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13266) );
  INV_X1 U16544 ( .A(DATAI_6_), .ZN(n21215) );
  NAND2_X1 U16545 ( .A1(n14263), .A2(n21215), .ZN(n13265) );
  INV_X1 U16546 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16803) );
  NAND2_X1 U16547 ( .A1(n14923), .A2(n16803), .ZN(n13264) );
  AND2_X1 U16548 ( .A1(n13265), .A2(n13264), .ZN(n14942) );
  NAND2_X1 U16549 ( .A1(n20426), .A2(n14942), .ZN(n13411) );
  NAND2_X1 U16550 ( .A1(n13266), .A2(n13411), .ZN(P1_U2958) );
  AOI22_X1 U16551 ( .A1(n20439), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20438), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n13269) );
  INV_X1 U16552 ( .A(DATAI_11_), .ZN(n13268) );
  NAND2_X1 U16553 ( .A1(n14923), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13267) );
  OAI21_X1 U16554 ( .B1(n14923), .B2(n13268), .A(n13267), .ZN(n14986) );
  NAND2_X1 U16555 ( .A1(n20426), .A2(n14986), .ZN(n13403) );
  NAND2_X1 U16556 ( .A1(n13269), .A2(n13403), .ZN(P1_U2963) );
  NAND2_X1 U16557 ( .A1(n13271), .A2(n13270), .ZN(n13278) );
  INV_X1 U16558 ( .A(n13272), .ZN(n13273) );
  NAND2_X1 U16559 ( .A1(n13273), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20051) );
  OAI211_X1 U16560 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n13273), .A(
        n20051), .B(n20196), .ZN(n13274) );
  INV_X1 U16561 ( .A(n13274), .ZN(n13275) );
  AOI21_X1 U16562 ( .B1(n13276), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13275), .ZN(n13277) );
  NAND3_X1 U16563 ( .A1(n13373), .A2(n13375), .A3(n13374), .ZN(n13372) );
  NAND2_X1 U16564 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19603), .ZN(
        n13285) );
  AND2_X1 U16565 ( .A1(n14549), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14342) );
  NAND2_X1 U16566 ( .A1(n13479), .A2(n14342), .ZN(n14341) );
  XOR2_X1 U16567 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14341), .Z(n13292)
         );
  INV_X1 U16568 ( .A(n13455), .ZN(n13287) );
  AOI21_X1 U16569 ( .B1(n13288), .B2(n14030), .A(n13287), .ZN(n19382) );
  NOR2_X1 U16570 ( .A1(n15449), .A2(n13289), .ZN(n13290) );
  AOI21_X1 U16571 ( .B1(n19382), .B2(n15449), .A(n13290), .ZN(n13291) );
  OAI21_X1 U16572 ( .B1(n13292), .B2(n15479), .A(n13291), .ZN(P2_U2882) );
  INV_X1 U16573 ( .A(n13293), .ZN(n13294) );
  AOI21_X1 U16574 ( .B1(n13294), .B2(n16416), .A(n13513), .ZN(n13295) );
  INV_X1 U16575 ( .A(n13296), .ZN(n13589) );
  NOR2_X1 U16576 ( .A1(n21050), .A2(n13297), .ZN(n13496) );
  NAND2_X1 U16577 ( .A1(n13589), .A2(n13496), .ZN(n13298) );
  INV_X1 U16578 ( .A(n13435), .ZN(n13314) );
  NAND2_X1 U16579 ( .A1(n13080), .A2(n13958), .ZN(n13519) );
  NAND2_X1 U16580 ( .A1(n13519), .A2(n10148), .ZN(n13301) );
  INV_X1 U16581 ( .A(n16182), .ZN(n13424) );
  NAND3_X1 U16582 ( .A1(n13301), .A2(n13424), .A3(n16416), .ZN(n13311) );
  NAND2_X1 U16583 ( .A1(n16159), .A2(n13302), .ZN(n13868) );
  AOI21_X1 U16584 ( .B1(n13303), .B2(n11900), .A(n14002), .ZN(n13304) );
  NAND2_X1 U16585 ( .A1(n13305), .A2(n13304), .ZN(n13346) );
  AND2_X1 U16586 ( .A1(n13306), .A2(n13346), .ZN(n13307) );
  NOR2_X1 U16587 ( .A1(n13080), .A2(n13307), .ZN(n13507) );
  OR2_X1 U16588 ( .A1(n13676), .A2(n13308), .ZN(n13343) );
  INV_X1 U16589 ( .A(n13343), .ZN(n13309) );
  NOR2_X1 U16590 ( .A1(n13507), .A2(n13309), .ZN(n13310) );
  OAI211_X1 U16591 ( .C1(n16159), .C2(n13311), .A(n13868), .B(n13310), .ZN(
        n13312) );
  INV_X1 U16592 ( .A(n13312), .ZN(n13313) );
  NAND2_X1 U16593 ( .A1(n13314), .A2(n13313), .ZN(n13587) );
  INV_X1 U16594 ( .A(n13587), .ZN(n16129) );
  NAND2_X1 U16595 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16421) );
  NOR2_X1 U16596 ( .A1(n21045), .A2(n16421), .ZN(n13593) );
  NAND2_X1 U16597 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13593), .ZN(n13315) );
  OAI21_X1 U16598 ( .B1(n16129), .B2(n20276), .A(n13315), .ZN(n13317) );
  AOI21_X1 U16599 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21045), .A(n13317), 
        .ZN(n15317) );
  INV_X1 U16600 ( .A(n15317), .ZN(n13320) );
  INV_X1 U16601 ( .A(n20583), .ZN(n13943) );
  OR2_X1 U16602 ( .A1(n12001), .A2(n13943), .ZN(n13316) );
  XNOR2_X1 U16603 ( .A(n13316), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20347) );
  NAND4_X1 U16604 ( .A1(n13317), .A2(n13367), .A3(n13589), .A4(n20347), .ZN(
        n13318) );
  OAI21_X1 U16605 ( .B1(n13320), .B2(n13319), .A(n13318), .ZN(P1_U3468) );
  NAND2_X1 U16606 ( .A1(n13322), .A2(n13321), .ZN(n13324) );
  AND2_X1 U16607 ( .A1(n13324), .A2(n10087), .ZN(n20213) );
  XNOR2_X1 U16608 ( .A(n20210), .B(n20213), .ZN(n13328) );
  NAND2_X1 U16609 ( .A1(n20222), .A2(n19409), .ZN(n13325) );
  OAI21_X1 U16610 ( .B1(n20222), .B2(n19409), .A(n13325), .ZN(n19489) );
  NOR2_X1 U16611 ( .A1(n20234), .A2(n19415), .ZN(n19496) );
  NOR2_X1 U16612 ( .A1(n19489), .A2(n19496), .ZN(n19488) );
  INV_X1 U16613 ( .A(n13325), .ZN(n13326) );
  NOR2_X1 U16614 ( .A1(n19488), .A2(n13326), .ZN(n13327) );
  NOR2_X1 U16615 ( .A1(n13327), .A2(n13328), .ZN(n19468) );
  AOI21_X1 U16616 ( .B1(n13328), .B2(n13327), .A(n19468), .ZN(n13340) );
  AND2_X1 U16617 ( .A1(n13329), .A2(n16659), .ZN(n13330) );
  INV_X1 U16618 ( .A(n10492), .ZN(n13334) );
  NAND2_X1 U16619 ( .A1(n19466), .A2(n13335), .ZN(n15558) );
  NAND2_X1 U16620 ( .A1(n19466), .A2(n13336), .ZN(n14117) );
  NAND2_X1 U16621 ( .A1(n15558), .A2(n14117), .ZN(n19459) );
  INV_X1 U16622 ( .A(n19466), .ZN(n19494) );
  AOI22_X1 U16623 ( .A1(n19459), .A2(n16484), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19494), .ZN(n13339) );
  INV_X1 U16624 ( .A(n20213), .ZN(n13337) );
  NAND2_X1 U16625 ( .A1(n13337), .A2(n19495), .ZN(n13338) );
  OAI211_X1 U16626 ( .C1(n13340), .C2(n19490), .A(n13339), .B(n13338), .ZN(
        P2_U2917) );
  INV_X1 U16627 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20760) );
  INV_X1 U16628 ( .A(n13572), .ZN(n13341) );
  AOI21_X1 U16629 ( .B1(n15312), .B2(n13341), .A(n15317), .ZN(n13371) );
  OAI21_X1 U16630 ( .B1(n13344), .B2(n13676), .A(n13343), .ZN(n13345) );
  INV_X1 U16631 ( .A(n13345), .ZN(n13347) );
  AND3_X1 U16632 ( .A1(n13348), .A2(n13347), .A3(n13346), .ZN(n13522) );
  NAND3_X1 U16633 ( .A1(n13349), .A2(n13521), .A3(n13528), .ZN(n13350) );
  NOR2_X1 U16634 ( .A1(n13350), .A2(n13300), .ZN(n13352) );
  AND3_X1 U16635 ( .A1(n13522), .A2(n13352), .A3(n13351), .ZN(n13353) );
  NAND2_X1 U16636 ( .A1(n13296), .A2(n13353), .ZN(n15305) );
  NOR2_X1 U16637 ( .A1(n13519), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15304) );
  NOR2_X1 U16638 ( .A1(n15302), .A2(n13354), .ZN(n13574) );
  INV_X1 U16639 ( .A(n13574), .ZN(n13355) );
  OAI22_X1 U16640 ( .A1(n13519), .A2(n15318), .B1(n13572), .B2(n13355), .ZN(
        n13356) );
  OAI21_X1 U16641 ( .B1(n15304), .B2(n13356), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13365) );
  NAND2_X1 U16642 ( .A1(n13525), .A2(n13357), .ZN(n13575) );
  NOR2_X1 U16643 ( .A1(n13358), .A2(n15318), .ZN(n13573) );
  XNOR2_X1 U16644 ( .A(n13573), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13360) );
  AOI22_X1 U16645 ( .A1(n13575), .A2(n13360), .B1(n13359), .B2(n13574), .ZN(
        n13364) );
  NOR2_X1 U16646 ( .A1(n13519), .A2(n13361), .ZN(n13571) );
  NAND2_X1 U16647 ( .A1(n13571), .A2(n13362), .ZN(n13363) );
  NAND3_X1 U16648 ( .A1(n13365), .A2(n13364), .A3(n13363), .ZN(n13366) );
  AOI21_X1 U16649 ( .B1(n13342), .B2(n15305), .A(n13366), .ZN(n13579) );
  INV_X1 U16650 ( .A(n13367), .ZN(n15315) );
  NOR2_X1 U16651 ( .A1(n13579), .A2(n15315), .ZN(n13368) );
  AOI21_X1 U16652 ( .B1(n15312), .B2(n13359), .A(n13368), .ZN(n13369) );
  OAI22_X1 U16653 ( .A1(n13371), .A2(n13370), .B1(n15317), .B2(n13369), .ZN(
        P1_U3469) );
  NAND2_X1 U16654 ( .A1(n13374), .A2(n13373), .ZN(n13377) );
  INV_X1 U16655 ( .A(n13375), .ZN(n13376) );
  INV_X1 U16656 ( .A(n16076), .ZN(n16678) );
  NAND2_X1 U16657 ( .A1(n13379), .A2(n16678), .ZN(n13390) );
  NAND2_X1 U16658 ( .A1(n16665), .A2(n16666), .ZN(n16080) );
  NOR2_X1 U16659 ( .A1(n13380), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16074) );
  INV_X1 U16660 ( .A(n16074), .ZN(n16070) );
  NAND2_X1 U16661 ( .A1(n10503), .A2(n13381), .ZN(n13382) );
  NAND2_X1 U16662 ( .A1(n13382), .A2(n9677), .ZN(n13383) );
  AOI21_X1 U16663 ( .B1(n16080), .B2(n16070), .A(n13383), .ZN(n13388) );
  NAND2_X1 U16664 ( .A1(n10508), .A2(n13384), .ZN(n13385) );
  NAND2_X1 U16665 ( .A1(n13385), .A2(n9677), .ZN(n16075) );
  INV_X1 U16666 ( .A(n13381), .ZN(n13386) );
  NAND2_X1 U16667 ( .A1(n10503), .A2(n13386), .ZN(n16073) );
  AND3_X1 U16668 ( .A1(n16075), .A2(n16070), .A3(n16073), .ZN(n13387) );
  MUX2_X1 U16669 ( .A(n13388), .B(n13387), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13389) );
  NAND2_X1 U16670 ( .A1(n13390), .A2(n13389), .ZN(n16677) );
  AOI22_X1 U16671 ( .A1(n19854), .A2(n20190), .B1(n20198), .B2(n16677), .ZN(
        n13392) );
  INV_X1 U16672 ( .A(n20192), .ZN(n20195) );
  NAND2_X1 U16673 ( .A1(n20195), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13391) );
  OAI21_X1 U16674 ( .B1(n13392), .B2(n20195), .A(n13391), .ZN(P2_U3596) );
  INV_X2 U16675 ( .A(n13393), .ZN(n20439) );
  AOI22_X1 U16676 ( .A1(n20439), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13396) );
  INV_X1 U16677 ( .A(DATAI_1_), .ZN(n21227) );
  NAND2_X1 U16678 ( .A1(n14263), .A2(n21227), .ZN(n13395) );
  INV_X1 U16679 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16813) );
  NAND2_X1 U16680 ( .A1(n14923), .A2(n16813), .ZN(n13394) );
  AND2_X1 U16681 ( .A1(n13395), .A2(n13394), .ZN(n14965) );
  NAND2_X1 U16682 ( .A1(n20426), .A2(n14965), .ZN(n13415) );
  NAND2_X1 U16683 ( .A1(n13396), .A2(n13415), .ZN(P1_U2938) );
  AOI22_X1 U16684 ( .A1(n20439), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13398) );
  NAND2_X1 U16685 ( .A1(n13398), .A2(n13397), .ZN(P1_U2940) );
  AOI22_X1 U16686 ( .A1(n20439), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13400) );
  INV_X1 U16687 ( .A(DATAI_9_), .ZN(n21228) );
  NAND2_X1 U16688 ( .A1(n14923), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13399) );
  OAI21_X1 U16689 ( .B1(n14923), .B2(n21228), .A(n13399), .ZN(n14933) );
  NAND2_X1 U16690 ( .A1(n20426), .A2(n14933), .ZN(n20430) );
  NAND2_X1 U16691 ( .A1(n13400), .A2(n20430), .ZN(P1_U2946) );
  AOI22_X1 U16692 ( .A1(n20439), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13402) );
  NAND2_X1 U16693 ( .A1(n13402), .A2(n13401), .ZN(P1_U2942) );
  AOI22_X1 U16694 ( .A1(n20439), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13404) );
  NAND2_X1 U16695 ( .A1(n13404), .A2(n13403), .ZN(P1_U2948) );
  AOI22_X1 U16696 ( .A1(n20439), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13407) );
  INV_X1 U16697 ( .A(DATAI_2_), .ZN(n13406) );
  NAND2_X1 U16698 ( .A1(n14923), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13405) );
  OAI21_X1 U16699 ( .B1(n14923), .B2(n13406), .A(n13405), .ZN(n14962) );
  NAND2_X1 U16700 ( .A1(n20426), .A2(n14962), .ZN(n13417) );
  NAND2_X1 U16701 ( .A1(n13407), .A2(n13417), .ZN(P1_U2939) );
  AOI22_X1 U16702 ( .A1(n20439), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13410) );
  INV_X1 U16703 ( .A(DATAI_0_), .ZN(n21208) );
  NAND2_X1 U16704 ( .A1(n14263), .A2(n21208), .ZN(n13409) );
  INV_X1 U16705 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16818) );
  NAND2_X1 U16706 ( .A1(n14923), .A2(n16818), .ZN(n13408) );
  AND2_X1 U16707 ( .A1(n13409), .A2(n13408), .ZN(n14971) );
  NAND2_X1 U16708 ( .A1(n20426), .A2(n14971), .ZN(n13413) );
  NAND2_X1 U16709 ( .A1(n13410), .A2(n13413), .ZN(P1_U2937) );
  AOI22_X1 U16710 ( .A1(n20439), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13412) );
  NAND2_X1 U16711 ( .A1(n13412), .A2(n13411), .ZN(P1_U2943) );
  AOI22_X1 U16712 ( .A1(n20439), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13414) );
  NAND2_X1 U16713 ( .A1(n13414), .A2(n13413), .ZN(P1_U2952) );
  AOI22_X1 U16714 ( .A1(n20439), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13416) );
  NAND2_X1 U16715 ( .A1(n13416), .A2(n13415), .ZN(P1_U2953) );
  AOI22_X1 U16716 ( .A1(n20439), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13418) );
  NAND2_X1 U16717 ( .A1(n13418), .A2(n13417), .ZN(P1_U2954) );
  AOI22_X1 U16718 ( .A1(n20439), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13420) );
  NAND2_X1 U16719 ( .A1(n13420), .A2(n13419), .ZN(P1_U2941) );
  AOI22_X1 U16720 ( .A1(n20439), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13422) );
  NAND2_X1 U16721 ( .A1(n13422), .A2(n13421), .ZN(P1_U2944) );
  INV_X1 U16722 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13428) );
  NAND2_X1 U16723 ( .A1(n13423), .A2(n13498), .ZN(n16152) );
  NAND2_X1 U16724 ( .A1(n13519), .A2(n16152), .ZN(n13425) );
  NAND3_X1 U16725 ( .A1(n13425), .A2(n13424), .A3(n13511), .ZN(n13426) );
  NAND2_X1 U16726 ( .A1(n20388), .A2(n13499), .ZN(n13787) );
  NOR2_X1 U16727 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16421), .ZN(n20414) );
  INV_X1 U16728 ( .A(n20414), .ZN(n21049) );
  NOR2_X4 U16729 ( .A1(n20388), .A2(n20400), .ZN(n20409) );
  AOI22_X1 U16730 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13427) );
  OAI21_X1 U16731 ( .B1(n13428), .B2(n13787), .A(n13427), .ZN(P1_U2913) );
  INV_X1 U16732 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U16733 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13429) );
  OAI21_X1 U16734 ( .B1(n13430), .B2(n13787), .A(n13429), .ZN(P1_U2907) );
  INV_X1 U16735 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13432) );
  AOI22_X1 U16736 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13431) );
  OAI21_X1 U16737 ( .B1(n13432), .B2(n13787), .A(n13431), .ZN(P1_U2911) );
  INV_X1 U16738 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U16739 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13433) );
  OAI21_X1 U16740 ( .B1(n13434), .B2(n13787), .A(n13433), .ZN(P1_U2909) );
  INV_X1 U16741 ( .A(n13875), .ZN(n14347) );
  NAND4_X1 U16742 ( .A1(n14347), .A2(n15338), .A3(n13511), .A4(n13967), .ZN(
        n13869) );
  OR2_X1 U16743 ( .A1(n13528), .A2(n13869), .ZN(n13436) );
  NAND2_X1 U16744 ( .A1(n14987), .A2(n13438), .ZN(n14989) );
  INV_X1 U16745 ( .A(n14971), .ZN(n13441) );
  NAND2_X2 U16746 ( .A1(n11880), .A2(n14987), .ZN(n14982) );
  XNOR2_X1 U16747 ( .A(n13440), .B(n13439), .ZN(n13919) );
  OAI222_X1 U16748 ( .A1(n14989), .A2(n13441), .B1(n14987), .B2(n12116), .C1(
        n14982), .C2(n13919), .ZN(P1_U2904) );
  INV_X1 U16749 ( .A(n14965), .ZN(n13445) );
  OR2_X1 U16750 ( .A1(n13443), .A2(n13442), .ZN(n13444) );
  AND2_X1 U16751 ( .A1(n13646), .A2(n13444), .ZN(n20372) );
  INV_X1 U16752 ( .A(n20372), .ZN(n13929) );
  OAI222_X1 U16753 ( .A1(n14989), .A2(n13445), .B1(n14987), .B2(n12108), .C1(
        n14982), .C2(n13929), .ZN(P1_U2903) );
  NAND2_X1 U16754 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13473) );
  NOR2_X1 U16755 ( .A1(n14341), .A2(n13473), .ZN(n13544) );
  XNOR2_X1 U16756 ( .A(n13544), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13450) );
  NOR2_X1 U16757 ( .A1(n13457), .A2(n13446), .ZN(n13447) );
  OR2_X1 U16758 ( .A1(n13695), .A2(n13447), .ZN(n16041) );
  INV_X1 U16759 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13448) );
  MUX2_X1 U16760 ( .A(n16041), .B(n13448), .S(n15448), .Z(n13449) );
  OAI21_X1 U16761 ( .B1(n13450), .B2(n15479), .A(n13449), .ZN(P2_U2880) );
  NOR2_X1 U16762 ( .A1(n14341), .A2(n13451), .ZN(n13453) );
  INV_X1 U16763 ( .A(n13544), .ZN(n13452) );
  OAI211_X1 U16764 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13453), .A(
        n13452), .B(n15470), .ZN(n13459) );
  AND2_X1 U16765 ( .A1(n13455), .A2(n13454), .ZN(n13456) );
  OR2_X1 U16766 ( .A1(n13457), .A2(n13456), .ZN(n16577) );
  INV_X1 U16767 ( .A(n16577), .ZN(n19371) );
  NAND2_X1 U16768 ( .A1(n19371), .A2(n15449), .ZN(n13458) );
  OAI211_X1 U16769 ( .C1(n15449), .C2(n10560), .A(n13459), .B(n13458), .ZN(
        P2_U2881) );
  XNOR2_X1 U16770 ( .A(n13460), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13543) );
  INV_X1 U16771 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13461) );
  OAI22_X1 U16772 ( .A1(n16260), .A2(n13462), .B1(n16406), .B2(n13461), .ZN(
        n13463) );
  AOI21_X1 U16773 ( .B1(n16285), .B2(n13462), .A(n13463), .ZN(n13465) );
  NAND2_X1 U16774 ( .A1(n20372), .A2(n16286), .ZN(n13464) );
  OAI211_X1 U16775 ( .C1(n13543), .C2(n20282), .A(n13465), .B(n13464), .ZN(
        P1_U2998) );
  NOR2_X1 U16776 ( .A1(n15302), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13466) );
  AOI21_X1 U16777 ( .B1(n20546), .B2(n15305), .A(n13466), .ZN(n16128) );
  OAI21_X1 U16778 ( .B1(n16128), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n16420), 
        .ZN(n13467) );
  INV_X1 U16779 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20455) );
  NOR2_X1 U16780 ( .A1(n16420), .A2(n20455), .ZN(n15310) );
  INV_X1 U16781 ( .A(n15310), .ZN(n15306) );
  AOI22_X1 U16782 ( .A1(n13467), .A2(n15306), .B1(n15312), .B2(n9955), .ZN(
        n13469) );
  INV_X1 U16783 ( .A(n13519), .ZN(n13468) );
  NAND2_X1 U16784 ( .A1(n13468), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16126) );
  OAI22_X1 U16785 ( .A1(n15317), .A2(n13469), .B1(n15315), .B2(n16126), .ZN(
        n13470) );
  AOI21_X1 U16786 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15317), .A(
        n13470), .ZN(n13471) );
  INV_X1 U16787 ( .A(n13471), .ZN(P1_U3474) );
  INV_X1 U16788 ( .A(n14549), .ZN(n13477) );
  NAND2_X1 U16789 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13472) );
  NOR2_X1 U16790 ( .A1(n13473), .A2(n13472), .ZN(n13474) );
  NAND3_X1 U16791 ( .A1(n13475), .A2(n13545), .A3(n13474), .ZN(n13476) );
  NOR2_X1 U16792 ( .A1(n13477), .A2(n13476), .ZN(n13478) );
  INV_X1 U16793 ( .A(n13481), .ZN(n13484) );
  INV_X1 U16794 ( .A(n13603), .ZN(n13482) );
  OAI211_X1 U16795 ( .C1(n13484), .C2(n13483), .A(n13482), .B(n15470), .ZN(
        n13488) );
  OR2_X1 U16796 ( .A1(n13485), .A2(n13547), .ZN(n13486) );
  AND2_X1 U16797 ( .A1(n13486), .A2(n13606), .ZN(n19350) );
  NAND2_X1 U16798 ( .A1(n19350), .A2(n15449), .ZN(n13487) );
  OAI211_X1 U16799 ( .C1(n15449), .C2(n13489), .A(n13488), .B(n13487), .ZN(
        P2_U2877) );
  OAI21_X1 U16800 ( .B1(n13491), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13490), .ZN(n20445) );
  OAI21_X1 U16801 ( .B1(n16291), .B2(n13492), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U16802 ( .A1(n16391), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20443) );
  OAI211_X1 U16803 ( .C1(n20445), .C2(n20282), .A(n13493), .B(n20443), .ZN(
        n13494) );
  INV_X1 U16804 ( .A(n13494), .ZN(n13495) );
  OAI21_X1 U16805 ( .B1(n13919), .B2(n16263), .A(n13495), .ZN(P1_U2999) );
  INV_X1 U16806 ( .A(n13496), .ZN(n13497) );
  AOI21_X1 U16807 ( .B1(n13958), .B2(n16182), .A(n13497), .ZN(n13504) );
  NAND2_X1 U16808 ( .A1(n13498), .A2(n16182), .ZN(n13673) );
  AND2_X1 U16809 ( .A1(n13673), .A2(n16416), .ZN(n13501) );
  NAND2_X1 U16810 ( .A1(n13499), .A2(n14267), .ZN(n13500) );
  AOI21_X1 U16811 ( .B1(n13300), .B2(n13501), .A(n13500), .ZN(n13502) );
  NOR2_X1 U16812 ( .A1(n16159), .A2(n13502), .ZN(n13503) );
  MUX2_X1 U16813 ( .A(n13504), .B(n13503), .S(n13941), .Z(n13505) );
  INV_X1 U16814 ( .A(n13505), .ZN(n13510) );
  INV_X1 U16815 ( .A(n13506), .ZN(n13508) );
  AOI21_X1 U16816 ( .B1(n16159), .B2(n13508), .A(n13507), .ZN(n13509) );
  NAND2_X1 U16817 ( .A1(n13510), .A2(n13509), .ZN(n13512) );
  AOI21_X1 U16818 ( .B1(n13515), .B2(n13514), .A(n13513), .ZN(n13516) );
  AND3_X1 U16819 ( .A1(n13517), .A2(n13516), .A3(n16140), .ZN(n13518) );
  AND4_X1 U16820 ( .A1(n13523), .A2(n13522), .A3(n13521), .A4(n13520), .ZN(
        n13524) );
  AND2_X2 U16821 ( .A1(n20453), .A2(n15149), .ZN(n16374) );
  NAND2_X1 U16822 ( .A1(n16374), .A2(n16371), .ZN(n15245) );
  INV_X1 U16823 ( .A(n15245), .ZN(n15282) );
  NOR2_X1 U16824 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16353), .ZN(
        n13562) );
  NOR3_X1 U16825 ( .A1(n15282), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13562), .ZN(n13539) );
  NAND2_X1 U16826 ( .A1(n13526), .A2(n15338), .ZN(n13527) );
  OR2_X1 U16827 ( .A1(n13528), .A2(n13527), .ZN(n13529) );
  AND2_X1 U16828 ( .A1(n16152), .A2(n13529), .ZN(n13530) );
  OR2_X1 U16829 ( .A1(n14656), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13534) );
  NAND3_X1 U16830 ( .A1(n13535), .A2(n13534), .A3(n13533), .ZN(n13555) );
  INV_X1 U16831 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13792) );
  OR2_X1 U16832 ( .A1(n14318), .A2(n13792), .ZN(n13537) );
  NAND2_X1 U16833 ( .A1(n14322), .A2(n13792), .ZN(n13536) );
  NAND2_X1 U16834 ( .A1(n13537), .A2(n13536), .ZN(n13789) );
  XNOR2_X1 U16835 ( .A(n13555), .B(n13789), .ZN(n13556) );
  XNOR2_X1 U16836 ( .A(n13556), .B(n9653), .ZN(n20359) );
  OAI22_X1 U16837 ( .A1(n16407), .A2(n20359), .B1(n13461), .B2(n16406), .ZN(
        n13538) );
  NOR2_X1 U16838 ( .A1(n13539), .A2(n13538), .ZN(n13542) );
  NOR2_X1 U16839 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16371), .ZN(
        n20442) );
  INV_X1 U16840 ( .A(n15149), .ZN(n16355) );
  NAND2_X1 U16841 ( .A1(n16355), .A2(n20455), .ZN(n20447) );
  NAND2_X1 U16842 ( .A1(n16406), .A2(n13540), .ZN(n20454) );
  NAND2_X1 U16843 ( .A1(n20447), .A2(n20454), .ZN(n15145) );
  OAI21_X1 U16844 ( .B1(n20442), .B2(n15145), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13541) );
  OAI211_X1 U16845 ( .C1(n13543), .C2(n20446), .A(n13542), .B(n13541), .ZN(
        P1_U3030) );
  NAND2_X1 U16846 ( .A1(n13544), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13699) );
  NOR2_X1 U16847 ( .A1(n13699), .A2(n13700), .ZN(n13698) );
  OAI211_X1 U16848 ( .C1(n13698), .C2(n13545), .A(n15470), .B(n13481), .ZN(
        n13551) );
  NAND2_X1 U16849 ( .A1(n13546), .A2(n13696), .ZN(n13549) );
  INV_X1 U16850 ( .A(n13547), .ZN(n13548) );
  NAND2_X1 U16851 ( .A1(n19360), .A2(n15449), .ZN(n13550) );
  OAI211_X1 U16852 ( .C1(n10570), .C2(n15449), .A(n13551), .B(n13550), .ZN(
        P2_U2878) );
  INV_X1 U16853 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15301) );
  NOR2_X1 U16854 ( .A1(n12683), .A2(n15301), .ZN(n15132) );
  OAI21_X1 U16855 ( .B1(n16374), .B2(n15132), .A(n15261), .ZN(n13554) );
  AND3_X1 U16856 ( .A1(n15147), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13553) );
  OAI21_X1 U16857 ( .B1(n13554), .B2(n13553), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13568) );
  AOI21_X1 U16858 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13817) );
  NAND2_X1 U16859 ( .A1(n15147), .A2(n13817), .ZN(n13729) );
  INV_X1 U16860 ( .A(n13729), .ZN(n13566) );
  AOI21_X1 U16861 ( .B1(n13556), .B2(n14652), .A(n13555), .ZN(n13560) );
  NOR2_X1 U16862 ( .A1(n14656), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13557) );
  NOR2_X1 U16863 ( .A1(n13558), .A2(n13557), .ZN(n13559) );
  NAND2_X1 U16864 ( .A1(n13560), .A2(n13559), .ZN(n13735) );
  OR2_X1 U16865 ( .A1(n13560), .A2(n13559), .ZN(n13561) );
  NAND2_X1 U16866 ( .A1(n13735), .A2(n13561), .ZN(n13932) );
  NAND3_X1 U16867 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16370), .A3(
        n12683), .ZN(n13564) );
  INV_X1 U16868 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20960) );
  NOR2_X1 U16869 ( .A1(n16406), .A2(n20960), .ZN(n13648) );
  INV_X1 U16870 ( .A(n13648), .ZN(n13563) );
  OAI211_X1 U16871 ( .C1(n16407), .C2(n13932), .A(n13564), .B(n13563), .ZN(
        n13565) );
  NOR2_X1 U16872 ( .A1(n13566), .A2(n13565), .ZN(n13567) );
  OAI211_X1 U16873 ( .C1(n13653), .C2(n20446), .A(n13568), .B(n13567), .ZN(
        P1_U3029) );
  NOR2_X1 U16874 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16420), .ZN(n13585) );
  INV_X1 U16875 ( .A(n13570), .ZN(n20460) );
  MUX2_X1 U16876 ( .A(n15304), .B(n13571), .S(n10154), .Z(n13577) );
  NOR2_X1 U16877 ( .A1(n13573), .A2(n13572), .ZN(n15313) );
  MUX2_X1 U16878 ( .A(n13575), .B(n13574), .S(n15313), .Z(n13576) );
  AOI211_X1 U16879 ( .C1(n20460), .C2(n15305), .A(n13577), .B(n13576), .ZN(
        n15316) );
  INV_X1 U16880 ( .A(n15316), .ZN(n13578) );
  MUX2_X1 U16881 ( .A(n15318), .B(n13578), .S(n13587), .Z(n16135) );
  AOI22_X1 U16882 ( .A1(n13585), .A2(n15318), .B1(n16420), .B2(n16135), .ZN(
        n13583) );
  OR2_X1 U16883 ( .A1(n13587), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13581) );
  NAND2_X1 U16884 ( .A1(n13587), .A2(n13579), .ZN(n13580) );
  AOI22_X1 U16885 ( .A1(n13585), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16420), .B2(n16125), .ZN(n13582) );
  NOR2_X1 U16886 ( .A1(n13583), .A2(n13582), .ZN(n16144) );
  INV_X1 U16887 ( .A(n13584), .ZN(n15300) );
  NAND2_X1 U16888 ( .A1(n16144), .A2(n15300), .ZN(n13592) );
  INV_X1 U16889 ( .A(n13585), .ZN(n13586) );
  OAI21_X1 U16890 ( .B1(n13587), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n13586), 
        .ZN(n13588) );
  NAND2_X1 U16891 ( .A1(n13588), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13591) );
  NAND3_X1 U16892 ( .A1(n20347), .A2(n13589), .A3(n16420), .ZN(n13590) );
  AND2_X1 U16893 ( .A1(n13591), .A2(n13590), .ZN(n16142) );
  NAND2_X1 U16894 ( .A1(n13592), .A2(n16142), .ZN(n13599) );
  OAI21_X1 U16895 ( .B1(n13599), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13593), .ZN(
        n13594) );
  NAND2_X1 U16896 ( .A1(n21042), .A2(n16420), .ZN(n21044) );
  NAND2_X1 U16897 ( .A1(n13594), .A2(n15326), .ZN(n21032) );
  NOR2_X1 U16898 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16420), .ZN(n21025) );
  NOR2_X1 U16899 ( .A1(n13570), .A2(n21025), .ZN(n13597) );
  AOI21_X1 U16900 ( .B1(n21021), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20883), 
        .ZN(n20551) );
  AND2_X1 U16901 ( .A1(n21021), .A2(n21030), .ZN(n20800) );
  MUX2_X1 U16902 ( .A(n20551), .B(n20800), .S(n20582), .Z(n13596) );
  OAI21_X1 U16903 ( .B1(n13597), .B2(n13596), .A(n21032), .ZN(n13598) );
  OAI21_X1 U16904 ( .B1(n12762), .B2(n21032), .A(n13598), .ZN(P1_U3476) );
  NOR2_X1 U16905 ( .A1(n13599), .A2(n16421), .ZN(n16147) );
  INV_X1 U16906 ( .A(n20546), .ZN(n13600) );
  OAI22_X1 U16907 ( .A1(n20518), .A2(n20883), .B1(n13600), .B2(n21025), .ZN(
        n13601) );
  OAI21_X1 U16908 ( .B1(n16147), .B2(n13601), .A(n21032), .ZN(n13602) );
  OAI21_X1 U16909 ( .B1(n21032), .B2(n20721), .A(n13602), .ZN(P1_U3478) );
  OAI211_X1 U16910 ( .C1(n13603), .C2(n13605), .A(n13604), .B(n15470), .ZN(
        n13611) );
  NAND2_X1 U16911 ( .A1(n13607), .A2(n13606), .ZN(n13609) );
  INV_X1 U16912 ( .A(n13809), .ZN(n13608) );
  AND2_X1 U16913 ( .A1(n13609), .A2(n13608), .ZN(n19340) );
  NAND2_X1 U16914 ( .A1(n19340), .A2(n15449), .ZN(n13610) );
  OAI211_X1 U16915 ( .C1(n15449), .C2(n10578), .A(n13611), .B(n13610), .ZN(
        P2_U2876) );
  NAND2_X1 U16916 ( .A1(n13661), .A2(n13614), .ZN(n13615) );
  AND2_X1 U16917 ( .A1(n13838), .A2(n13615), .ZN(n20355) );
  INV_X1 U16918 ( .A(n20355), .ZN(n13877) );
  INV_X1 U16919 ( .A(n14989), .ZN(n14980) );
  AOI22_X1 U16920 ( .A1(n14980), .A2(n15337), .B1(P1_EAX_REG_4__SCAN_IN), .B2(
        n14979), .ZN(n13616) );
  OAI21_X1 U16921 ( .B1(n13877), .B2(n14982), .A(n13616), .ZN(P1_U2900) );
  NAND2_X1 U16922 ( .A1(n9658), .A2(n13617), .ZN(n13618) );
  XNOR2_X1 U16923 ( .A(n15726), .B(n13618), .ZN(n13627) );
  XOR2_X1 U16924 ( .A(n13620), .B(n13619), .Z(n19463) );
  NAND2_X1 U16925 ( .A1(n19463), .A2(n19420), .ZN(n13625) );
  AOI22_X1 U16926 ( .A1(n13621), .A2(n12839), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19406), .ZN(n13622) );
  OAI211_X1 U16927 ( .C1(n10567), .C2(n19416), .A(n13622), .B(n19333), .ZN(
        n13623) );
  AOI21_X1 U16928 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19431), .A(
        n13623), .ZN(n13624) );
  OAI211_X1 U16929 ( .C1(n16041), .C2(n19389), .A(n13625), .B(n13624), .ZN(
        n13626) );
  AOI21_X1 U16930 ( .B1(n13627), .B2(n19411), .A(n13626), .ZN(n13628) );
  INV_X1 U16931 ( .A(n13628), .ZN(P2_U2848) );
  NAND2_X1 U16932 ( .A1(n9658), .A2(n13629), .ZN(n13630) );
  XNOR2_X1 U16933 ( .A(n13985), .B(n13630), .ZN(n13644) );
  INV_X1 U16934 ( .A(n19428), .ZN(n19390) );
  OR2_X1 U16935 ( .A1(n13632), .A2(n13631), .ZN(n13634) );
  NAND2_X1 U16936 ( .A1(n13634), .A2(n13633), .ZN(n20206) );
  INV_X1 U16937 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20136) );
  OAI22_X1 U16938 ( .A1(n19418), .A2(n13635), .B1(n13983), .B2(n19386), .ZN(
        n13636) );
  AOI21_X1 U16939 ( .B1(n19402), .B2(P2_REIP_REG_3__SCAN_IN), .A(n13636), .ZN(
        n13639) );
  NAND2_X1 U16940 ( .A1(n12839), .A2(n10026), .ZN(n13638) );
  OAI211_X1 U16941 ( .C1(n20206), .C2(n19408), .A(n13639), .B(n13638), .ZN(
        n13640) );
  INV_X1 U16942 ( .A(n13640), .ZN(n13642) );
  NAND2_X1 U16943 ( .A1(n13379), .A2(n19425), .ZN(n13641) );
  OAI211_X1 U16944 ( .C1(n20204), .C2(n19390), .A(n13642), .B(n13641), .ZN(
        n13643) );
  AOI21_X1 U16945 ( .B1(n13644), .B2(n19411), .A(n13643), .ZN(n13645) );
  INV_X1 U16946 ( .A(n13645), .ZN(P2_U2852) );
  OAI21_X1 U16947 ( .B1(n9696), .B2(n12120), .A(n13657), .ZN(n13930) );
  INV_X1 U16948 ( .A(n13930), .ZN(n13651) );
  AOI21_X1 U16949 ( .B1(n16291), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13648), .ZN(n13649) );
  OAI21_X1 U16950 ( .B1(n16299), .B2(n13687), .A(n13649), .ZN(n13650) );
  AOI21_X1 U16951 ( .B1(n13651), .B2(n16286), .A(n13650), .ZN(n13652) );
  OAI21_X1 U16952 ( .B1(n20282), .B2(n13653), .A(n13652), .ZN(P1_U2997) );
  XNOR2_X1 U16953 ( .A(n13655), .B(n13654), .ZN(n13740) );
  INV_X1 U16954 ( .A(n13656), .ZN(n13659) );
  NAND3_X1 U16955 ( .A1(n13659), .A2(n13658), .A3(n13657), .ZN(n13660) );
  NAND2_X1 U16956 ( .A1(n13661), .A2(n13660), .ZN(n13880) );
  INV_X1 U16957 ( .A(n13880), .ZN(n13664) );
  INV_X1 U16958 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20963) );
  NOR2_X1 U16959 ( .A1(n16406), .A2(n20963), .ZN(n13737) );
  AOI21_X1 U16960 ( .B1(n16291), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13737), .ZN(n13662) );
  OAI21_X1 U16961 ( .B1(n16299), .B2(n13802), .A(n13662), .ZN(n13663) );
  AOI21_X1 U16962 ( .B1(n13664), .B2(n16286), .A(n13663), .ZN(n13665) );
  OAI21_X1 U16963 ( .B1(n13740), .B2(n20282), .A(n13665), .ZN(P1_U2996) );
  AND2_X1 U16964 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21045), .ZN(n13666) );
  NOR2_X1 U16965 ( .A1(n20760), .A2(n21044), .ZN(n16150) );
  AOI22_X1 U16966 ( .A1(n13667), .A2(n13666), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16150), .ZN(n13668) );
  AND2_X1 U16967 ( .A1(n16406), .A2(n13668), .ZN(n13669) );
  NOR2_X1 U16968 ( .A1(n13685), .A2(n16420), .ZN(n13670) );
  NAND2_X1 U16969 ( .A1(n14864), .A2(n13671), .ZN(n20371) );
  INV_X1 U16970 ( .A(n20371), .ZN(n13808) );
  NOR2_X1 U16971 ( .A1(n14002), .A2(n21042), .ZN(n13672) );
  AND2_X1 U16972 ( .A1(n16416), .A2(n21172), .ZN(n16151) );
  AND2_X1 U16973 ( .A1(n13673), .A2(n16151), .ZN(n13681) );
  INV_X1 U16974 ( .A(n14099), .ZN(n13674) );
  NOR2_X1 U16975 ( .A1(n13674), .A2(n13461), .ZN(n20367) );
  NAND2_X1 U16976 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20367), .ZN(n14078) );
  AND2_X1 U16977 ( .A1(n14812), .A2(n14078), .ZN(n13804) );
  NAND2_X1 U16978 ( .A1(n13805), .A2(n20960), .ZN(n13675) );
  NAND2_X1 U16979 ( .A1(n13804), .A2(n13675), .ZN(n13692) );
  NOR2_X1 U16980 ( .A1(n13676), .A2(n21042), .ZN(n13677) );
  AND2_X1 U16981 ( .A1(n14099), .A2(n13677), .ZN(n20363) );
  AOI22_X1 U16982 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20348), .B1(
        n20363), .B2(n20460), .ZN(n13691) );
  AND2_X1 U16983 ( .A1(n13958), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13680) );
  INV_X1 U16984 ( .A(n13680), .ZN(n13678) );
  NOR2_X1 U16985 ( .A1(n13678), .A2(n16151), .ZN(n13679) );
  INV_X1 U16986 ( .A(n13932), .ZN(n13684) );
  NOR2_X1 U16987 ( .A1(n13681), .A2(n13680), .ZN(n13682) );
  AOI22_X1 U16988 ( .A1(n20362), .A2(n13684), .B1(n20360), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13690) );
  AND2_X1 U16989 ( .A1(n13685), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13686) );
  INV_X1 U16990 ( .A(n13687), .ZN(n13688) );
  NAND2_X1 U16991 ( .A1(n20349), .A2(n13688), .ZN(n13689) );
  AND4_X1 U16992 ( .A1(n13692), .A2(n13691), .A3(n13690), .A4(n13689), .ZN(
        n13693) );
  OAI21_X1 U16993 ( .B1(n13808), .B2(n13930), .A(n13693), .ZN(P1_U2838) );
  OR2_X1 U16994 ( .A1(n13695), .A2(n13694), .ZN(n13697) );
  AND2_X1 U16995 ( .A1(n13697), .A2(n13696), .ZN(n16644) );
  INV_X1 U16996 ( .A(n16644), .ZN(n13918) );
  NOR2_X1 U16997 ( .A1(n13918), .A2(n15448), .ZN(n13702) );
  AOI211_X1 U16998 ( .C1(n13700), .C2(n13699), .A(n15479), .B(n13698), .ZN(
        n13701) );
  AOI211_X1 U16999 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n15448), .A(n13702), .B(
        n13701), .ZN(n13703) );
  INV_X1 U17000 ( .A(n13703), .ZN(P2_U2879) );
  XNOR2_X1 U17001 ( .A(n13705), .B(n13704), .ZN(n13754) );
  INV_X1 U17002 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n13706) );
  NOR2_X1 U17003 ( .A1(n16406), .A2(n13706), .ZN(n13751) );
  NOR2_X1 U17004 ( .A1(n16260), .A2(n13707), .ZN(n13708) );
  AOI211_X1 U17005 ( .C1(n16285), .C2(n20350), .A(n13751), .B(n13708), .ZN(
        n13710) );
  NAND2_X1 U17006 ( .A1(n20355), .A2(n16286), .ZN(n13709) );
  OAI211_X1 U17007 ( .C1(n13754), .C2(n20282), .A(n13710), .B(n13709), .ZN(
        P1_U2995) );
  INV_X1 U17008 ( .A(n14959), .ZN(n13711) );
  OAI222_X1 U17009 ( .A1(n13880), .A2(n14982), .B1(n14989), .B2(n13711), .C1(
        n14987), .C2(n12125), .ZN(P1_U2901) );
  INV_X1 U17010 ( .A(n14962), .ZN(n13712) );
  OAI222_X1 U17011 ( .A1(n13930), .A2(n14982), .B1(n14989), .B2(n13712), .C1(
        n20412), .C2(n14987), .ZN(P1_U2902) );
  AND2_X1 U17012 ( .A1(n20204), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19794) );
  NAND2_X1 U17013 ( .A1(n19794), .A2(n13723), .ZN(n13713) );
  NAND3_X1 U17014 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20209), .A3(
        n20229), .ZN(n19710) );
  NAND2_X1 U17015 ( .A1(n13713), .A2(n19710), .ZN(n13716) );
  NOR2_X1 U17016 ( .A1(n20239), .A2(n19710), .ZN(n19763) );
  INV_X1 U17017 ( .A(n19763), .ZN(n13714) );
  OAI21_X1 U17018 ( .B1(n13719), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13714), 
        .ZN(n13715) );
  MUX2_X1 U17019 ( .A(n13716), .B(n13715), .S(n20202), .Z(n13717) );
  NAND2_X1 U17020 ( .A1(n13717), .A2(n20053), .ZN(n19753) );
  INV_X1 U17021 ( .A(n19753), .ZN(n19739) );
  INV_X1 U17022 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13728) );
  NOR2_X2 U17023 ( .A1(n19504), .A2(n19764), .ZN(n20047) );
  INV_X1 U17024 ( .A(n19710), .ZN(n13718) );
  NAND2_X1 U17025 ( .A1(n13718), .A2(n20196), .ZN(n13722) );
  INV_X1 U17026 ( .A(n13719), .ZN(n13720) );
  OAI21_X1 U17027 ( .B1(n13720), .B2(n9804), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13721) );
  NAND2_X1 U17028 ( .A1(n13722), .A2(n13721), .ZN(n19752) );
  INV_X1 U17029 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16772) );
  INV_X1 U17030 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18546) );
  OAI22_X2 U17031 ( .A1(n16772), .A2(n19611), .B1(n18546), .B2(n19609), .ZN(
        n20055) );
  INV_X1 U17032 ( .A(n20055), .ZN(n13725) );
  AOI22_X2 U17033 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19608), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19607), .ZN(n20058) );
  INV_X1 U17034 ( .A(n20058), .ZN(n19621) );
  AOI22_X1 U17035 ( .A1(n19771), .A2(n19621), .B1(n20046), .B2(n9804), .ZN(
        n13724) );
  OAI21_X1 U17036 ( .B1(n19748), .B2(n13725), .A(n13724), .ZN(n13726) );
  AOI21_X1 U17037 ( .B1(n20047), .B2(n19752), .A(n13726), .ZN(n13727) );
  OAI21_X1 U17038 ( .B1(n19739), .B2(n13728), .A(n13727), .ZN(P2_U3088) );
  OAI211_X1 U17039 ( .C1(n16374), .C2(n15132), .A(n15261), .B(n13729), .ZN(
        n13744) );
  NOR2_X1 U17040 ( .A1(n15147), .A2(n15281), .ZN(n15263) );
  NOR2_X1 U17041 ( .A1(n13817), .A2(n15263), .ZN(n13820) );
  AOI22_X1 U17042 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13744), .B1(
        n13820), .B2(n13741), .ZN(n13739) );
  NAND2_X1 U17043 ( .A1(n14318), .A2(n13741), .ZN(n13730) );
  OAI211_X1 U17044 ( .C1(n9653), .C2(P1_EBX_REG_3__SCAN_IN), .A(n13730), .B(
        n14291), .ZN(n13733) );
  INV_X1 U17045 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13731) );
  NAND2_X1 U17046 ( .A1(n14322), .A2(n13731), .ZN(n13732) );
  AND2_X1 U17047 ( .A1(n13733), .A2(n13732), .ZN(n13734) );
  NAND2_X1 U17048 ( .A1(n13735), .A2(n13734), .ZN(n13736) );
  AND2_X1 U17049 ( .A1(n13749), .A2(n13736), .ZN(n13878) );
  AOI21_X1 U17050 ( .B1(n20451), .B2(n13878), .A(n13737), .ZN(n13738) );
  OAI211_X1 U17051 ( .C1(n20446), .C2(n13740), .A(n13739), .B(n13738), .ZN(
        P1_U3028) );
  NOR2_X1 U17052 ( .A1(n13742), .A2(n13741), .ZN(n15133) );
  AOI21_X1 U17053 ( .B1(n13742), .B2(n13741), .A(n15133), .ZN(n13743) );
  AOI22_X1 U17054 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13744), .B1(
        n13820), .B2(n13743), .ZN(n13753) );
  INV_X1 U17055 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13745) );
  NAND2_X1 U17056 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13746) );
  OAI211_X1 U17057 ( .C1(n9653), .C2(P1_EBX_REG_4__SCAN_IN), .A(n14318), .B(
        n13746), .ZN(n13747) );
  NAND2_X1 U17058 ( .A1(n13748), .A2(n13747), .ZN(n13750) );
  AOI21_X1 U17059 ( .B1(n13750), .B2(n13749), .A(n16403), .ZN(n20345) );
  AOI21_X1 U17060 ( .B1(n20451), .B2(n20345), .A(n13751), .ZN(n13752) );
  OAI211_X1 U17061 ( .C1(n20446), .C2(n13754), .A(n13753), .B(n13752), .ZN(
        P1_U3027) );
  NAND2_X1 U17062 ( .A1(n19794), .A2(n19819), .ZN(n13755) );
  NOR2_X1 U17063 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19675) );
  NAND2_X1 U17064 ( .A1(n19675), .A2(n20229), .ZN(n19565) );
  NAND2_X1 U17065 ( .A1(n13755), .A2(n19565), .ZN(n13759) );
  OR2_X1 U17066 ( .A1(n13760), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13757) );
  NAND2_X1 U17067 ( .A1(n20229), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19853) );
  INV_X1 U17068 ( .A(n19675), .ZN(n19673) );
  NOR2_X1 U17069 ( .A1(n19853), .A2(n19673), .ZN(n19637) );
  NOR2_X1 U17070 ( .A1(n19637), .A2(n20196), .ZN(n13756) );
  AOI21_X1 U17071 ( .B1(n13757), .B2(n13756), .A(n19764), .ZN(n13758) );
  NAND2_X1 U17072 ( .A1(n13759), .A2(n13758), .ZN(n19640) );
  INV_X1 U17073 ( .A(n19640), .ZN(n19625) );
  INV_X1 U17074 ( .A(n13760), .ZN(n13761) );
  OAI21_X1 U17075 ( .B1(n13761), .B2(n19637), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13762) );
  OAI21_X1 U17076 ( .B1(n19565), .B2(n20202), .A(n13762), .ZN(n19638) );
  NOR2_X2 U17077 ( .A1(n19480), .A2(n19764), .ZN(n20078) );
  NOR2_X2 U17078 ( .A1(n10486), .A2(n19596), .ZN(n20077) );
  INV_X1 U17079 ( .A(n20077), .ZN(n19873) );
  INV_X1 U17080 ( .A(n19637), .ZN(n13764) );
  NAND2_X1 U17081 ( .A1(n19819), .A2(n19788), .ZN(n19643) );
  INV_X1 U17082 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16779) );
  INV_X1 U17083 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18565) );
  AOI22_X1 U17084 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19607), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19608), .ZN(n20082) );
  INV_X1 U17085 ( .A(n20082), .ZN(n20025) );
  AOI22_X1 U17086 ( .A1(n19669), .A2(n20079), .B1(n19639), .B2(n20025), .ZN(
        n13763) );
  OAI21_X1 U17087 ( .B1(n19873), .B2(n13764), .A(n13763), .ZN(n13765) );
  AOI21_X1 U17088 ( .B1(n19638), .B2(n20078), .A(n13765), .ZN(n13766) );
  OAI21_X1 U17089 ( .B1(n19625), .B2(n13767), .A(n13766), .ZN(P2_U3060) );
  AOI22_X1 U17090 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20400), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20409), .ZN(n13768) );
  OAI21_X1 U17091 ( .B1(n12662), .B2(n13787), .A(n13768), .ZN(P1_U2906) );
  INV_X1 U17092 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13770) );
  AOI22_X1 U17093 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13769) );
  OAI21_X1 U17094 ( .B1(n13770), .B2(n13787), .A(n13769), .ZN(P1_U2908) );
  INV_X1 U17095 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13772) );
  AOI22_X1 U17096 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13771) );
  OAI21_X1 U17097 ( .B1(n13772), .B2(n13787), .A(n13771), .ZN(P1_U2915) );
  INV_X1 U17098 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13774) );
  AOI22_X1 U17099 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13773) );
  OAI21_X1 U17100 ( .B1(n13774), .B2(n13787), .A(n13773), .ZN(P1_U2916) );
  INV_X1 U17101 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13776) );
  AOI22_X1 U17102 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13775) );
  OAI21_X1 U17103 ( .B1(n13776), .B2(n13787), .A(n13775), .ZN(P1_U2918) );
  AOI22_X1 U17104 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13777) );
  OAI21_X1 U17105 ( .B1(n14956), .B2(n13787), .A(n13777), .ZN(P1_U2917) );
  INV_X1 U17106 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13779) );
  AOI22_X1 U17107 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13778) );
  OAI21_X1 U17108 ( .B1(n13779), .B2(n13787), .A(n13778), .ZN(P1_U2920) );
  INV_X1 U17109 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13781) );
  AOI22_X1 U17110 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13780) );
  OAI21_X1 U17111 ( .B1(n13781), .B2(n13787), .A(n13780), .ZN(P1_U2919) );
  INV_X1 U17112 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13783) );
  AOI22_X1 U17113 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13782) );
  OAI21_X1 U17114 ( .B1(n13783), .B2(n13787), .A(n13782), .ZN(P1_U2910) );
  INV_X1 U17115 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13785) );
  AOI22_X1 U17116 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13784) );
  OAI21_X1 U17117 ( .B1(n13785), .B2(n13787), .A(n13784), .ZN(P1_U2912) );
  INV_X1 U17118 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U17119 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13786) );
  OAI21_X1 U17120 ( .B1(n13788), .B2(n13787), .A(n13786), .ZN(P1_U2914) );
  INV_X1 U17121 ( .A(n13789), .ZN(n13791) );
  OR2_X1 U17122 ( .A1(n14656), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13790) );
  AND2_X1 U17123 ( .A1(n13791), .A2(n13790), .ZN(n20450) );
  INV_X1 U17124 ( .A(n20450), .ZN(n13920) );
  OAI22_X1 U17125 ( .A1(n13792), .A2(n20325), .B1(n20320), .B2(n13920), .ZN(
        n13793) );
  AOI21_X1 U17126 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n14812), .A(n13793), .ZN(
        n13797) );
  AOI21_X1 U17127 ( .B1(n20365), .B2(n20375), .A(n13794), .ZN(n13795) );
  AOI21_X1 U17128 ( .B1(n20363), .B2(n20546), .A(n13795), .ZN(n13796) );
  OAI211_X1 U17129 ( .C1(n13808), .C2(n13919), .A(n13797), .B(n13796), .ZN(
        P1_U2840) );
  INV_X1 U17130 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13798) );
  NOR2_X1 U17131 ( .A1(n20365), .A2(n13798), .ZN(n13799) );
  AOI21_X1 U17132 ( .B1(n20363), .B2(n13342), .A(n13799), .ZN(n13801) );
  AOI22_X1 U17133 ( .A1(n13878), .A2(n20362), .B1(n20360), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13800) );
  OAI211_X1 U17134 ( .C1(n13802), .C2(n20375), .A(n13801), .B(n13800), .ZN(
        n13803) );
  AOI21_X1 U17135 ( .B1(n13804), .B2(P1_REIP_REG_3__SCAN_IN), .A(n13803), .ZN(
        n13807) );
  NAND2_X1 U17136 ( .A1(n20344), .A2(n20963), .ZN(n13806) );
  OAI211_X1 U17137 ( .C1(n13808), .C2(n13880), .A(n13807), .B(n13806), .ZN(
        P1_U2837) );
  XNOR2_X1 U17138 ( .A(n13604), .B(n13846), .ZN(n13813) );
  OR2_X1 U17139 ( .A1(n13810), .A2(n13809), .ZN(n13811) );
  AND2_X1 U17140 ( .A1(n13849), .A2(n13811), .ZN(n16532) );
  INV_X1 U17141 ( .A(n16532), .ZN(n16612) );
  MUX2_X1 U17142 ( .A(n16612), .B(n10584), .S(n15448), .Z(n13812) );
  OAI21_X1 U17143 ( .B1(n13813), .B2(n15479), .A(n13812), .ZN(P2_U2875) );
  XNOR2_X1 U17144 ( .A(n13815), .B(n13814), .ZN(n13844) );
  NAND2_X1 U17145 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15133), .ZN(
        n13816) );
  NOR2_X1 U17146 ( .A1(n13817), .A2(n13816), .ZN(n15258) );
  OAI21_X1 U17147 ( .B1(n15258), .B2(n16371), .A(n15261), .ZN(n16376) );
  INV_X1 U17148 ( .A(n16376), .ZN(n13818) );
  OAI221_X1 U17149 ( .B1(n16374), .B2(n15133), .C1(n16374), .C2(n15132), .A(
        n13818), .ZN(n15279) );
  INV_X1 U17150 ( .A(n15133), .ZN(n13819) );
  NOR2_X1 U17151 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13819), .ZN(
        n15280) );
  AOI22_X1 U17152 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15279), .B1(
        n15280), .B2(n13820), .ZN(n13824) );
  MUX2_X1 U17153 ( .A(n14291), .B(n14318), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n13822) );
  NAND2_X1 U17154 ( .A1(n9653), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13821) );
  NAND2_X1 U17155 ( .A1(n13822), .A2(n13821), .ZN(n16402) );
  INV_X1 U17156 ( .A(n16402), .ZN(n14084) );
  XNOR2_X1 U17157 ( .A(n16403), .B(n14084), .ZN(n20331) );
  INV_X1 U17158 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20966) );
  NOR2_X1 U17159 ( .A1(n16406), .A2(n20966), .ZN(n13840) );
  AOI21_X1 U17160 ( .B1(n20451), .B2(n20331), .A(n13840), .ZN(n13823) );
  OAI211_X1 U17161 ( .C1(n20446), .C2(n13844), .A(n13824), .B(n13823), .ZN(
        P1_U3026) );
  OR2_X1 U17162 ( .A1(n13851), .A2(n13825), .ZN(n13827) );
  AND2_X1 U17163 ( .A1(n13827), .A2(n13826), .ZN(n16599) );
  INV_X1 U17164 ( .A(n16599), .ZN(n14046) );
  INV_X1 U17165 ( .A(n13933), .ZN(n13833) );
  OAI211_X1 U17166 ( .C1(n10221), .C2(n13834), .A(n13833), .B(n15470), .ZN(
        n13836) );
  NAND2_X1 U17167 ( .A1(n15448), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13835) );
  OAI211_X1 U17168 ( .C1(n14046), .C2(n15448), .A(n13836), .B(n13835), .ZN(
        P2_U2873) );
  NAND2_X1 U17169 ( .A1(n13838), .A2(n13837), .ZN(n13839) );
  AND2_X1 U17170 ( .A1(n14016), .A2(n13839), .ZN(n20338) );
  AOI21_X1 U17171 ( .B1(n16291), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13840), .ZN(n13841) );
  OAI21_X1 U17172 ( .B1(n16299), .B2(n20332), .A(n13841), .ZN(n13842) );
  AOI21_X1 U17173 ( .B1(n20338), .B2(n16286), .A(n13842), .ZN(n13843) );
  OAI21_X1 U17174 ( .B1(n13844), .B2(n20282), .A(n13843), .ZN(P1_U2994) );
  OAI21_X1 U17175 ( .B1(n13604), .B2(n13846), .A(n13845), .ZN(n13847) );
  NAND3_X1 U17176 ( .A1(n13847), .A2(n15470), .A3(n13832), .ZN(n13853) );
  AND2_X1 U17177 ( .A1(n13849), .A2(n13848), .ZN(n13850) );
  OR2_X1 U17178 ( .A1(n13851), .A2(n13850), .ZN(n19329) );
  INV_X1 U17179 ( .A(n19329), .ZN(n16517) );
  NAND2_X1 U17180 ( .A1(n16517), .A2(n15449), .ZN(n13852) );
  OAI211_X1 U17181 ( .C1(n10590), .C2(n15449), .A(n13853), .B(n13852), .ZN(
        P2_U2874) );
  NOR2_X2 U17182 ( .A1(n20003), .A2(n19974), .ZN(n19999) );
  NOR2_X2 U17183 ( .A1(n19970), .A2(n20197), .ZN(n19965) );
  OAI21_X1 U17184 ( .B1(n19999), .B2(n19965), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13860) );
  NOR2_X1 U17185 ( .A1(n13855), .A2(n13854), .ZN(n19708) );
  NAND2_X1 U17186 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19708), .ZN(
        n13861) );
  NAND3_X1 U17187 ( .A1(n20229), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19973) );
  NOR2_X1 U17188 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19973), .ZN(
        n19963) );
  INV_X1 U17189 ( .A(n19963), .ZN(n13856) );
  AND2_X1 U17190 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13856), .ZN(n13857) );
  NAND2_X1 U17191 ( .A1(n13858), .A2(n13857), .ZN(n13863) );
  OAI211_X1 U17192 ( .C1(n19963), .C2(n20205), .A(n13863), .B(n20053), .ZN(
        n13859) );
  INV_X1 U17193 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13866) );
  AOI22_X1 U17194 ( .A1(n19965), .A2(n20055), .B1(n19999), .B2(n19621), .ZN(
        n13865) );
  OAI21_X1 U17195 ( .B1(n13861), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19761), 
        .ZN(n13862) );
  AND2_X1 U17196 ( .A1(n13863), .A2(n13862), .ZN(n19964) );
  AOI22_X1 U17197 ( .A1(n19964), .A2(n20047), .B1(n20046), .B2(n19963), .ZN(
        n13864) );
  OAI211_X1 U17198 ( .C1(n19969), .C2(n13866), .A(n13865), .B(n13864), .ZN(
        P2_U3144) );
  INV_X1 U17199 ( .A(n14950), .ZN(n13867) );
  INV_X1 U17200 ( .A(n20338), .ZN(n13882) );
  OAI222_X1 U17201 ( .A1(n14989), .A2(n13867), .B1(n14987), .B2(n12144), .C1(
        n14982), .C2(n13882), .ZN(P1_U2899) );
  INV_X1 U17202 ( .A(n13869), .ZN(n13872) );
  NAND4_X1 U17203 ( .A1(n14652), .A2(n13872), .A3(n13871), .A4(n13870), .ZN(
        n13873) );
  AOI22_X1 U17204 ( .A1(n20382), .A2(n20345), .B1(n14902), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13876) );
  OAI21_X1 U17205 ( .B1(n13877), .B2(n14914), .A(n13876), .ZN(P1_U2868) );
  AOI22_X1 U17206 ( .A1(n20382), .A2(n13878), .B1(n14902), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13879) );
  OAI21_X1 U17207 ( .B1(n13880), .B2(n14914), .A(n13879), .ZN(P1_U2869) );
  AOI22_X1 U17208 ( .A1(n20382), .A2(n20331), .B1(n14902), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n13881) );
  OAI21_X1 U17209 ( .B1(n13882), .B2(n14914), .A(n13881), .ZN(P1_U2867) );
  NOR2_X1 U17210 ( .A1(n19393), .A2(n13883), .ZN(n13884) );
  XNOR2_X1 U17211 ( .A(n13884), .B(n16538), .ZN(n13894) );
  INV_X1 U17212 ( .A(n13885), .ZN(n13886) );
  AOI22_X1 U17213 ( .A1(n13886), .A2(n12839), .B1(n19431), .B2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13887) );
  OAI21_X1 U17214 ( .B1(n19418), .B2(n10584), .A(n13887), .ZN(n13888) );
  AOI211_X1 U17215 ( .C1(n19402), .C2(P2_REIP_REG_12__SCAN_IN), .A(n16616), 
        .B(n13888), .ZN(n13892) );
  AOI21_X1 U17216 ( .B1(n13890), .B2(n16006), .A(n13889), .ZN(n19448) );
  NAND2_X1 U17217 ( .A1(n19420), .A2(n19448), .ZN(n13891) );
  OAI211_X1 U17218 ( .C1(n16612), .C2(n19389), .A(n13892), .B(n13891), .ZN(
        n13893) );
  AOI21_X1 U17219 ( .B1(n13894), .B2(n19411), .A(n13893), .ZN(n13895) );
  INV_X1 U17220 ( .A(n13895), .ZN(P2_U2843) );
  NOR2_X1 U17221 ( .A1(n19393), .A2(n16068), .ZN(n13896) );
  XNOR2_X1 U17222 ( .A(n13896), .B(n14644), .ZN(n13897) );
  NAND2_X1 U17223 ( .A1(n13897), .A2(n19411), .ZN(n13905) );
  INV_X1 U17224 ( .A(n13898), .ZN(n13900) );
  AOI22_X1 U17225 ( .A1(n19402), .A2(P2_REIP_REG_2__SCAN_IN), .B1(n19406), 
        .B2(P2_EBX_REG_2__SCAN_IN), .ZN(n13899) );
  OAI21_X1 U17226 ( .B1(n13900), .B2(n19423), .A(n13899), .ZN(n13902) );
  OAI22_X1 U17227 ( .A1(n20213), .A2(n19408), .B1(n10534), .B2(n19386), .ZN(
        n13901) );
  AOI211_X1 U17228 ( .C1(n19425), .C2(n13903), .A(n13902), .B(n13901), .ZN(
        n13904) );
  OAI211_X1 U17229 ( .C1(n19390), .C2(n20210), .A(n13905), .B(n13904), .ZN(
        P2_U2853) );
  NOR2_X1 U17230 ( .A1(n19393), .A2(n13906), .ZN(n13907) );
  XNOR2_X1 U17231 ( .A(n13907), .B(n16576), .ZN(n13908) );
  NAND2_X1 U17232 ( .A1(n13908), .A2(n19411), .ZN(n13917) );
  AOI21_X1 U17233 ( .B1(n13910), .B2(n13909), .A(n16025), .ZN(n19458) );
  AOI22_X1 U17234 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19431), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19406), .ZN(n13911) );
  OAI211_X1 U17235 ( .C1(n19416), .C2(n13912), .A(n13911), .B(n19333), .ZN(
        n13915) );
  NOR2_X1 U17236 ( .A1(n13913), .A2(n19423), .ZN(n13914) );
  AOI211_X1 U17237 ( .C1(n19420), .C2(n19458), .A(n13915), .B(n13914), .ZN(
        n13916) );
  OAI211_X1 U17238 ( .C1(n13918), .C2(n19389), .A(n13917), .B(n13916), .ZN(
        P2_U2847) );
  OAI222_X1 U17239 ( .A1(n14916), .A2(n13920), .B1(n20387), .B2(n13792), .C1(
        n14884), .C2(n13919), .ZN(P1_U2872) );
  INV_X1 U17240 ( .A(n13023), .ZN(n13922) );
  NAND2_X1 U17241 ( .A1(n13922), .A2(n13921), .ZN(n16680) );
  MUX2_X1 U17242 ( .A(n10503), .B(n16680), .S(n13923), .Z(n13924) );
  AOI21_X1 U17243 ( .B1(n13050), .B2(n16678), .A(n13924), .ZN(n16683) );
  OAI21_X1 U17244 ( .B1(n16683), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n10598), 
        .ZN(n13926) );
  OAI221_X1 U17245 ( .B1(n19393), .B2(n19426), .C1(n9658), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(P2_STATE2_REG_1__SCAN_IN), .ZN(
        n20187) );
  AOI22_X1 U17246 ( .A1(n13926), .A2(n20187), .B1(n13925), .B2(n20190), .ZN(
        n13928) );
  NAND2_X1 U17247 ( .A1(n20195), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13927) );
  OAI21_X1 U17248 ( .B1(n13928), .B2(n20195), .A(n13927), .ZN(P2_U3601) );
  OAI222_X1 U17249 ( .A1(n20359), .A2(n14916), .B1(n13532), .B2(n20387), .C1(
        n13929), .C2(n14884), .ZN(P1_U2871) );
  INV_X1 U17250 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13931) );
  OAI222_X1 U17251 ( .A1(n13932), .A2(n14916), .B1(n13931), .B2(n20387), .C1(
        n13930), .C2(n14884), .ZN(P1_U2870) );
  OAI211_X1 U17252 ( .C1(n13933), .C2(n13934), .A(n14065), .B(n15470), .ZN(
        n13939) );
  OR2_X1 U17253 ( .A1(n13936), .A2(n13935), .ZN(n13937) );
  AND2_X1 U17254 ( .A1(n14069), .A2(n13937), .ZN(n19314) );
  NAND2_X1 U17255 ( .A1(n19314), .A2(n15449), .ZN(n13938) );
  OAI211_X1 U17256 ( .C1(n10599), .C2(n15449), .A(n13939), .B(n13938), .ZN(
        P2_U2872) );
  NAND3_X1 U17257 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20692), .ZN(n15324) );
  NOR2_X1 U17258 ( .A1(n20721), .A2(n15324), .ZN(n14003) );
  INV_X1 U17259 ( .A(n14003), .ZN(n15353) );
  NOR2_X2 U17260 ( .A1(n15339), .A2(n13941), .ZN(n20902) );
  INV_X1 U17261 ( .A(n20902), .ZN(n13953) );
  INV_X1 U17262 ( .A(n15324), .ZN(n13948) );
  OR2_X1 U17263 ( .A1(n13570), .A2(n13943), .ZN(n20876) );
  OR2_X1 U17264 ( .A1(n20876), .A2(n13944), .ZN(n13945) );
  AND2_X1 U17265 ( .A1(n13945), .A2(n15353), .ZN(n13947) );
  OAI211_X1 U17266 ( .C1(n21022), .C2(n21172), .A(n20889), .B(n13947), .ZN(
        n13946) );
  OAI211_X1 U17267 ( .C1(n20889), .C2(n13948), .A(n20888), .B(n13946), .ZN(
        n15346) );
  NAND2_X1 U17268 ( .A1(n15346), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13952) );
  NOR2_X2 U17269 ( .A1(n21022), .A2(n20728), .ZN(n20870) );
  INV_X1 U17270 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n19582) );
  INV_X1 U17271 ( .A(DATAI_18_), .ZN(n21209) );
  OAI22_X1 U17272 ( .A1(n19582), .A2(n15341), .B1(n21209), .B2(n15340), .ZN(
        n20771) );
  INV_X1 U17273 ( .A(n20518), .ZN(n15322) );
  INV_X1 U17274 ( .A(n20835), .ZN(n15348) );
  INV_X1 U17275 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16768) );
  INV_X1 U17276 ( .A(DATAI_26_), .ZN(n21083) );
  OAI22_X1 U17277 ( .A1(n16768), .A2(n15341), .B1(n21083), .B2(n15340), .ZN(
        n20903) );
  NAND2_X1 U17278 ( .A1(n20464), .A2(n14962), .ZN(n20774) );
  INV_X1 U17279 ( .A(n13947), .ZN(n13949) );
  AOI22_X1 U17280 ( .A1(n13949), .A2(n20889), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13948), .ZN(n15347) );
  OAI22_X1 U17281 ( .A1(n15348), .A2(n9812), .B1(n20774), .B2(n15347), .ZN(
        n13950) );
  AOI21_X1 U17282 ( .B1(n20870), .B2(n20771), .A(n13950), .ZN(n13951) );
  OAI211_X1 U17283 ( .C1(n15353), .C2(n13953), .A(n13952), .B(n13951), .ZN(
        P1_U3139) );
  NAND2_X1 U17284 ( .A1(n13968), .A2(n13954), .ZN(n20476) );
  NAND2_X1 U17285 ( .A1(n15346), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13957) );
  INV_X1 U17286 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16781) );
  INV_X1 U17287 ( .A(DATAI_19_), .ZN(n21231) );
  INV_X1 U17288 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19586) );
  INV_X1 U17289 ( .A(DATAI_27_), .ZN(n21191) );
  OAI22_X1 U17290 ( .A1(n19586), .A2(n15341), .B1(n21191), .B2(n15340), .ZN(
        n20857) );
  INV_X1 U17291 ( .A(n20857), .ZN(n20912) );
  NAND2_X1 U17292 ( .A1(n20464), .A2(n14959), .ZN(n20777) );
  OAI22_X1 U17293 ( .A1(n15348), .A2(n20912), .B1(n15347), .B2(n20777), .ZN(
        n13955) );
  AOI21_X1 U17294 ( .B1(n20870), .B2(n20909), .A(n13955), .ZN(n13956) );
  OAI211_X1 U17295 ( .C1(n15353), .C2(n20476), .A(n13957), .B(n13956), .ZN(
        P1_U3140) );
  NAND2_X1 U17296 ( .A1(n13968), .A2(n13958), .ZN(n20471) );
  NAND2_X1 U17297 ( .A1(n15346), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13963) );
  INV_X1 U17298 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n19576) );
  INV_X1 U17299 ( .A(DATAI_17_), .ZN(n13959) );
  OAI22_X1 U17300 ( .A1(n19576), .A2(n15341), .B1(n13959), .B2(n15340), .ZN(
        n20823) );
  INV_X1 U17301 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16770) );
  INV_X1 U17302 ( .A(DATAI_25_), .ZN(n13960) );
  OAI22_X1 U17303 ( .A1(n16770), .A2(n15341), .B1(n13960), .B2(n15340), .ZN(
        n20897) );
  NAND2_X1 U17304 ( .A1(n20464), .A2(n14965), .ZN(n20770) );
  OAI22_X1 U17305 ( .A1(n15348), .A2(n9810), .B1(n15347), .B2(n20770), .ZN(
        n13961) );
  AOI21_X1 U17306 ( .B1(n20870), .B2(n20823), .A(n13961), .ZN(n13962) );
  OAI211_X1 U17307 ( .C1(n15353), .C2(n20471), .A(n13963), .B(n13962), .ZN(
        P1_U3138) );
  NAND2_X1 U17308 ( .A1(n13968), .A2(n14265), .ZN(n20481) );
  NAND2_X1 U17309 ( .A1(n15346), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13966) );
  INV_X1 U17310 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19595) );
  INV_X1 U17311 ( .A(DATAI_21_), .ZN(n21171) );
  OAI22_X1 U17312 ( .A1(n19595), .A2(n15341), .B1(n21171), .B2(n15340), .ZN(
        n20828) );
  INV_X1 U17313 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16763) );
  INV_X1 U17314 ( .A(DATAI_29_), .ZN(n21160) );
  INV_X1 U17315 ( .A(n20921), .ZN(n20831) );
  NAND2_X1 U17316 ( .A1(n20464), .A2(n14950), .ZN(n20784) );
  OAI22_X1 U17317 ( .A1(n15348), .A2(n20831), .B1(n15347), .B2(n20784), .ZN(
        n13964) );
  AOI21_X1 U17318 ( .B1(n20870), .B2(n20828), .A(n13964), .ZN(n13965) );
  OAI211_X1 U17319 ( .C1(n15353), .C2(n20481), .A(n13966), .B(n13965), .ZN(
        P1_U3142) );
  NAND2_X1 U17320 ( .A1(n13968), .A2(n13967), .ZN(n20484) );
  NAND2_X1 U17321 ( .A1(n15346), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13972) );
  INV_X1 U17322 ( .A(DATAI_22_), .ZN(n13969) );
  INV_X1 U17323 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16776) );
  OAI22_X1 U17324 ( .A1(n13969), .A2(n15340), .B1(n16776), .B2(n15341), .ZN(
        n20832) );
  INV_X1 U17325 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19601) );
  INV_X1 U17326 ( .A(DATAI_30_), .ZN(n21069) );
  OAI22_X1 U17327 ( .A1(n19601), .A2(n15341), .B1(n21069), .B2(n15340), .ZN(
        n20927) );
  NAND2_X1 U17328 ( .A1(n20464), .A2(n14942), .ZN(n20787) );
  OAI22_X1 U17329 ( .A1(n15348), .A2(n9808), .B1(n15347), .B2(n20787), .ZN(
        n13970) );
  AOI21_X1 U17330 ( .B1(n20870), .B2(n20832), .A(n13970), .ZN(n13971) );
  OAI211_X1 U17331 ( .C1(n15353), .C2(n20484), .A(n13972), .B(n13971), .ZN(
        P1_U3143) );
  INV_X1 U17332 ( .A(n15346), .ZN(n14007) );
  INV_X1 U17333 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13976) );
  NOR2_X2 U17334 ( .A1(n15339), .A2(n14347), .ZN(n20933) );
  INV_X1 U17335 ( .A(DATAI_23_), .ZN(n21061) );
  INV_X1 U17336 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16774) );
  OAI22_X1 U17337 ( .A1(n21061), .A2(n15340), .B1(n16774), .B2(n15341), .ZN(
        n20937) );
  INV_X1 U17338 ( .A(DATAI_31_), .ZN(n21222) );
  INV_X1 U17339 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19612) );
  AOI22_X1 U17340 ( .A1(n20870), .A2(n20937), .B1(n20835), .B2(n20869), .ZN(
        n13973) );
  OAI21_X1 U17341 ( .B1(n20793), .B2(n15347), .A(n13973), .ZN(n13974) );
  AOI21_X1 U17342 ( .B1(n14003), .B2(n20933), .A(n13974), .ZN(n13975) );
  OAI21_X1 U17343 ( .B1(n14007), .B2(n13976), .A(n13975), .ZN(P1_U3144) );
  NAND2_X1 U17344 ( .A1(n13978), .A2(n13977), .ZN(n13980) );
  XNOR2_X1 U17345 ( .A(n13980), .B(n13979), .ZN(n14000) );
  XOR2_X1 U17346 ( .A(n13982), .B(n13981), .Z(n13998) );
  OAI22_X1 U17347 ( .A1(n16593), .A2(n13983), .B1(n20136), .B2(n19333), .ZN(
        n13984) );
  AOI21_X1 U17348 ( .B1(n16583), .B2(n13985), .A(n13984), .ZN(n13986) );
  OAI21_X1 U17349 ( .B1(n11339), .B2(n19559), .A(n13986), .ZN(n13987) );
  AOI21_X1 U17350 ( .B1(n13998), .B2(n19554), .A(n13987), .ZN(n13988) );
  OAI21_X1 U17351 ( .B1(n14000), .B2(n16586), .A(n13988), .ZN(P2_U3011) );
  NOR2_X1 U17352 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14625), .ZN(
        n15734) );
  INV_X1 U17353 ( .A(n15734), .ZN(n14623) );
  NAND2_X1 U17354 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14625), .ZN(
        n14624) );
  INV_X1 U17355 ( .A(n14624), .ZN(n13989) );
  OR2_X1 U17356 ( .A1(n15940), .A2(n13989), .ZN(n13990) );
  AND2_X1 U17357 ( .A1(n13990), .A2(n14629), .ZN(n15736) );
  OAI21_X1 U17358 ( .B1(n15944), .B2(n14623), .A(n15736), .ZN(n16038) );
  OR2_X1 U17359 ( .A1(n15944), .A2(n15734), .ZN(n13992) );
  OR2_X1 U17360 ( .A1(n15940), .A2(n14624), .ZN(n13991) );
  NAND2_X1 U17361 ( .A1(n13992), .A2(n13991), .ZN(n15751) );
  INV_X1 U17362 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15732) );
  NOR2_X1 U17363 ( .A1(n20136), .A2(n19333), .ZN(n13993) );
  AOI21_X1 U17364 ( .B1(n15751), .B2(n15732), .A(n13993), .ZN(n13994) );
  OAI21_X1 U17365 ( .B1(n20206), .B2(n16624), .A(n13994), .ZN(n13995) );
  AOI21_X1 U17366 ( .B1(n16038), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13995), .ZN(n13996) );
  OAI21_X1 U17367 ( .B1(n11339), .B2(n16629), .A(n13996), .ZN(n13997) );
  AOI21_X1 U17368 ( .B1(n13998), .B2(n16646), .A(n13997), .ZN(n13999) );
  OAI21_X1 U17369 ( .B1(n14000), .B2(n16651), .A(n13999), .ZN(P2_U3043) );
  INV_X1 U17370 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14006) );
  INV_X1 U17371 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16785) );
  INV_X1 U17372 ( .A(DATAI_16_), .ZN(n21224) );
  OAI22_X1 U17373 ( .A1(n16785), .A2(n15341), .B1(n21224), .B2(n15340), .ZN(
        n20757) );
  INV_X1 U17374 ( .A(DATAI_24_), .ZN(n21214) );
  OAI22_X1 U17375 ( .A1(n21214), .A2(n15340), .B1(n16772), .B2(n15341), .ZN(
        n20891) );
  NAND2_X1 U17376 ( .A1(n20464), .A2(n14971), .ZN(n20767) );
  OAI22_X1 U17377 ( .A1(n15348), .A2(n9806), .B1(n20767), .B2(n15347), .ZN(
        n14001) );
  AOI21_X1 U17378 ( .B1(n20870), .B2(n20757), .A(n14001), .ZN(n14005) );
  NOR2_X2 U17379 ( .A1(n15339), .A2(n14002), .ZN(n20881) );
  NAND2_X1 U17380 ( .A1(n20881), .A2(n14003), .ZN(n14004) );
  OAI211_X1 U17381 ( .C1(n14007), .C2(n14006), .A(n14005), .B(n14004), .ZN(
        P1_U3137) );
  AOI21_X1 U17382 ( .B1(n14105), .B2(n14009), .A(n14010), .ZN(n14011) );
  OR2_X1 U17383 ( .A1(n14008), .A2(n14011), .ZN(n15129) );
  INV_X1 U17384 ( .A(DATAI_8_), .ZN(n21166) );
  NAND2_X1 U17385 ( .A1(n14923), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14012) );
  OAI21_X1 U17386 ( .B1(n14923), .B2(n21166), .A(n14012), .ZN(n20417) );
  AOI22_X1 U17387 ( .A1(n14980), .A2(n20417), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14979), .ZN(n14013) );
  OAI21_X1 U17388 ( .B1(n15129), .B2(n14982), .A(n14013), .ZN(P1_U2896) );
  XNOR2_X1 U17389 ( .A(n14015), .B(n14014), .ZN(n16411) );
  AOI21_X1 U17390 ( .B1(n14017), .B2(n14016), .A(n14105), .ZN(n20384) );
  AOI22_X1 U17391 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n14018) );
  OAI21_X1 U17392 ( .B1(n16299), .B2(n20330), .A(n14018), .ZN(n14019) );
  AOI21_X1 U17393 ( .B1(n20384), .B2(n16286), .A(n14019), .ZN(n14020) );
  OAI21_X1 U17394 ( .B1(n20282), .B2(n16411), .A(n14020), .ZN(P1_U2993) );
  INV_X1 U17395 ( .A(n14942), .ZN(n14022) );
  INV_X1 U17396 ( .A(n20384), .ZN(n14021) );
  OAI222_X1 U17397 ( .A1(n14989), .A2(n14022), .B1(n14987), .B2(n12153), .C1(
        n14982), .C2(n14021), .ZN(P1_U2898) );
  NAND2_X1 U17398 ( .A1(n14024), .A2(n14023), .ZN(n14025) );
  XNOR2_X1 U17399 ( .A(n14025), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19555) );
  INV_X1 U17400 ( .A(n19555), .ZN(n14039) );
  XNOR2_X1 U17401 ( .A(n14026), .B(n10302), .ZN(n19553) );
  NAND2_X1 U17402 ( .A1(n14028), .A2(n14027), .ZN(n14029) );
  NAND2_X1 U17403 ( .A1(n14030), .A2(n14029), .ZN(n19558) );
  NAND2_X1 U17404 ( .A1(n14031), .A2(n13633), .ZN(n14033) );
  INV_X1 U17405 ( .A(n14130), .ZN(n14032) );
  AND2_X1 U17406 ( .A1(n14033), .A2(n14032), .ZN(n19474) );
  NAND2_X1 U17407 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15751), .ZN(
        n16056) );
  INV_X1 U17408 ( .A(n16609), .ZN(n15741) );
  AOI21_X1 U17409 ( .B1(n15732), .B2(n15741), .A(n16038), .ZN(n14131) );
  INV_X1 U17410 ( .A(n19333), .ZN(n16616) );
  NAND2_X1 U17411 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n16616), .ZN(n14034) );
  OAI221_X1 U17412 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16056), .C1(
        n14127), .C2(n14131), .A(n14034), .ZN(n14035) );
  AOI21_X1 U17413 ( .B1(n16643), .B2(n19474), .A(n14035), .ZN(n14036) );
  OAI21_X1 U17414 ( .B1(n16629), .B2(n19558), .A(n14036), .ZN(n14037) );
  AOI21_X1 U17415 ( .B1(n19553), .B2(n16600), .A(n14037), .ZN(n14038) );
  OAI21_X1 U17416 ( .B1(n16630), .B2(n14039), .A(n14038), .ZN(P2_U3042) );
  INV_X1 U17417 ( .A(n14040), .ZN(n14051) );
  NOR2_X1 U17418 ( .A1(n19393), .A2(n19319), .ZN(n14041) );
  XNOR2_X1 U17419 ( .A(n14041), .B(n16513), .ZN(n14042) );
  NAND2_X1 U17420 ( .A1(n14042), .A2(n19411), .ZN(n14050) );
  AOI21_X1 U17421 ( .B1(n14043), .B2(n15987), .A(n15969), .ZN(n19443) );
  AOI22_X1 U17422 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19431), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19406), .ZN(n14044) );
  OAI211_X1 U17423 ( .C1(n19416), .C2(n14045), .A(n14044), .B(n19364), .ZN(
        n14048) );
  NOR2_X1 U17424 ( .A1(n14046), .A2(n19389), .ZN(n14047) );
  AOI211_X1 U17425 ( .C1(n19420), .C2(n19443), .A(n14048), .B(n14047), .ZN(
        n14049) );
  OAI211_X1 U17426 ( .C1(n19423), .C2(n14051), .A(n14050), .B(n14049), .ZN(
        P2_U2841) );
  INV_X1 U17427 ( .A(n14065), .ZN(n14067) );
  AOI22_X1 U17428 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n10744), .B1(
        n10779), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U17429 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U17430 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14053) );
  AOI22_X1 U17431 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14052) );
  NAND4_X1 U17432 ( .A1(n14055), .A2(n14054), .A3(n14053), .A4(n14052), .ZN(
        n14064) );
  AOI22_X1 U17433 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U17434 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14061) );
  INV_X1 U17435 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14057) );
  NAND2_X1 U17436 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n14437), .ZN(
        n14056) );
  OAI21_X1 U17437 ( .B1(n14440), .B2(n14057), .A(n14056), .ZN(n14058) );
  AOI21_X1 U17438 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n14058), .ZN(n14060) );
  NAND2_X1 U17439 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14059) );
  NAND4_X1 U17440 ( .A1(n14062), .A2(n14061), .A3(n14060), .A4(n14059), .ZN(
        n14063) );
  OR2_X1 U17441 ( .A1(n14064), .A2(n14063), .ZN(n14066) );
  OAI21_X1 U17442 ( .B1(n14067), .B2(n14066), .A(n10224), .ZN(n14123) );
  INV_X1 U17443 ( .A(n15474), .ZN(n14068) );
  AOI21_X1 U17444 ( .B1(n14070), .B2(n14069), .A(n14068), .ZN(n19301) );
  NOR2_X1 U17445 ( .A1(n15449), .A2(n14071), .ZN(n14072) );
  AOI21_X1 U17446 ( .B1(n19301), .B2(n15449), .A(n14072), .ZN(n14073) );
  OAI21_X1 U17447 ( .B1(n14123), .B2(n15479), .A(n14073), .ZN(P2_U2871) );
  NOR2_X1 U17448 ( .A1(n14008), .A2(n14075), .ZN(n14076) );
  OR2_X1 U17449 ( .A1(n14074), .A2(n14076), .ZN(n15118) );
  NAND3_X1 U17450 ( .A1(n20344), .A2(P1_REIP_REG_4__SCAN_IN), .A3(
        P1_REIP_REG_3__SCAN_IN), .ZN(n20343) );
  NAND4_X1 U17451 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14077)
         );
  INV_X1 U17452 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20972) );
  INV_X1 U17453 ( .A(n14077), .ZN(n14080) );
  NAND2_X1 U17454 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .ZN(n14079) );
  NOR2_X1 U17455 ( .A1(n14079), .A2(n14078), .ZN(n20305) );
  NAND2_X1 U17456 ( .A1(n14080), .A2(n20305), .ZN(n14327) );
  NAND2_X1 U17457 ( .A1(n14327), .A2(n14812), .ZN(n20299) );
  NOR2_X1 U17458 ( .A1(n20299), .A2(n20972), .ZN(n14103) );
  INV_X1 U17459 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20386) );
  NAND2_X1 U17460 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14081) );
  OAI211_X1 U17461 ( .C1(n9653), .C2(P1_EBX_REG_6__SCAN_IN), .A(n14318), .B(
        n14081), .ZN(n14082) );
  NAND2_X1 U17462 ( .A1(n14083), .A2(n14082), .ZN(n16400) );
  NOR2_X1 U17463 ( .A1(n14084), .A2(n16400), .ZN(n14085) );
  MUX2_X1 U17464 ( .A(n14291), .B(n14318), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n14087) );
  NAND2_X1 U17465 ( .A1(n9653), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14086) );
  NAND2_X1 U17466 ( .A1(n14087), .A2(n14086), .ZN(n15287) );
  INV_X1 U17467 ( .A(n15287), .ZN(n14091) );
  INV_X1 U17468 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n20379) );
  NAND2_X1 U17469 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14088) );
  OAI211_X1 U17470 ( .C1(n9653), .C2(P1_EBX_REG_8__SCAN_IN), .A(n14318), .B(
        n14088), .ZN(n14089) );
  NAND2_X1 U17471 ( .A1(n14090), .A2(n14089), .ZN(n15288) );
  NOR2_X1 U17472 ( .A1(n14091), .A2(n15288), .ZN(n14092) );
  NAND2_X1 U17473 ( .A1(n16405), .A2(n14092), .ZN(n15290) );
  MUX2_X1 U17474 ( .A(n14291), .B(n14318), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n14095) );
  NAND2_X1 U17475 ( .A1(n9653), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14094) );
  AND2_X1 U17476 ( .A1(n14095), .A2(n14094), .ZN(n14096) );
  NAND2_X1 U17477 ( .A1(n15290), .A2(n14096), .ZN(n14097) );
  NAND2_X1 U17478 ( .A1(n14170), .A2(n14097), .ZN(n15272) );
  INV_X1 U17479 ( .A(n15272), .ZN(n14098) );
  AOI22_X1 U17480 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n20360), .B1(n20362), .B2(
        n14098), .ZN(n14101) );
  NAND3_X1 U17481 ( .A1(n20889), .A2(n16420), .A3(n14099), .ZN(n20308) );
  AOI21_X1 U17482 ( .B1(n20348), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20346), .ZN(n14100) );
  OAI211_X1 U17483 ( .C1(n15120), .C2(n20375), .A(n14101), .B(n14100), .ZN(
        n14102) );
  AOI211_X1 U17484 ( .C1(n16235), .C2(n20972), .A(n14103), .B(n14102), .ZN(
        n14104) );
  OAI21_X1 U17485 ( .B1(n14864), .B2(n15118), .A(n14104), .ZN(P1_U2831) );
  XOR2_X1 U17486 ( .A(n14105), .B(n14009), .Z(n20316) );
  INV_X1 U17487 ( .A(n20316), .ZN(n14143) );
  INV_X1 U17488 ( .A(n14939), .ZN(n14106) );
  OAI222_X1 U17489 ( .A1(n14982), .A2(n14143), .B1(n14989), .B2(n14106), .C1(
        n14987), .C2(n12077), .ZN(P1_U2897) );
  OAI21_X1 U17490 ( .B1(n14074), .B2(n14108), .A(n14107), .ZN(n16242) );
  INV_X1 U17491 ( .A(DATAI_10_), .ZN(n21175) );
  NAND2_X1 U17492 ( .A1(n14923), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14109) );
  OAI21_X1 U17493 ( .B1(n14923), .B2(n21175), .A(n14109), .ZN(n20419) );
  AOI22_X1 U17494 ( .A1(n14980), .A2(n20419), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14979), .ZN(n14110) );
  OAI21_X1 U17495 ( .B1(n16242), .B2(n14982), .A(n14110), .ZN(P1_U2894) );
  INV_X1 U17496 ( .A(n14933), .ZN(n14112) );
  OAI222_X1 U17497 ( .A1(n15118), .A2(n14982), .B1(n14989), .B2(n14112), .C1(
        n14111), .C2(n14987), .ZN(P1_U2895) );
  OAI21_X1 U17498 ( .B1(n14114), .B2(n14113), .A(n9685), .ZN(n19302) );
  INV_X1 U17499 ( .A(n19302), .ZN(n14121) );
  OAI22_X1 U17500 ( .A1(n15558), .A2(n19504), .B1(n19466), .B2(n14115), .ZN(
        n14120) );
  NOR2_X1 U17501 ( .A1(n14117), .A2(n14611), .ZN(n19436) );
  INV_X1 U17502 ( .A(n19436), .ZN(n15561) );
  NOR2_X1 U17503 ( .A1(n14117), .A2(n14116), .ZN(n19438) );
  INV_X1 U17504 ( .A(n19438), .ZN(n15560) );
  INV_X1 U17505 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n14118) );
  OAI22_X1 U17506 ( .A1(n15561), .A2(n16785), .B1(n15560), .B2(n14118), .ZN(
        n14119) );
  AOI211_X1 U17507 ( .C1(n19495), .C2(n14121), .A(n14120), .B(n14119), .ZN(
        n14122) );
  OAI21_X1 U17508 ( .B1(n14123), .B2(n19490), .A(n14122), .ZN(P2_U2903) );
  XNOR2_X1 U17509 ( .A(n14124), .B(n14125), .ZN(n16587) );
  NAND2_X1 U17510 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16057) );
  INV_X1 U17511 ( .A(n16057), .ZN(n14126) );
  AOI211_X1 U17512 ( .C1(n14128), .C2(n14127), .A(n14126), .B(n16056), .ZN(
        n14135) );
  OAI21_X1 U17513 ( .B1(n14130), .B2(n14129), .A(n16052), .ZN(n19472) );
  INV_X1 U17514 ( .A(n14131), .ZN(n14132) );
  INV_X1 U17515 ( .A(n19333), .ZN(n15989) );
  AOI22_X1 U17516 ( .A1(n14132), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n15989), .B2(P2_REIP_REG_5__SCAN_IN), .ZN(n14133) );
  OAI21_X1 U17517 ( .B1(n19472), .B2(n16624), .A(n14133), .ZN(n14134) );
  AOI211_X1 U17518 ( .C1(n19382), .C2(n16645), .A(n14135), .B(n14134), .ZN(
        n14141) );
  AND2_X1 U17519 ( .A1(n14137), .A2(n14136), .ZN(n14138) );
  OAI22_X1 U17520 ( .A1(n11657), .A2(n10278), .B1(n14139), .B2(n14138), .ZN(
        n16585) );
  OR2_X1 U17521 ( .A1(n16585), .A2(n16630), .ZN(n14140) );
  OAI211_X1 U17522 ( .C1(n16587), .C2(n16651), .A(n14141), .B(n14140), .ZN(
        P2_U3041) );
  INV_X1 U17523 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14142) );
  OAI222_X1 U17524 ( .A1(n15272), .A2(n14916), .B1(n20387), .B2(n14142), .C1(
        n14884), .C2(n15118), .ZN(P1_U2863) );
  INV_X1 U17525 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14144) );
  XNOR2_X1 U17526 ( .A(n16405), .B(n15287), .ZN(n20312) );
  OAI222_X1 U17527 ( .A1(n14144), .A2(n20387), .B1(n14916), .B2(n20312), .C1(
        n14914), .C2(n14143), .ZN(P1_U2865) );
  AOI22_X1 U17528 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10779), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U17529 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U17530 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U17531 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14145) );
  NAND4_X1 U17532 ( .A1(n14148), .A2(n14147), .A3(n14146), .A4(n14145), .ZN(
        n14157) );
  AOI22_X1 U17533 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14155) );
  AOI22_X1 U17534 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14154) );
  NAND2_X1 U17535 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14437), .ZN(
        n14149) );
  OAI21_X1 U17536 ( .B1(n14440), .B2(n14150), .A(n14149), .ZN(n14151) );
  AOI21_X1 U17537 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n14151), .ZN(n14153) );
  NAND2_X1 U17538 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n14152) );
  NAND4_X1 U17539 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        n14156) );
  OR2_X1 U17540 ( .A1(n14157), .A2(n14156), .ZN(n14159) );
  INV_X1 U17541 ( .A(n14363), .ZN(n15468) );
  OAI21_X1 U17542 ( .B1(n14158), .B2(n14159), .A(n15468), .ZN(n15480) );
  INV_X1 U17543 ( .A(n14160), .ZN(n14161) );
  XNOR2_X1 U17544 ( .A(n14161), .B(n9685), .ZN(n19293) );
  OAI22_X1 U17545 ( .A1(n15558), .A2(n19578), .B1(n14162), .B2(n19466), .ZN(
        n14165) );
  INV_X1 U17546 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14163) );
  OAI22_X1 U17547 ( .A1(n15561), .A2(n19576), .B1(n15560), .B2(n14163), .ZN(
        n14164) );
  AOI211_X1 U17548 ( .C1(n19495), .C2(n19293), .A(n14165), .B(n14164), .ZN(
        n14166) );
  OAI21_X1 U17549 ( .B1(n15480), .B2(n19490), .A(n14166), .ZN(P2_U2902) );
  INV_X1 U17550 ( .A(n14167), .ZN(n14168) );
  OAI21_X1 U17551 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n14656), .A(
        n14168), .ZN(n14169) );
  NAND2_X1 U17552 ( .A1(n14170), .A2(n14169), .ZN(n14171) );
  NAND2_X1 U17553 ( .A1(n14908), .A2(n14171), .ZN(n16236) );
  INV_X1 U17554 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14172) );
  OAI222_X1 U17555 ( .A1(n16236), .A2(n14916), .B1(n14172), .B2(n20387), .C1(
        n16242), .C2(n14884), .ZN(P1_U2862) );
  AND2_X1 U17556 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17302) );
  INV_X1 U17557 ( .A(n18991), .ZN(n16108) );
  INV_X1 U17558 ( .A(n19206), .ZN(n19044) );
  NAND2_X1 U17559 ( .A1(n17711), .A2(n9669), .ZN(n17585) );
  INV_X2 U17560 ( .A(n17583), .ZN(n17578) );
  INV_X1 U17561 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17265) );
  INV_X1 U17562 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16975) );
  INV_X1 U17563 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17343) );
  INV_X1 U17564 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17357) );
  INV_X1 U17565 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17400) );
  INV_X1 U17566 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17054) );
  INV_X1 U17567 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17464) );
  AND2_X1 U17568 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17575) );
  NAND2_X1 U17569 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17575), .ZN(n17570) );
  INV_X1 U17570 ( .A(n17570), .ZN(n14175) );
  NAND4_X1 U17571 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17581), .A4(n14175), .ZN(n17564) );
  NAND4_X1 U17572 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_7__SCAN_IN), .ZN(n14176) );
  NOR2_X1 U17573 ( .A1(n17564), .A2(n14176), .ZN(n14177) );
  NAND4_X1 U17574 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n14177), .ZN(n17495) );
  INV_X1 U17575 ( .A(n17495), .ZN(n17465) );
  NAND2_X1 U17576 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17444), .ZN(n17417) );
  NOR2_X2 U17577 ( .A1(n17054), .A2(n17417), .ZN(n17415) );
  NAND2_X1 U17578 ( .A1(n17711), .A2(n17372), .ZN(n17344) );
  NOR2_X2 U17579 ( .A1(n17343), .A2(n17344), .ZN(n17327) );
  NAND2_X1 U17580 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17327), .ZN(n17321) );
  NOR2_X2 U17581 ( .A1(n16975), .A2(n17321), .ZN(n17326) );
  NAND2_X1 U17582 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17326), .ZN(n17312) );
  NOR2_X2 U17583 ( .A1(n17265), .A2(n17312), .ZN(n17317) );
  NAND2_X1 U17584 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17317), .ZN(n17308) );
  NAND2_X1 U17585 ( .A1(n17578), .A2(n17308), .ZN(n17306) );
  OAI21_X1 U17586 ( .B1(n17302), .B2(n17585), .A(n17306), .ZN(n17303) );
  AOI22_X1 U17587 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14178) );
  OAI21_X1 U17588 ( .B1(n17500), .B2(n16085), .A(n14178), .ZN(n14188) );
  AOI22_X1 U17589 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14186) );
  OAI22_X1 U17590 ( .A1(n9652), .A2(n17347), .B1(n10316), .B2(n14179), .ZN(
        n14184) );
  AOI22_X1 U17591 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14182) );
  AOI22_X1 U17592 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14181) );
  AOI22_X1 U17593 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14180) );
  NAND3_X1 U17594 ( .A1(n14182), .A2(n14181), .A3(n14180), .ZN(n14183) );
  AOI211_X1 U17595 ( .C1(n17497), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n14184), .B(n14183), .ZN(n14185) );
  OAI211_X1 U17596 ( .C1(n17274), .C2(n18796), .A(n14186), .B(n14185), .ZN(
        n14187) );
  AOI211_X1 U17597 ( .C1(n17540), .C2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n14188), .B(n14187), .ZN(n14257) );
  AOI22_X1 U17598 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14189) );
  OAI21_X1 U17599 ( .B1(n17500), .B2(n17486), .A(n14189), .ZN(n14200) );
  AOI22_X1 U17600 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14197) );
  OAI22_X1 U17601 ( .A1(n17274), .A2(n18790), .B1(n11036), .B2(n14190), .ZN(
        n14195) );
  AOI22_X1 U17602 ( .A1(n14248), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14193) );
  AOI22_X1 U17603 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14192) );
  AOI22_X1 U17604 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14191) );
  NAND3_X1 U17605 ( .A1(n14193), .A2(n14192), .A3(n14191), .ZN(n14194) );
  AOI211_X1 U17606 ( .C1(n9670), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n14195), .B(n14194), .ZN(n14196) );
  OAI211_X1 U17607 ( .C1(n14198), .C2(n18760), .A(n14197), .B(n14196), .ZN(
        n14199) );
  AOI211_X1 U17608 ( .C1(n9647), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n14200), .B(n14199), .ZN(n17309) );
  AOI22_X1 U17609 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14201) );
  OAI21_X1 U17610 ( .B1(n14202), .B2(n10316), .A(n14201), .ZN(n14213) );
  AOI22_X1 U17611 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9651), .ZN(n14210) );
  INV_X1 U17612 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17523) );
  AOI22_X1 U17613 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17541), .ZN(n14203) );
  OAI21_X1 U17614 ( .B1(n17523), .B2(n10314), .A(n14203), .ZN(n14208) );
  AOI22_X1 U17615 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17544), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n9648), .ZN(n14205) );
  AOI22_X1 U17616 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17501), .ZN(n14204) );
  OAI211_X1 U17617 ( .C1(n14206), .C2(n17526), .A(n14205), .B(n14204), .ZN(
        n14207) );
  AOI211_X1 U17618 ( .C1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .C2(n17433), .A(
        n14208), .B(n14207), .ZN(n14209) );
  OAI211_X1 U17619 ( .C1(n17468), .C2(n14211), .A(n14210), .B(n14209), .ZN(
        n14212) );
  AOI211_X1 U17620 ( .C1(n9647), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n14213), .B(n14212), .ZN(n17318) );
  AOI22_X1 U17621 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14223) );
  AOI22_X1 U17622 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14222) );
  AOI22_X1 U17623 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14221) );
  OAI22_X1 U17624 ( .A1(n17274), .A2(n18782), .B1(n11036), .B2(n17419), .ZN(
        n14219) );
  AOI22_X1 U17625 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14217) );
  AOI22_X1 U17626 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14216) );
  AOI22_X1 U17627 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14215) );
  NAND2_X1 U17628 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14214) );
  NAND4_X1 U17629 ( .A1(n14217), .A2(n14216), .A3(n14215), .A4(n14214), .ZN(
        n14218) );
  AOI211_X1 U17630 ( .C1(n17544), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n14219), .B(n14218), .ZN(n14220) );
  NAND4_X1 U17631 ( .A1(n14223), .A2(n14222), .A3(n14221), .A4(n14220), .ZN(
        n17323) );
  AOI22_X1 U17632 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14233) );
  AOI22_X1 U17633 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14224) );
  OAI21_X1 U17634 ( .B1(n17388), .B2(n17282), .A(n14224), .ZN(n14231) );
  OAI22_X1 U17635 ( .A1(n9652), .A2(n18590), .B1(n17526), .B2(n17442), .ZN(
        n14225) );
  AOI21_X1 U17636 ( .B1(n17497), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n14225), .ZN(n14229) );
  AOI22_X1 U17637 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14228) );
  AOI22_X1 U17638 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U17639 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14226) );
  NAND4_X1 U17640 ( .A1(n14229), .A2(n14228), .A3(n14227), .A4(n14226), .ZN(
        n14230) );
  AOI211_X1 U17641 ( .C1(n17544), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n14231), .B(n14230), .ZN(n14232) );
  OAI211_X1 U17642 ( .C1(n11021), .C2(n14234), .A(n14233), .B(n14232), .ZN(
        n17324) );
  NAND2_X1 U17643 ( .A1(n17323), .A2(n17324), .ZN(n17322) );
  NOR2_X1 U17644 ( .A1(n17318), .A2(n17322), .ZN(n17315) );
  AOI22_X1 U17645 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14245) );
  AOI22_X1 U17646 ( .A1(n14248), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14235) );
  OAI21_X1 U17647 ( .B1(n17500), .B2(n17498), .A(n14235), .ZN(n14243) );
  AOI22_X1 U17648 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U17649 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14237) );
  AOI22_X1 U17650 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14236) );
  OAI211_X1 U17651 ( .C1(n11036), .C2(n14238), .A(n14237), .B(n14236), .ZN(
        n14239) );
  AOI21_X1 U17652 ( .B1(n9641), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(n14239), .ZN(n14240) );
  OAI211_X1 U17653 ( .C1(n17526), .C2(n17499), .A(n14241), .B(n14240), .ZN(
        n14242) );
  AOI211_X1 U17654 ( .C1(n17497), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n14243), .B(n14242), .ZN(n14244) );
  OAI211_X1 U17655 ( .C1(n9709), .C2(n18560), .A(n14245), .B(n14244), .ZN(
        n17314) );
  NAND2_X1 U17656 ( .A1(n17315), .A2(n17314), .ZN(n17313) );
  NOR2_X1 U17657 ( .A1(n17309), .A2(n17313), .ZN(n17609) );
  AOI22_X1 U17658 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14256) );
  INV_X1 U17659 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U17660 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9649), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14247) );
  AOI22_X1 U17661 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14246) );
  OAI211_X1 U17662 ( .C1(n17526), .C2(n17470), .A(n14247), .B(n14246), .ZN(
        n14254) );
  AOI22_X1 U17663 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14252) );
  AOI22_X1 U17664 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14251) );
  AOI22_X1 U17665 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U17666 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n14249) );
  NAND4_X1 U17667 ( .A1(n14252), .A2(n14251), .A3(n14250), .A4(n14249), .ZN(
        n14253) );
  AOI211_X1 U17668 ( .C1(n9641), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n14254), .B(n14253), .ZN(n14255) );
  OAI211_X1 U17669 ( .C1(n9652), .C2(n17361), .A(n14256), .B(n14255), .ZN(
        n17608) );
  NAND2_X1 U17670 ( .A1(n17609), .A2(n17608), .ZN(n17607) );
  NOR2_X1 U17671 ( .A1(n14257), .A2(n17607), .ZN(n17300) );
  AOI21_X1 U17672 ( .B1(n14257), .B2(n17607), .A(n17300), .ZN(n17604) );
  AOI22_X1 U17673 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17303), .B1(n17583), 
        .B2(n17604), .ZN(n14260) );
  INV_X1 U17674 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14258) );
  INV_X1 U17675 ( .A(n17308), .ZN(n17311) );
  NAND3_X1 U17676 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14258), .A3(n17311), 
        .ZN(n14259) );
  NAND2_X1 U17677 ( .A1(n14260), .A2(n14259), .ZN(P3_U2675) );
  NOR2_X1 U17678 ( .A1(n14267), .A2(n14263), .ZN(n14264) );
  NAND2_X1 U17679 ( .A1(n14987), .A2(n14264), .ZN(n14957) );
  AOI22_X1 U17680 ( .A1(n14969), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14979), .ZN(n14270) );
  NOR3_X4 U17681 ( .A1(n14979), .A2(n14347), .A3(n14265), .ZN(n14972) );
  INV_X1 U17682 ( .A(DATAI_12_), .ZN(n21077) );
  NAND2_X1 U17683 ( .A1(n14923), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14266) );
  OAI21_X1 U17684 ( .B1(n14923), .B2(n21077), .A(n14266), .ZN(n20421) );
  NOR3_X1 U17685 ( .A1(n14979), .A2(n14923), .A3(n14267), .ZN(n14268) );
  AOI22_X1 U17686 ( .A1(n14972), .A2(n20421), .B1(n14970), .B2(DATAI_28_), 
        .ZN(n14269) );
  OAI211_X1 U17687 ( .C1(n15003), .C2(n14982), .A(n14270), .B(n14269), .ZN(
        P1_U2876) );
  MUX2_X1 U17688 ( .A(n14291), .B(n14318), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n14272) );
  NAND2_X1 U17689 ( .A1(n9653), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14271) );
  AND2_X1 U17690 ( .A1(n14272), .A2(n14271), .ZN(n14907) );
  NOR2_X1 U17691 ( .A1(n14656), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14273) );
  NOR2_X1 U17692 ( .A1(n14274), .A2(n14273), .ZN(n14855) );
  NAND2_X1 U17693 ( .A1(n14910), .A2(n14855), .ZN(n14900) );
  NAND2_X1 U17694 ( .A1(n14318), .A2(n16357), .ZN(n14275) );
  OAI211_X1 U17695 ( .C1(n9653), .C2(P1_EBX_REG_13__SCAN_IN), .A(n14275), .B(
        n14291), .ZN(n14277) );
  INV_X1 U17696 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n16217) );
  NAND2_X1 U17697 ( .A1(n14322), .A2(n16217), .ZN(n14276) );
  AND2_X1 U17698 ( .A1(n14277), .A2(n14276), .ZN(n14899) );
  INV_X1 U17699 ( .A(n14278), .ZN(n14279) );
  OAI21_X1 U17700 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14656), .A(
        n14279), .ZN(n14840) );
  NAND2_X1 U17701 ( .A1(n14318), .A2(n14280), .ZN(n14281) );
  OAI211_X1 U17702 ( .C1(n9653), .C2(P1_EBX_REG_15__SCAN_IN), .A(n14281), .B(
        n14291), .ZN(n14284) );
  INV_X1 U17703 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14282) );
  NAND2_X1 U17704 ( .A1(n14322), .A2(n14282), .ZN(n14283) );
  NAND2_X1 U17705 ( .A1(n14284), .A2(n14283), .ZN(n14826) );
  INV_X1 U17706 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14285) );
  NAND2_X1 U17707 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14286) );
  OAI211_X1 U17708 ( .C1(n9653), .C2(P1_EBX_REG_16__SCAN_IN), .A(n14318), .B(
        n14286), .ZN(n14287) );
  AND2_X1 U17709 ( .A1(n14288), .A2(n14287), .ZN(n14814) );
  NOR2_X1 U17710 ( .A1(n14656), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14289) );
  NOR2_X1 U17711 ( .A1(n14290), .A2(n14289), .ZN(n14797) );
  MUX2_X1 U17712 ( .A(n14291), .B(n14318), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14293) );
  NAND2_X1 U17713 ( .A1(n9653), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14292) );
  NAND2_X1 U17714 ( .A1(n14293), .A2(n14292), .ZN(n14889) );
  NAND2_X1 U17715 ( .A1(n14797), .A2(n14889), .ZN(n14294) );
  NAND2_X1 U17716 ( .A1(n14318), .A2(n15220), .ZN(n14295) );
  OAI211_X1 U17717 ( .C1(n9653), .C2(P1_EBX_REG_19__SCAN_IN), .A(n14295), .B(
        n14291), .ZN(n14297) );
  INV_X1 U17718 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14880) );
  NAND2_X1 U17719 ( .A1(n14322), .A2(n14880), .ZN(n14296) );
  AND2_X1 U17720 ( .A1(n14297), .A2(n14296), .ZN(n14785) );
  NOR2_X2 U17721 ( .A1(n9707), .A2(n14785), .ZN(n14786) );
  INV_X1 U17722 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14877) );
  NAND2_X1 U17723 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14298) );
  OAI211_X1 U17724 ( .C1(n9653), .C2(P1_EBX_REG_20__SCAN_IN), .A(n14318), .B(
        n14298), .ZN(n14299) );
  AND2_X1 U17725 ( .A1(n14300), .A2(n14299), .ZN(n14774) );
  NAND2_X1 U17726 ( .A1(n14318), .A2(n14301), .ZN(n14302) );
  OAI211_X1 U17727 ( .C1(n9653), .C2(P1_EBX_REG_21__SCAN_IN), .A(n14302), .B(
        n14291), .ZN(n14304) );
  INV_X1 U17728 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n16248) );
  NAND2_X1 U17729 ( .A1(n14322), .A2(n16248), .ZN(n14303) );
  AND2_X1 U17730 ( .A1(n14304), .A2(n14303), .ZN(n16170) );
  INV_X1 U17731 ( .A(n14305), .ZN(n14306) );
  OAI21_X1 U17732 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n14656), .A(
        n14306), .ZN(n14761) );
  MUX2_X1 U17733 ( .A(n14291), .B(n14318), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n14308) );
  NAND2_X1 U17734 ( .A1(n9653), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14307) );
  AND2_X1 U17735 ( .A1(n14308), .A2(n14307), .ZN(n14750) );
  NOR2_X2 U17736 ( .A1(n14762), .A2(n14750), .ZN(n14749) );
  NOR2_X1 U17737 ( .A1(n14656), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14309) );
  NOR2_X1 U17738 ( .A1(n14310), .A2(n14309), .ZN(n14737) );
  NAND2_X1 U17739 ( .A1(n14749), .A2(n14737), .ZN(n14739) );
  NAND2_X1 U17740 ( .A1(n14318), .A2(n15205), .ZN(n14311) );
  OAI211_X1 U17741 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n9653), .A(n14311), .B(
        n14291), .ZN(n14314) );
  INV_X1 U17742 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U17743 ( .A1(n14322), .A2(n14312), .ZN(n14313) );
  AND2_X1 U17744 ( .A1(n14314), .A2(n14313), .ZN(n14723) );
  INV_X1 U17745 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14871) );
  NAND2_X1 U17746 ( .A1(n14291), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14315) );
  OAI211_X1 U17747 ( .C1(n9653), .C2(P1_EBX_REG_26__SCAN_IN), .A(n14318), .B(
        n14315), .ZN(n14316) );
  NAND2_X1 U17748 ( .A1(n14317), .A2(n14316), .ZN(n14709) );
  NAND2_X1 U17749 ( .A1(n14318), .A2(n15190), .ZN(n14319) );
  OAI211_X1 U17750 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n9653), .A(n14319), .B(
        n14291), .ZN(n14321) );
  INV_X1 U17751 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14870) );
  NAND2_X1 U17752 ( .A1(n14322), .A2(n14870), .ZN(n14320) );
  NAND2_X1 U17753 ( .A1(n14321), .A2(n14320), .ZN(n14696) );
  NOR2_X1 U17754 ( .A1(n14656), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14323) );
  NOR2_X1 U17755 ( .A1(n14324), .A2(n14323), .ZN(n14325) );
  OR2_X1 U17756 ( .A1(n14698), .A2(n14325), .ZN(n14326) );
  NAND2_X1 U17757 ( .A1(n14683), .A2(n14326), .ZN(n15179) );
  INV_X1 U17758 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14334) );
  OAI222_X1 U17759 ( .A1(n15179), .A2(n14916), .B1(n14334), .B2(n20387), .C1(
        n15003), .C2(n14884), .ZN(P1_U2844) );
  INV_X1 U17760 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21079) );
  AND2_X1 U17761 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14337) );
  INV_X1 U17762 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20983) );
  NAND2_X1 U17763 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14330) );
  NAND2_X1 U17764 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14859) );
  INV_X1 U17765 ( .A(n14859), .ZN(n14329) );
  NAND2_X1 U17766 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14328) );
  NOR2_X1 U17767 ( .A1(n14328), .A2(n14327), .ZN(n14858) );
  NAND4_X1 U17768 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n14329), .A4(n14858), .ZN(n14811) );
  NOR3_X1 U17769 ( .A1(n20983), .A2(n14330), .A3(n14811), .ZN(n14784) );
  AND4_X1 U17770 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .A4(n14784), .ZN(n14759) );
  AND2_X1 U17771 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n14759), .ZN(n14331) );
  AND2_X1 U17772 ( .A1(n14337), .A2(n14331), .ZN(n14725) );
  NAND4_X1 U17773 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_24__SCAN_IN), .A4(n14725), .ZN(n14700) );
  NOR2_X1 U17774 ( .A1(n21079), .A2(n14700), .ZN(n14332) );
  AOI21_X1 U17775 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14332), .A(n20307), 
        .ZN(n14688) );
  AOI22_X1 U17776 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20348), .B1(
        n20349), .B2(n15006), .ZN(n14333) );
  OAI21_X1 U17777 ( .B1(n20325), .B2(n14334), .A(n14333), .ZN(n14336) );
  NOR2_X1 U17778 ( .A1(n15179), .A2(n20320), .ZN(n14335) );
  AOI211_X1 U17779 ( .C1(n14688), .C2(P1_REIP_REG_28__SCAN_IN), .A(n14336), 
        .B(n14335), .ZN(n14340) );
  INV_X1 U17780 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20979) );
  NAND3_X1 U17781 ( .A1(n16235), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n16234) );
  NOR2_X2 U17782 ( .A1(n16234), .A2(n14859), .ZN(n16221) );
  NAND3_X1 U17783 ( .A1(n14804), .A2(P1_REIP_REG_19__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n14773) );
  INV_X1 U17784 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20990) );
  NAND2_X1 U17785 ( .A1(n16207), .A2(n14337), .ZN(n14753) );
  INV_X1 U17786 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20995) );
  NAND2_X1 U17787 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14338) );
  NOR2_X1 U17788 ( .A1(n14742), .A2(n14338), .ZN(n14717) );
  NAND3_X1 U17789 ( .A1(n14705), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n21079), 
        .ZN(n14339) );
  OAI211_X1 U17790 ( .C1(n15003), .C2(n14864), .A(n14340), .B(n14339), .ZN(
        P1_U2812) );
  OAI21_X1 U17791 ( .B1(n13479), .B2(n14342), .A(n14341), .ZN(n19476) );
  MUX2_X1 U17792 ( .A(n14343), .B(n19558), .S(n15449), .Z(n14344) );
  OAI21_X1 U17793 ( .B1(n19476), .B2(n15479), .A(n14344), .ZN(P2_U2883) );
  NOR2_X1 U17794 ( .A1(n11339), .A2(n15448), .ZN(n14345) );
  AOI21_X1 U17795 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n15448), .A(n14345), .ZN(
        n14346) );
  OAI21_X1 U17796 ( .B1(n20204), .B2(n15479), .A(n14346), .ZN(P2_U2884) );
  NAND2_X1 U17797 ( .A1(n10293), .A2(n14651), .ZN(n14349) );
  AOI22_X1 U17798 ( .A1(n14970), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14979), .ZN(n14348) );
  OAI211_X1 U17799 ( .C1(n14957), .C2(n19612), .A(n14349), .B(n14348), .ZN(
        P1_U2873) );
  AOI22_X1 U17800 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10779), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14353) );
  AOI22_X1 U17801 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14352) );
  AOI22_X1 U17802 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14351) );
  AOI22_X1 U17803 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14350) );
  NAND4_X1 U17804 ( .A1(n14353), .A2(n14352), .A3(n14351), .A4(n14350), .ZN(
        n14362) );
  AOI22_X1 U17805 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U17806 ( .A1(n9643), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14359) );
  INV_X1 U17807 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14355) );
  NAND2_X1 U17808 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14437), .ZN(
        n14354) );
  OAI21_X1 U17809 ( .B1(n14440), .B2(n14355), .A(n14354), .ZN(n14356) );
  AOI21_X1 U17810 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n14356), .ZN(n14358) );
  NAND2_X1 U17811 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n14357) );
  NAND4_X1 U17812 ( .A1(n14360), .A2(n14359), .A3(n14358), .A4(n14357), .ZN(
        n14361) );
  OR2_X1 U17813 ( .A1(n14362), .A2(n14361), .ZN(n15467) );
  AND2_X2 U17814 ( .A1(n14363), .A2(n15467), .ZN(n15460) );
  AOI22_X1 U17815 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10779), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14367) );
  AOI22_X1 U17816 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U17817 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14365) );
  AOI22_X1 U17818 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14364) );
  NAND4_X1 U17819 ( .A1(n14367), .A2(n14366), .A3(n14365), .A4(n14364), .ZN(
        n14376) );
  AOI22_X1 U17820 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14374) );
  AOI22_X1 U17821 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14373) );
  NAND2_X1 U17822 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14437), .ZN(
        n14368) );
  OAI21_X1 U17823 ( .B1(n14440), .B2(n14369), .A(n14368), .ZN(n14370) );
  AOI21_X1 U17824 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n14370), .ZN(n14372) );
  NAND2_X1 U17825 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n14371) );
  NAND4_X1 U17826 ( .A1(n14374), .A2(n14373), .A3(n14372), .A4(n14371), .ZN(
        n14375) );
  OR2_X1 U17827 ( .A1(n14376), .A2(n14375), .ZN(n15461) );
  AOI22_X1 U17828 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10779), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14380) );
  AOI22_X1 U17829 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14379) );
  AOI22_X1 U17830 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14378) );
  AOI22_X1 U17831 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n14448), .B1(
        n10701), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14377) );
  NAND4_X1 U17832 ( .A1(n14380), .A2(n14379), .A3(n14378), .A4(n14377), .ZN(
        n14389) );
  AOI22_X1 U17833 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U17834 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14386) );
  INV_X1 U17835 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14382) );
  NAND2_X1 U17836 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14437), .ZN(
        n14381) );
  OAI21_X1 U17837 ( .B1(n14440), .B2(n14382), .A(n14381), .ZN(n14383) );
  AOI21_X1 U17838 ( .B1(n14406), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n14383), .ZN(n14385) );
  NAND2_X1 U17839 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n14384) );
  NAND4_X1 U17840 ( .A1(n14387), .A2(n14386), .A3(n14385), .A4(n14384), .ZN(
        n14388) );
  NOR2_X1 U17841 ( .A1(n14389), .A2(n14388), .ZN(n15456) );
  INV_X1 U17842 ( .A(n9642), .ZN(n14393) );
  AOI22_X1 U17843 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14392) );
  NAND2_X1 U17844 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14391) );
  OAI211_X1 U17845 ( .C1(n13451), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        n14405) );
  AOI22_X1 U17846 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10779), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U17847 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14396) );
  AOI22_X1 U17848 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14395) );
  AOI22_X1 U17849 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14394) );
  NAND4_X1 U17850 ( .A1(n14397), .A2(n14396), .A3(n14395), .A4(n14394), .ZN(
        n14404) );
  INV_X1 U17851 ( .A(n14398), .ZN(n14402) );
  AOI22_X1 U17852 ( .A1(n14407), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__5__SCAN_IN), .B2(n14437), .ZN(n14400) );
  NAND2_X1 U17853 ( .A1(n14406), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14399) );
  OAI211_X1 U17854 ( .C1(n14402), .C2(n14401), .A(n14400), .B(n14399), .ZN(
        n14403) );
  NOR3_X1 U17855 ( .A1(n14405), .A2(n14404), .A3(n14403), .ZN(n15446) );
  INV_X1 U17856 ( .A(n14406), .ZN(n14410) );
  AOI22_X1 U17857 ( .A1(n14407), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n14437), .ZN(n14408) );
  OAI21_X1 U17858 ( .B1(n14410), .B2(n14409), .A(n14408), .ZN(n14411) );
  AOI21_X1 U17859 ( .B1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n14398), .A(
        n14411), .ZN(n14419) );
  AOI22_X1 U17860 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U17861 ( .A1(n9642), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U17862 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10779), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14415) );
  AOI22_X1 U17863 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14414) );
  AOI22_X1 U17864 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U17865 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14412) );
  AND4_X1 U17866 ( .A1(n14415), .A2(n14414), .A3(n14413), .A4(n14412), .ZN(
        n14416) );
  NAND4_X1 U17867 ( .A1(n14419), .A2(n14418), .A3(n14417), .A4(n14416), .ZN(
        n15443) );
  NAND2_X1 U17868 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14423) );
  NAND2_X1 U17869 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14422) );
  NAND2_X1 U17870 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14421) );
  NAND2_X1 U17871 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n14420) );
  AND4_X1 U17872 ( .A1(n14423), .A2(n14422), .A3(n14421), .A4(n14420), .ZN(
        n14426) );
  AOI22_X1 U17873 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14425) );
  AOI22_X1 U17874 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9671), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14424) );
  XNOR2_X1 U17875 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14591) );
  NAND4_X1 U17876 ( .A1(n14426), .A2(n14425), .A3(n14424), .A4(n14591), .ZN(
        n14435) );
  NAND2_X1 U17877 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n14430) );
  NAND2_X1 U17878 ( .A1(n14595), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14429) );
  NAND2_X1 U17879 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n14428) );
  NAND2_X1 U17880 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n14427) );
  AND4_X1 U17881 ( .A1(n14430), .A2(n14429), .A3(n14428), .A4(n14427), .ZN(
        n14433) );
  INV_X1 U17882 ( .A(n14591), .ZN(n14598) );
  AOI22_X1 U17883 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U17884 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14431) );
  NAND4_X1 U17885 ( .A1(n14433), .A2(n14598), .A3(n14432), .A4(n14431), .ZN(
        n14434) );
  NAND2_X1 U17886 ( .A1(n14435), .A2(n14434), .ZN(n14481) );
  NOR2_X1 U17887 ( .A1(n10493), .A2(n14481), .ZN(n14455) );
  AOI22_X1 U17888 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n9640), .B1(
        n14406), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14445) );
  INV_X1 U17889 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14439) );
  NAND2_X1 U17890 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14437), .ZN(
        n14438) );
  OAI21_X1 U17891 ( .B1(n14440), .B2(n14439), .A(n14438), .ZN(n14441) );
  AOI21_X1 U17892 ( .B1(n9642), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(n14441), .ZN(n14444) );
  AOI22_X1 U17893 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10779), .B1(
        n10744), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14443) );
  NAND2_X1 U17894 ( .A1(n14398), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n14442) );
  NAND4_X1 U17895 ( .A1(n14445), .A2(n14444), .A3(n14443), .A4(n14442), .ZN(
        n14454) );
  AOI22_X1 U17896 ( .A1(n10766), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14452) );
  AOI22_X1 U17897 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10743), .B1(
        n14446), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U17898 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10720), .B1(
        n10700), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14450) );
  AOI22_X1 U17899 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10701), .B1(
        n14448), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14449) );
  NAND4_X1 U17900 ( .A1(n14452), .A2(n14451), .A3(n14450), .A4(n14449), .ZN(
        n14453) );
  NOR2_X1 U17901 ( .A1(n14454), .A2(n14453), .ZN(n14476) );
  XNOR2_X1 U17902 ( .A(n14455), .B(n14476), .ZN(n14483) );
  INV_X1 U17903 ( .A(n14483), .ZN(n14456) );
  INV_X1 U17904 ( .A(n14481), .ZN(n14477) );
  NAND2_X1 U17905 ( .A1(n10493), .A2(n14477), .ZN(n15438) );
  INV_X1 U17906 ( .A(n14457), .ZN(n14458) );
  AOI22_X1 U17907 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U17908 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n14462) );
  NAND2_X1 U17909 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14461) );
  NAND2_X1 U17910 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14460) );
  NAND2_X1 U17911 ( .A1(n9671), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14459) );
  AND4_X1 U17912 ( .A1(n14462), .A2(n14461), .A3(n14460), .A4(n14459), .ZN(
        n14464) );
  AOI22_X1 U17913 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14463) );
  NAND4_X1 U17914 ( .A1(n14465), .A2(n14464), .A3(n14463), .A4(n14591), .ZN(
        n14475) );
  AOI22_X1 U17915 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14473) );
  NAND2_X1 U17916 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n14470) );
  NAND2_X1 U17917 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14469) );
  NAND2_X1 U17918 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14468) );
  NAND2_X1 U17919 ( .A1(n9671), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14467) );
  AND4_X1 U17920 ( .A1(n14470), .A2(n14469), .A3(n14468), .A4(n14467), .ZN(
        n14472) );
  AOI22_X1 U17921 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14471) );
  NAND4_X1 U17922 ( .A1(n14473), .A2(n14472), .A3(n14471), .A4(n14598), .ZN(
        n14474) );
  NAND2_X1 U17923 ( .A1(n14475), .A2(n14474), .ZN(n14484) );
  INV_X1 U17924 ( .A(n14476), .ZN(n14478) );
  NAND2_X1 U17925 ( .A1(n14478), .A2(n14477), .ZN(n14485) );
  XOR2_X1 U17926 ( .A(n14484), .B(n14485), .Z(n14479) );
  NAND2_X1 U17927 ( .A1(n14479), .A2(n14549), .ZN(n15428) );
  INV_X1 U17928 ( .A(n14484), .ZN(n14480) );
  NAND2_X1 U17929 ( .A1(n10493), .A2(n14480), .ZN(n15430) );
  NOR2_X1 U17930 ( .A1(n15430), .A2(n14481), .ZN(n14482) );
  NOR2_X1 U17931 ( .A1(n14485), .A2(n14484), .ZN(n14502) );
  AOI22_X1 U17932 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14492) );
  NAND2_X1 U17933 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14489) );
  NAND2_X1 U17934 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14488) );
  NAND2_X1 U17935 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14487) );
  NAND2_X1 U17936 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14486) );
  AND4_X1 U17937 ( .A1(n14489), .A2(n14488), .A3(n14487), .A4(n14486), .ZN(
        n14491) );
  AOI22_X1 U17938 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14490) );
  NAND4_X1 U17939 ( .A1(n14492), .A2(n14491), .A3(n14490), .A4(n14591), .ZN(
        n14501) );
  AOI22_X1 U17940 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14499) );
  NAND2_X1 U17941 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n14496) );
  NAND2_X1 U17942 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14495) );
  NAND2_X1 U17943 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14494) );
  NAND2_X1 U17944 ( .A1(n9671), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14493) );
  AND4_X1 U17945 ( .A1(n14496), .A2(n14495), .A3(n14494), .A4(n14493), .ZN(
        n14498) );
  AOI22_X1 U17946 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14497) );
  NAND4_X1 U17947 ( .A1(n14499), .A2(n14498), .A3(n14497), .A4(n14598), .ZN(
        n14500) );
  AND2_X1 U17948 ( .A1(n14501), .A2(n14500), .ZN(n14503) );
  NAND2_X1 U17949 ( .A1(n14502), .A2(n14503), .ZN(n14546) );
  OAI211_X1 U17950 ( .C1(n14502), .C2(n14503), .A(n14546), .B(n14549), .ZN(
        n14506) );
  INV_X1 U17951 ( .A(n14503), .ZN(n14504) );
  NOR2_X1 U17952 ( .A1(n16700), .A2(n14504), .ZN(n15424) );
  AOI22_X1 U17953 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14515) );
  NAND2_X1 U17954 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n14512) );
  NAND2_X1 U17955 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14511) );
  NAND2_X1 U17956 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14510) );
  NAND2_X1 U17957 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14509) );
  AND4_X1 U17958 ( .A1(n14512), .A2(n14511), .A3(n14510), .A4(n14509), .ZN(
        n14514) );
  AOI22_X1 U17959 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14513) );
  NAND4_X1 U17960 ( .A1(n14515), .A2(n14514), .A3(n14513), .A4(n14591), .ZN(
        n14524) );
  AOI22_X1 U17961 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14522) );
  NAND2_X1 U17962 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n14519) );
  NAND2_X1 U17963 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14518) );
  NAND2_X1 U17964 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14517) );
  NAND2_X1 U17965 ( .A1(n9671), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14516) );
  AND4_X1 U17966 ( .A1(n14519), .A2(n14518), .A3(n14517), .A4(n14516), .ZN(
        n14521) );
  AOI22_X1 U17967 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14520) );
  NAND4_X1 U17968 ( .A1(n14522), .A2(n14521), .A3(n14520), .A4(n14598), .ZN(
        n14523) );
  AND2_X1 U17969 ( .A1(n14524), .A2(n14523), .ZN(n14544) );
  XNOR2_X1 U17970 ( .A(n14546), .B(n14544), .ZN(n14525) );
  NAND2_X1 U17971 ( .A1(n10493), .A2(n14544), .ZN(n15419) );
  AOI22_X1 U17972 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U17973 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14531) );
  NAND2_X1 U17974 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14530) );
  NAND2_X1 U17975 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14529) );
  NAND2_X1 U17976 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14528) );
  AND4_X1 U17977 ( .A1(n14531), .A2(n14530), .A3(n14529), .A4(n14528), .ZN(
        n14533) );
  AOI22_X1 U17978 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14532) );
  NAND4_X1 U17979 ( .A1(n14534), .A2(n14533), .A3(n14532), .A4(n14591), .ZN(
        n14543) );
  AOI22_X1 U17980 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14541) );
  NAND2_X1 U17981 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n14538) );
  NAND2_X1 U17982 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14537) );
  NAND2_X1 U17983 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14536) );
  NAND2_X1 U17984 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14535) );
  AND4_X1 U17985 ( .A1(n14538), .A2(n14537), .A3(n14536), .A4(n14535), .ZN(
        n14540) );
  AOI22_X1 U17986 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14539) );
  NAND4_X1 U17987 ( .A1(n14541), .A2(n14540), .A3(n14539), .A4(n14598), .ZN(
        n14542) );
  NAND2_X1 U17988 ( .A1(n14543), .A2(n14542), .ZN(n14547) );
  INV_X1 U17989 ( .A(n14547), .ZN(n14554) );
  INV_X1 U17990 ( .A(n14544), .ZN(n14545) );
  OR2_X1 U17991 ( .A1(n14546), .A2(n14545), .ZN(n14548) );
  INV_X1 U17992 ( .A(n14548), .ZN(n14550) );
  OR2_X1 U17993 ( .A1(n14548), .A2(n14547), .ZN(n15395) );
  OAI211_X1 U17994 ( .C1(n14554), .C2(n14550), .A(n15395), .B(n14549), .ZN(
        n14551) );
  OR2_X2 U17995 ( .A1(n14552), .A2(n14551), .ZN(n15396) );
  NAND2_X1 U17996 ( .A1(n10493), .A2(n14554), .ZN(n15409) );
  AOI22_X1 U17997 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14561) );
  NAND2_X1 U17998 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14558) );
  NAND2_X1 U17999 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14557) );
  NAND2_X1 U18000 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14556) );
  NAND2_X1 U18001 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14555) );
  AND4_X1 U18002 ( .A1(n14558), .A2(n14557), .A3(n14556), .A4(n14555), .ZN(
        n14560) );
  AOI22_X1 U18003 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14559) );
  NAND4_X1 U18004 ( .A1(n14561), .A2(n14560), .A3(n14559), .A4(n14591), .ZN(
        n14570) );
  AOI22_X1 U18005 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14568) );
  NAND2_X1 U18006 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n14565) );
  NAND2_X1 U18007 ( .A1(n14600), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14564) );
  NAND2_X1 U18008 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14563) );
  NAND2_X1 U18009 ( .A1(n9671), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14562) );
  AND4_X1 U18010 ( .A1(n14565), .A2(n14564), .A3(n14563), .A4(n14562), .ZN(
        n14567) );
  AOI22_X1 U18011 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14566) );
  NAND4_X1 U18012 ( .A1(n14568), .A2(n14567), .A3(n14566), .A4(n14598), .ZN(
        n14569) );
  AND2_X1 U18013 ( .A1(n14570), .A2(n14569), .ZN(n15397) );
  NAND2_X1 U18014 ( .A1(n16700), .A2(n15397), .ZN(n14571) );
  NOR2_X1 U18015 ( .A1(n15395), .A2(n14571), .ZN(n14586) );
  AOI22_X1 U18016 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14573) );
  AOI22_X1 U18017 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14572) );
  AND2_X1 U18018 ( .A1(n14573), .A2(n14572), .ZN(n14576) );
  AOI22_X1 U18019 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14577), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14575) );
  AOI22_X1 U18020 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14574) );
  NAND4_X1 U18021 ( .A1(n14576), .A2(n14575), .A3(n14574), .A4(n14591), .ZN(
        n14584) );
  AOI22_X1 U18022 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14579) );
  AOI22_X1 U18023 ( .A1(n14577), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14578) );
  AND2_X1 U18024 ( .A1(n14579), .A2(n14578), .ZN(n14582) );
  AOI22_X1 U18025 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14581) );
  AOI22_X1 U18026 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14580) );
  NAND4_X1 U18027 ( .A1(n14582), .A2(n14598), .A3(n14581), .A4(n14580), .ZN(
        n14583) );
  AND2_X1 U18028 ( .A1(n14584), .A2(n14583), .ZN(n14585) );
  NAND2_X1 U18029 ( .A1(n14586), .A2(n14585), .ZN(n14587) );
  OAI21_X1 U18030 ( .B1(n14586), .B2(n14585), .A(n14587), .ZN(n15392) );
  INV_X1 U18031 ( .A(n14587), .ZN(n14588) );
  AOI22_X1 U18032 ( .A1(n9660), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14590) );
  AOI22_X1 U18033 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14589) );
  NAND2_X1 U18034 ( .A1(n14590), .A2(n14589), .ZN(n14608) );
  AOI22_X1 U18035 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14577), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14593) );
  AOI22_X1 U18036 ( .A1(n14594), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14595), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14592) );
  NAND3_X1 U18037 ( .A1(n14593), .A2(n14592), .A3(n14591), .ZN(n14607) );
  AOI22_X1 U18038 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14594), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14599) );
  AOI22_X1 U18039 ( .A1(n14596), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9674), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14597) );
  NAND3_X1 U18040 ( .A1(n14599), .A2(n14598), .A3(n14597), .ZN(n14606) );
  AOI22_X1 U18041 ( .A1(n9661), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14600), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14604) );
  AOI22_X1 U18042 ( .A1(n14602), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9671), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14603) );
  NAND2_X1 U18043 ( .A1(n14604), .A2(n14603), .ZN(n14605) );
  OAI22_X1 U18044 ( .A1(n14608), .A2(n14607), .B1(n14606), .B2(n14605), .ZN(
        n14609) );
  XNOR2_X1 U18045 ( .A(n14610), .B(n14609), .ZN(n14622) );
  INV_X1 U18046 ( .A(n15768), .ZN(n14617) );
  NAND2_X1 U18047 ( .A1(n14611), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14613) );
  INV_X1 U18048 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16788) );
  OR2_X1 U18049 ( .A1(n14611), .A2(n16788), .ZN(n14612) );
  NAND2_X1 U18050 ( .A1(n14613), .A2(n14612), .ZN(n19546) );
  INV_X1 U18051 ( .A(n19546), .ZN(n14615) );
  INV_X1 U18052 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14614) );
  OAI22_X1 U18053 ( .A1(n15558), .A2(n14615), .B1(n19466), .B2(n14614), .ZN(
        n14616) );
  AOI21_X1 U18054 ( .B1(n14617), .B2(n19495), .A(n14616), .ZN(n14619) );
  AOI22_X1 U18055 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19436), .B1(n19438), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n14618) );
  OAI211_X1 U18056 ( .C1(n14622), .C2(n19490), .A(n14619), .B(n14618), .ZN(
        P2_U2889) );
  NAND2_X1 U18057 ( .A1(n15766), .A2(n15449), .ZN(n14621) );
  NAND2_X1 U18058 ( .A1(n15448), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14620) );
  OAI211_X1 U18059 ( .C1(n14622), .C2(n15479), .A(n14621), .B(n14620), .ZN(
        P2_U2857) );
  AOI21_X1 U18060 ( .B1(n14623), .B2(n14624), .A(n15944), .ZN(n14640) );
  INV_X1 U18061 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14628) );
  OR2_X1 U18062 ( .A1(n19333), .A2(n10535), .ZN(n14643) );
  OAI21_X1 U18063 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14625), .A(
        n14624), .ZN(n14626) );
  OR2_X1 U18064 ( .A1(n15940), .A2(n14626), .ZN(n14627) );
  OAI211_X1 U18065 ( .C1(n14629), .C2(n14628), .A(n14643), .B(n14627), .ZN(
        n14630) );
  INV_X1 U18066 ( .A(n14630), .ZN(n14635) );
  INV_X1 U18067 ( .A(n14631), .ZN(n14632) );
  XNOR2_X1 U18068 ( .A(n14633), .B(n14632), .ZN(n14646) );
  NAND2_X1 U18069 ( .A1(n14646), .A2(n16646), .ZN(n14634) );
  OAI211_X1 U18070 ( .C1(n20213), .C2(n16624), .A(n14635), .B(n14634), .ZN(
        n14639) );
  NAND2_X1 U18071 ( .A1(n14637), .A2(n14636), .ZN(n14647) );
  AND3_X1 U18072 ( .A1(n14648), .A2(n16600), .A3(n14647), .ZN(n14638) );
  NOR3_X1 U18073 ( .A1(n14640), .A2(n14639), .A3(n14638), .ZN(n14641) );
  OAI21_X1 U18074 ( .B1(n9675), .B2(n16629), .A(n14641), .ZN(P2_U3044) );
  NAND2_X1 U18075 ( .A1(n19551), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14642) );
  OAI211_X1 U18076 ( .C1(n19564), .C2(n14644), .A(n14643), .B(n14642), .ZN(
        n14645) );
  AOI21_X1 U18077 ( .B1(n19554), .B2(n14646), .A(n14645), .ZN(n14650) );
  NAND3_X1 U18078 ( .A1(n14648), .A2(n19552), .A3(n14647), .ZN(n14649) );
  OAI211_X1 U18079 ( .C1(n19559), .C2(n9675), .A(n14650), .B(n14649), .ZN(
        P2_U3012) );
  INV_X1 U18080 ( .A(n14651), .ZN(n14666) );
  OR2_X1 U18081 ( .A1(n14656), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14654) );
  INV_X1 U18082 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14869) );
  NAND2_X1 U18083 ( .A1(n14652), .A2(n14869), .ZN(n14653) );
  AND2_X1 U18084 ( .A1(n14654), .A2(n14653), .ZN(n14668) );
  NOR2_X1 U18085 ( .A1(n14291), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14655) );
  AOI21_X1 U18086 ( .B1(n14668), .B2(n14291), .A(n14655), .ZN(n14682) );
  NOR2_X1 U18087 ( .A1(n14685), .A2(n14291), .ZN(n14667) );
  AOI22_X1 U18088 ( .A1(n14656), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n9653), .ZN(n14659) );
  NOR2_X1 U18089 ( .A1(n14667), .A2(n14659), .ZN(n14660) );
  INV_X1 U18090 ( .A(n14685), .ZN(n14657) );
  AOI22_X1 U18091 ( .A1(n14656), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n9653), .ZN(n14669) );
  NOR2_X1 U18092 ( .A1(n14657), .A2(n14669), .ZN(n14658) );
  MUX2_X1 U18093 ( .A(n14660), .B(n14659), .S(n14658), .Z(n15140) );
  NAND2_X1 U18094 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14662) );
  AOI21_X1 U18095 ( .B1(n14662), .B2(n14812), .A(n14688), .ZN(n14674) );
  AOI22_X1 U18096 ( .A1(n20360), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20348), .ZN(n14661) );
  OAI21_X1 U18097 ( .B1(n14674), .B2(n21165), .A(n14661), .ZN(n14664) );
  NOR3_X1 U18098 ( .A1(n14673), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14662), 
        .ZN(n14663) );
  AOI211_X1 U18099 ( .C1(n20362), .C2(n15140), .A(n14664), .B(n14663), .ZN(
        n14665) );
  OAI21_X1 U18100 ( .B1(n14666), .B2(n14864), .A(n14665), .ZN(P1_U2809) );
  AOI21_X1 U18101 ( .B1(n10129), .B2(n14668), .A(n14667), .ZN(n14670) );
  XNOR2_X1 U18102 ( .A(n14670), .B(n14669), .ZN(n14867) );
  INV_X1 U18103 ( .A(n14867), .ZN(n15161) );
  INV_X1 U18104 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14868) );
  AOI22_X1 U18105 ( .A1(n14671), .A2(n20349), .B1(n20348), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14672) );
  OAI21_X1 U18106 ( .B1(n20325), .B2(n14868), .A(n14672), .ZN(n14677) );
  NOR2_X1 U18107 ( .A1(n14675), .A2(n14674), .ZN(n14676) );
  AOI211_X1 U18108 ( .C1(n15161), .C2(n20362), .A(n14677), .B(n14676), .ZN(
        n14678) );
  INV_X1 U18109 ( .A(n14996), .ZN(n14926) );
  INV_X1 U18110 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21094) );
  AND2_X1 U18111 ( .A1(n14683), .A2(n14682), .ZN(n14684) );
  OR2_X1 U18112 ( .A1(n14685), .A2(n14684), .ZN(n15173) );
  OAI22_X1 U18113 ( .A1(n14686), .A2(n20365), .B1(n20375), .B2(n14994), .ZN(
        n14687) );
  AOI21_X1 U18114 ( .B1(n20360), .B2(P1_EBX_REG_29__SCAN_IN), .A(n14687), .ZN(
        n14690) );
  NAND2_X1 U18115 ( .A1(n14688), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14689) );
  OAI211_X1 U18116 ( .C1(n15173), .C2(n20320), .A(n14690), .B(n14689), .ZN(
        n14691) );
  AOI21_X1 U18117 ( .B1(n14692), .B2(n21094), .A(n14691), .ZN(n14693) );
  OAI21_X1 U18118 ( .B1(n14926), .B2(n14864), .A(n14693), .ZN(P1_U2811) );
  AOI21_X1 U18119 ( .B1(n14695), .B2(n14707), .A(n14694), .ZN(n15016) );
  INV_X1 U18120 ( .A(n15016), .ZN(n14929) );
  INV_X1 U18121 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21163) );
  NOR2_X1 U18122 ( .A1(n14710), .A2(n14696), .ZN(n14697) );
  OR2_X1 U18123 ( .A1(n14698), .A2(n14697), .ZN(n15186) );
  OAI22_X1 U18124 ( .A1(n14699), .A2(n20365), .B1(n20375), .B2(n15014), .ZN(
        n14702) );
  NAND2_X1 U18125 ( .A1(n14812), .A2(n14700), .ZN(n14714) );
  NOR2_X1 U18126 ( .A1(n14714), .A2(n21163), .ZN(n14701) );
  AOI211_X1 U18127 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n20360), .A(n14702), .B(
        n14701), .ZN(n14703) );
  OAI21_X1 U18128 ( .B1(n15186), .B2(n20320), .A(n14703), .ZN(n14704) );
  AOI21_X1 U18129 ( .B1(n14705), .B2(n21163), .A(n14704), .ZN(n14706) );
  OAI21_X1 U18130 ( .B1(n14929), .B2(n14864), .A(n14706), .ZN(P1_U2813) );
  AOI21_X1 U18131 ( .B1(n14708), .B2(n14721), .A(n10243), .ZN(n15027) );
  INV_X1 U18132 ( .A(n15027), .ZN(n14932) );
  AND2_X1 U18133 ( .A1(n9706), .A2(n14709), .ZN(n14711) );
  OR2_X1 U18134 ( .A1(n14711), .A2(n14710), .ZN(n15200) );
  INV_X1 U18135 ( .A(n15200), .ZN(n14716) );
  INV_X1 U18136 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21000) );
  AOI22_X1 U18137 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20348), .B1(
        n20349), .B2(n15023), .ZN(n14713) );
  NAND2_X1 U18138 ( .A1(n20360), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14712) );
  OAI211_X1 U18139 ( .C1(n14714), .C2(n21000), .A(n14713), .B(n14712), .ZN(
        n14715) );
  AOI21_X1 U18140 ( .B1(n14716), .B2(n20362), .A(n14715), .ZN(n14719) );
  NAND2_X1 U18141 ( .A1(n14717), .A2(n21000), .ZN(n14718) );
  OAI211_X1 U18142 ( .C1(n14932), .C2(n14864), .A(n14719), .B(n14718), .ZN(
        P1_U2814) );
  XNOR2_X1 U18143 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14733) );
  AOI21_X1 U18144 ( .B1(n14722), .B2(n14735), .A(n12542), .ZN(n15034) );
  NAND2_X1 U18145 ( .A1(n15034), .A2(n20328), .ZN(n14732) );
  NAND2_X1 U18146 ( .A1(n14739), .A2(n14723), .ZN(n14724) );
  AND2_X1 U18147 ( .A1(n9706), .A2(n14724), .ZN(n15209) );
  INV_X1 U18148 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21187) );
  INV_X1 U18149 ( .A(n14725), .ZN(n14726) );
  NAND2_X1 U18150 ( .A1(n14812), .A2(n14726), .ZN(n14752) );
  OAI22_X1 U18151 ( .A1(n14727), .A2(n20365), .B1(n20375), .B2(n15032), .ZN(
        n14728) );
  AOI21_X1 U18152 ( .B1(n20360), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14728), .ZN(
        n14729) );
  OAI21_X1 U18153 ( .B1(n21187), .B2(n14752), .A(n14729), .ZN(n14730) );
  AOI21_X1 U18154 ( .B1(n15209), .B2(n20362), .A(n14730), .ZN(n14731) );
  OAI211_X1 U18155 ( .C1(n14742), .C2(n14733), .A(n14732), .B(n14731), .ZN(
        P1_U2815) );
  OAI21_X1 U18156 ( .B1(n14734), .B2(n14736), .A(n14735), .ZN(n15039) );
  OR2_X1 U18157 ( .A1(n14749), .A2(n14737), .ZN(n14738) );
  AND2_X1 U18158 ( .A1(n14739), .A2(n14738), .ZN(n16305) );
  INV_X1 U18159 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21169) );
  AOI22_X1 U18160 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20348), .B1(
        n20349), .B2(n15042), .ZN(n14741) );
  NAND2_X1 U18161 ( .A1(n20360), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14740) );
  OAI211_X1 U18162 ( .C1(n14752), .C2(n21169), .A(n14741), .B(n14740), .ZN(
        n14744) );
  NOR2_X1 U18163 ( .A1(n14742), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14743) );
  AOI211_X1 U18164 ( .C1(n16305), .C2(n20362), .A(n14744), .B(n14743), .ZN(
        n14745) );
  OAI21_X1 U18165 ( .B1(n15039), .B2(n14864), .A(n14745), .ZN(P1_U2816) );
  INV_X1 U18166 ( .A(n14734), .ZN(n14747) );
  OAI21_X1 U18167 ( .B1(n14748), .B2(n14746), .A(n14747), .ZN(n15047) );
  AOI21_X1 U18168 ( .B1(n14750), .B2(n14762), .A(n14749), .ZN(n15213) );
  INV_X1 U18169 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14874) );
  AOI22_X1 U18170 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20348), .B1(
        n20349), .B2(n15050), .ZN(n14751) );
  OAI21_X1 U18171 ( .B1(n20325), .B2(n14874), .A(n14751), .ZN(n14755) );
  AOI21_X1 U18172 ( .B1(n14753), .B2(n20995), .A(n14752), .ZN(n14754) );
  AOI211_X1 U18173 ( .C1(n15213), .C2(n20362), .A(n14755), .B(n14754), .ZN(
        n14756) );
  OAI21_X1 U18174 ( .B1(n15047), .B2(n14864), .A(n14756), .ZN(P1_U2817) );
  INV_X1 U18175 ( .A(n16207), .ZN(n14769) );
  XNOR2_X1 U18176 ( .A(P1_REIP_REG_22__SCAN_IN), .B(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14768) );
  AOI21_X1 U18177 ( .B1(n14758), .B2(n14757), .A(n14746), .ZN(n15059) );
  NAND2_X1 U18178 ( .A1(n15059), .A2(n20328), .ZN(n14767) );
  NOR2_X1 U18179 ( .A1(n20307), .A2(n14759), .ZN(n16206) );
  INV_X1 U18180 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14876) );
  AOI22_X1 U18181 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20348), .B1(
        n20349), .B2(n15055), .ZN(n14760) );
  OAI21_X1 U18182 ( .B1(n20325), .B2(n14876), .A(n14760), .ZN(n14765) );
  OAI21_X1 U18183 ( .B1(n16169), .B2(n16170), .A(n14761), .ZN(n14763) );
  NAND2_X1 U18184 ( .A1(n14763), .A2(n14762), .ZN(n16314) );
  NOR2_X1 U18185 ( .A1(n16314), .A2(n20320), .ZN(n14764) );
  AOI211_X1 U18186 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n16206), .A(n14765), 
        .B(n14764), .ZN(n14766) );
  OAI211_X1 U18187 ( .C1(n14769), .C2(n14768), .A(n14767), .B(n14766), .ZN(
        P1_U2818) );
  OAI21_X1 U18188 ( .B1(n14770), .B2(n14772), .A(n14947), .ZN(n16255) );
  NAND2_X1 U18189 ( .A1(n20990), .A2(n14773), .ZN(n14779) );
  OR2_X1 U18190 ( .A1(n14786), .A2(n14774), .ZN(n14775) );
  AND2_X1 U18191 ( .A1(n16169), .A2(n14775), .ZN(n16193) );
  NAND2_X1 U18192 ( .A1(n16193), .A2(n20362), .ZN(n14777) );
  AOI22_X1 U18193 ( .A1(n20348), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n20349), .B2(n16257), .ZN(n14776) );
  OAI211_X1 U18194 ( .C1(n14877), .C2(n20325), .A(n14777), .B(n14776), .ZN(
        n14778) );
  AOI21_X1 U18195 ( .B1(n16206), .B2(n14779), .A(n14778), .ZN(n14780) );
  OAI21_X1 U18196 ( .B1(n16255), .B2(n14864), .A(n14780), .ZN(P1_U2820) );
  NOR2_X1 U18197 ( .A1(n9711), .A2(n14781), .ZN(n14782) );
  OR2_X1 U18198 ( .A1(n14770), .A2(n14782), .ZN(n16264) );
  NAND2_X1 U18199 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14783) );
  OAI211_X1 U18200 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(P1_REIP_REG_18__SCAN_IN), .A(n14804), .B(n14783), .ZN(n14795) );
  NOR2_X1 U18201 ( .A1(n14784), .A2(n20307), .ZN(n16211) );
  AND2_X1 U18202 ( .A1(n9707), .A2(n14785), .ZN(n14787) );
  OR2_X1 U18203 ( .A1(n14787), .A2(n14786), .ZN(n15223) );
  NAND2_X1 U18204 ( .A1(n20348), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14790) );
  NAND2_X1 U18205 ( .A1(n20349), .A2(n14788), .ZN(n14789) );
  AND3_X1 U18206 ( .A1(n14790), .A2(n14789), .A3(n20308), .ZN(n14792) );
  NAND2_X1 U18207 ( .A1(n20360), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n14791) );
  OAI211_X1 U18208 ( .C1(n15223), .C2(n20320), .A(n14792), .B(n14791), .ZN(
        n14793) );
  AOI21_X1 U18209 ( .B1(n16211), .B2(P1_REIP_REG_19__SCAN_IN), .A(n14793), 
        .ZN(n14794) );
  OAI211_X1 U18210 ( .C1(n16264), .C2(n14864), .A(n14795), .B(n14794), .ZN(
        P1_U2821) );
  INV_X1 U18211 ( .A(n14889), .ZN(n14796) );
  NOR2_X1 U18212 ( .A1(n9753), .A2(n14796), .ZN(n14798) );
  OAI21_X1 U18213 ( .B1(n14798), .B2(n14797), .A(n9707), .ZN(n16323) );
  AOI21_X1 U18214 ( .B1(n14800), .B2(n14799), .A(n9711), .ZN(n14883) );
  NAND2_X1 U18215 ( .A1(n14883), .A2(n20328), .ZN(n14806) );
  INV_X1 U18216 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20987) );
  AOI22_X1 U18217 ( .A1(n20360), .A2(P1_EBX_REG_18__SCAN_IN), .B1(n20349), 
        .B2(n15066), .ZN(n14801) );
  OAI211_X1 U18218 ( .C1(n20365), .C2(n14802), .A(n14801), .B(n20308), .ZN(
        n14803) );
  AOI221_X1 U18219 ( .B1(n14804), .B2(n20987), .C1(n16211), .C2(
        P1_REIP_REG_18__SCAN_IN), .A(n14803), .ZN(n14805) );
  OAI211_X1 U18220 ( .C1(n20320), .C2(n16323), .A(n14806), .B(n14805), .ZN(
        P1_U2822) );
  NAND2_X1 U18221 ( .A1(n14849), .A2(n14808), .ZN(n14824) );
  AOI21_X1 U18222 ( .B1(n14810), .B2(n14824), .A(n10231), .ZN(n15078) );
  NAND2_X1 U18223 ( .A1(n14812), .A2(n14811), .ZN(n14843) );
  INV_X1 U18224 ( .A(n14843), .ZN(n14833) );
  XNOR2_X1 U18225 ( .A(P1_REIP_REG_16__SCAN_IN), .B(n10076), .ZN(n14813) );
  AOI22_X1 U18226 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n14833), .B1(n9755), 
        .B2(n14813), .ZN(n14820) );
  AOI21_X1 U18227 ( .B1(n20348), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20346), .ZN(n14819) );
  OR2_X1 U18228 ( .A1(n14828), .A2(n14814), .ZN(n14815) );
  AND2_X1 U18229 ( .A1(n9753), .A2(n14815), .ZN(n16331) );
  AOI22_X1 U18230 ( .A1(n16331), .A2(n20362), .B1(n20360), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14818) );
  INV_X1 U18231 ( .A(n15076), .ZN(n14816) );
  NAND2_X1 U18232 ( .A1(n20349), .A2(n14816), .ZN(n14817) );
  NAND4_X1 U18233 ( .A1(n14820), .A2(n14819), .A3(n14818), .A4(n14817), .ZN(
        n14821) );
  AOI21_X1 U18234 ( .B1(n15078), .B2(n20328), .A(n14821), .ZN(n14822) );
  INV_X1 U18235 ( .A(n14822), .ZN(P1_U2824) );
  AND2_X1 U18236 ( .A1(n14849), .A2(n14823), .ZN(n14837) );
  INV_X1 U18237 ( .A(n16280), .ZN(n14831) );
  NOR2_X1 U18238 ( .A1(n14839), .A2(n14826), .ZN(n14827) );
  OR2_X1 U18239 ( .A1(n14828), .A2(n14827), .ZN(n16338) );
  INV_X1 U18240 ( .A(n16338), .ZN(n14892) );
  AOI22_X1 U18241 ( .A1(n14892), .A2(n20362), .B1(n20360), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14830) );
  AOI21_X1 U18242 ( .B1(n20348), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20346), .ZN(n14829) );
  OAI211_X1 U18243 ( .C1(n20375), .C2(n14831), .A(n14830), .B(n14829), .ZN(
        n14832) );
  AOI21_X1 U18244 ( .B1(n14833), .B2(P1_REIP_REG_15__SCAN_IN), .A(n14832), 
        .ZN(n14835) );
  NAND2_X1 U18245 ( .A1(n9755), .A2(n10076), .ZN(n14834) );
  OAI211_X1 U18246 ( .C1(n16279), .C2(n14864), .A(n14835), .B(n14834), .ZN(
        P1_U2825) );
  NAND2_X1 U18247 ( .A1(n14849), .A2(n14836), .ZN(n14895) );
  AOI21_X1 U18248 ( .B1(n14838), .B2(n14895), .A(n14837), .ZN(n15088) );
  INV_X1 U18249 ( .A(n15088), .ZN(n14978) );
  INV_X1 U18250 ( .A(n15086), .ZN(n14847) );
  INV_X1 U18251 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14842) );
  AOI21_X1 U18252 ( .B1(n14840), .B2(n10309), .A(n14839), .ZN(n16348) );
  AOI22_X1 U18253 ( .A1(n20362), .A2(n16348), .B1(n20360), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14841) );
  OAI211_X1 U18254 ( .C1(n20365), .C2(n14842), .A(n14841), .B(n20308), .ZN(
        n14846) );
  AOI21_X1 U18255 ( .B1(n20979), .B2(n14844), .A(n14843), .ZN(n14845) );
  AOI211_X1 U18256 ( .C1(n20349), .C2(n14847), .A(n14846), .B(n14845), .ZN(
        n14848) );
  OAI21_X1 U18257 ( .B1(n14978), .B2(n14864), .A(n14848), .ZN(P1_U2826) );
  NAND2_X1 U18258 ( .A1(n14849), .A2(n14851), .ZN(n14897) );
  INV_X1 U18259 ( .A(n14851), .ZN(n14853) );
  NAND3_X1 U18260 ( .A1(n14850), .A2(n14853), .A3(n14852), .ZN(n14854) );
  NAND2_X1 U18261 ( .A1(n14897), .A2(n14854), .ZN(n15110) );
  INV_X1 U18262 ( .A(n15106), .ZN(n14862) );
  INV_X1 U18263 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14857) );
  OAI21_X1 U18264 ( .B1(n14910), .B2(n14855), .A(n14900), .ZN(n14906) );
  INV_X1 U18265 ( .A(n14906), .ZN(n16369) );
  AOI22_X1 U18266 ( .A1(n20362), .A2(n16369), .B1(n20360), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n14856) );
  OAI211_X1 U18267 ( .C1(n20365), .C2(n14857), .A(n14856), .B(n20308), .ZN(
        n14861) );
  INV_X1 U18268 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20977) );
  INV_X1 U18269 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20975) );
  OR2_X1 U18270 ( .A1(n14858), .A2(n20307), .ZN(n16226) );
  INV_X1 U18271 ( .A(n16226), .ZN(n16241) );
  AOI21_X1 U18272 ( .B1(n20366), .B2(n14859), .A(n16241), .ZN(n16225) );
  AOI221_X1 U18273 ( .B1(n16234), .B2(n20977), .C1(n20975), .C2(n20977), .A(
        n16225), .ZN(n14860) );
  AOI211_X1 U18274 ( .C1(n20349), .C2(n14862), .A(n14861), .B(n14860), .ZN(
        n14863) );
  OAI21_X1 U18275 ( .B1(n14864), .B2(n15110), .A(n14863), .ZN(P1_U2828) );
  INV_X1 U18276 ( .A(n15140), .ZN(n14866) );
  INV_X1 U18277 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14865) );
  OAI22_X1 U18278 ( .A1(n14866), .A2(n14916), .B1(n14865), .B2(n20387), .ZN(
        P1_U2841) );
  OAI222_X1 U18279 ( .A1(n14914), .A2(n14921), .B1(n20387), .B2(n14868), .C1(
        n14867), .C2(n14916), .ZN(P1_U2842) );
  OAI222_X1 U18280 ( .A1(n15173), .A2(n14916), .B1(n14869), .B2(n20387), .C1(
        n14926), .C2(n14884), .ZN(P1_U2843) );
  OAI222_X1 U18281 ( .A1(n15186), .A2(n14916), .B1(n14870), .B2(n20387), .C1(
        n14929), .C2(n14884), .ZN(P1_U2845) );
  OAI222_X1 U18282 ( .A1(n15200), .A2(n14916), .B1(n14871), .B2(n20387), .C1(
        n14932), .C2(n14884), .ZN(P1_U2846) );
  INV_X1 U18283 ( .A(n15034), .ZN(n14936) );
  AOI22_X1 U18284 ( .A1(n15209), .A2(n20382), .B1(n14902), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14872) );
  OAI21_X1 U18285 ( .B1(n14936), .B2(n14914), .A(n14872), .ZN(P1_U2847) );
  AOI22_X1 U18286 ( .A1(n16305), .A2(n20382), .B1(n14902), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n14873) );
  OAI21_X1 U18287 ( .B1(n15039), .B2(n14914), .A(n14873), .ZN(P1_U2848) );
  INV_X1 U18288 ( .A(n15213), .ZN(n14875) );
  OAI222_X1 U18289 ( .A1(n14875), .A2(n14916), .B1(n14874), .B2(n20387), .C1(
        n15047), .C2(n14884), .ZN(P1_U2849) );
  INV_X1 U18290 ( .A(n15059), .ZN(n14945) );
  OAI222_X1 U18291 ( .A1(n16314), .A2(n14916), .B1(n14876), .B2(n20387), .C1(
        n14945), .C2(n14884), .ZN(P1_U2850) );
  NOR2_X1 U18292 ( .A1(n20387), .A2(n14877), .ZN(n14878) );
  AOI21_X1 U18293 ( .B1(n16193), .B2(n20382), .A(n14878), .ZN(n14879) );
  OAI21_X1 U18294 ( .B1(n16255), .B2(n14914), .A(n14879), .ZN(P1_U2852) );
  OAI22_X1 U18295 ( .A1(n15223), .A2(n14916), .B1(n14880), .B2(n20387), .ZN(
        n14881) );
  INV_X1 U18296 ( .A(n14881), .ZN(n14882) );
  OAI21_X1 U18297 ( .B1(n16264), .B2(n14914), .A(n14882), .ZN(P1_U2853) );
  INV_X1 U18298 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14885) );
  INV_X1 U18299 ( .A(n14883), .ZN(n15068) );
  OAI222_X1 U18300 ( .A1(n16323), .A2(n14916), .B1(n14885), .B2(n20387), .C1(
        n15068), .C2(n14884), .ZN(P1_U2854) );
  INV_X1 U18301 ( .A(n14799), .ZN(n14886) );
  AOI21_X1 U18302 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n16270) );
  INV_X1 U18303 ( .A(n16270), .ZN(n14968) );
  XNOR2_X1 U18304 ( .A(n9753), .B(n14889), .ZN(n16210) );
  AOI22_X1 U18305 ( .A1(n16210), .A2(n20382), .B1(n14902), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n14890) );
  OAI21_X1 U18306 ( .B1(n14968), .B2(n14914), .A(n14890), .ZN(P1_U2855) );
  INV_X1 U18307 ( .A(n15078), .ZN(n14975) );
  AOI22_X1 U18308 ( .A1(n16331), .A2(n20382), .B1(n14902), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14891) );
  OAI21_X1 U18309 ( .B1(n14975), .B2(n14914), .A(n14891), .ZN(P1_U2856) );
  AOI22_X1 U18310 ( .A1(n14892), .A2(n20382), .B1(n14902), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14893) );
  OAI21_X1 U18311 ( .B1(n16279), .B2(n14914), .A(n14893), .ZN(P1_U2857) );
  AOI22_X1 U18312 ( .A1(n16348), .A2(n20382), .B1(n14902), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14894) );
  OAI21_X1 U18313 ( .B1(n14978), .B2(n14914), .A(n14894), .ZN(P1_U2858) );
  INV_X1 U18314 ( .A(n14895), .ZN(n14896) );
  AOI21_X1 U18315 ( .B1(n14898), .B2(n14897), .A(n14896), .ZN(n16222) );
  INV_X1 U18316 ( .A(n16222), .ZN(n14983) );
  NAND2_X1 U18317 ( .A1(n14900), .A2(n14899), .ZN(n14901) );
  NAND2_X1 U18318 ( .A1(n10309), .A2(n14901), .ZN(n16359) );
  INV_X1 U18319 ( .A(n16359), .ZN(n14903) );
  AOI22_X1 U18320 ( .A1(n20382), .A2(n14903), .B1(n14902), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14904) );
  OAI21_X1 U18321 ( .B1(n14983), .B2(n14914), .A(n14904), .ZN(P1_U2859) );
  INV_X1 U18322 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14905) );
  OAI222_X1 U18323 ( .A1(n14906), .A2(n14916), .B1(n14905), .B2(n20387), .C1(
        n14914), .C2(n15110), .ZN(P1_U2860) );
  AND2_X1 U18324 ( .A1(n14908), .A2(n14907), .ZN(n14909) );
  NOR2_X1 U18325 ( .A1(n14910), .A2(n14909), .ZN(n16386) );
  INV_X1 U18326 ( .A(n16386), .ZN(n16227) );
  INV_X1 U18327 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14915) );
  OR2_X1 U18328 ( .A1(n14912), .A2(n14911), .ZN(n14913) );
  AND2_X1 U18329 ( .A1(n14850), .A2(n14913), .ZN(n16231) );
  INV_X1 U18330 ( .A(n16231), .ZN(n14990) );
  OAI222_X1 U18331 ( .A1(n16227), .A2(n14916), .B1(n20387), .B2(n14915), .C1(
        n14914), .C2(n14990), .ZN(P1_U2861) );
  AOI22_X1 U18332 ( .A1(n14969), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14979), .ZN(n14920) );
  INV_X1 U18333 ( .A(DATAI_14_), .ZN(n14918) );
  NAND2_X1 U18334 ( .A1(n14923), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14917) );
  OAI21_X1 U18335 ( .B1(n14923), .B2(n14918), .A(n14917), .ZN(n20425) );
  AOI22_X1 U18336 ( .A1(n14972), .A2(n20425), .B1(n14970), .B2(DATAI_30_), 
        .ZN(n14919) );
  OAI211_X1 U18337 ( .C1(n14921), .C2(n14982), .A(n14920), .B(n14919), .ZN(
        P1_U2874) );
  AOI22_X1 U18338 ( .A1(n14969), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14979), .ZN(n14925) );
  INV_X1 U18339 ( .A(DATAI_13_), .ZN(n21206) );
  NAND2_X1 U18340 ( .A1(n14923), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14922) );
  OAI21_X1 U18341 ( .B1(n14923), .B2(n21206), .A(n14922), .ZN(n20423) );
  AOI22_X1 U18342 ( .A1(n14972), .A2(n20423), .B1(n14970), .B2(DATAI_29_), 
        .ZN(n14924) );
  OAI211_X1 U18343 ( .C1(n14926), .C2(n14982), .A(n14925), .B(n14924), .ZN(
        P1_U2875) );
  AOI22_X1 U18344 ( .A1(n14969), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14979), .ZN(n14928) );
  AOI22_X1 U18345 ( .A1(n14972), .A2(n14986), .B1(n14970), .B2(DATAI_27_), 
        .ZN(n14927) );
  OAI211_X1 U18346 ( .C1(n14929), .C2(n14982), .A(n14928), .B(n14927), .ZN(
        P1_U2877) );
  AOI22_X1 U18347 ( .A1(n14969), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14979), .ZN(n14931) );
  AOI22_X1 U18348 ( .A1(n14972), .A2(n20419), .B1(n14970), .B2(DATAI_26_), 
        .ZN(n14930) );
  OAI211_X1 U18349 ( .C1(n14932), .C2(n14982), .A(n14931), .B(n14930), .ZN(
        P1_U2878) );
  AOI22_X1 U18350 ( .A1(n14969), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14979), .ZN(n14935) );
  AOI22_X1 U18351 ( .A1(n14972), .A2(n14933), .B1(n14970), .B2(DATAI_25_), 
        .ZN(n14934) );
  OAI211_X1 U18352 ( .C1(n14936), .C2(n14982), .A(n14935), .B(n14934), .ZN(
        P1_U2879) );
  AOI22_X1 U18353 ( .A1(n14969), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14979), .ZN(n14938) );
  AOI22_X1 U18354 ( .A1(n14972), .A2(n20417), .B1(n14970), .B2(DATAI_24_), 
        .ZN(n14937) );
  OAI211_X1 U18355 ( .C1(n15039), .C2(n14982), .A(n14938), .B(n14937), .ZN(
        P1_U2880) );
  AOI22_X1 U18356 ( .A1(n14969), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14979), .ZN(n14941) );
  AOI22_X1 U18357 ( .A1(n14972), .A2(n14939), .B1(n14970), .B2(DATAI_23_), 
        .ZN(n14940) );
  OAI211_X1 U18358 ( .C1(n15047), .C2(n14982), .A(n14941), .B(n14940), .ZN(
        P1_U2881) );
  AOI22_X1 U18359 ( .A1(n14969), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14979), .ZN(n14944) );
  AOI22_X1 U18360 ( .A1(n14972), .A2(n14942), .B1(n14970), .B2(DATAI_22_), 
        .ZN(n14943) );
  OAI211_X1 U18361 ( .C1(n14945), .C2(n14982), .A(n14944), .B(n14943), .ZN(
        P1_U2882) );
  INV_X1 U18362 ( .A(n14757), .ZN(n14946) );
  AOI21_X1 U18363 ( .B1(n14948), .B2(n14947), .A(n14946), .ZN(n16250) );
  INV_X1 U18364 ( .A(n16250), .ZN(n14953) );
  OAI22_X1 U18365 ( .A1(n14957), .A2(n19595), .B1(n13772), .B2(n14987), .ZN(
        n14949) );
  INV_X1 U18366 ( .A(n14949), .ZN(n14952) );
  AOI22_X1 U18367 ( .A1(n14972), .A2(n14950), .B1(n14970), .B2(DATAI_21_), 
        .ZN(n14951) );
  OAI211_X1 U18368 ( .C1(n14953), .C2(n14982), .A(n14952), .B(n14951), .ZN(
        P1_U2883) );
  AOI22_X1 U18369 ( .A1(n14969), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14979), .ZN(n14955) );
  AOI22_X1 U18370 ( .A1(n14972), .A2(n15337), .B1(n14970), .B2(DATAI_20_), 
        .ZN(n14954) );
  OAI211_X1 U18371 ( .C1(n16255), .C2(n14982), .A(n14955), .B(n14954), .ZN(
        P1_U2884) );
  OAI22_X1 U18372 ( .A1(n14957), .A2(n16781), .B1(n14956), .B2(n14987), .ZN(
        n14958) );
  INV_X1 U18373 ( .A(n14958), .ZN(n14961) );
  AOI22_X1 U18374 ( .A1(n14972), .A2(n14959), .B1(n14970), .B2(DATAI_19_), 
        .ZN(n14960) );
  OAI211_X1 U18375 ( .C1(n16264), .C2(n14982), .A(n14961), .B(n14960), .ZN(
        P1_U2885) );
  AOI22_X1 U18376 ( .A1(n14969), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14979), .ZN(n14964) );
  AOI22_X1 U18377 ( .A1(n14972), .A2(n14962), .B1(n14970), .B2(DATAI_18_), 
        .ZN(n14963) );
  OAI211_X1 U18378 ( .C1(n15068), .C2(n14982), .A(n14964), .B(n14963), .ZN(
        P1_U2886) );
  AOI22_X1 U18379 ( .A1(n14969), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14979), .ZN(n14967) );
  AOI22_X1 U18380 ( .A1(n14972), .A2(n14965), .B1(n14970), .B2(DATAI_17_), 
        .ZN(n14966) );
  OAI211_X1 U18381 ( .C1(n14968), .C2(n14982), .A(n14967), .B(n14966), .ZN(
        P1_U2887) );
  AOI22_X1 U18382 ( .A1(n14969), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14979), .ZN(n14974) );
  AOI22_X1 U18383 ( .A1(n14972), .A2(n14971), .B1(n14970), .B2(DATAI_16_), 
        .ZN(n14973) );
  OAI211_X1 U18384 ( .C1(n14975), .C2(n14982), .A(n14974), .B(n14973), .ZN(
        P1_U2888) );
  OAI222_X1 U18385 ( .A1(n16279), .A2(n14982), .B1(n14989), .B2(n14976), .C1(
        n14987), .C2(n12239), .ZN(P1_U2889) );
  AOI22_X1 U18386 ( .A1(n14980), .A2(n20425), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14979), .ZN(n14977) );
  OAI21_X1 U18387 ( .B1(n14978), .B2(n14982), .A(n14977), .ZN(P1_U2890) );
  AOI22_X1 U18388 ( .A1(n14980), .A2(n20423), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14979), .ZN(n14981) );
  OAI21_X1 U18389 ( .B1(n14983), .B2(n14982), .A(n14981), .ZN(P1_U2891) );
  INV_X1 U18390 ( .A(n20421), .ZN(n14985) );
  OAI222_X1 U18391 ( .A1(n15110), .A2(n14982), .B1(n14989), .B2(n14985), .C1(
        n14984), .C2(n14987), .ZN(P1_U2892) );
  INV_X1 U18392 ( .A(n14986), .ZN(n14988) );
  OAI222_X1 U18393 ( .A1(n14990), .A2(n14982), .B1(n14989), .B2(n14988), .C1(
        n20397), .C2(n14987), .ZN(P1_U2893) );
  XNOR2_X1 U18394 ( .A(n15224), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14991) );
  XNOR2_X1 U18395 ( .A(n14992), .B(n14991), .ZN(n15177) );
  NOR2_X1 U18396 ( .A1(n16406), .A2(n21094), .ZN(n15170) );
  AOI21_X1 U18397 ( .B1(n16291), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15170), .ZN(n14993) );
  OAI21_X1 U18398 ( .B1(n16299), .B2(n14994), .A(n14993), .ZN(n14995) );
  AOI21_X1 U18399 ( .B1(n14996), .B2(n16286), .A(n14995), .ZN(n14997) );
  OAI21_X1 U18400 ( .B1(n15177), .B2(n20282), .A(n14997), .ZN(P1_U2970) );
  INV_X1 U18401 ( .A(n15045), .ZN(n14998) );
  OAI21_X1 U18402 ( .B1(n14998), .B2(n15151), .A(n15036), .ZN(n15000) );
  NAND2_X1 U18403 ( .A1(n16391), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15178) );
  OAI21_X1 U18404 ( .B1(n16260), .B2(n15002), .A(n15178), .ZN(n15005) );
  NOR2_X1 U18405 ( .A1(n15003), .A2(n16263), .ZN(n15004) );
  AOI211_X2 U18406 ( .C1(n16285), .C2(n15006), .A(n15005), .B(n15004), .ZN(
        n15007) );
  MUX2_X1 U18407 ( .A(n15009), .B(n15008), .S(n16163), .Z(n15011) );
  NOR2_X1 U18408 ( .A1(n15011), .A2(n15010), .ZN(n15012) );
  XNOR2_X1 U18409 ( .A(n15012), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15194) );
  NOR2_X1 U18410 ( .A1(n16406), .A2(n21163), .ZN(n15188) );
  AOI21_X1 U18411 ( .B1(n16291), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15188), .ZN(n15013) );
  OAI21_X1 U18412 ( .B1(n16299), .B2(n15014), .A(n15013), .ZN(n15015) );
  AOI21_X1 U18413 ( .B1(n15016), .B2(n16286), .A(n15015), .ZN(n15017) );
  OAI21_X1 U18414 ( .B1(n20282), .B2(n15194), .A(n15017), .ZN(P1_U2972) );
  NOR2_X1 U18415 ( .A1(n15018), .A2(n15151), .ZN(n15020) );
  OAI21_X1 U18416 ( .B1(n15021), .B2(n15020), .A(n15019), .ZN(n15022) );
  XOR2_X1 U18417 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15022), .Z(
        n15204) );
  INV_X1 U18418 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15025) );
  NAND2_X1 U18419 ( .A1(n16285), .A2(n15023), .ZN(n15024) );
  NAND2_X1 U18420 ( .A1(n16391), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15198) );
  OAI211_X1 U18421 ( .C1(n16260), .C2(n15025), .A(n15024), .B(n15198), .ZN(
        n15026) );
  AOI21_X1 U18422 ( .B1(n15027), .B2(n16286), .A(n15026), .ZN(n15028) );
  OAI21_X1 U18423 ( .B1(n20282), .B2(n15204), .A(n15028), .ZN(P1_U2973) );
  MUX2_X1 U18424 ( .A(n15018), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .S(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n15029) );
  OAI211_X1 U18425 ( .C1(n16302), .C2(n15045), .A(n15036), .B(n15029), .ZN(
        n15030) );
  XNOR2_X1 U18426 ( .A(n15030), .B(n15205), .ZN(n15212) );
  NOR2_X1 U18427 ( .A1(n16406), .A2(n21187), .ZN(n15208) );
  AOI21_X1 U18428 ( .B1(n16291), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15208), .ZN(n15031) );
  OAI21_X1 U18429 ( .B1(n16299), .B2(n15032), .A(n15031), .ZN(n15033) );
  AOI21_X1 U18430 ( .B1(n15034), .B2(n16286), .A(n15033), .ZN(n15035) );
  OAI21_X1 U18431 ( .B1(n20282), .B2(n15212), .A(n15035), .ZN(P1_U2974) );
  XNOR2_X1 U18432 ( .A(n15227), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15044) );
  NAND3_X1 U18433 ( .A1(n15036), .A2(n15044), .A3(n15019), .ZN(n15037) );
  XNOR2_X1 U18434 ( .A(n15037), .B(n16301), .ZN(n16304) );
  OAI22_X1 U18435 ( .A1(n16260), .A2(n15038), .B1(n16406), .B2(n21169), .ZN(
        n15041) );
  NOR2_X1 U18436 ( .A1(n15039), .A2(n16263), .ZN(n15040) );
  AOI211_X1 U18437 ( .C1(n16285), .C2(n15042), .A(n15041), .B(n15040), .ZN(
        n15043) );
  OAI21_X1 U18438 ( .B1(n20282), .B2(n16304), .A(n15043), .ZN(P1_U2975) );
  XNOR2_X1 U18439 ( .A(n15045), .B(n15044), .ZN(n15219) );
  NAND2_X1 U18440 ( .A1(n16391), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15215) );
  OAI21_X1 U18441 ( .B1(n16260), .B2(n15046), .A(n15215), .ZN(n15049) );
  NOR2_X1 U18442 ( .A1(n15047), .A2(n16263), .ZN(n15048) );
  AOI211_X1 U18443 ( .C1(n16285), .C2(n15050), .A(n15049), .B(n15048), .ZN(
        n15051) );
  OAI21_X1 U18444 ( .B1(n15219), .B2(n20282), .A(n15051), .ZN(P1_U2976) );
  NAND2_X1 U18445 ( .A1(n15053), .A2(n15052), .ZN(n15054) );
  XOR2_X1 U18446 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15054), .Z(
        n16313) );
  INV_X1 U18447 ( .A(n15055), .ZN(n15057) );
  AOI22_X1 U18448 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15056) );
  OAI21_X1 U18449 ( .B1(n16299), .B2(n15057), .A(n15056), .ZN(n15058) );
  AOI21_X1 U18450 ( .B1(n15059), .B2(n16286), .A(n15058), .ZN(n15060) );
  OAI21_X1 U18451 ( .B1(n20282), .B2(n16313), .A(n15060), .ZN(P1_U2977) );
  OAI22_X1 U18452 ( .A1(n16260), .A2(n14802), .B1(n16406), .B2(n20987), .ZN(
        n15065) );
  OAI21_X1 U18453 ( .B1(n15063), .B2(n15062), .A(n15061), .ZN(n16322) );
  NOR2_X1 U18454 ( .A1(n16322), .A2(n20282), .ZN(n15064) );
  AOI211_X1 U18455 ( .C1(n16285), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15067) );
  OAI21_X1 U18456 ( .B1(n15068), .B2(n16263), .A(n15067), .ZN(P1_U2981) );
  INV_X1 U18457 ( .A(n15092), .ZN(n15070) );
  OAI21_X1 U18458 ( .B1(n15069), .B2(n15071), .A(n15070), .ZN(n16274) );
  OAI21_X1 U18459 ( .B1(n16274), .B2(n15072), .A(n16275), .ZN(n15073) );
  XOR2_X1 U18460 ( .A(n15074), .B(n15073), .Z(n16330) );
  AOI22_X1 U18461 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15075) );
  OAI21_X1 U18462 ( .B1(n16299), .B2(n15076), .A(n15075), .ZN(n15077) );
  AOI21_X1 U18463 ( .B1(n15078), .B2(n16286), .A(n15077), .ZN(n15079) );
  OAI21_X1 U18464 ( .B1(n20282), .B2(n16330), .A(n15079), .ZN(P1_U2983) );
  INV_X1 U18465 ( .A(n15069), .ZN(n15252) );
  NOR2_X1 U18466 ( .A1(n15252), .A2(n15092), .ZN(n15237) );
  NAND2_X1 U18467 ( .A1(n15080), .A2(n15102), .ZN(n15082) );
  OAI21_X1 U18468 ( .B1(n15237), .B2(n15082), .A(n15081), .ZN(n15084) );
  XNOR2_X1 U18469 ( .A(n15018), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15083) );
  XNOR2_X1 U18470 ( .A(n15084), .B(n15083), .ZN(n16349) );
  INV_X1 U18471 ( .A(n16349), .ZN(n15090) );
  AOI22_X1 U18472 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15085) );
  OAI21_X1 U18473 ( .B1(n16299), .B2(n15086), .A(n15085), .ZN(n15087) );
  AOI21_X1 U18474 ( .B1(n15088), .B2(n16286), .A(n15087), .ZN(n15089) );
  OAI21_X1 U18475 ( .B1(n15090), .B2(n20282), .A(n15089), .ZN(P1_U2985) );
  NOR2_X1 U18476 ( .A1(n15069), .A2(n15091), .ZN(n15099) );
  OAI21_X1 U18477 ( .B1(n15099), .B2(n15092), .A(n15102), .ZN(n15094) );
  XNOR2_X1 U18478 ( .A(n15094), .B(n15093), .ZN(n16360) );
  AOI22_X1 U18479 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n15095) );
  OAI21_X1 U18480 ( .B1(n16299), .B2(n15096), .A(n15095), .ZN(n15097) );
  AOI21_X1 U18481 ( .B1(n16222), .B2(n16286), .A(n15097), .ZN(n15098) );
  OAI21_X1 U18482 ( .B1(n20282), .B2(n16360), .A(n15098), .ZN(P1_U2986) );
  INV_X1 U18483 ( .A(n15099), .ZN(n15101) );
  NAND2_X1 U18484 ( .A1(n15101), .A2(n15100), .ZN(n15105) );
  NAND2_X1 U18485 ( .A1(n15103), .A2(n15102), .ZN(n15104) );
  XNOR2_X1 U18486 ( .A(n15105), .B(n15104), .ZN(n16379) );
  INV_X1 U18487 ( .A(n20282), .ZN(n16296) );
  NAND2_X1 U18488 ( .A1(n16379), .A2(n16296), .ZN(n15109) );
  NOR2_X1 U18489 ( .A1(n16406), .A2(n20977), .ZN(n16368) );
  NOR2_X1 U18490 ( .A1(n16299), .A2(n15106), .ZN(n15107) );
  AOI211_X1 U18491 ( .C1(n16291), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16368), .B(n15107), .ZN(n15108) );
  OAI211_X1 U18492 ( .C1(n16263), .C2(n15110), .A(n15109), .B(n15108), .ZN(
        P1_U2987) );
  NOR3_X1 U18493 ( .A1(n15069), .A2(n15018), .A3(n15266), .ZN(n15255) );
  NOR3_X1 U18494 ( .A1(n15251), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15224), .ZN(n15111) );
  NOR2_X1 U18495 ( .A1(n15255), .A2(n15111), .ZN(n15112) );
  XNOR2_X1 U18496 ( .A(n15112), .B(n16389), .ZN(n16384) );
  AOI22_X1 U18497 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15113) );
  OAI21_X1 U18498 ( .B1(n16299), .B2(n16229), .A(n15113), .ZN(n15114) );
  AOI21_X1 U18499 ( .B1(n16231), .B2(n16286), .A(n15114), .ZN(n15115) );
  OAI21_X1 U18500 ( .B1(n16384), .B2(n20282), .A(n15115), .ZN(P1_U2988) );
  XNOR2_X1 U18501 ( .A(n15227), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15116) );
  XNOR2_X1 U18502 ( .A(n15117), .B(n15116), .ZN(n15278) );
  INV_X1 U18503 ( .A(n15118), .ZN(n15122) );
  AOI22_X1 U18504 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n15119) );
  OAI21_X1 U18505 ( .B1(n16299), .B2(n15120), .A(n15119), .ZN(n15121) );
  AOI21_X1 U18506 ( .B1(n15122), .B2(n16286), .A(n15121), .ZN(n15123) );
  OAI21_X1 U18507 ( .B1(n15278), .B2(n20282), .A(n15123), .ZN(P1_U2990) );
  XOR2_X1 U18508 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n15124), .Z(
        n15125) );
  XNOR2_X1 U18509 ( .A(n15126), .B(n15125), .ZN(n15295) );
  INV_X1 U18510 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U18511 ( .A1(n16406), .A2(n15127), .ZN(n15292) );
  AND2_X1 U18512 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15128) );
  AOI211_X1 U18513 ( .C1(n16285), .C2(n20301), .A(n15292), .B(n15128), .ZN(
        n15131) );
  NAND2_X1 U18514 ( .A1(n20377), .A2(n16286), .ZN(n15130) );
  OAI211_X1 U18515 ( .C1(n15295), .C2(n20282), .A(n15131), .B(n15130), .ZN(
        P1_U2991) );
  NAND2_X1 U18516 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16311) );
  INV_X1 U18517 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15226) );
  NAND3_X1 U18518 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15141) );
  INV_X1 U18519 ( .A(n15141), .ZN(n15246) );
  INV_X1 U18520 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15284) );
  INV_X1 U18521 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15283) );
  NOR3_X1 U18522 ( .A1(n15284), .A2(n15283), .A3(n16414), .ZN(n15257) );
  NOR2_X1 U18523 ( .A1(n15266), .A2(n15275), .ZN(n16346) );
  NAND2_X1 U18524 ( .A1(n15257), .A2(n16346), .ZN(n15134) );
  NOR2_X1 U18525 ( .A1(n16389), .A2(n15134), .ZN(n16372) );
  NAND3_X1 U18526 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15258), .A3(
        n16372), .ZN(n16358) );
  NOR2_X1 U18527 ( .A1(n16357), .A2(n16358), .ZN(n15244) );
  NAND3_X1 U18528 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15133), .A3(
        n15132), .ZN(n15260) );
  NOR2_X1 U18529 ( .A1(n15134), .A2(n15260), .ZN(n16373) );
  NAND3_X1 U18530 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n16373), .ZN(n16367) );
  NOR2_X1 U18531 ( .A1(n16357), .A2(n16367), .ZN(n15241) );
  AOI22_X1 U18532 ( .A1(n15147), .A2(n15244), .B1(n15241), .B2(n16370), .ZN(
        n15135) );
  INV_X1 U18533 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16347) );
  NOR2_X1 U18534 ( .A1(n15135), .A2(n16347), .ZN(n16334) );
  NAND2_X1 U18535 ( .A1(n15246), .A2(n16334), .ZN(n16328) );
  NOR2_X1 U18536 ( .A1(n15226), .A2(n16328), .ZN(n16186) );
  NAND2_X1 U18537 ( .A1(n16167), .A2(n16186), .ZN(n16320) );
  INV_X1 U18538 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15196) );
  NOR2_X1 U18539 ( .A1(n15151), .A2(n15196), .ZN(n15136) );
  INV_X1 U18540 ( .A(n15182), .ZN(n15169) );
  NAND3_X1 U18541 ( .A1(n15191), .A2(n15169), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15162) );
  NOR3_X1 U18542 ( .A1(n15162), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15137), .ZN(n15138) );
  AOI211_X1 U18543 ( .C1(n20451), .C2(n15140), .A(n15139), .B(n15138), .ZN(
        n15157) );
  NOR3_X1 U18544 ( .A1(n15226), .A2(n16347), .A3(n15141), .ZN(n15142) );
  NAND2_X1 U18545 ( .A1(n15244), .A2(n15142), .ZN(n15144) );
  AOI21_X1 U18546 ( .B1(n15142), .B2(n15241), .A(n16374), .ZN(n15143) );
  NOR2_X1 U18547 ( .A1(n15145), .A2(n15245), .ZN(n15146) );
  AOI21_X1 U18548 ( .B1(n16167), .B2(n16195), .A(n15146), .ZN(n16312) );
  AOI21_X1 U18549 ( .B1(n15245), .B2(n16311), .A(n16312), .ZN(n15216) );
  NAND2_X1 U18550 ( .A1(n15147), .A2(n16302), .ZN(n15148) );
  NAND2_X1 U18551 ( .A1(n15216), .A2(n15148), .ZN(n16300) );
  NOR2_X1 U18552 ( .A1(n15149), .A2(n15195), .ZN(n15150) );
  OR2_X1 U18553 ( .A1(n16300), .A2(n15150), .ZN(n15155) );
  INV_X1 U18554 ( .A(n15151), .ZN(n15197) );
  OAI22_X1 U18555 ( .A1(n15197), .A2(n20453), .B1(n16371), .B2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15152) );
  NOR2_X1 U18556 ( .A1(n15155), .A2(n15152), .ZN(n15206) );
  NAND2_X1 U18557 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15153) );
  NAND2_X1 U18558 ( .A1(n15245), .A2(n15153), .ZN(n15154) );
  NAND2_X1 U18559 ( .A1(n15206), .A2(n15154), .ZN(n15189) );
  AOI21_X1 U18560 ( .B1(n15182), .B2(n15245), .A(n15189), .ZN(n15168) );
  OAI211_X1 U18561 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15282), .A(
        n15168), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15163) );
  OAI211_X1 U18562 ( .C1(n15245), .C2(n15155), .A(n15163), .B(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15156) );
  OAI211_X1 U18563 ( .C1(n15158), .C2(n20446), .A(n15157), .B(n15156), .ZN(
        P1_U3000) );
  INV_X1 U18564 ( .A(n15159), .ZN(n15160) );
  AOI21_X1 U18565 ( .B1(n15161), .B2(n20451), .A(n15160), .ZN(n15166) );
  INV_X1 U18566 ( .A(n15162), .ZN(n15164) );
  OAI21_X1 U18567 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15164), .A(
        n15163), .ZN(n15165) );
  OAI211_X1 U18568 ( .C1(n15167), .C2(n20446), .A(n15166), .B(n15165), .ZN(
        P1_U3001) );
  INV_X1 U18569 ( .A(n15168), .ZN(n15175) );
  NAND3_X1 U18570 ( .A1(n15191), .A2(n15169), .A3(n12846), .ZN(n15172) );
  INV_X1 U18571 ( .A(n15170), .ZN(n15171) );
  OAI211_X1 U18572 ( .C1(n16407), .C2(n15173), .A(n15172), .B(n15171), .ZN(
        n15174) );
  AOI21_X1 U18573 ( .B1(n15175), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15174), .ZN(n15176) );
  OAI21_X1 U18574 ( .B1(n15177), .B2(n20446), .A(n15176), .ZN(P1_U3002) );
  OAI21_X1 U18575 ( .B1(n15179), .B2(n16407), .A(n15178), .ZN(n15180) );
  AOI21_X1 U18576 ( .B1(n15189), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15180), .ZN(n15184) );
  NAND3_X1 U18577 ( .A1(n15191), .A2(n15182), .A3(n15181), .ZN(n15183) );
  OAI211_X1 U18578 ( .C1(n15185), .C2(n20446), .A(n15184), .B(n15183), .ZN(
        P1_U3003) );
  NOR2_X1 U18579 ( .A1(n15186), .A2(n16407), .ZN(n15187) );
  AOI211_X1 U18580 ( .C1(n15189), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15188), .B(n15187), .ZN(n15193) );
  NAND2_X1 U18581 ( .A1(n15191), .A2(n15190), .ZN(n15192) );
  OAI211_X1 U18582 ( .C1(n15194), .C2(n20446), .A(n15193), .B(n15192), .ZN(
        P1_U3004) );
  NAND3_X1 U18583 ( .A1(n16303), .A2(n15195), .A3(n15205), .ZN(n15210) );
  NAND2_X1 U18584 ( .A1(n15210), .A2(n15206), .ZN(n15202) );
  NAND3_X1 U18585 ( .A1(n16303), .A2(n15197), .A3(n15196), .ZN(n15199) );
  OAI211_X1 U18586 ( .C1(n16407), .C2(n15200), .A(n15199), .B(n15198), .ZN(
        n15201) );
  AOI21_X1 U18587 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15202), .A(
        n15201), .ZN(n15203) );
  OAI21_X1 U18588 ( .B1(n15204), .B2(n20446), .A(n15203), .ZN(P1_U3005) );
  NOR2_X1 U18589 ( .A1(n15206), .A2(n15205), .ZN(n15207) );
  AOI211_X1 U18590 ( .C1(n20451), .C2(n15209), .A(n15208), .B(n15207), .ZN(
        n15211) );
  OAI211_X1 U18591 ( .C1(n15212), .C2(n20446), .A(n15211), .B(n15210), .ZN(
        P1_U3006) );
  NAND2_X1 U18592 ( .A1(n15213), .A2(n20451), .ZN(n15214) );
  OAI211_X1 U18593 ( .C1(n15216), .C2(n16302), .A(n15215), .B(n15214), .ZN(
        n15217) );
  AOI21_X1 U18594 ( .B1(n16303), .B2(n16302), .A(n15217), .ZN(n15218) );
  OAI21_X1 U18595 ( .B1(n15219), .B2(n20446), .A(n15218), .ZN(P1_U3008) );
  OR2_X1 U18596 ( .A1(n16195), .A2(n15220), .ZN(n15222) );
  NAND2_X1 U18597 ( .A1(n16391), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15221) );
  OAI211_X1 U18598 ( .C1(n16407), .C2(n15223), .A(n15222), .B(n15221), .ZN(
        n15233) );
  NAND2_X1 U18599 ( .A1(n15227), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16187) );
  NOR2_X1 U18600 ( .A1(n15224), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16166) );
  INV_X1 U18601 ( .A(n16187), .ZN(n15225) );
  OR2_X1 U18602 ( .A1(n16166), .A2(n15225), .ZN(n15229) );
  OR2_X1 U18603 ( .A1(n15227), .A2(n15226), .ZN(n15228) );
  NAND2_X1 U18604 ( .A1(n15061), .A2(n15228), .ZN(n16164) );
  MUX2_X1 U18605 ( .A(n16187), .B(n15229), .S(n16164), .Z(n15231) );
  INV_X1 U18606 ( .A(n16166), .ZN(n15230) );
  AND2_X1 U18607 ( .A1(n15231), .A2(n16189), .ZN(n16262) );
  NOR2_X1 U18608 ( .A1(n16262), .A2(n20446), .ZN(n15232) );
  AOI211_X1 U18609 ( .C1(n16186), .C2(n15220), .A(n15233), .B(n15232), .ZN(
        n15234) );
  INV_X1 U18610 ( .A(n15234), .ZN(P1_U3012) );
  AOI21_X1 U18611 ( .B1(n15237), .B2(n15236), .A(n15235), .ZN(n15239) );
  NOR2_X1 U18612 ( .A1(n15239), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15238) );
  MUX2_X1 U18613 ( .A(n15239), .B(n15238), .S(n16163), .Z(n15240) );
  XNOR2_X1 U18614 ( .A(n15240), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16273) );
  AOI22_X1 U18615 ( .A1(n16210), .A2(n20451), .B1(n16391), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n15250) );
  OAI21_X1 U18616 ( .B1(n16374), .B2(n15241), .A(n15261), .ZN(n15242) );
  INV_X1 U18617 ( .A(n15242), .ZN(n15243) );
  OAI21_X1 U18618 ( .B1(n15244), .B2(n16371), .A(n15243), .ZN(n16363) );
  AOI21_X1 U18619 ( .B1(n16347), .B2(n15245), .A(n16363), .ZN(n16329) );
  OAI21_X1 U18620 ( .B1(n15282), .B2(n15246), .A(n16329), .ZN(n16321) );
  NAND2_X1 U18621 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16333) );
  INV_X1 U18622 ( .A(n16334), .ZN(n16344) );
  OAI21_X1 U18623 ( .B1(n16333), .B2(n16344), .A(n15247), .ZN(n15248) );
  NAND2_X1 U18624 ( .A1(n16321), .A2(n15248), .ZN(n15249) );
  OAI211_X1 U18625 ( .C1(n16273), .C2(n20446), .A(n15250), .B(n15249), .ZN(
        P1_U3014) );
  XNOR2_X1 U18626 ( .A(n15251), .B(n15266), .ZN(n15254) );
  NOR2_X1 U18627 ( .A1(n15252), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15253) );
  MUX2_X1 U18628 ( .A(n15254), .B(n15253), .S(n15227), .Z(n15256) );
  OR2_X1 U18629 ( .A1(n15256), .A2(n15255), .ZN(n16290) );
  INV_X1 U18630 ( .A(n16374), .ZN(n15259) );
  INV_X1 U18631 ( .A(n15257), .ZN(n15265) );
  INV_X1 U18632 ( .A(n15258), .ZN(n15264) );
  AOI211_X1 U18633 ( .C1(n15260), .C2(n15259), .A(n15265), .B(n15264), .ZN(
        n15262) );
  OAI21_X1 U18634 ( .B1(n15282), .B2(n15262), .A(n15261), .ZN(n15274) );
  NOR2_X1 U18635 ( .A1(n15264), .A2(n15263), .ZN(n16399) );
  INV_X1 U18636 ( .A(n16399), .ZN(n16383) );
  NOR2_X1 U18637 ( .A1(n15265), .A2(n16383), .ZN(n16345) );
  AOI21_X1 U18638 ( .B1(n15266), .B2(n15275), .A(n16346), .ZN(n15267) );
  AOI22_X1 U18639 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15274), .B1(
        n16345), .B2(n15267), .ZN(n15271) );
  INV_X1 U18640 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15268) );
  OAI22_X1 U18641 ( .A1(n16407), .A2(n16236), .B1(n16406), .B2(n15268), .ZN(
        n15269) );
  INV_X1 U18642 ( .A(n15269), .ZN(n15270) );
  OAI211_X1 U18643 ( .C1(n16290), .C2(n20446), .A(n15271), .B(n15270), .ZN(
        P1_U3021) );
  OAI22_X1 U18644 ( .A1(n16407), .A2(n15272), .B1(n20972), .B2(n16406), .ZN(
        n15273) );
  AOI21_X1 U18645 ( .B1(n15274), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15273), .ZN(n15277) );
  NAND2_X1 U18646 ( .A1(n16345), .A2(n15275), .ZN(n15276) );
  OAI211_X1 U18647 ( .C1(n15278), .C2(n20446), .A(n15277), .B(n15276), .ZN(
        P1_U3022) );
  AOI21_X1 U18648 ( .B1(n15281), .B2(n15280), .A(n15279), .ZN(n16415) );
  OAI21_X1 U18649 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15282), .A(
        n16415), .ZN(n16395) );
  AOI211_X1 U18650 ( .C1(n15284), .C2(n15283), .A(n16414), .B(n16383), .ZN(
        n15286) );
  NAND2_X1 U18651 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15285) );
  AOI22_X1 U18652 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16395), .B1(
        n15286), .B2(n15285), .ZN(n15294) );
  NAND2_X1 U18653 ( .A1(n16405), .A2(n15287), .ZN(n15289) );
  NAND2_X1 U18654 ( .A1(n15289), .A2(n15288), .ZN(n15291) );
  AND2_X1 U18655 ( .A1(n15291), .A2(n15290), .ZN(n20376) );
  AOI21_X1 U18656 ( .B1(n20451), .B2(n20376), .A(n15292), .ZN(n15293) );
  OAI211_X1 U18657 ( .C1(n20446), .C2(n15295), .A(n15294), .B(n15293), .ZN(
        P1_U3023) );
  OAI21_X1 U18658 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21021), .A(n20551), 
        .ZN(n15297) );
  OAI21_X1 U18659 ( .B1(n21025), .B2(n20693), .A(n15297), .ZN(n15298) );
  MUX2_X1 U18660 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15298), .S(
        n21032), .Z(P1_U3477) );
  INV_X1 U18661 ( .A(n15312), .ZN(n15308) );
  INV_X1 U18662 ( .A(n13358), .ZN(n15299) );
  NAND2_X1 U18663 ( .A1(n15300), .A2(n15299), .ZN(n15307) );
  AOI22_X1 U18664 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n15301), .B2(n12852), .ZN(
        n15311) );
  NOR2_X1 U18665 ( .A1(n15302), .A2(n15307), .ZN(n15303) );
  AOI211_X1 U18666 ( .C1(n11995), .C2(n15305), .A(n15304), .B(n15303), .ZN(
        n16130) );
  OAI222_X1 U18667 ( .A1(n15308), .A2(n15307), .B1(n15311), .B2(n15306), .C1(
        n15315), .C2(n16130), .ZN(n15309) );
  MUX2_X1 U18668 ( .A(n15309), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15317), .Z(P1_U3473) );
  AOI22_X1 U18669 ( .A1(n15313), .A2(n15312), .B1(n15311), .B2(n15310), .ZN(
        n15314) );
  OAI21_X1 U18670 ( .B1(n15316), .B2(n15315), .A(n15314), .ZN(n15319) );
  MUX2_X1 U18671 ( .A(n15319), .B(n15318), .S(n15317), .Z(P1_U3472) );
  NOR2_X1 U18672 ( .A1(n20835), .A2(n20883), .ZN(n15323) );
  INV_X1 U18673 ( .A(n15320), .ZN(n15321) );
  NOR2_X1 U18674 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20883), .ZN(n20725) );
  AOI21_X1 U18675 ( .B1(n15323), .B2(n20841), .A(n20725), .ZN(n15327) );
  OR2_X1 U18676 ( .A1(n20876), .A2(n11995), .ZN(n15328) );
  NAND2_X1 U18677 ( .A1(n20461), .A2(n20753), .ZN(n20694) );
  NAND2_X1 U18678 ( .A1(n15325), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20845) );
  OAI22_X1 U18679 ( .A1(n15327), .A2(n15328), .B1(n20694), .B2(n20845), .ZN(
        n20837) );
  INV_X1 U18680 ( .A(n20837), .ZN(n15345) );
  NOR2_X1 U18681 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15324), .ZN(
        n20836) );
  NOR2_X1 U18682 ( .A1(n15325), .A2(n21042), .ZN(n20755) );
  INV_X1 U18683 ( .A(n15327), .ZN(n15329) );
  AOI22_X1 U18684 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20694), .B1(n15329), 
        .B2(n15328), .ZN(n15330) );
  OAI211_X1 U18685 ( .C1(n20836), .C2(n20760), .A(n20849), .B(n15330), .ZN(
        n20838) );
  AOI22_X1 U18686 ( .A1(n20835), .A2(n20757), .B1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n20838), .ZN(n15331) );
  OAI21_X1 U18687 ( .B1(n20841), .B2(n9806), .A(n15331), .ZN(n15332) );
  AOI21_X1 U18688 ( .B1(n20836), .B2(n20881), .A(n15332), .ZN(n15333) );
  OAI21_X1 U18689 ( .B1(n15345), .B2(n20767), .A(n15333), .ZN(P1_U3129) );
  AOI22_X1 U18690 ( .A1(n20835), .A2(n20771), .B1(
        P1_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n20838), .ZN(n15334) );
  OAI21_X1 U18691 ( .B1(n20841), .B2(n9812), .A(n15334), .ZN(n15335) );
  AOI21_X1 U18692 ( .B1(n20836), .B2(n20902), .A(n15335), .ZN(n15336) );
  OAI21_X1 U18693 ( .B1(n15345), .B2(n20774), .A(n15336), .ZN(P1_U3131) );
  NAND2_X1 U18694 ( .A1(n20464), .A2(n15337), .ZN(n20781) );
  NOR2_X2 U18695 ( .A1(n15339), .A2(n15338), .ZN(n20914) );
  INV_X1 U18696 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16765) );
  INV_X1 U18697 ( .A(DATAI_28_), .ZN(n21068) );
  INV_X1 U18698 ( .A(n20915), .ZN(n20739) );
  INV_X1 U18699 ( .A(DATAI_20_), .ZN(n21225) );
  OAI22_X1 U18700 ( .A1(n16779), .A2(n15341), .B1(n21225), .B2(n15340), .ZN(
        n20778) );
  AOI22_X1 U18701 ( .A1(n20835), .A2(n20778), .B1(
        P1_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n20838), .ZN(n15342) );
  OAI21_X1 U18702 ( .B1(n20841), .B2(n20739), .A(n15342), .ZN(n15343) );
  AOI21_X1 U18703 ( .B1(n20836), .B2(n20914), .A(n15343), .ZN(n15344) );
  OAI21_X1 U18704 ( .B1(n15345), .B2(n20781), .A(n15344), .ZN(P1_U3133) );
  INV_X1 U18705 ( .A(n20914), .ZN(n15352) );
  NAND2_X1 U18706 ( .A1(n15346), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n15351) );
  OAI22_X1 U18707 ( .A1(n15348), .A2(n20739), .B1(n20781), .B2(n15347), .ZN(
        n15349) );
  AOI21_X1 U18708 ( .B1(n20870), .B2(n20778), .A(n15349), .ZN(n15350) );
  OAI211_X1 U18709 ( .C1(n15353), .C2(n15352), .A(n15351), .B(n15350), .ZN(
        P1_U3141) );
  OR2_X1 U18710 ( .A1(n15399), .A2(n15354), .ZN(n15355) );
  NAND2_X1 U18711 ( .A1(n15356), .A2(n15355), .ZN(n15777) );
  OR2_X1 U18712 ( .A1(n15488), .A2(n15357), .ZN(n15358) );
  NAND2_X1 U18713 ( .A1(n12826), .A2(n15358), .ZN(n15779) );
  AOI22_X1 U18714 ( .A1(n15359), .A2(n12839), .B1(P2_REIP_REG_29__SCAN_IN), 
        .B2(n19402), .ZN(n15361) );
  AOI22_X1 U18715 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19406), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19431), .ZN(n15360) );
  OAI211_X1 U18716 ( .C1(n15779), .C2(n19408), .A(n15361), .B(n15360), .ZN(
        n15364) );
  AOI211_X1 U18717 ( .C1(n9771), .C2(n15627), .A(n15365), .B(n19394), .ZN(
        n15366) );
  INV_X1 U18718 ( .A(n15366), .ZN(n15375) );
  OR2_X1 U18719 ( .A1(n15433), .A2(n15367), .ZN(n15368) );
  AND2_X1 U18720 ( .A1(n15415), .A2(n15368), .ZN(n15837) );
  OR2_X1 U18721 ( .A1(n15527), .A2(n15369), .ZN(n15370) );
  NAND2_X1 U18722 ( .A1(n15511), .A2(n15370), .ZN(n15835) );
  AOI22_X1 U18723 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19431), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19406), .ZN(n15372) );
  NAND2_X1 U18724 ( .A1(n19402), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15371) );
  OAI211_X1 U18725 ( .C1(n19408), .C2(n15835), .A(n15372), .B(n15371), .ZN(
        n15373) );
  AOI21_X1 U18726 ( .B1(n15837), .B2(n19425), .A(n15373), .ZN(n15374) );
  OAI211_X1 U18727 ( .C1(n19423), .C2(n15376), .A(n15375), .B(n15374), .ZN(
        P2_U2830) );
  NOR2_X1 U18728 ( .A1(n19289), .A2(n19393), .ZN(n15377) );
  XNOR2_X1 U18729 ( .A(n15377), .B(n15697), .ZN(n15378) );
  NAND2_X1 U18730 ( .A1(n15378), .A2(n19411), .ZN(n15389) );
  OR2_X1 U18731 ( .A1(n15381), .A2(n15380), .ZN(n15382) );
  AND2_X1 U18732 ( .A1(n15379), .A2(n15382), .ZN(n16486) );
  AOI22_X1 U18733 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19431), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19406), .ZN(n15383) );
  OAI211_X1 U18734 ( .C1(n19416), .C2(n15696), .A(n15383), .B(n19364), .ZN(
        n15387) );
  OAI21_X1 U18735 ( .B1(n15475), .B2(n15385), .A(n15384), .ZN(n15929) );
  NOR2_X1 U18736 ( .A1(n15929), .A2(n19389), .ZN(n15386) );
  AOI211_X1 U18737 ( .C1(n19420), .C2(n16486), .A(n15387), .B(n15386), .ZN(
        n15388) );
  OAI211_X1 U18738 ( .C1(n19423), .C2(n15390), .A(n15389), .B(n15388), .ZN(
        P2_U2837) );
  MUX2_X1 U18739 ( .A(n15757), .B(P2_EBX_REG_31__SCAN_IN), .S(n15448), .Z(
        P2_U2856) );
  NAND2_X1 U18740 ( .A1(n15391), .A2(n15392), .ZN(n15481) );
  NAND3_X1 U18741 ( .A1(n9715), .A2(n15470), .A3(n15481), .ZN(n15394) );
  NAND2_X1 U18742 ( .A1(n15448), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15393) );
  OAI211_X1 U18743 ( .C1(n15777), .C2(n15448), .A(n15394), .B(n15393), .ZN(
        P2_U2858) );
  NAND2_X1 U18744 ( .A1(n15396), .A2(n15395), .ZN(n15398) );
  XNOR2_X1 U18745 ( .A(n15398), .B(n15397), .ZN(n15497) );
  INV_X1 U18746 ( .A(n15399), .ZN(n15402) );
  OR2_X1 U18747 ( .A1(n15406), .A2(n15400), .ZN(n15401) );
  NOR2_X1 U18748 ( .A1(n16423), .A2(n15448), .ZN(n15403) );
  AOI21_X1 U18749 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15448), .A(n15403), .ZN(
        n15404) );
  OAI21_X1 U18750 ( .B1(n15497), .B2(n15479), .A(n15404), .ZN(P2_U2859) );
  AND2_X1 U18751 ( .A1(n15413), .A2(n15405), .ZN(n15407) );
  OR2_X1 U18752 ( .A1(n15407), .A2(n15406), .ZN(n16442) );
  AOI21_X1 U18753 ( .B1(n15410), .B2(n15409), .A(n15408), .ZN(n15498) );
  NAND2_X1 U18754 ( .A1(n15498), .A2(n15470), .ZN(n15412) );
  NAND2_X1 U18755 ( .A1(n15448), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15411) );
  OAI211_X1 U18756 ( .C1(n16442), .C2(n15448), .A(n15412), .B(n15411), .ZN(
        P2_U2860) );
  INV_X1 U18757 ( .A(n15413), .ZN(n15414) );
  AOI21_X1 U18758 ( .B1(n15416), .B2(n15415), .A(n15414), .ZN(n16455) );
  INV_X1 U18759 ( .A(n16455), .ZN(n15827) );
  AOI21_X1 U18760 ( .B1(n15417), .B2(n15419), .A(n15418), .ZN(n15509) );
  NAND2_X1 U18761 ( .A1(n15509), .A2(n15470), .ZN(n15421) );
  NAND2_X1 U18762 ( .A1(n15448), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15420) );
  OAI211_X1 U18763 ( .C1(n15827), .C2(n15448), .A(n15421), .B(n15420), .ZN(
        P2_U2861) );
  OAI21_X1 U18764 ( .B1(n15422), .B2(n15424), .A(n15423), .ZN(n15524) );
  NAND2_X1 U18765 ( .A1(n15448), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15426) );
  NAND2_X1 U18766 ( .A1(n15837), .A2(n15449), .ZN(n15425) );
  OAI211_X1 U18767 ( .C1(n15524), .C2(n15479), .A(n15426), .B(n15425), .ZN(
        P2_U2862) );
  AOI21_X1 U18768 ( .B1(n9768), .B2(n15428), .A(n15427), .ZN(n15429) );
  XOR2_X1 U18769 ( .A(n15430), .B(n15429), .Z(n15532) );
  AND2_X1 U18770 ( .A1(n15432), .A2(n15431), .ZN(n15434) );
  OR2_X1 U18771 ( .A1(n15434), .A2(n15433), .ZN(n16469) );
  NOR2_X1 U18772 ( .A1(n16469), .A2(n15448), .ZN(n15435) );
  AOI21_X1 U18773 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15448), .A(n15435), .ZN(
        n15436) );
  OAI21_X1 U18774 ( .B1(n15532), .B2(n15479), .A(n15436), .ZN(P2_U2863) );
  AOI21_X1 U18775 ( .B1(n15439), .B2(n15438), .A(n15437), .ZN(n15533) );
  NAND2_X1 U18776 ( .A1(n15533), .A2(n15470), .ZN(n15441) );
  NAND2_X1 U18777 ( .A1(n15448), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15440) );
  OAI211_X1 U18778 ( .C1(n15862), .C2(n15448), .A(n15441), .B(n15440), .ZN(
        P2_U2864) );
  OAI21_X1 U18779 ( .B1(n15442), .B2(n15443), .A(n14457), .ZN(n15547) );
  NAND2_X1 U18780 ( .A1(n15448), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15445) );
  NAND2_X1 U18781 ( .A1(n16492), .A2(n15449), .ZN(n15444) );
  OAI211_X1 U18782 ( .C1(n15547), .C2(n15479), .A(n15445), .B(n15444), .ZN(
        P2_U2865) );
  AOI21_X1 U18783 ( .B1(n15446), .B2(n9680), .A(n15442), .ZN(n15447) );
  INV_X1 U18784 ( .A(n15447), .ZN(n15554) );
  NAND2_X1 U18785 ( .A1(n15448), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U18786 ( .A1(n15891), .A2(n15449), .ZN(n15450) );
  OAI211_X1 U18787 ( .C1(n15554), .C2(n15479), .A(n15451), .B(n15450), .ZN(
        P2_U2866) );
  NAND2_X1 U18788 ( .A1(n15464), .A2(n15452), .ZN(n15453) );
  NAND2_X1 U18789 ( .A1(n15454), .A2(n15453), .ZN(n15911) );
  NAND2_X1 U18790 ( .A1(n15455), .A2(n15456), .ZN(n15457) );
  AND2_X1 U18791 ( .A1(n9680), .A2(n15457), .ZN(n16480) );
  NAND2_X1 U18792 ( .A1(n16480), .A2(n15470), .ZN(n15459) );
  NAND2_X1 U18793 ( .A1(n15448), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15458) );
  OAI211_X1 U18794 ( .C1(n15911), .C2(n15448), .A(n15459), .B(n15458), .ZN(
        P2_U2867) );
  OAI21_X1 U18795 ( .B1(n15460), .B2(n15461), .A(n15455), .ZN(n15565) );
  NAND2_X1 U18796 ( .A1(n15384), .A2(n15462), .ZN(n15463) );
  NAND2_X1 U18797 ( .A1(n15464), .A2(n15463), .ZN(n19273) );
  NOR2_X1 U18798 ( .A1(n19273), .A2(n15448), .ZN(n15465) );
  AOI21_X1 U18799 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15448), .A(n15465), .ZN(
        n15466) );
  OAI21_X1 U18800 ( .B1(n15565), .B2(n15479), .A(n15466), .ZN(P2_U2868) );
  INV_X1 U18801 ( .A(n15467), .ZN(n15469) );
  AOI21_X1 U18802 ( .B1(n15469), .B2(n15468), .A(n15460), .ZN(n16487) );
  NAND2_X1 U18803 ( .A1(n16487), .A2(n15470), .ZN(n15472) );
  NAND2_X1 U18804 ( .A1(n15448), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15471) );
  OAI211_X1 U18805 ( .C1(n15929), .C2(n15448), .A(n15472), .B(n15471), .ZN(
        P2_U2869) );
  AND2_X1 U18806 ( .A1(n15474), .A2(n15473), .ZN(n15476) );
  OR2_X1 U18807 ( .A1(n15476), .A2(n15475), .ZN(n19286) );
  NOR2_X1 U18808 ( .A1(n19286), .A2(n15448), .ZN(n15477) );
  AOI21_X1 U18809 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15448), .A(n15477), .ZN(
        n15478) );
  OAI21_X1 U18810 ( .B1(n15480), .B2(n15479), .A(n15478), .ZN(P2_U2870) );
  NAND3_X1 U18811 ( .A1(n9715), .A2(n19497), .A3(n15481), .ZN(n15487) );
  INV_X1 U18812 ( .A(n15779), .ZN(n15484) );
  OAI22_X1 U18813 ( .A1(n15558), .A2(n19446), .B1(n19466), .B2(n15482), .ZN(
        n15483) );
  AOI21_X1 U18814 ( .B1(n19495), .B2(n15484), .A(n15483), .ZN(n15486) );
  AOI22_X1 U18815 ( .A1(n19436), .A2(BUF1_REG_29__SCAN_IN), .B1(n19438), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15485) );
  NAND3_X1 U18816 ( .A1(n15487), .A2(n15486), .A3(n15485), .ZN(P2_U2890) );
  INV_X1 U18817 ( .A(n15488), .ZN(n15491) );
  NAND2_X1 U18818 ( .A1(n15501), .A2(n15489), .ZN(n15490) );
  NAND2_X1 U18819 ( .A1(n15491), .A2(n15490), .ZN(n16422) );
  INV_X1 U18820 ( .A(n16422), .ZN(n15494) );
  OAI22_X1 U18821 ( .A1(n15558), .A2(n19449), .B1(n19466), .B2(n15492), .ZN(
        n15493) );
  AOI21_X1 U18822 ( .B1(n15494), .B2(n19495), .A(n15493), .ZN(n15496) );
  AOI22_X1 U18823 ( .A1(n19436), .A2(BUF1_REG_28__SCAN_IN), .B1(n19438), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15495) );
  OAI211_X1 U18824 ( .C1(n15497), .C2(n19490), .A(n15496), .B(n15495), .ZN(
        P2_U2891) );
  INV_X1 U18825 ( .A(n15498), .ZN(n15508) );
  NAND2_X1 U18826 ( .A1(n15513), .A2(n15499), .ZN(n15500) );
  NAND2_X1 U18827 ( .A1(n15501), .A2(n15500), .ZN(n16449) );
  INV_X1 U18828 ( .A(n16449), .ZN(n15506) );
  OAI22_X1 U18829 ( .A1(n15558), .A2(n19451), .B1(n19466), .B2(n15502), .ZN(
        n15505) );
  INV_X1 U18830 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15503) );
  OAI22_X1 U18831 ( .A1(n15561), .A2(n19586), .B1(n15560), .B2(n15503), .ZN(
        n15504) );
  AOI211_X1 U18832 ( .C1(n19495), .C2(n15506), .A(n15505), .B(n15504), .ZN(
        n15507) );
  OAI21_X1 U18833 ( .B1(n15508), .B2(n19490), .A(n15507), .ZN(P2_U2892) );
  NAND2_X1 U18834 ( .A1(n15509), .A2(n19497), .ZN(n15517) );
  INV_X1 U18835 ( .A(n15558), .ZN(n16485) );
  AOI22_X1 U18836 ( .A1(n16485), .A2(n19453), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19494), .ZN(n15516) );
  AOI22_X1 U18837 ( .A1(n19436), .A2(BUF1_REG_26__SCAN_IN), .B1(n19438), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15515) );
  NAND2_X1 U18838 ( .A1(n15511), .A2(n15510), .ZN(n15512) );
  AND2_X1 U18839 ( .A1(n15513), .A2(n15512), .ZN(n16462) );
  NAND2_X1 U18840 ( .A1(n19495), .A2(n16462), .ZN(n15514) );
  NAND4_X1 U18841 ( .A1(n15517), .A2(n15516), .A3(n15515), .A4(n15514), .ZN(
        P2_U2893) );
  INV_X1 U18842 ( .A(n15835), .ZN(n15522) );
  OAI22_X1 U18843 ( .A1(n15558), .A2(n19456), .B1(n19466), .B2(n15518), .ZN(
        n15521) );
  INV_X1 U18844 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n15519) );
  OAI22_X1 U18845 ( .A1(n15561), .A2(n16770), .B1(n15560), .B2(n15519), .ZN(
        n15520) );
  AOI211_X1 U18846 ( .C1(n19495), .C2(n15522), .A(n15521), .B(n15520), .ZN(
        n15523) );
  OAI21_X1 U18847 ( .B1(n15524), .B2(n19490), .A(n15523), .ZN(P2_U2894) );
  AND2_X1 U18848 ( .A1(n9777), .A2(n15525), .ZN(n15526) );
  NOR2_X1 U18849 ( .A1(n15527), .A2(n15526), .ZN(n16467) );
  INV_X1 U18850 ( .A(n19460), .ZN(n15528) );
  OAI22_X1 U18851 ( .A1(n15558), .A2(n15528), .B1(n19466), .B2(n13245), .ZN(
        n15529) );
  AOI21_X1 U18852 ( .B1(n19495), .B2(n16467), .A(n15529), .ZN(n15531) );
  AOI22_X1 U18853 ( .A1(n19436), .A2(BUF1_REG_24__SCAN_IN), .B1(n19438), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n15530) );
  OAI211_X1 U18854 ( .C1(n15532), .C2(n19490), .A(n15531), .B(n15530), .ZN(
        P2_U2895) );
  INV_X1 U18855 ( .A(n15533), .ZN(n15540) );
  INV_X1 U18856 ( .A(n15859), .ZN(n15538) );
  OAI22_X1 U18857 ( .A1(n15558), .A2(n19616), .B1(n15534), .B2(n19466), .ZN(
        n15537) );
  INV_X1 U18858 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15535) );
  OAI22_X1 U18859 ( .A1(n15561), .A2(n16774), .B1(n15560), .B2(n15535), .ZN(
        n15536) );
  AOI211_X1 U18860 ( .C1(n19495), .C2(n15538), .A(n15537), .B(n15536), .ZN(
        n15539) );
  OAI21_X1 U18861 ( .B1(n15540), .B2(n19490), .A(n15539), .ZN(P2_U2896) );
  INV_X1 U18862 ( .A(n15878), .ZN(n15545) );
  OAI22_X1 U18863 ( .A1(n15558), .A2(n19604), .B1(n19466), .B2(n15541), .ZN(
        n15544) );
  INV_X1 U18864 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n15542) );
  OAI22_X1 U18865 ( .A1(n15561), .A2(n16776), .B1(n15560), .B2(n15542), .ZN(
        n15543) );
  AOI211_X1 U18866 ( .C1(n19495), .C2(n15545), .A(n15544), .B(n15543), .ZN(
        n15546) );
  OAI21_X1 U18867 ( .B1(n15547), .B2(n19490), .A(n15546), .ZN(P2_U2897) );
  INV_X1 U18868 ( .A(n15886), .ZN(n15552) );
  OAI22_X1 U18869 ( .A1(n15558), .A2(n19598), .B1(n15548), .B2(n19466), .ZN(
        n15551) );
  AOI22_X1 U18870 ( .A1(n19436), .A2(BUF1_REG_21__SCAN_IN), .B1(n19438), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15549) );
  INV_X1 U18871 ( .A(n15549), .ZN(n15550) );
  AOI211_X1 U18872 ( .C1(n15552), .C2(n19495), .A(n15551), .B(n15550), .ZN(
        n15553) );
  OAI21_X1 U18873 ( .B1(n15554), .B2(n19490), .A(n15553), .ZN(P2_U2898) );
  NAND2_X1 U18874 ( .A1(n15379), .A2(n15555), .ZN(n15556) );
  NAND2_X1 U18875 ( .A1(n15905), .A2(n15556), .ZN(n19280) );
  INV_X1 U18876 ( .A(n19280), .ZN(n15918) );
  OAI22_X1 U18877 ( .A1(n15558), .A2(n19587), .B1(n15557), .B2(n19466), .ZN(
        n15563) );
  INV_X1 U18878 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15559) );
  OAI22_X1 U18879 ( .A1(n15561), .A2(n16781), .B1(n15560), .B2(n15559), .ZN(
        n15562) );
  AOI211_X1 U18880 ( .C1(n19495), .C2(n15918), .A(n15563), .B(n15562), .ZN(
        n15564) );
  OAI21_X1 U18881 ( .B1(n15565), .B2(n19490), .A(n15564), .ZN(P2_U2900) );
  NAND2_X1 U18882 ( .A1(n15566), .A2(n15581), .ZN(n15571) );
  INV_X1 U18883 ( .A(n15567), .ZN(n15568) );
  NOR2_X1 U18884 ( .A1(n15569), .A2(n15568), .ZN(n15570) );
  XNOR2_X1 U18885 ( .A(n15571), .B(n15570), .ZN(n15775) );
  XOR2_X1 U18886 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15584), .Z(
        n15773) );
  INV_X1 U18887 ( .A(n15573), .ZN(n15575) );
  NOR2_X1 U18888 ( .A1(n19364), .A2(n20174), .ZN(n15767) );
  AOI21_X1 U18889 ( .B1(n19551), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15767), .ZN(n15574) );
  INV_X1 U18890 ( .A(n15577), .ZN(n15578) );
  AOI21_X1 U18891 ( .B1(n15773), .B2(n19554), .A(n15578), .ZN(n15579) );
  OAI21_X1 U18892 ( .B1(n15775), .B2(n16586), .A(n15579), .ZN(P2_U2984) );
  NAND2_X1 U18893 ( .A1(n15581), .A2(n15580), .ZN(n15583) );
  XOR2_X1 U18894 ( .A(n15583), .B(n15582), .Z(n15791) );
  OR2_X1 U18895 ( .A1(n19333), .A2(n20171), .ZN(n15778) );
  OAI21_X1 U18896 ( .B1(n16593), .B2(n15586), .A(n15778), .ZN(n15587) );
  AOI21_X1 U18897 ( .B1(n16583), .B2(n15588), .A(n15587), .ZN(n15589) );
  OAI21_X1 U18898 ( .B1(n15777), .B2(n19559), .A(n15589), .ZN(n15590) );
  AOI21_X1 U18899 ( .B1(n15789), .B2(n19554), .A(n15590), .ZN(n15591) );
  OAI21_X1 U18900 ( .B1(n15791), .B2(n16586), .A(n15591), .ZN(P2_U2985) );
  NAND2_X1 U18901 ( .A1(n15593), .A2(n15592), .ZN(n15594) );
  INV_X1 U18902 ( .A(n15594), .ZN(n15596) );
  XNOR2_X1 U18903 ( .A(n15594), .B(n15595), .ZN(n15605) );
  NAND2_X1 U18904 ( .A1(n15605), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15805) );
  OAI21_X1 U18905 ( .B1(n15596), .B2(n15595), .A(n15805), .ZN(n15599) );
  XNOR2_X1 U18906 ( .A(n15597), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15598) );
  XNOR2_X1 U18907 ( .A(n15599), .B(n15598), .ZN(n15803) );
  NOR2_X1 U18908 ( .A1(n19364), .A2(n20169), .ZN(n15793) );
  NOR2_X1 U18909 ( .A1(n19564), .A2(n15600), .ZN(n15601) );
  AOI211_X1 U18910 ( .C1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n19551), .A(
        n15793), .B(n15601), .ZN(n15602) );
  OAI21_X1 U18911 ( .B1(n16423), .B2(n19559), .A(n15602), .ZN(n15603) );
  AOI21_X1 U18912 ( .B1(n15801), .B2(n19554), .A(n15603), .ZN(n15604) );
  OAI21_X1 U18913 ( .B1(n15803), .B2(n16586), .A(n15604), .ZN(P2_U2986) );
  NAND2_X1 U18914 ( .A1(n15619), .A2(n15783), .ZN(n15804) );
  NAND2_X1 U18915 ( .A1(n15804), .A2(n19554), .ZN(n15611) );
  OR2_X1 U18916 ( .A1(n15605), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15806) );
  NAND3_X1 U18917 ( .A1(n15806), .A2(n15805), .A3(n19552), .ZN(n15610) );
  OR2_X1 U18918 ( .A1(n19364), .A2(n20168), .ZN(n15807) );
  OAI21_X1 U18919 ( .B1(n16593), .B2(n15606), .A(n15807), .ZN(n15608) );
  NOR2_X1 U18920 ( .A1(n16442), .A2(n19559), .ZN(n15607) );
  AOI211_X1 U18921 ( .C1(n16583), .C2(n16445), .A(n15608), .B(n15607), .ZN(
        n15609) );
  OAI211_X1 U18922 ( .C1(n15817), .C2(n15611), .A(n15610), .B(n15609), .ZN(
        P2_U2987) );
  NOR2_X1 U18923 ( .A1(n15612), .A2(n15624), .ZN(n15613) );
  XOR2_X1 U18924 ( .A(n15614), .B(n15613), .Z(n15832) );
  NOR2_X1 U18925 ( .A1(n19364), .A2(n15615), .ZN(n15824) );
  AOI21_X1 U18926 ( .B1(n19551), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15824), .ZN(n15616) );
  OAI21_X1 U18927 ( .B1(n19564), .B2(n15617), .A(n15616), .ZN(n15621) );
  NOR2_X1 U18928 ( .A1(n15818), .A2(n16584), .ZN(n15620) );
  OAI21_X1 U18929 ( .B1(n15832), .B2(n16586), .A(n15622), .ZN(P2_U2988) );
  NOR2_X1 U18930 ( .A1(n15624), .A2(n15623), .ZN(n15626) );
  XOR2_X1 U18931 ( .A(n15626), .B(n15625), .Z(n15845) );
  NAND2_X1 U18932 ( .A1(n16583), .A2(n15627), .ZN(n15628) );
  OR2_X1 U18933 ( .A1(n19333), .A2(n20164), .ZN(n15834) );
  OAI211_X1 U18934 ( .C1(n15629), .C2(n16593), .A(n15628), .B(n15834), .ZN(
        n15632) );
  INV_X1 U18935 ( .A(n15630), .ZN(n15637) );
  NOR2_X1 U18936 ( .A1(n15637), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15833) );
  NOR3_X1 U18937 ( .A1(n15833), .A2(n15618), .A3(n16584), .ZN(n15631) );
  AOI211_X1 U18938 ( .C1(n16589), .C2(n15837), .A(n15632), .B(n15631), .ZN(
        n15633) );
  OAI21_X1 U18939 ( .B1(n16586), .B2(n15845), .A(n15633), .ZN(P2_U2989) );
  XNOR2_X1 U18940 ( .A(n15634), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15635) );
  XNOR2_X1 U18941 ( .A(n15636), .B(n15635), .ZN(n15854) );
  AOI21_X1 U18942 ( .B1(n15819), .B2(n9946), .A(n15637), .ZN(n15852) );
  NOR2_X1 U18943 ( .A1(n19364), .A2(n20162), .ZN(n15848) );
  AOI21_X1 U18944 ( .B1(n19551), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15848), .ZN(n15639) );
  NAND2_X1 U18945 ( .A1(n16583), .A2(n16473), .ZN(n15638) );
  OAI211_X1 U18946 ( .C1(n16469), .C2(n19559), .A(n15639), .B(n15638), .ZN(
        n15640) );
  AOI21_X1 U18947 ( .B1(n15852), .B2(n19554), .A(n15640), .ZN(n15641) );
  OAI21_X1 U18948 ( .B1(n15854), .B2(n16586), .A(n15641), .ZN(P2_U2990) );
  XNOR2_X1 U18949 ( .A(n15643), .B(n15642), .ZN(n15867) );
  AOI21_X1 U18950 ( .B1(n15855), .B2(n15868), .A(n15644), .ZN(n15865) );
  OR2_X1 U18951 ( .A1(n19333), .A2(n20160), .ZN(n15857) );
  OAI21_X1 U18952 ( .B1(n16593), .B2(n15645), .A(n15857), .ZN(n15646) );
  AOI21_X1 U18953 ( .B1(n16583), .B2(n15647), .A(n15646), .ZN(n15648) );
  OAI21_X1 U18954 ( .B1(n15862), .B2(n19559), .A(n15648), .ZN(n15649) );
  AOI21_X1 U18955 ( .B1(n15865), .B2(n19554), .A(n15649), .ZN(n15650) );
  OAI21_X1 U18956 ( .B1(n15867), .B2(n16586), .A(n15650), .ZN(P2_U2991) );
  NAND2_X1 U18957 ( .A1(n15652), .A2(n15651), .ZN(n15663) );
  NAND2_X1 U18958 ( .A1(n16523), .A2(n16521), .ZN(n16525) );
  NAND2_X1 U18959 ( .A1(n15656), .A2(n15655), .ZN(n15703) );
  INV_X1 U18960 ( .A(n15656), .ZN(n15657) );
  NOR2_X1 U18961 ( .A1(n15660), .A2(n15659), .ZN(n15673) );
  INV_X1 U18962 ( .A(n15660), .ZN(n15661) );
  NAND2_X1 U18963 ( .A1(n15672), .A2(n15661), .ZN(n15662) );
  XOR2_X1 U18964 ( .A(n15663), .B(n15662), .Z(n15897) );
  NAND2_X1 U18965 ( .A1(n16583), .A2(n15664), .ZN(n15665) );
  NAND2_X1 U18966 ( .A1(n15989), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15887) );
  OAI211_X1 U18967 ( .C1(n15666), .C2(n16593), .A(n15665), .B(n15887), .ZN(
        n15670) );
  NAND2_X1 U18968 ( .A1(n15667), .A2(n10199), .ZN(n15668) );
  NAND2_X1 U18969 ( .A1(n15869), .A2(n15668), .ZN(n15885) );
  NOR2_X1 U18970 ( .A1(n15885), .A2(n16584), .ZN(n15669) );
  AOI211_X1 U18971 ( .C1(n16589), .C2(n15891), .A(n15670), .B(n15669), .ZN(
        n15671) );
  OAI21_X1 U18972 ( .B1(n15897), .B2(n16586), .A(n15671), .ZN(P2_U2993) );
  OAI21_X1 U18973 ( .B1(n9692), .B2(n15673), .A(n15672), .ZN(n15916) );
  INV_X1 U18974 ( .A(n15911), .ZN(n19259) );
  NOR2_X1 U18975 ( .A1(n19364), .A2(n15674), .ZN(n15908) );
  AOI21_X1 U18976 ( .B1(n19551), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15908), .ZN(n15675) );
  OAI21_X1 U18977 ( .B1(n19564), .B2(n15676), .A(n15675), .ZN(n15679) );
  OAI21_X1 U18978 ( .B1(n15677), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15667), .ZN(n15898) );
  NOR2_X1 U18979 ( .A1(n15898), .A2(n16584), .ZN(n15678) );
  AOI211_X1 U18980 ( .C1(n16589), .C2(n19259), .A(n15679), .B(n15678), .ZN(
        n15680) );
  OAI21_X1 U18981 ( .B1(n15916), .B2(n16586), .A(n15680), .ZN(P2_U2994) );
  INV_X1 U18982 ( .A(n15683), .ZN(n15689) );
  AND2_X1 U18983 ( .A1(n15694), .A2(n15899), .ZN(n15684) );
  NOR2_X1 U18984 ( .A1(n15677), .A2(n15684), .ZN(n15925) );
  NAND2_X1 U18985 ( .A1(n19270), .A2(n16583), .ZN(n15686) );
  NOR2_X1 U18986 ( .A1(n19364), .A2(n20154), .ZN(n15917) );
  AOI21_X1 U18987 ( .B1(n19551), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15917), .ZN(n15685) );
  OAI211_X1 U18988 ( .C1(n19273), .C2(n19559), .A(n15686), .B(n15685), .ZN(
        n15687) );
  AOI21_X1 U18989 ( .B1(n15925), .B2(n19554), .A(n15687), .ZN(n15688) );
  OAI21_X1 U18990 ( .B1(n15927), .B2(n16586), .A(n15688), .ZN(P2_U2995) );
  NOR2_X1 U18991 ( .A1(n15690), .A2(n15689), .ZN(n15691) );
  XNOR2_X1 U18992 ( .A(n15692), .B(n15691), .ZN(n15939) );
  NAND2_X1 U18993 ( .A1(n16024), .A2(n15693), .ZN(n15710) );
  INV_X1 U18994 ( .A(n15694), .ZN(n15695) );
  AOI21_X1 U18995 ( .B1(n15934), .B2(n15710), .A(n15695), .ZN(n15937) );
  NOR2_X1 U18996 ( .A1(n19333), .A2(n15696), .ZN(n15931) );
  NOR2_X1 U18997 ( .A1(n15697), .A2(n19564), .ZN(n15698) );
  AOI211_X1 U18998 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19551), .A(
        n15931), .B(n15698), .ZN(n15699) );
  OAI21_X1 U18999 ( .B1(n19559), .B2(n15929), .A(n15699), .ZN(n15700) );
  AOI21_X1 U19000 ( .B1(n15937), .B2(n19554), .A(n15700), .ZN(n15701) );
  OAI21_X1 U19001 ( .B1(n15939), .B2(n16586), .A(n15701), .ZN(P2_U2996) );
  AOI21_X1 U19002 ( .B1(n15704), .B2(n15703), .A(n15702), .ZN(n15953) );
  INV_X1 U19003 ( .A(n19286), .ZN(n15708) );
  NOR2_X1 U19004 ( .A1(n20151), .A2(n19333), .ZN(n15707) );
  INV_X1 U19005 ( .A(n19291), .ZN(n19283) );
  OAI22_X1 U19006 ( .A1(n16593), .A2(n15705), .B1(n19564), .B2(n19283), .ZN(
        n15706) );
  AOI211_X1 U19007 ( .C1(n16589), .C2(n15708), .A(n15707), .B(n15706), .ZN(
        n15712) );
  INV_X1 U19008 ( .A(n15709), .ZN(n15941) );
  NAND2_X1 U19009 ( .A1(n16508), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15979) );
  NOR2_X1 U19010 ( .A1(n15979), .A2(n15958), .ZN(n15943) );
  OAI211_X1 U19011 ( .C1(n15943), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19554), .B(n15710), .ZN(n15711) );
  OAI211_X1 U19012 ( .C1(n15953), .C2(n16586), .A(n15712), .B(n15711), .ZN(
        P2_U2997) );
  XNOR2_X1 U19013 ( .A(n15714), .B(n15713), .ZN(n15961) );
  INV_X1 U19014 ( .A(n19300), .ZN(n15715) );
  NAND2_X1 U19015 ( .A1(n16583), .A2(n15715), .ZN(n15716) );
  NAND2_X1 U19016 ( .A1(n15989), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15954) );
  OAI211_X1 U19017 ( .C1(n10321), .C2(n16593), .A(n15716), .B(n15954), .ZN(
        n15718) );
  AOI211_X1 U19018 ( .C1(n15958), .C2(n15979), .A(n16584), .B(n15943), .ZN(
        n15717) );
  AOI211_X1 U19019 ( .C1(n16589), .C2(n19301), .A(n15718), .B(n15717), .ZN(
        n15719) );
  OAI21_X1 U19020 ( .B1(n16586), .B2(n15961), .A(n15719), .ZN(P2_U2998) );
  INV_X1 U19021 ( .A(n16015), .ZN(n15722) );
  NOR2_X1 U19022 ( .A1(n15722), .A2(n15721), .ZN(n15723) );
  XNOR2_X1 U19023 ( .A(n15720), .B(n15723), .ZN(n16046) );
  OAI22_X1 U19024 ( .A1(n16593), .A2(n15725), .B1(n10567), .B2(n19333), .ZN(
        n15728) );
  AND2_X1 U19025 ( .A1(n16583), .A2(n15726), .ZN(n15727) );
  NOR2_X1 U19026 ( .A1(n15728), .A2(n15727), .ZN(n15729) );
  OAI21_X1 U19027 ( .B1(n16041), .B2(n19559), .A(n15729), .ZN(n15730) );
  AOI21_X1 U19028 ( .B1(n16035), .B2(n19554), .A(n15730), .ZN(n15731) );
  OAI21_X1 U19029 ( .B1(n16046), .B2(n16586), .A(n15731), .ZN(P2_U3007) );
  NOR3_X1 U19030 ( .A1(n15732), .A2(n16055), .A3(n16057), .ZN(n16036) );
  INV_X1 U19031 ( .A(n16036), .ZN(n15733) );
  NAND2_X1 U19032 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16636) );
  NOR3_X1 U19033 ( .A1(n15734), .A2(n15733), .A3(n16636), .ZN(n15735) );
  OR2_X1 U19034 ( .A1(n16609), .A2(n15735), .ZN(n15737) );
  AND2_X1 U19035 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15738) );
  AND2_X1 U19036 ( .A1(n15903), .A2(n15738), .ZN(n15752) );
  AND2_X1 U19037 ( .A1(n15752), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15739) );
  OR2_X1 U19038 ( .A1(n16609), .A2(n15739), .ZN(n15740) );
  AND2_X1 U19039 ( .A1(n16608), .A2(n15740), .ZN(n15893) );
  NOR2_X1 U19040 ( .A1(n15855), .A2(n15882), .ZN(n15753) );
  INV_X1 U19041 ( .A(n15753), .ZN(n15856) );
  AOI21_X1 U19042 ( .B1(n15741), .B2(n15856), .A(n15819), .ZN(n15742) );
  NAND2_X1 U19043 ( .A1(n15893), .A2(n15742), .ZN(n15846) );
  NAND2_X1 U19044 ( .A1(n16608), .A2(n16609), .ZN(n15745) );
  NAND2_X1 U19045 ( .A1(n15846), .A2(n15745), .ZN(n15841) );
  NAND2_X1 U19046 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15743) );
  NAND2_X1 U19047 ( .A1(n15745), .A2(n15743), .ZN(n15744) );
  AND2_X1 U19048 ( .A1(n15841), .A2(n15744), .ZN(n15776) );
  NAND2_X1 U19049 ( .A1(n15745), .A2(n15763), .ZN(n15746) );
  NAND2_X1 U19050 ( .A1(n15776), .A2(n15746), .ZN(n15769) );
  NOR2_X1 U19051 ( .A1(n16609), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15747) );
  OAI21_X1 U19052 ( .B1(n15769), .B2(n15747), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15750) );
  INV_X1 U19053 ( .A(n15748), .ZN(n15749) );
  OAI211_X1 U19054 ( .C1(n19435), .C2(n16624), .A(n15750), .B(n15749), .ZN(
        n15756) );
  NAND2_X1 U19055 ( .A1(n16036), .A2(n15751), .ZN(n16638) );
  NAND2_X1 U19056 ( .A1(n16597), .A2(n15752), .ZN(n15888) );
  NOR2_X1 U19057 ( .A1(n10199), .A2(n15888), .ZN(n15873) );
  NAND2_X1 U19058 ( .A1(n15873), .A2(n15753), .ZN(n15823) );
  INV_X1 U19059 ( .A(n15823), .ZN(n15847) );
  NAND2_X1 U19060 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15822) );
  INV_X1 U19061 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15821) );
  NOR2_X1 U19062 ( .A1(n15822), .A2(n15821), .ZN(n15754) );
  NAND2_X1 U19063 ( .A1(n15847), .A2(n15754), .ZN(n15782) );
  NOR4_X1 U19064 ( .A1(n15782), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15764), .A4(n15763), .ZN(n15755) );
  AOI211_X1 U19065 ( .C1(n16645), .C2(n15757), .A(n15756), .B(n15755), .ZN(
        n15761) );
  INV_X1 U19066 ( .A(n15758), .ZN(n15759) );
  NAND2_X1 U19067 ( .A1(n15759), .A2(n16646), .ZN(n15760) );
  INV_X1 U19068 ( .A(n15763), .ZN(n15765) );
  NAND2_X1 U19069 ( .A1(n15765), .A2(n15764), .ZN(n15771) );
  NAND2_X1 U19070 ( .A1(n15766), .A2(n16645), .ZN(n15770) );
  AOI21_X1 U19071 ( .B1(n15773), .B2(n16646), .A(n15772), .ZN(n15774) );
  OAI21_X1 U19072 ( .B1(n15775), .B2(n16651), .A(n15774), .ZN(P2_U3016) );
  NOR2_X1 U19073 ( .A1(n15782), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15813) );
  INV_X1 U19074 ( .A(n15776), .ZN(n15809) );
  NOR2_X1 U19075 ( .A1(n15813), .A2(n15809), .ZN(n15797) );
  INV_X1 U19076 ( .A(n15777), .ZN(n15781) );
  OAI21_X1 U19077 ( .B1(n16624), .B2(n15779), .A(n15778), .ZN(n15780) );
  AOI21_X1 U19078 ( .B1(n15781), .B2(n16645), .A(n15780), .ZN(n15786) );
  INV_X1 U19079 ( .A(n15782), .ZN(n15795) );
  OAI21_X1 U19080 ( .B1(n15783), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15784) );
  OAI211_X1 U19081 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n15795), .B(n15784), .ZN(
        n15785) );
  OAI211_X1 U19082 ( .C1(n15797), .C2(n15787), .A(n15786), .B(n15785), .ZN(
        n15788) );
  AOI21_X1 U19083 ( .B1(n15789), .B2(n16646), .A(n15788), .ZN(n15790) );
  OAI21_X1 U19084 ( .B1(n15791), .B2(n16651), .A(n15790), .ZN(P2_U3017) );
  INV_X1 U19085 ( .A(n16423), .ZN(n15794) );
  NOR2_X1 U19086 ( .A1(n16624), .A2(n16422), .ZN(n15792) );
  AOI211_X1 U19087 ( .C1(n15794), .C2(n16645), .A(n15793), .B(n15792), .ZN(
        n15799) );
  NAND3_X1 U19088 ( .A1(n15795), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15796), .ZN(n15798) );
  NAND3_X1 U19089 ( .A1(n15799), .A2(n15798), .A3(n10300), .ZN(n15800) );
  OAI21_X1 U19090 ( .B1(n15803), .B2(n16651), .A(n15802), .ZN(P2_U3018) );
  NAND2_X1 U19091 ( .A1(n15804), .A2(n16646), .ZN(n15816) );
  NAND3_X1 U19092 ( .A1(n15806), .A2(n15805), .A3(n16600), .ZN(n15815) );
  OAI21_X1 U19093 ( .B1(n16624), .B2(n16449), .A(n15807), .ZN(n15808) );
  INV_X1 U19094 ( .A(n15808), .ZN(n15811) );
  NAND2_X1 U19095 ( .A1(n15809), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15810) );
  OAI211_X1 U19096 ( .C1(n16442), .C2(n16629), .A(n15811), .B(n15810), .ZN(
        n15812) );
  NOR2_X1 U19097 ( .A1(n15813), .A2(n15812), .ZN(n15814) );
  OAI211_X1 U19098 ( .C1(n15817), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        P2_U3019) );
  INV_X1 U19099 ( .A(n15818), .ZN(n15830) );
  NOR2_X1 U19100 ( .A1(n15819), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15820) );
  NAND2_X1 U19101 ( .A1(n15847), .A2(n15820), .ZN(n15839) );
  AOI21_X1 U19102 ( .B1(n15839), .B2(n15841), .A(n15821), .ZN(n15829) );
  OR3_X1 U19103 ( .A1(n15823), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15822), .ZN(n15826) );
  AOI21_X1 U19104 ( .B1(n16643), .B2(n16462), .A(n15824), .ZN(n15825) );
  OAI211_X1 U19105 ( .C1(n15827), .C2(n16629), .A(n15826), .B(n15825), .ZN(
        n15828) );
  AOI211_X1 U19106 ( .C1(n15830), .C2(n16646), .A(n15829), .B(n15828), .ZN(
        n15831) );
  OAI21_X1 U19107 ( .B1(n15832), .B2(n16651), .A(n15831), .ZN(P2_U3020) );
  NOR3_X1 U19108 ( .A1(n15833), .A2(n15618), .A3(n16630), .ZN(n15843) );
  OAI21_X1 U19109 ( .B1(n16624), .B2(n15835), .A(n15834), .ZN(n15836) );
  AOI21_X1 U19110 ( .B1(n15837), .B2(n16645), .A(n15836), .ZN(n15838) );
  OAI211_X1 U19111 ( .C1(n15841), .C2(n15840), .A(n15839), .B(n15838), .ZN(
        n15842) );
  NOR2_X1 U19112 ( .A1(n15843), .A2(n15842), .ZN(n15844) );
  OAI21_X1 U19113 ( .B1(n16651), .B2(n15845), .A(n15844), .ZN(P2_U3021) );
  OAI21_X1 U19114 ( .B1(n15847), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15846), .ZN(n15850) );
  AOI21_X1 U19115 ( .B1(n16643), .B2(n16467), .A(n15848), .ZN(n15849) );
  OAI211_X1 U19116 ( .C1(n16629), .C2(n16469), .A(n15850), .B(n15849), .ZN(
        n15851) );
  AOI21_X1 U19117 ( .B1(n15852), .B2(n16646), .A(n15851), .ZN(n15853) );
  OAI21_X1 U19118 ( .B1(n15854), .B2(n16651), .A(n15853), .ZN(P2_U3022) );
  NOR2_X1 U19119 ( .A1(n15893), .A2(n15855), .ZN(n15864) );
  OAI211_X1 U19120 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15873), .B(n15856), .ZN(
        n15858) );
  OAI211_X1 U19121 ( .C1(n16624), .C2(n15859), .A(n15858), .B(n15857), .ZN(
        n15860) );
  INV_X1 U19122 ( .A(n15860), .ZN(n15861) );
  OAI21_X1 U19123 ( .B1(n15862), .B2(n16629), .A(n15861), .ZN(n15863) );
  AOI211_X1 U19124 ( .C1(n15865), .C2(n16646), .A(n15864), .B(n15863), .ZN(
        n15866) );
  OAI21_X1 U19125 ( .B1(n15867), .B2(n16651), .A(n15866), .ZN(P2_U3023) );
  NOR2_X1 U19126 ( .A1(n15871), .A2(n9761), .ZN(n15872) );
  XNOR2_X1 U19127 ( .A(n15870), .B(n15872), .ZN(n16493) );
  NAND2_X1 U19128 ( .A1(n16493), .A2(n16600), .ZN(n15881) );
  NOR2_X1 U19129 ( .A1(n10965), .A2(n19364), .ZN(n15876) );
  INV_X1 U19130 ( .A(n15873), .ZN(n15874) );
  NOR2_X1 U19131 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15874), .ZN(
        n15875) );
  NOR2_X1 U19132 ( .A1(n15876), .A2(n15875), .ZN(n15877) );
  OAI21_X1 U19133 ( .B1(n16624), .B2(n15878), .A(n15877), .ZN(n15879) );
  AOI21_X1 U19134 ( .B1(n16492), .B2(n16645), .A(n15879), .ZN(n15880) );
  OAI211_X1 U19135 ( .C1(n15893), .C2(n15882), .A(n15881), .B(n15880), .ZN(
        n15883) );
  AOI21_X1 U19136 ( .B1(n16491), .B2(n16646), .A(n15883), .ZN(n15884) );
  INV_X1 U19137 ( .A(n15884), .ZN(P2_U3024) );
  INV_X1 U19138 ( .A(n15885), .ZN(n15895) );
  NOR2_X1 U19139 ( .A1(n16624), .A2(n15886), .ZN(n15890) );
  OAI21_X1 U19140 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15888), .A(
        n15887), .ZN(n15889) );
  AOI211_X1 U19141 ( .C1(n15891), .C2(n16645), .A(n15890), .B(n15889), .ZN(
        n15892) );
  OAI21_X1 U19142 ( .B1(n15893), .B2(n10199), .A(n15892), .ZN(n15894) );
  AOI21_X1 U19143 ( .B1(n15895), .B2(n16646), .A(n15894), .ZN(n15896) );
  OAI21_X1 U19144 ( .B1(n15897), .B2(n16651), .A(n15896), .ZN(P2_U3025) );
  INV_X1 U19145 ( .A(n15898), .ZN(n15914) );
  AND2_X1 U19146 ( .A1(n15903), .A2(n15899), .ZN(n15900) );
  NAND2_X1 U19147 ( .A1(n16597), .A2(n15900), .ZN(n15923) );
  OR2_X1 U19148 ( .A1(n16609), .A2(n15903), .ZN(n15901) );
  AND2_X1 U19149 ( .A1(n16608), .A2(n15901), .ZN(n15935) );
  AOI21_X1 U19150 ( .B1(n15923), .B2(n15935), .A(n15902), .ZN(n15913) );
  NAND4_X1 U19151 ( .A1(n16597), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15903), .A4(n15902), .ZN(n15910) );
  AND2_X1 U19152 ( .A1(n15905), .A2(n15904), .ZN(n15906) );
  NOR2_X1 U19153 ( .A1(n15907), .A2(n15906), .ZN(n19258) );
  AOI21_X1 U19154 ( .B1(n16643), .B2(n19258), .A(n15908), .ZN(n15909) );
  OAI211_X1 U19155 ( .C1(n15911), .C2(n16629), .A(n15910), .B(n15909), .ZN(
        n15912) );
  AOI211_X1 U19156 ( .C1(n15914), .C2(n16646), .A(n15913), .B(n15912), .ZN(
        n15915) );
  OAI21_X1 U19157 ( .B1(n15916), .B2(n16651), .A(n15915), .ZN(P2_U3026) );
  INV_X1 U19158 ( .A(n15935), .ZN(n15921) );
  AOI21_X1 U19159 ( .B1(n16643), .B2(n15918), .A(n15917), .ZN(n15919) );
  OAI21_X1 U19160 ( .B1(n16629), .B2(n19273), .A(n15919), .ZN(n15920) );
  AOI21_X1 U19161 ( .B1(n15921), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15920), .ZN(n15922) );
  NAND2_X1 U19162 ( .A1(n15923), .A2(n15922), .ZN(n15924) );
  AOI21_X1 U19163 ( .B1(n15925), .B2(n16646), .A(n15924), .ZN(n15926) );
  OAI21_X1 U19164 ( .B1(n15927), .B2(n16651), .A(n15926), .ZN(P2_U3027) );
  AND2_X1 U19165 ( .A1(n16597), .A2(n15941), .ZN(n15978) );
  NAND4_X1 U19166 ( .A1(n15978), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15928), .A4(n15934), .ZN(n15933) );
  NOR2_X1 U19167 ( .A1(n16629), .A2(n15929), .ZN(n15930) );
  AOI211_X1 U19168 ( .C1(n16643), .C2(n16486), .A(n15931), .B(n15930), .ZN(
        n15932) );
  OAI211_X1 U19169 ( .C1(n15935), .C2(n15934), .A(n15933), .B(n15932), .ZN(
        n15936) );
  AOI21_X1 U19170 ( .B1(n15937), .B2(n16646), .A(n15936), .ZN(n15938) );
  OAI21_X1 U19171 ( .B1(n15939), .B2(n16651), .A(n15938), .ZN(P2_U3028) );
  INV_X1 U19172 ( .A(n15940), .ZN(n15945) );
  OR2_X1 U19173 ( .A1(n16609), .A2(n15941), .ZN(n15942) );
  NAND2_X1 U19174 ( .A1(n16608), .A2(n15942), .ZN(n15967) );
  OAI21_X1 U19175 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16609), .A(
        n15956), .ZN(n15951) );
  AOI21_X1 U19176 ( .B1(n16508), .B2(n16646), .A(n15978), .ZN(n15946) );
  NOR2_X1 U19177 ( .A1(n15946), .A2(n15977), .ZN(n15959) );
  NAND3_X1 U19178 ( .A1(n15959), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15947), .ZN(n15949) );
  AOI22_X1 U19179 ( .A1(n16643), .A2(n19293), .B1(P2_REIP_REG_17__SCAN_IN), 
        .B2(n16616), .ZN(n15948) );
  OAI211_X1 U19180 ( .C1(n19286), .C2(n16629), .A(n15949), .B(n15948), .ZN(
        n15950) );
  AOI21_X1 U19181 ( .B1(n15951), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15950), .ZN(n15952) );
  OAI21_X1 U19182 ( .B1(n15953), .B2(n16651), .A(n15952), .ZN(P2_U3029) );
  NAND2_X1 U19183 ( .A1(n16645), .A2(n19301), .ZN(n15955) );
  OAI211_X1 U19184 ( .C1(n16624), .C2(n19302), .A(n15955), .B(n15954), .ZN(
        n15957) );
  OAI21_X1 U19185 ( .B1(n16651), .B2(n15961), .A(n15960), .ZN(P2_U3030) );
  INV_X1 U19186 ( .A(n15962), .ZN(n15964) );
  NOR2_X1 U19187 ( .A1(n15964), .A2(n15963), .ZN(n15965) );
  XNOR2_X1 U19188 ( .A(n15966), .B(n15965), .ZN(n16498) );
  INV_X1 U19189 ( .A(n19314), .ZN(n15975) );
  NAND2_X1 U19190 ( .A1(n15967), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15974) );
  INV_X1 U19191 ( .A(n14113), .ZN(n15968) );
  OAI21_X1 U19192 ( .B1(n15970), .B2(n15969), .A(n15968), .ZN(n19442) );
  INV_X1 U19193 ( .A(n19442), .ZN(n15972) );
  NOR2_X1 U19194 ( .A1(n10948), .A2(n19364), .ZN(n15971) );
  AOI21_X1 U19195 ( .B1(n16643), .B2(n15972), .A(n15971), .ZN(n15973) );
  OAI211_X1 U19196 ( .C1(n16629), .C2(n15975), .A(n15974), .B(n15973), .ZN(
        n15976) );
  AOI21_X1 U19197 ( .B1(n15978), .B2(n15977), .A(n15976), .ZN(n15981) );
  OAI21_X1 U19198 ( .B1(n16508), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15979), .ZN(n16497) );
  OR2_X1 U19199 ( .A1(n16497), .A2(n16630), .ZN(n15980) );
  OAI211_X1 U19200 ( .C1(n16498), .C2(n16651), .A(n15981), .B(n15980), .ZN(
        P2_U3031) );
  NAND2_X1 U19201 ( .A1(n15983), .A2(n15982), .ZN(n15984) );
  XOR2_X1 U19202 ( .A(n15984), .B(n9721), .Z(n16514) );
  NAND2_X1 U19203 ( .A1(n16024), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16545) );
  NOR2_X1 U19204 ( .A1(n16545), .A2(n16001), .ZN(n15996) );
  NAND2_X1 U19205 ( .A1(n15996), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16531) );
  INV_X1 U19206 ( .A(n16531), .ZN(n15985) );
  NAND2_X1 U19207 ( .A1(n16024), .A2(n16594), .ZN(n16509) );
  OAI21_X1 U19208 ( .B1(n15985), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16509), .ZN(n16515) );
  INV_X1 U19209 ( .A(n16515), .ZN(n15994) );
  NAND2_X1 U19210 ( .A1(n16610), .A2(n16597), .ZN(n15986) );
  NOR2_X1 U19211 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15986), .ZN(
        n16603) );
  NAND3_X1 U19212 ( .A1(n16610), .A2(n16597), .A3(n16528), .ZN(n16618) );
  OAI211_X1 U19213 ( .C1(n16610), .C2(n16609), .A(n16608), .B(n16618), .ZN(
        n16602) );
  AOI22_X1 U19214 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16603), .B1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16602), .ZN(n15992) );
  OAI21_X1 U19215 ( .B1(n15988), .B2(n13889), .A(n15987), .ZN(n19447) );
  INV_X1 U19216 ( .A(n19447), .ZN(n15990) );
  AOI22_X1 U19217 ( .A1(n16643), .A2(n15990), .B1(n15989), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n15991) );
  OAI211_X1 U19218 ( .C1(n16629), .C2(n19329), .A(n15992), .B(n15991), .ZN(
        n15993) );
  AOI21_X1 U19219 ( .B1(n15994), .B2(n16646), .A(n15993), .ZN(n15995) );
  OAI21_X1 U19220 ( .B1(n16651), .B2(n16514), .A(n15995), .ZN(P2_U3033) );
  NOR2_X1 U19221 ( .A1(n16545), .A2(n11519), .ZN(n16546) );
  INV_X1 U19222 ( .A(n15996), .ZN(n16529) );
  OAI21_X1 U19223 ( .B1(n16546), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16529), .ZN(n16540) );
  NOR2_X1 U19224 ( .A1(n15998), .A2(n10273), .ZN(n15999) );
  XNOR2_X1 U19225 ( .A(n16000), .B(n15999), .ZN(n16539) );
  OAI21_X1 U19226 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16609), .A(
        n16608), .ZN(n16627) );
  INV_X1 U19227 ( .A(n16001), .ZN(n16002) );
  NAND2_X1 U19228 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16597), .ZN(
        n16623) );
  AOI211_X1 U19229 ( .C1(n11519), .C2(n16003), .A(n16002), .B(n16623), .ZN(
        n16005) );
  NOR2_X1 U19230 ( .A1(n10888), .A2(n19364), .ZN(n16004) );
  AOI211_X1 U19231 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16627), .A(
        n16005), .B(n16004), .ZN(n16011) );
  OAI21_X1 U19232 ( .B1(n16008), .B2(n16007), .A(n16006), .ZN(n19452) );
  INV_X1 U19233 ( .A(n19452), .ZN(n16009) );
  AOI22_X1 U19234 ( .A1(n16643), .A2(n16009), .B1(n16645), .B2(n19340), .ZN(
        n16010) );
  OAI211_X1 U19235 ( .C1(n16539), .C2(n16651), .A(n16011), .B(n16010), .ZN(
        n16012) );
  INV_X1 U19236 ( .A(n16012), .ZN(n16013) );
  OAI21_X1 U19237 ( .B1(n16540), .B2(n16630), .A(n16013), .ZN(P2_U3035) );
  NAND2_X1 U19238 ( .A1(n16014), .A2(n16015), .ZN(n16567) );
  INV_X1 U19239 ( .A(n16565), .ZN(n16017) );
  INV_X1 U19240 ( .A(n16016), .ZN(n16566) );
  AOI21_X1 U19241 ( .B1(n16567), .B2(n16017), .A(n16566), .ZN(n16021) );
  NAND2_X1 U19242 ( .A1(n16021), .A2(n16019), .ZN(n16549) );
  INV_X1 U19243 ( .A(n16548), .ZN(n16018) );
  OR2_X1 U19244 ( .A1(n16549), .A2(n16018), .ZN(n16023) );
  AND2_X1 U19245 ( .A1(n16019), .A2(n16548), .ZN(n16020) );
  OR2_X1 U19246 ( .A1(n16021), .A2(n16020), .ZN(n16022) );
  NAND2_X1 U19247 ( .A1(n16023), .A2(n16022), .ZN(n16559) );
  OAI21_X1 U19248 ( .B1(n16024), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16545), .ZN(n16560) );
  OR2_X1 U19249 ( .A1(n16560), .A2(n16630), .ZN(n16034) );
  OAI21_X1 U19250 ( .B1(n16026), .B2(n16025), .A(n16622), .ZN(n19457) );
  INV_X1 U19251 ( .A(n19457), .ZN(n16028) );
  NOR2_X1 U19252 ( .A1(n10855), .A2(n19364), .ZN(n16027) );
  AOI21_X1 U19253 ( .B1(n16643), .B2(n16028), .A(n16027), .ZN(n16030) );
  NAND2_X1 U19254 ( .A1(n16645), .A2(n19360), .ZN(n16029) );
  OAI211_X1 U19255 ( .C1(n16608), .C2(n16032), .A(n16030), .B(n16029), .ZN(
        n16031) );
  AOI21_X1 U19256 ( .B1(n16597), .B2(n16032), .A(n16031), .ZN(n16033) );
  OAI211_X1 U19257 ( .C1(n16651), .C2(n16559), .A(n16034), .B(n16033), .ZN(
        P2_U3037) );
  NAND2_X1 U19258 ( .A1(n16035), .A2(n16646), .ZN(n16045) );
  NOR2_X1 U19259 ( .A1(n16609), .A2(n16036), .ZN(n16037) );
  NOR2_X1 U19260 ( .A1(n16038), .A2(n16037), .ZN(n16640) );
  NAND2_X1 U19261 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n16616), .ZN(n16039) );
  OAI221_X1 U19262 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16638), .C1(
        n16040), .C2(n16640), .A(n16039), .ZN(n16043) );
  NOR2_X1 U19263 ( .A1(n16041), .A2(n16629), .ZN(n16042) );
  AOI211_X1 U19264 ( .C1(n19463), .C2(n16643), .A(n16043), .B(n16042), .ZN(
        n16044) );
  OAI211_X1 U19265 ( .C1(n16046), .C2(n16651), .A(n16045), .B(n16044), .ZN(
        P2_U3039) );
  XOR2_X1 U19266 ( .A(n16048), .B(n16047), .Z(n16580) );
  INV_X1 U19267 ( .A(n16580), .ZN(n16067) );
  INV_X1 U19268 ( .A(n16049), .ZN(n16051) );
  NAND3_X1 U19269 ( .A1(n16052), .A2(n16051), .A3(n16050), .ZN(n16053) );
  NAND2_X1 U19270 ( .A1(n16054), .A2(n16053), .ZN(n19465) );
  OAI22_X1 U19271 ( .A1(n16640), .A2(n16055), .B1(n16624), .B2(n19465), .ZN(
        n16061) );
  NOR3_X1 U19272 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16057), .A3(
        n16056), .ZN(n16060) );
  NOR2_X1 U19273 ( .A1(n19333), .A2(n16058), .ZN(n16059) );
  OR3_X1 U19274 ( .A1(n16061), .A2(n16060), .A3(n16059), .ZN(n16065) );
  OAI21_X1 U19275 ( .B1(n16063), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16062), .ZN(n16578) );
  NOR2_X1 U19276 ( .A1(n16578), .A2(n16630), .ZN(n16064) );
  AOI211_X1 U19277 ( .C1(n19371), .C2(n16645), .A(n16065), .B(n16064), .ZN(
        n16066) );
  OAI21_X1 U19278 ( .B1(n16651), .B2(n16067), .A(n16066), .ZN(P2_U3040) );
  INV_X1 U19279 ( .A(n20190), .ZN(n16081) );
  AOI211_X1 U19280 ( .C1(n19426), .C2(n16069), .A(n19393), .B(n16068), .ZN(
        n19412) );
  AOI21_X1 U19281 ( .B1(n19393), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19412), .ZN(n20188) );
  NAND2_X1 U19282 ( .A1(n9677), .A2(n16070), .ZN(n16079) );
  OAI22_X1 U19283 ( .A1(n16075), .A2(n16074), .B1(n16073), .B2(n16072), .ZN(
        n16078) );
  NOR2_X1 U19284 ( .A1(n9675), .A2(n16076), .ZN(n16077) );
  AOI211_X1 U19285 ( .C1(n16080), .C2(n16079), .A(n16078), .B(n16077), .ZN(
        n16652) );
  OAI222_X1 U19286 ( .A1(n20210), .A2(n16081), .B1(n20188), .B2(n20187), .C1(
        n19233), .C2(n16652), .ZN(n16082) );
  MUX2_X1 U19287 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16082), .S(
        n20192), .Z(P2_U3599) );
  INV_X1 U19288 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16084) );
  AOI22_X1 U19289 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16083) );
  OAI21_X1 U19290 ( .B1(n10316), .B2(n16084), .A(n16083), .ZN(n16094) );
  AOI22_X1 U19291 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17545), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16092) );
  OAI22_X1 U19292 ( .A1(n9652), .A2(n16085), .B1(n11180), .B2(n17347), .ZN(
        n16090) );
  AOI22_X1 U19293 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16088) );
  AOI22_X1 U19294 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16087) );
  AOI22_X1 U19295 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16086) );
  NAND3_X1 U19296 ( .A1(n16088), .A2(n16087), .A3(n16086), .ZN(n16089) );
  AOI211_X1 U19297 ( .C1(n9647), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n16090), .B(n16089), .ZN(n16091) );
  OAI211_X1 U19298 ( .C1(n10314), .C2(n18576), .A(n16092), .B(n16091), .ZN(
        n16093) );
  AOI211_X1 U19299 ( .C1(n17450), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n16094), .B(n16093), .ZN(n17681) );
  OAI211_X1 U19300 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n17482), .A(n17460), .B(
        n17578), .ZN(n16095) );
  OAI21_X1 U19301 ( .B1(n17681), .B2(n17578), .A(n16095), .ZN(P3_U2690) );
  NOR2_X1 U19302 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19160), .ZN(
        n18532) );
  NAND3_X1 U19303 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19158)
         );
  INV_X1 U19304 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17196) );
  OAI21_X1 U19305 ( .B1(n19026), .B2(n19167), .A(n17196), .ZN(n16111) );
  NOR2_X1 U19306 ( .A1(n9651), .A2(n16111), .ZN(n18531) );
  INV_X1 U19307 ( .A(n18905), .ZN(n18656) );
  INV_X1 U19308 ( .A(n19158), .ZN(n16096) );
  NAND2_X1 U19309 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n16096), .ZN(n16110) );
  OAI211_X1 U19310 ( .C1(n19158), .C2(n18531), .A(n18656), .B(n16110), .ZN(
        n18539) );
  INV_X1 U19311 ( .A(n18539), .ZN(n18535) );
  NOR2_X1 U19312 ( .A1(n18532), .A2(n18535), .ZN(n16098) );
  INV_X1 U19313 ( .A(n18853), .ZN(n18902) );
  INV_X1 U19314 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19010) );
  OAI22_X1 U19315 ( .A1(n18166), .A2(n19205), .B1(n19010), .B2(n19160), .ZN(
        n16101) );
  NAND3_X1 U19316 ( .A1(n19012), .A2(n18539), .A3(n16101), .ZN(n16097) );
  OAI221_X1 U19317 ( .B1(n19012), .B2(n16098), .C1(n19012), .C2(n18902), .A(
        n16097), .ZN(P3_U2864) );
  NAND2_X1 U19318 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18724) );
  NOR2_X1 U19319 ( .A1(n18166), .A2(n19205), .ZN(n16100) );
  INV_X1 U19320 ( .A(n16098), .ZN(n16099) );
  AOI221_X1 U19321 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18724), .C1(n16100), 
        .C2(n18724), .A(n16099), .ZN(n18538) );
  OAI221_X1 U19322 ( .B1(n18853), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18853), .C2(n16101), .A(n18539), .ZN(n18536) );
  AOI22_X1 U19323 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18538), .B1(
        n18536), .B2(n19030), .ZN(P3_U2865) );
  NAND2_X1 U19324 ( .A1(n18986), .A2(n19213), .ZN(n16106) );
  OAI21_X1 U19325 ( .B1(n16104), .B2(n19046), .A(n16103), .ZN(n17745) );
  OAI21_X1 U19326 ( .B1(n16106), .B2(n17745), .A(n16105), .ZN(n16107) );
  NAND2_X1 U19327 ( .A1(n19052), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18543) );
  OAI211_X1 U19328 ( .C1(n19044), .C2(n19029), .A(n18543), .B(n16110), .ZN(
        n19189) );
  INV_X1 U19329 ( .A(n16111), .ZN(n16112) );
  NOR2_X1 U19330 ( .A1(n16112), .A2(n19014), .ZN(n18994) );
  NAND3_X1 U19331 ( .A1(n19189), .A2(n19223), .A3(n18994), .ZN(n16113) );
  OAI21_X1 U19332 ( .B1(n19189), .B2(n17196), .A(n16113), .ZN(P3_U3284) );
  AOI21_X1 U19333 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16114), .A(
        n16115), .ZN(n16743) );
  INV_X1 U19334 ( .A(n18431), .ZN(n18372) );
  NAND2_X1 U19335 ( .A1(n16173), .A2(n18220), .ZN(n16725) );
  INV_X1 U19336 ( .A(n16724), .ZN(n16116) );
  AOI22_X1 U19337 ( .A1(n18372), .A2(n16725), .B1(n18527), .B2(n16116), .ZN(
        n16177) );
  OAI21_X1 U19338 ( .B1(n18382), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16117), .ZN(n16749) );
  AOI22_X1 U19339 ( .A1(n18521), .A2(n16749), .B1(n18515), .B2(n17852), .ZN(
        n16118) );
  NAND3_X1 U19340 ( .A1(n16177), .A2(n16118), .A3(n18511), .ZN(n16123) );
  INV_X1 U19341 ( .A(n18527), .ZN(n18518) );
  OAI21_X1 U19342 ( .B1(n18518), .B2(n18218), .A(n16119), .ZN(n16120) );
  AOI21_X1 U19343 ( .B1(n18220), .B2(n18372), .A(n16120), .ZN(n16181) );
  NOR2_X1 U19344 ( .A1(n16181), .A2(n16729), .ZN(n16122) );
  AOI22_X1 U19345 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16123), .B1(
        n16122), .B2(n16121), .ZN(n16124) );
  NAND2_X1 U19346 ( .A1(n18483), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16739) );
  OAI211_X1 U19347 ( .C1(n16743), .C2(n21258), .A(n16124), .B(n16739), .ZN(
        P3_U2833) );
  INV_X1 U19348 ( .A(n16125), .ZN(n16137) );
  AND2_X1 U19349 ( .A1(n16126), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16127) );
  AND2_X1 U19350 ( .A1(n16128), .A2(n16127), .ZN(n16133) );
  AOI211_X1 U19351 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16133), .A(
        n16130), .B(n16129), .ZN(n16131) );
  INV_X1 U19352 ( .A(n16131), .ZN(n16132) );
  OAI21_X1 U19353 ( .B1(n16133), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16132), .ZN(n16134) );
  AOI222_X1 U19354 ( .A1(n12762), .A2(n16135), .B1(n12762), .B2(n16134), .C1(
        n16135), .C2(n16134), .ZN(n16136) );
  AOI222_X1 U19355 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16137), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16136), .C1(n16137), 
        .C2(n16136), .ZN(n16146) );
  OAI21_X1 U19356 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n16138), .ZN(n16139) );
  NAND4_X1 U19357 ( .A1(n16142), .A2(n16141), .A3(n16140), .A4(n16139), .ZN(
        n16143) );
  OR2_X1 U19358 ( .A1(n16144), .A2(n16143), .ZN(n16145) );
  AOI21_X1 U19359 ( .B1(n16146), .B2(n20456), .A(n16145), .ZN(n16156) );
  INV_X1 U19360 ( .A(n16156), .ZN(n16148) );
  AOI21_X1 U19361 ( .B1(n16149), .B2(n16148), .A(n16147), .ZN(n16162) );
  INV_X1 U19362 ( .A(n16150), .ZN(n16158) );
  NAND3_X1 U19363 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21050), .A3(n21045), 
        .ZN(n16155) );
  INV_X1 U19364 ( .A(n16151), .ZN(n16153) );
  NOR3_X1 U19365 ( .A1(n16153), .A2(n16182), .A3(n16152), .ZN(n16154) );
  AOI21_X1 U19366 ( .B1(n16155), .B2(n20944), .A(n16154), .ZN(n16417) );
  OAI221_X1 U19367 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n16156), 
        .A(n16417), .ZN(n16157) );
  OAI211_X1 U19368 ( .C1(n16416), .C2(P1_STATE2_REG_2__SCAN_IN), .A(n16158), 
        .B(n20945), .ZN(n16419) );
  INV_X1 U19369 ( .A(n16419), .ZN(n16161) );
  OAI21_X1 U19370 ( .B1(n16159), .B2(n16158), .A(n16157), .ZN(n16160) );
  AOI22_X1 U19371 ( .A1(n16162), .A2(n16161), .B1(n21045), .B2(n16160), .ZN(
        P1_U3161) );
  AOI22_X1 U19372 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n16312), .B1(
        n16391), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n16172) );
  OAI22_X1 U19373 ( .A1(n16164), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16163), .B2(n15061), .ZN(n16165) );
  OAI21_X1 U19374 ( .B1(n16167), .B2(n16166), .A(n16165), .ZN(n16168) );
  XNOR2_X1 U19375 ( .A(n16168), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16249) );
  XOR2_X1 U19376 ( .A(n16170), .B(n16169), .Z(n16246) );
  AOI22_X1 U19377 ( .A1(n16249), .A2(n16394), .B1(n20451), .B2(n16246), .ZN(
        n16171) );
  OAI211_X1 U19378 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n16320), .A(
        n16172), .B(n16171), .ZN(P1_U3010) );
  NAND2_X1 U19379 ( .A1(n16173), .A2(n16176), .ZN(n16728) );
  AOI21_X1 U19380 ( .B1(n16175), .B2(n16176), .A(n16174), .ZN(n16723) );
  AOI21_X1 U19381 ( .B1(n16178), .B2(n16177), .A(n16176), .ZN(n16179) );
  AOI21_X1 U19382 ( .B1(n9631), .B2(n16723), .A(n16179), .ZN(n16180) );
  NAND2_X1 U19383 ( .A1(n18483), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16720) );
  OAI211_X1 U19384 ( .C1(n16181), .C2(n16728), .A(n16180), .B(n16720), .ZN(
        P3_U2832) );
  INV_X1 U19385 ( .A(HOLD), .ZN(n21190) );
  NAND2_X1 U19386 ( .A1(n11877), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20952) );
  INV_X1 U19387 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21188) );
  NOR2_X1 U19388 ( .A1(n13206), .A2(n21188), .ZN(n20950) );
  NAND2_X1 U19389 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21050), .ZN(n20953) );
  INV_X1 U19390 ( .A(n20953), .ZN(n20951) );
  AOI221_X1 U19391 ( .B1(n21190), .B2(n20950), .C1(n11877), .C2(n20950), .A(
        n20951), .ZN(n16183) );
  OAI211_X1 U19392 ( .C1(n21190), .C2(n20952), .A(n16183), .B(n16182), .ZN(
        P1_U3195) );
  AND2_X1 U19393 ( .A1(n20409), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AND3_X1 U19394 ( .A1(n16186), .A2(n16185), .A3(n16184), .ZN(n16192) );
  OR2_X1 U19395 ( .A1(n15061), .A2(n16187), .ZN(n16188) );
  NAND2_X1 U19396 ( .A1(n16189), .A2(n16188), .ZN(n16190) );
  XNOR2_X1 U19397 ( .A(n16190), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16254) );
  NOR2_X1 U19398 ( .A1(n16254), .A2(n20446), .ZN(n16191) );
  AOI211_X1 U19399 ( .C1(n20451), .C2(n16193), .A(n16192), .B(n16191), .ZN(
        n16194) );
  NAND2_X1 U19400 ( .A1(n16391), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16258) );
  OAI211_X1 U19401 ( .C1(n16195), .C2(n12753), .A(n16194), .B(n16258), .ZN(
        P1_U3011) );
  INV_X1 U19402 ( .A(n16196), .ZN(n16705) );
  NOR3_X1 U19403 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16197) );
  NOR3_X1 U19404 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20256), .A3(n20257), 
        .ZN(n16697) );
  OR2_X1 U19405 ( .A1(n16197), .A2(n16697), .ZN(n20108) );
  NOR3_X1 U19406 ( .A1(n16705), .A2(n16699), .A3(n20108), .ZN(P2_U3178) );
  INV_X1 U19407 ( .A(n16699), .ZN(n16713) );
  OAI221_X1 U19408 ( .B1(n11632), .B2(n16713), .C1(n20243), .C2(n16713), .A(
        n19764), .ZN(n20238) );
  NOR2_X1 U19409 ( .A1(n16198), .A2(n20238), .ZN(P2_U3047) );
  NOR3_X1 U19410 ( .A1(n16199), .A2(n18545), .A3(n18551), .ZN(n16200) );
  NAND2_X1 U19411 ( .A1(n17711), .A2(n17586), .ZN(n17589) );
  INV_X1 U19412 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17817) );
  AOI22_X1 U19413 ( .A1(n17741), .A2(BUF2_REG_0__SCAN_IN), .B1(n17730), .B2(
        n18205), .ZN(n16203) );
  OAI221_X1 U19414 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17589), .C1(n17817), 
        .C2(n17586), .A(n16203), .ZN(P3_U2735) );
  INV_X1 U19415 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20992) );
  AOI22_X1 U19416 ( .A1(n20360), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20348), .ZN(n16204) );
  OAI21_X1 U19417 ( .B1(n16253), .B2(n20375), .A(n16204), .ZN(n16205) );
  AOI221_X1 U19418 ( .B1(n16207), .B2(n20992), .C1(n16206), .C2(
        P1_REIP_REG_21__SCAN_IN), .A(n16205), .ZN(n16209) );
  AOI22_X1 U19419 ( .A1(n16250), .A2(n20328), .B1(n20362), .B2(n16246), .ZN(
        n16208) );
  NAND2_X1 U19420 ( .A1(n16209), .A2(n16208), .ZN(P1_U2819) );
  AOI22_X1 U19421 ( .A1(n20360), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20348), .ZN(n16215) );
  AOI21_X1 U19422 ( .B1(n20349), .B2(n16269), .A(n20346), .ZN(n16214) );
  AOI22_X1 U19423 ( .A1(n16270), .A2(n20328), .B1(n20362), .B2(n16210), .ZN(
        n16213) );
  OAI21_X1 U19424 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n9769), .A(n16211), .ZN(
        n16212) );
  NAND4_X1 U19425 ( .A1(n16215), .A2(n16214), .A3(n16213), .A4(n16212), .ZN(
        P1_U2823) );
  OAI21_X1 U19426 ( .B1(n20365), .B2(n16216), .A(n20308), .ZN(n16219) );
  OAI22_X1 U19427 ( .A1(n16217), .A2(n20325), .B1(n20320), .B2(n16359), .ZN(
        n16218) );
  AOI211_X1 U19428 ( .C1(n16220), .C2(n20349), .A(n16219), .B(n16218), .ZN(
        n16224) );
  AOI22_X1 U19429 ( .A1(n16222), .A2(n20328), .B1(n10074), .B2(n16221), .ZN(
        n16223) );
  OAI211_X1 U19430 ( .C1(n16225), .C2(n10074), .A(n16224), .B(n16223), .ZN(
        P1_U2827) );
  OAI222_X1 U19431 ( .A1(n16227), .A2(n20320), .B1(n20325), .B2(n14915), .C1(
        n20975), .C2(n16226), .ZN(n16228) );
  AOI211_X1 U19432 ( .C1(n20348), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20346), .B(n16228), .ZN(n16233) );
  INV_X1 U19433 ( .A(n16229), .ZN(n16230) );
  AOI22_X1 U19434 ( .A1(n16231), .A2(n20328), .B1(n20349), .B2(n16230), .ZN(
        n16232) );
  OAI211_X1 U19435 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n16234), .A(n16233), 
        .B(n16232), .ZN(P1_U2829) );
  NAND2_X1 U19436 ( .A1(n16235), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16245) );
  INV_X1 U19437 ( .A(n16236), .ZN(n16237) );
  AOI22_X1 U19438 ( .A1(n20362), .A2(n16237), .B1(n20360), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n16238) );
  OAI211_X1 U19439 ( .C1(n20365), .C2(n16239), .A(n16238), .B(n20308), .ZN(
        n16240) );
  AOI21_X1 U19440 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n16241), .A(n16240), 
        .ZN(n16244) );
  INV_X1 U19441 ( .A(n16242), .ZN(n16287) );
  AOI22_X1 U19442 ( .A1(n16287), .A2(n20328), .B1(n20349), .B2(n16284), .ZN(
        n16243) );
  OAI211_X1 U19443 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n16245), .A(n16244), 
        .B(n16243), .ZN(P1_U2830) );
  AOI22_X1 U19444 ( .A1(n16250), .A2(n20383), .B1(n20382), .B2(n16246), .ZN(
        n16247) );
  OAI21_X1 U19445 ( .B1(n20387), .B2(n16248), .A(n16247), .ZN(P1_U2851) );
  AOI22_X1 U19446 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n16252) );
  AOI22_X1 U19447 ( .A1(n16250), .A2(n16286), .B1(n16296), .B2(n16249), .ZN(
        n16251) );
  OAI211_X1 U19448 ( .C1(n16299), .C2(n16253), .A(n16252), .B(n16251), .ZN(
        P1_U2978) );
  OAI22_X1 U19449 ( .A1(n16255), .A2(n16263), .B1(n20282), .B2(n16254), .ZN(
        n16256) );
  AOI21_X1 U19450 ( .B1(n16285), .B2(n16257), .A(n16256), .ZN(n16259) );
  OAI211_X1 U19451 ( .C1(n16261), .C2(n16260), .A(n16259), .B(n16258), .ZN(
        P1_U2979) );
  AOI22_X1 U19452 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16267) );
  OAI22_X1 U19453 ( .A1(n16264), .A2(n16263), .B1(n16262), .B2(n20282), .ZN(
        n16265) );
  INV_X1 U19454 ( .A(n16265), .ZN(n16266) );
  OAI211_X1 U19455 ( .C1(n16299), .C2(n16268), .A(n16267), .B(n16266), .ZN(
        P1_U2980) );
  AOI22_X1 U19456 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16272) );
  AOI22_X1 U19457 ( .A1(n16270), .A2(n16286), .B1(n16269), .B2(n16285), .ZN(
        n16271) );
  OAI211_X1 U19458 ( .C1(n20282), .C2(n16273), .A(n16272), .B(n16271), .ZN(
        P1_U2982) );
  NOR2_X1 U19459 ( .A1(n16274), .A2(n9950), .ZN(n16278) );
  NAND2_X1 U19460 ( .A1(n16276), .A2(n16275), .ZN(n16277) );
  XNOR2_X1 U19461 ( .A(n16278), .B(n16277), .ZN(n16339) );
  AOI22_X1 U19462 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16283) );
  INV_X1 U19463 ( .A(n16279), .ZN(n16281) );
  AOI22_X1 U19464 ( .A1(n16281), .A2(n16286), .B1(n16285), .B2(n16280), .ZN(
        n16282) );
  OAI211_X1 U19465 ( .C1(n16339), .C2(n20282), .A(n16283), .B(n16282), .ZN(
        P1_U2984) );
  AOI22_X1 U19466 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n16289) );
  AOI22_X1 U19467 ( .A1(n16287), .A2(n16286), .B1(n16285), .B2(n16284), .ZN(
        n16288) );
  OAI211_X1 U19468 ( .C1(n20282), .C2(n16290), .A(n16289), .B(n16288), .ZN(
        P1_U2989) );
  AOI22_X1 U19469 ( .A1(n16291), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16391), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16298) );
  NAND2_X1 U19470 ( .A1(n16293), .A2(n16292), .ZN(n16294) );
  XNOR2_X1 U19471 ( .A(n16295), .B(n16294), .ZN(n16393) );
  AOI22_X1 U19472 ( .A1(n16393), .A2(n16296), .B1(n20316), .B2(n16286), .ZN(
        n16297) );
  OAI211_X1 U19473 ( .C1(n16299), .C2(n20319), .A(n16298), .B(n16297), .ZN(
        P1_U2992) );
  AOI211_X1 U19474 ( .C1(n16370), .C2(n16302), .A(n16301), .B(n16300), .ZN(
        n16310) );
  AOI21_X1 U19475 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16303), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16309) );
  INV_X1 U19476 ( .A(n16304), .ZN(n16306) );
  AOI22_X1 U19477 ( .A1(n16306), .A2(n16394), .B1(n20451), .B2(n16305), .ZN(
        n16308) );
  NAND2_X1 U19478 ( .A1(n16391), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16307) );
  OAI211_X1 U19479 ( .C1(n16310), .C2(n16309), .A(n16308), .B(n16307), .ZN(
        P1_U3007) );
  OAI21_X1 U19480 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16311), .ZN(n16319) );
  AOI22_X1 U19481 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16312), .B1(
        n16391), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16318) );
  INV_X1 U19482 ( .A(n16313), .ZN(n16316) );
  INV_X1 U19483 ( .A(n16314), .ZN(n16315) );
  AOI22_X1 U19484 ( .A1(n16316), .A2(n16394), .B1(n20451), .B2(n16315), .ZN(
        n16317) );
  OAI211_X1 U19485 ( .C1(n16320), .C2(n16319), .A(n16318), .B(n16317), .ZN(
        P1_U3009) );
  AOI22_X1 U19486 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16321), .B1(
        n16391), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n16327) );
  INV_X1 U19487 ( .A(n16322), .ZN(n16325) );
  INV_X1 U19488 ( .A(n16323), .ZN(n16324) );
  AOI22_X1 U19489 ( .A1(n16325), .A2(n16394), .B1(n20451), .B2(n16324), .ZN(
        n16326) );
  OAI211_X1 U19490 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n16328), .A(
        n16327), .B(n16326), .ZN(P1_U3013) );
  INV_X1 U19491 ( .A(n16329), .ZN(n16342) );
  AOI22_X1 U19492 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16342), .B1(
        n16391), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16337) );
  INV_X1 U19493 ( .A(n16330), .ZN(n16332) );
  AOI22_X1 U19494 ( .A1(n16332), .A2(n16394), .B1(n20451), .B2(n16331), .ZN(
        n16336) );
  OAI211_X1 U19495 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16334), .B(n16333), .ZN(
        n16335) );
  NAND3_X1 U19496 ( .A1(n16337), .A2(n16336), .A3(n16335), .ZN(P1_U3015) );
  NOR2_X1 U19497 ( .A1(n16406), .A2(n10076), .ZN(n16341) );
  OAI22_X1 U19498 ( .A1(n16339), .A2(n20446), .B1(n16407), .B2(n16338), .ZN(
        n16340) );
  AOI211_X1 U19499 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16342), .A(
        n16341), .B(n16340), .ZN(n16343) );
  OAI21_X1 U19500 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16344), .A(
        n16343), .ZN(P1_U3016) );
  NAND2_X1 U19501 ( .A1(n16346), .A2(n16345), .ZN(n16390) );
  NAND4_X1 U19502 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n16347), .ZN(n16352) );
  AOI22_X1 U19503 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16363), .B1(
        n16391), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16351) );
  AOI22_X1 U19504 ( .A1(n16349), .A2(n16394), .B1(n20451), .B2(n16348), .ZN(
        n16350) );
  OAI211_X1 U19505 ( .C1(n16390), .C2(n16352), .A(n16351), .B(n16350), .ZN(
        P1_U3017) );
  NAND2_X1 U19506 ( .A1(n16353), .A2(n16357), .ZN(n16366) );
  INV_X1 U19507 ( .A(n16367), .ZN(n16354) );
  NAND3_X1 U19508 ( .A1(n16355), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n16354), .ZN(n16356) );
  OAI211_X1 U19509 ( .C1(n16371), .C2(n16358), .A(n16357), .B(n16356), .ZN(
        n16362) );
  OAI22_X1 U19510 ( .A1(n16360), .A2(n20446), .B1(n16407), .B2(n16359), .ZN(
        n16361) );
  AOI21_X1 U19511 ( .B1(n16363), .B2(n16362), .A(n16361), .ZN(n16365) );
  NAND2_X1 U19512 ( .A1(n16391), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16364) );
  OAI211_X1 U19513 ( .C1(n16367), .C2(n16366), .A(n16365), .B(n16364), .ZN(
        P1_U3018) );
  NAND2_X1 U19514 ( .A1(n16372), .A2(n12745), .ZN(n16382) );
  AOI21_X1 U19515 ( .B1(n20451), .B2(n16369), .A(n16368), .ZN(n16381) );
  INV_X1 U19516 ( .A(n16370), .ZN(n16377) );
  OAI22_X1 U19517 ( .A1(n16374), .A2(n16373), .B1(n16372), .B2(n16371), .ZN(
        n16375) );
  NOR2_X1 U19518 ( .A1(n16376), .A2(n16375), .ZN(n16388) );
  OAI21_X1 U19519 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16377), .A(
        n16388), .ZN(n16378) );
  AOI22_X1 U19520 ( .A1(n16379), .A2(n16394), .B1(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16378), .ZN(n16380) );
  OAI211_X1 U19521 ( .C1(n16383), .C2(n16382), .A(n16381), .B(n16380), .ZN(
        P1_U3019) );
  INV_X1 U19522 ( .A(n16384), .ZN(n16385) );
  AOI222_X1 U19523 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n16391), .B1(n20451), 
        .B2(n16386), .C1(n16394), .C2(n16385), .ZN(n16387) );
  OAI221_X1 U19524 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16390), 
        .C1(n16389), .C2(n16388), .A(n16387), .ZN(P1_U3020) );
  NAND2_X1 U19525 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16399), .ZN(
        n16398) );
  INV_X1 U19526 ( .A(n20312), .ZN(n16392) );
  AOI22_X1 U19527 ( .A1(n20451), .A2(n16392), .B1(n16391), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16397) );
  AOI22_X1 U19528 ( .A1(n16395), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16394), .B2(n16393), .ZN(n16396) );
  OAI211_X1 U19529 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16398), .A(
        n16397), .B(n16396), .ZN(P1_U3024) );
  NAND2_X1 U19530 ( .A1(n16399), .A2(n16414), .ZN(n16410) );
  INV_X1 U19531 ( .A(n16400), .ZN(n16401) );
  AOI21_X1 U19532 ( .B1(n16403), .B2(n16402), .A(n16401), .ZN(n16404) );
  OR2_X1 U19533 ( .A1(n16405), .A2(n16404), .ZN(n20380) );
  INV_X1 U19534 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20968) );
  OAI22_X1 U19535 ( .A1(n16407), .A2(n20380), .B1(n20968), .B2(n16406), .ZN(
        n16408) );
  INV_X1 U19536 ( .A(n16408), .ZN(n16409) );
  OAI211_X1 U19537 ( .C1(n16411), .C2(n20446), .A(n16410), .B(n16409), .ZN(
        n16412) );
  INV_X1 U19538 ( .A(n16412), .ZN(n16413) );
  OAI21_X1 U19539 ( .B1(n16415), .B2(n16414), .A(n16413), .ZN(P1_U3025) );
  OAI221_X1 U19540 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n21045), .C2(n16416), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20946) );
  AOI21_X1 U19541 ( .B1(n16421), .B2(n20946), .A(n16417), .ZN(n16418) );
  AOI21_X1 U19542 ( .B1(n16420), .B2(n16419), .A(n16418), .ZN(P1_U3162) );
  OAI22_X1 U19543 ( .A1(n20945), .A2(n20760), .B1(n21045), .B2(n16421), .ZN(
        P1_U3466) );
  AOI22_X1 U19544 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19406), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19431), .ZN(n16433) );
  OAI22_X1 U19545 ( .A1(n16423), .A2(n19389), .B1(n16422), .B2(n19408), .ZN(
        n16431) );
  AOI211_X1 U19546 ( .C1(n16426), .C2(n16425), .A(n16424), .B(n19394), .ZN(
        n16430) );
  INV_X1 U19547 ( .A(n16427), .ZN(n16428) );
  OAI22_X1 U19548 ( .A1(n16428), .A2(n19423), .B1(n20169), .B2(n19416), .ZN(
        n16429) );
  NOR3_X1 U19549 ( .A1(n16431), .A2(n16430), .A3(n16429), .ZN(n16432) );
  NAND2_X1 U19550 ( .A1(n16433), .A2(n16432), .ZN(P2_U2827) );
  INV_X1 U19551 ( .A(n16434), .ZN(n16436) );
  OAI211_X1 U19552 ( .C1(n16437), .C2(n16436), .A(n16435), .B(n12839), .ZN(
        n16441) );
  AOI22_X1 U19553 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19406), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19431), .ZN(n16438) );
  OAI21_X1 U19554 ( .B1(n19416), .B2(n20168), .A(n16438), .ZN(n16439) );
  INV_X1 U19555 ( .A(n16439), .ZN(n16440) );
  OAI211_X1 U19556 ( .C1(n19389), .C2(n16442), .A(n16441), .B(n16440), .ZN(
        n16447) );
  AOI211_X1 U19557 ( .C1(n16445), .C2(n16444), .A(n16443), .B(n19394), .ZN(
        n16446) );
  NOR2_X1 U19558 ( .A1(n16447), .A2(n16446), .ZN(n16448) );
  OAI21_X1 U19559 ( .B1(n16449), .B2(n19408), .A(n16448), .ZN(P2_U2828) );
  AOI211_X1 U19560 ( .C1(n16452), .C2(n16451), .A(n16450), .B(n19394), .ZN(
        n16461) );
  OAI211_X1 U19561 ( .C1(n16454), .C2(n11012), .A(n16453), .B(n12839), .ZN(
        n16459) );
  AOI22_X1 U19562 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19406), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19402), .ZN(n16458) );
  NAND2_X1 U19563 ( .A1(n16455), .A2(n19425), .ZN(n16457) );
  NAND2_X1 U19564 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19431), .ZN(
        n16456) );
  NAND4_X1 U19565 ( .A1(n16459), .A2(n16458), .A3(n16457), .A4(n16456), .ZN(
        n16460) );
  AOI211_X1 U19566 ( .C1(n19420), .C2(n16462), .A(n16461), .B(n16460), .ZN(
        n16463) );
  INV_X1 U19567 ( .A(n16463), .ZN(P2_U2829) );
  AOI22_X1 U19568 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19431), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19402), .ZN(n16478) );
  INV_X1 U19569 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16464) );
  OAI22_X1 U19570 ( .A1(n16465), .A2(n19423), .B1(n19418), .B2(n16464), .ZN(
        n16466) );
  INV_X1 U19571 ( .A(n16466), .ZN(n16477) );
  INV_X1 U19572 ( .A(n16467), .ZN(n16468) );
  OAI22_X1 U19573 ( .A1(n16469), .A2(n19389), .B1(n19408), .B2(n16468), .ZN(
        n16470) );
  INV_X1 U19574 ( .A(n16470), .ZN(n16476) );
  AOI21_X1 U19575 ( .B1(n16473), .B2(n16472), .A(n16471), .ZN(n16474) );
  NAND2_X1 U19576 ( .A1(n19411), .A2(n16474), .ZN(n16475) );
  NAND4_X1 U19577 ( .A1(n16478), .A2(n16477), .A3(n16476), .A4(n16475), .ZN(
        P2_U2831) );
  AOI22_X1 U19578 ( .A1(n16485), .A2(n16479), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19494), .ZN(n16483) );
  AOI22_X1 U19579 ( .A1(n19438), .A2(BUF2_REG_20__SCAN_IN), .B1(n19436), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U19580 ( .A1(n16480), .A2(n19497), .B1(n19495), .B2(n19258), .ZN(
        n16481) );
  NAND3_X1 U19581 ( .A1(n16483), .A2(n16482), .A3(n16481), .ZN(P2_U2899) );
  AOI22_X1 U19582 ( .A1(n16485), .A2(n16484), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19494), .ZN(n16490) );
  AOI22_X1 U19583 ( .A1(n19438), .A2(BUF2_REG_18__SCAN_IN), .B1(n19436), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U19584 ( .A1(n16487), .A2(n19497), .B1(n19495), .B2(n16486), .ZN(
        n16488) );
  NAND3_X1 U19585 ( .A1(n16490), .A2(n16489), .A3(n16488), .ZN(P2_U2901) );
  AOI22_X1 U19586 ( .A1(n19551), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n16616), .ZN(n16495) );
  AOI222_X1 U19587 ( .A1(n16493), .A2(n19552), .B1(n16589), .B2(n16492), .C1(
        n19554), .C2(n16491), .ZN(n16494) );
  OAI211_X1 U19588 ( .C1(n19564), .C2(n16496), .A(n16495), .B(n16494), .ZN(
        P2_U2992) );
  AOI22_X1 U19589 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n16616), .B1(n16583), 
        .B2(n19313), .ZN(n16501) );
  OAI22_X1 U19590 ( .A1(n16498), .A2(n16586), .B1(n16584), .B2(n16497), .ZN(
        n16499) );
  AOI21_X1 U19591 ( .B1(n16589), .B2(n19314), .A(n16499), .ZN(n16500) );
  OAI211_X1 U19592 ( .C1(n16593), .C2(n16502), .A(n16501), .B(n16500), .ZN(
        P2_U2999) );
  AOI22_X1 U19593 ( .A1(n19551), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n16616), .ZN(n16512) );
  INV_X1 U19594 ( .A(n16503), .ZN(n16505) );
  NOR2_X1 U19595 ( .A1(n16505), .A2(n16504), .ZN(n16506) );
  XNOR2_X1 U19596 ( .A(n16507), .B(n16506), .ZN(n16601) );
  AOI21_X1 U19597 ( .B1(n16510), .B2(n16509), .A(n16508), .ZN(n16598) );
  AOI222_X1 U19598 ( .A1(n16601), .A2(n19552), .B1(n16589), .B2(n16599), .C1(
        n19554), .C2(n16598), .ZN(n16511) );
  OAI211_X1 U19599 ( .C1(n19564), .C2(n16513), .A(n16512), .B(n16511), .ZN(
        P2_U3000) );
  AOI22_X1 U19600 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n16616), .B1(n16583), 
        .B2(n19327), .ZN(n16519) );
  OAI22_X1 U19601 ( .A1(n16515), .A2(n16584), .B1(n16586), .B2(n16514), .ZN(
        n16516) );
  AOI21_X1 U19602 ( .B1(n16589), .B2(n16517), .A(n16516), .ZN(n16518) );
  OAI211_X1 U19603 ( .C1(n16593), .C2(n16520), .A(n16519), .B(n16518), .ZN(
        P2_U3001) );
  AOI22_X1 U19604 ( .A1(n19551), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n16616), .ZN(n16537) );
  NAND2_X1 U19605 ( .A1(n9721), .A2(n16521), .ZN(n16527) );
  INV_X1 U19606 ( .A(n16522), .ZN(n16524) );
  OAI21_X1 U19607 ( .B1(n16525), .B2(n16524), .A(n16523), .ZN(n16526) );
  NAND2_X1 U19608 ( .A1(n16527), .A2(n16526), .ZN(n16613) );
  NAND2_X1 U19609 ( .A1(n16529), .A2(n16528), .ZN(n16530) );
  NAND2_X1 U19610 ( .A1(n16615), .A2(n19554), .ZN(n16534) );
  NAND2_X1 U19611 ( .A1(n16589), .A2(n16532), .ZN(n16533) );
  OAI211_X1 U19612 ( .C1(n16613), .C2(n16586), .A(n16534), .B(n16533), .ZN(
        n16535) );
  INV_X1 U19613 ( .A(n16535), .ZN(n16536) );
  OAI211_X1 U19614 ( .C1(n19564), .C2(n16538), .A(n16537), .B(n16536), .ZN(
        P2_U3002) );
  AOI22_X1 U19615 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n16616), .B1(n16583), 
        .B2(n19339), .ZN(n16543) );
  OAI22_X1 U19616 ( .A1(n16540), .A2(n16584), .B1(n16539), .B2(n16586), .ZN(
        n16541) );
  AOI21_X1 U19617 ( .B1(n16589), .B2(n19340), .A(n16541), .ZN(n16542) );
  OAI211_X1 U19618 ( .C1(n16593), .C2(n16544), .A(n16543), .B(n16542), .ZN(
        P2_U3003) );
  AOI22_X1 U19619 ( .A1(n19551), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n16616), .ZN(n16558) );
  AND2_X1 U19620 ( .A1(n16545), .A2(n11519), .ZN(n16547) );
  OR2_X1 U19621 ( .A1(n16547), .A2(n16546), .ZN(n16631) );
  NAND2_X1 U19622 ( .A1(n16549), .A2(n16548), .ZN(n16553) );
  AND2_X1 U19623 ( .A1(n16551), .A2(n16550), .ZN(n16552) );
  XNOR2_X1 U19624 ( .A(n16553), .B(n16552), .ZN(n16635) );
  OR2_X1 U19625 ( .A1(n16635), .A2(n16586), .ZN(n16555) );
  NAND2_X1 U19626 ( .A1(n16589), .A2(n19350), .ZN(n16554) );
  OAI211_X1 U19627 ( .C1(n16631), .C2(n16584), .A(n16555), .B(n16554), .ZN(
        n16556) );
  INV_X1 U19628 ( .A(n16556), .ZN(n16557) );
  OAI211_X1 U19629 ( .C1(n19564), .C2(n19348), .A(n16558), .B(n16557), .ZN(
        P2_U3004) );
  AOI22_X1 U19630 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n16616), .B1(n16583), 
        .B2(n19359), .ZN(n16563) );
  OAI22_X1 U19631 ( .A1(n16560), .A2(n16584), .B1(n16586), .B2(n16559), .ZN(
        n16561) );
  AOI21_X1 U19632 ( .B1(n16589), .B2(n19360), .A(n16561), .ZN(n16562) );
  OAI211_X1 U19633 ( .C1(n16593), .C2(n16564), .A(n16563), .B(n16562), .ZN(
        P2_U3005) );
  AOI22_X1 U19634 ( .A1(n19551), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n16616), .ZN(n16575) );
  NOR2_X1 U19635 ( .A1(n16566), .A2(n16565), .ZN(n16568) );
  XOR2_X1 U19636 ( .A(n16568), .B(n16567), .Z(n16650) );
  INV_X1 U19637 ( .A(n16650), .ZN(n16573) );
  NAND2_X1 U19638 ( .A1(n16570), .A2(n16569), .ZN(n16571) );
  AND2_X1 U19639 ( .A1(n16572), .A2(n16571), .ZN(n16647) );
  AOI222_X1 U19640 ( .A1(n19552), .A2(n16573), .B1(n16647), .B2(n19554), .C1(
        n16589), .C2(n16644), .ZN(n16574) );
  OAI211_X1 U19641 ( .C1(n19564), .C2(n16576), .A(n16575), .B(n16574), .ZN(
        P2_U3006) );
  AOI22_X1 U19642 ( .A1(n19551), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n16616), .ZN(n16582) );
  OAI22_X1 U19643 ( .A1(n16578), .A2(n16584), .B1(n19559), .B2(n16577), .ZN(
        n16579) );
  AOI21_X1 U19644 ( .B1(n19552), .B2(n16580), .A(n16579), .ZN(n16581) );
  OAI211_X1 U19645 ( .C1(n19564), .C2(n19369), .A(n16582), .B(n16581), .ZN(
        P2_U3008) );
  AOI22_X1 U19646 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n16616), .B1(n16583), 
        .B2(n19381), .ZN(n16591) );
  OAI22_X1 U19647 ( .A1(n16587), .A2(n16586), .B1(n16585), .B2(n16584), .ZN(
        n16588) );
  AOI21_X1 U19648 ( .B1(n16589), .B2(n19382), .A(n16588), .ZN(n16590) );
  OAI211_X1 U19649 ( .C1(n16593), .C2(n16592), .A(n16591), .B(n16590), .ZN(
        P2_U3009) );
  INV_X1 U19650 ( .A(n16594), .ZN(n16595) );
  NOR2_X1 U19651 ( .A1(n16595), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16596) );
  AOI22_X1 U19652 ( .A1(n16597), .A2(n16596), .B1(n16643), .B2(n19443), .ZN(
        n16607) );
  AOI222_X1 U19653 ( .A1(n16601), .A2(n16600), .B1(n16645), .B2(n16599), .C1(
        n16646), .C2(n16598), .ZN(n16606) );
  NAND2_X1 U19654 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n16616), .ZN(n16605) );
  OAI21_X1 U19655 ( .B1(n16603), .B2(n16602), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16604) );
  NAND4_X1 U19656 ( .A1(n16607), .A2(n16606), .A3(n16605), .A4(n16604), .ZN(
        P2_U3032) );
  OAI21_X1 U19657 ( .B1(n16610), .B2(n16609), .A(n16608), .ZN(n16611) );
  AOI22_X1 U19658 ( .A1(n16611), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16643), .B2(n19448), .ZN(n16620) );
  OAI22_X1 U19659 ( .A1(n16613), .A2(n16651), .B1(n16629), .B2(n16612), .ZN(
        n16614) );
  AOI21_X1 U19660 ( .B1(n16646), .B2(n16615), .A(n16614), .ZN(n16619) );
  NAND2_X1 U19661 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n16616), .ZN(n16617) );
  NAND4_X1 U19662 ( .A1(n16620), .A2(n16619), .A3(n16618), .A4(n16617), .ZN(
        P2_U3034) );
  NOR2_X1 U19663 ( .A1(n10577), .A2(n19333), .ZN(n16626) );
  XNOR2_X1 U19664 ( .A(n16622), .B(n16621), .ZN(n19455) );
  OAI22_X1 U19665 ( .A1(n16624), .A2(n19455), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16623), .ZN(n16625) );
  AOI211_X1 U19666 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16627), .A(
        n16626), .B(n16625), .ZN(n16634) );
  INV_X1 U19667 ( .A(n19350), .ZN(n16628) );
  OAI22_X1 U19668 ( .A1(n16631), .A2(n16630), .B1(n16629), .B2(n16628), .ZN(
        n16632) );
  INV_X1 U19669 ( .A(n16632), .ZN(n16633) );
  OAI211_X1 U19670 ( .C1(n16635), .C2(n16651), .A(n16634), .B(n16633), .ZN(
        P2_U3036) );
  NOR2_X1 U19671 ( .A1(n19364), .A2(n13912), .ZN(n16642) );
  OAI21_X1 U19672 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16636), .ZN(n16637) );
  OAI22_X1 U19673 ( .A1(n16640), .A2(n16639), .B1(n16638), .B2(n16637), .ZN(
        n16641) );
  AOI211_X1 U19674 ( .C1(n19458), .C2(n16643), .A(n16642), .B(n16641), .ZN(
        n16649) );
  AOI22_X1 U19675 ( .A1(n16647), .A2(n16646), .B1(n16645), .B2(n16644), .ZN(
        n16648) );
  OAI211_X1 U19676 ( .C1(n16651), .C2(n16650), .A(n16649), .B(n16648), .ZN(
        P2_U3038) );
  MUX2_X1 U19677 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16677), .S(
        n16685), .Z(n16696) );
  MUX2_X1 U19678 ( .A(n16653), .B(n16652), .S(n16685), .Z(n16676) );
  INV_X1 U19679 ( .A(n16676), .ZN(n16695) );
  INV_X1 U19680 ( .A(n16654), .ZN(n16657) );
  NOR3_X1 U19681 ( .A1(n16657), .A2(n16656), .A3(n16655), .ZN(n19238) );
  OAI21_X1 U19682 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19238), .ZN(n16661) );
  NAND3_X1 U19683 ( .A1(n10484), .A2(n16659), .A3(n16658), .ZN(n16660) );
  OAI211_X1 U19684 ( .C1(n16663), .C2(n16662), .A(n16661), .B(n16660), .ZN(
        n16673) );
  INV_X1 U19685 ( .A(n16664), .ZN(n16671) );
  OR2_X1 U19686 ( .A1(n16668), .A2(n16665), .ZN(n16670) );
  INV_X1 U19687 ( .A(n16666), .ZN(n16667) );
  NAND2_X1 U19688 ( .A1(n16668), .A2(n16667), .ZN(n16669) );
  OAI211_X1 U19689 ( .C1(n16672), .C2(n16671), .A(n16670), .B(n16669), .ZN(
        n20242) );
  NOR2_X1 U19690 ( .A1(n16673), .A2(n20242), .ZN(n16674) );
  OAI21_X1 U19691 ( .B1(n16675), .B2(n16685), .A(n16674), .ZN(n16694) );
  NOR2_X1 U19692 ( .A1(n16676), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16690) );
  AOI22_X1 U19693 ( .A1(n16690), .A2(n20219), .B1(n16696), .B2(n20209), .ZN(
        n16692) );
  INV_X1 U19694 ( .A(n16677), .ZN(n16688) );
  NAND2_X1 U19695 ( .A1(n9644), .A2(n16678), .ZN(n16682) );
  MUX2_X1 U19696 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n20194), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n16679) );
  AOI22_X1 U19697 ( .A1(n16680), .A2(n16679), .B1(n20194), .B2(n10503), .ZN(
        n16681) );
  NAND2_X1 U19698 ( .A1(n16682), .A2(n16681), .ZN(n20191) );
  NAND2_X1 U19699 ( .A1(n20191), .A2(n20229), .ZN(n16684) );
  NAND3_X1 U19700 ( .A1(n16684), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        n16683), .ZN(n16686) );
  OAI211_X1 U19701 ( .C1(n20229), .C2(n20191), .A(n16686), .B(n16685), .ZN(
        n16687) );
  AOI21_X1 U19702 ( .B1(n16688), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16687), .ZN(n16689) );
  OAI21_X1 U19703 ( .B1(n16690), .B2(n20219), .A(n16689), .ZN(n16691) );
  AOI21_X1 U19704 ( .B1(n16692), .B2(n16691), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16693) );
  AOI211_X1 U19705 ( .C1(n16696), .C2(n16695), .A(n16694), .B(n16693), .ZN(
        n16711) );
  AOI211_X1 U19706 ( .C1(n20243), .C2(n16699), .A(n16698), .B(n16697), .ZN(
        n16710) );
  NOR3_X1 U19707 ( .A1(n10672), .A2(n16701), .A3(n16700), .ZN(n16703) );
  INV_X1 U19708 ( .A(n20252), .ZN(n16702) );
  NOR3_X1 U19709 ( .A1(n16703), .A2(n16702), .A3(n19761), .ZN(n16707) );
  INV_X1 U19710 ( .A(n16707), .ZN(n16704) );
  NOR2_X1 U19711 ( .A1(n16704), .A2(n20257), .ZN(n20110) );
  AOI21_X1 U19712 ( .B1(n20190), .B2(n16705), .A(n20110), .ZN(n16708) );
  AOI21_X1 U19713 ( .B1(n16711), .B2(n10598), .A(n20256), .ZN(n16706) );
  INV_X1 U19714 ( .A(n16706), .ZN(n20109) );
  NAND2_X1 U19715 ( .A1(n20109), .A2(n16707), .ZN(n20111) );
  NAND2_X1 U19716 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20111), .ZN(n16712) );
  OAI21_X1 U19717 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16708), .A(n16712), 
        .ZN(n16709) );
  OAI211_X1 U19718 ( .C1(n16711), .C2(n19237), .A(n16710), .B(n16709), .ZN(
        P2_U3176) );
  INV_X1 U19719 ( .A(n16712), .ZN(n16714) );
  OAI21_X1 U19720 ( .B1(n16714), .B2(n20205), .A(n16713), .ZN(P2_U3593) );
  INV_X1 U19721 ( .A(n11318), .ZN(n18081) );
  NAND2_X1 U19722 ( .A1(n18213), .A2(n18021), .ZN(n17886) );
  INV_X1 U19723 ( .A(n17886), .ZN(n17931) );
  NAND2_X1 U19724 ( .A1(n16715), .A2(n17931), .ZN(n17874) );
  AOI21_X1 U19725 ( .B1(n16718), .B2(n16717), .A(n16716), .ZN(n16722) );
  OAI21_X1 U19726 ( .B1(n16731), .B2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16719), .ZN(n16901) );
  OAI21_X1 U19727 ( .B1(n18063), .B2(n16901), .A(n16720), .ZN(n16721) );
  NOR2_X1 U19728 ( .A1(n16724), .A2(n18211), .ZN(n16741) );
  INV_X1 U19729 ( .A(n18058), .ZN(n18119) );
  AND2_X1 U19730 ( .A1(n16725), .A2(n18119), .ZN(n16730) );
  OAI21_X1 U19731 ( .B1(n16741), .B2(n16730), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16726) );
  OAI211_X1 U19732 ( .C1(n16728), .C2(n17874), .A(n16727), .B(n16726), .ZN(
        P3_U2800) );
  NOR2_X1 U19733 ( .A1(n18218), .A2(n16729), .ZN(n16748) );
  INV_X1 U19734 ( .A(n18220), .ZN(n17864) );
  NOR2_X1 U19735 ( .A1(n16729), .A2(n17864), .ZN(n16747) );
  OAI21_X1 U19736 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16747), .A(
        n16730), .ZN(n16738) );
  INV_X1 U19737 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16732) );
  AOI21_X1 U19738 ( .B1(n16732), .B2(n16884), .A(n16731), .ZN(n16910) );
  OAI21_X1 U19739 ( .B1(n17970), .B2(n16733), .A(n16910), .ZN(n16737) );
  OAI221_X1 U19740 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16735), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18932), .A(n16734), .ZN(
        n16736) );
  NAND4_X1 U19741 ( .A1(n16739), .A2(n16738), .A3(n16737), .A4(n16736), .ZN(
        n16740) );
  AOI221_X1 U19742 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16741), 
        .C1(n16748), .C2(n16741), .A(n16740), .ZN(n16742) );
  OAI21_X1 U19743 ( .B1(n16743), .B2(n18122), .A(n16742), .ZN(P3_U2801) );
  NAND2_X1 U19744 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16744), .ZN(
        n17870) );
  NAND2_X1 U19745 ( .A1(n10177), .A2(n18354), .ZN(n16752) );
  NOR2_X1 U19746 ( .A1(n18987), .A2(n16746), .ZN(n18272) );
  OAI22_X1 U19747 ( .A1(n16748), .A2(n18501), .B1(n16747), .B2(n18401), .ZN(
        n16750) );
  INV_X1 U19748 ( .A(n18343), .ZN(n18271) );
  OAI22_X1 U19749 ( .A1(n18501), .A2(n18273), .B1(n18271), .B2(n18401), .ZN(
        n18314) );
  INV_X1 U19750 ( .A(n18212), .ZN(n18317) );
  OAI22_X1 U19751 ( .A1(n19023), .A2(n18253), .B1(n18317), .B2(n18491), .ZN(
        n18238) );
  NOR2_X1 U19752 ( .A1(n18293), .A2(n18276), .ZN(n18270) );
  NAND2_X1 U19753 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18270), .ZN(
        n18264) );
  NOR2_X1 U19754 ( .A1(n17887), .A2(n18264), .ZN(n18231) );
  NAND2_X1 U19755 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18231), .ZN(
        n18221) );
  NOR4_X1 U19756 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n11149), .A3(
        n18510), .A4(n18221), .ZN(n16753) );
  NAND3_X1 U19757 ( .A1(n16754), .A2(n18525), .A3(n17856), .ZN(n16756) );
  NAND3_X1 U19758 ( .A1(n17857), .A2(n17869), .A3(n9631), .ZN(n16755) );
  NAND3_X1 U19759 ( .A1(n16757), .A2(n16756), .A3(n16755), .ZN(P3_U2834) );
  NOR3_X1 U19760 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16759) );
  NOR4_X1 U19761 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16758) );
  NAND4_X1 U19762 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16759), .A3(n16758), .A4(
        U215), .ZN(U213) );
  INV_X1 U19763 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19505) );
  INV_X2 U19764 ( .A(U214), .ZN(n16814) );
  INV_X1 U19765 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16852) );
  OAI222_X1 U19766 ( .A1(U212), .A2(n19505), .B1(n16817), .B2(n19612), .C1(
        U214), .C2(n16852), .ZN(U216) );
  INV_X1 U19767 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16761) );
  INV_X1 U19768 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19510) );
  OAI222_X1 U19769 ( .A1(U214), .A2(n16761), .B1(n16817), .B2(n19601), .C1(
        U212), .C2(n19510), .ZN(U217) );
  INV_X2 U19770 ( .A(U212), .ZN(n16815) );
  AOI22_X1 U19771 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16814), .ZN(n16762) );
  OAI21_X1 U19772 ( .B1(n16763), .B2(n16817), .A(n16762), .ZN(U218) );
  AOI22_X1 U19773 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16814), .ZN(n16764) );
  OAI21_X1 U19774 ( .B1(n16765), .B2(n16817), .A(n16764), .ZN(U219) );
  AOI22_X1 U19775 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16814), .ZN(n16766) );
  OAI21_X1 U19776 ( .B1(n19586), .B2(n16817), .A(n16766), .ZN(U220) );
  AOI22_X1 U19777 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16814), .ZN(n16767) );
  OAI21_X1 U19778 ( .B1(n16768), .B2(n16817), .A(n16767), .ZN(U221) );
  AOI22_X1 U19779 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16814), .ZN(n16769) );
  OAI21_X1 U19780 ( .B1(n16770), .B2(n16817), .A(n16769), .ZN(U222) );
  AOI22_X1 U19781 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16814), .ZN(n16771) );
  OAI21_X1 U19782 ( .B1(n16772), .B2(n16817), .A(n16771), .ZN(U223) );
  AOI22_X1 U19783 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16814), .ZN(n16773) );
  OAI21_X1 U19784 ( .B1(n16774), .B2(n16817), .A(n16773), .ZN(U224) );
  AOI22_X1 U19785 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16814), .ZN(n16775) );
  OAI21_X1 U19786 ( .B1(n16776), .B2(n16817), .A(n16775), .ZN(U225) );
  AOI22_X1 U19787 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16814), .ZN(n16777) );
  OAI21_X1 U19788 ( .B1(n19595), .B2(n16817), .A(n16777), .ZN(U226) );
  AOI22_X1 U19789 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16814), .ZN(n16778) );
  OAI21_X1 U19790 ( .B1(n16779), .B2(n16817), .A(n16778), .ZN(U227) );
  AOI22_X1 U19791 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16814), .ZN(n16780) );
  OAI21_X1 U19792 ( .B1(n16781), .B2(n16817), .A(n16780), .ZN(U228) );
  AOI22_X1 U19793 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16814), .ZN(n16782) );
  OAI21_X1 U19794 ( .B1(n19582), .B2(n16817), .A(n16782), .ZN(U229) );
  AOI22_X1 U19795 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16814), .ZN(n16783) );
  OAI21_X1 U19796 ( .B1(n19576), .B2(n16817), .A(n16783), .ZN(U230) );
  AOI22_X1 U19797 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16814), .ZN(n16784) );
  OAI21_X1 U19798 ( .B1(n16785), .B2(n16817), .A(n16784), .ZN(U231) );
  AOI22_X1 U19799 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16814), .ZN(n16786) );
  OAI21_X1 U19800 ( .B1(n13249), .B2(n16817), .A(n16786), .ZN(U232) );
  AOI22_X1 U19801 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16814), .ZN(n16787) );
  OAI21_X1 U19802 ( .B1(n16788), .B2(n16817), .A(n16787), .ZN(U233) );
  AOI22_X1 U19803 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16814), .ZN(n16789) );
  OAI21_X1 U19804 ( .B1(n16790), .B2(n16817), .A(n16789), .ZN(U234) );
  AOI22_X1 U19805 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16814), .ZN(n16791) );
  OAI21_X1 U19806 ( .B1(n16792), .B2(n16817), .A(n16791), .ZN(U235) );
  AOI22_X1 U19807 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16814), .ZN(n16793) );
  OAI21_X1 U19808 ( .B1(n12993), .B2(n16817), .A(n16793), .ZN(U236) );
  AOI22_X1 U19809 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16814), .ZN(n16794) );
  OAI21_X1 U19810 ( .B1(n16795), .B2(n16817), .A(n16794), .ZN(U237) );
  AOI22_X1 U19811 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16814), .ZN(n16796) );
  OAI21_X1 U19812 ( .B1(n16797), .B2(n16817), .A(n16796), .ZN(U238) );
  AOI22_X1 U19813 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16814), .ZN(n16798) );
  OAI21_X1 U19814 ( .B1(n16799), .B2(n16817), .A(n16798), .ZN(U239) );
  INV_X1 U19815 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16801) );
  AOI22_X1 U19816 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16814), .ZN(n16800) );
  OAI21_X1 U19817 ( .B1(n16801), .B2(n16817), .A(n16800), .ZN(U240) );
  AOI22_X1 U19818 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16814), .ZN(n16802) );
  OAI21_X1 U19819 ( .B1(n16803), .B2(n16817), .A(n16802), .ZN(U241) );
  AOI22_X1 U19820 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16814), .ZN(n16804) );
  OAI21_X1 U19821 ( .B1(n16805), .B2(n16817), .A(n16804), .ZN(U242) );
  AOI22_X1 U19822 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16814), .ZN(n16806) );
  OAI21_X1 U19823 ( .B1(n16807), .B2(n16817), .A(n16806), .ZN(U243) );
  INV_X1 U19824 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16809) );
  AOI22_X1 U19825 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16814), .ZN(n16808) );
  OAI21_X1 U19826 ( .B1(n16809), .B2(n16817), .A(n16808), .ZN(U244) );
  AOI22_X1 U19827 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16814), .ZN(n16810) );
  OAI21_X1 U19828 ( .B1(n16811), .B2(n16817), .A(n16810), .ZN(U245) );
  AOI22_X1 U19829 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16814), .ZN(n16812) );
  OAI21_X1 U19830 ( .B1(n16813), .B2(n16817), .A(n16812), .ZN(U246) );
  AOI22_X1 U19831 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16815), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16814), .ZN(n16816) );
  OAI21_X1 U19832 ( .B1(n16818), .B2(n16817), .A(n16816), .ZN(U247) );
  OAI22_X1 U19833 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16850), .ZN(n16819) );
  INV_X1 U19834 ( .A(n16819), .ZN(U251) );
  OAI22_X1 U19835 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16850), .ZN(n16820) );
  INV_X1 U19836 ( .A(n16820), .ZN(U252) );
  INV_X1 U19837 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16821) );
  AOI22_X1 U19838 ( .A1(n16845), .A2(n16821), .B1(n18556), .B2(U215), .ZN(U253) );
  OAI22_X1 U19839 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16850), .ZN(n16822) );
  INV_X1 U19840 ( .A(n16822), .ZN(U254) );
  INV_X1 U19841 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16823) );
  INV_X1 U19842 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18566) );
  AOI22_X1 U19843 ( .A1(n16850), .A2(n16823), .B1(n18566), .B2(U215), .ZN(U255) );
  INV_X1 U19844 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16824) );
  INV_X1 U19845 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18572) );
  AOI22_X1 U19846 ( .A1(n16850), .A2(n16824), .B1(n18572), .B2(U215), .ZN(U256) );
  INV_X1 U19847 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16825) );
  INV_X1 U19848 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18577) );
  AOI22_X1 U19849 ( .A1(n16850), .A2(n16825), .B1(n18577), .B2(U215), .ZN(U257) );
  INV_X1 U19850 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16826) );
  INV_X1 U19851 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18583) );
  AOI22_X1 U19852 ( .A1(n16845), .A2(n16826), .B1(n18583), .B2(U215), .ZN(U258) );
  INV_X1 U19853 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16827) );
  INV_X1 U19854 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17710) );
  AOI22_X1 U19855 ( .A1(n16850), .A2(n16827), .B1(n17710), .B2(U215), .ZN(U259) );
  INV_X1 U19856 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16828) );
  INV_X1 U19857 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U19858 ( .A1(n16850), .A2(n16828), .B1(n17704), .B2(U215), .ZN(U260) );
  INV_X1 U19859 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16829) );
  INV_X1 U19860 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17698) );
  AOI22_X1 U19861 ( .A1(n16845), .A2(n16829), .B1(n17698), .B2(U215), .ZN(U261) );
  INV_X1 U19862 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16830) );
  INV_X1 U19863 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17693) );
  AOI22_X1 U19864 ( .A1(n16845), .A2(n16830), .B1(n17693), .B2(U215), .ZN(U262) );
  INV_X1 U19865 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16831) );
  INV_X1 U19866 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17689) );
  AOI22_X1 U19867 ( .A1(n16850), .A2(n16831), .B1(n17689), .B2(U215), .ZN(U263) );
  INV_X1 U19868 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16832) );
  INV_X1 U19869 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17684) );
  AOI22_X1 U19870 ( .A1(n16845), .A2(n16832), .B1(n17684), .B2(U215), .ZN(U264) );
  OAI22_X1 U19871 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16850), .ZN(n16833) );
  INV_X1 U19872 ( .A(n16833), .ZN(U265) );
  OAI22_X1 U19873 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16850), .ZN(n16834) );
  INV_X1 U19874 ( .A(n16834), .ZN(U266) );
  OAI22_X1 U19875 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16850), .ZN(n16835) );
  INV_X1 U19876 ( .A(n16835), .ZN(U267) );
  INV_X1 U19877 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16836) );
  AOI22_X1 U19878 ( .A1(n16850), .A2(n16836), .B1(n14163), .B2(U215), .ZN(U268) );
  INV_X1 U19879 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16837) );
  INV_X1 U19880 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19581) );
  AOI22_X1 U19881 ( .A1(n16845), .A2(n16837), .B1(n19581), .B2(U215), .ZN(U269) );
  OAI22_X1 U19882 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16850), .ZN(n16838) );
  INV_X1 U19883 ( .A(n16838), .ZN(U270) );
  INV_X1 U19884 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16839) );
  AOI22_X1 U19885 ( .A1(n16845), .A2(n16839), .B1(n18565), .B2(U215), .ZN(U271) );
  INV_X1 U19886 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16840) );
  INV_X1 U19887 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19594) );
  AOI22_X1 U19888 ( .A1(n16850), .A2(n16840), .B1(n19594), .B2(U215), .ZN(U272) );
  INV_X1 U19889 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16841) );
  AOI22_X1 U19890 ( .A1(n16850), .A2(n16841), .B1(n15542), .B2(U215), .ZN(U273) );
  OAI22_X1 U19891 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16845), .ZN(n16842) );
  INV_X1 U19892 ( .A(n16842), .ZN(U274) );
  INV_X1 U19893 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16843) );
  AOI22_X1 U19894 ( .A1(n16850), .A2(n16843), .B1(n18546), .B2(U215), .ZN(U275) );
  OAI22_X1 U19895 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16845), .ZN(n16844) );
  INV_X1 U19896 ( .A(n16844), .ZN(U276) );
  OAI22_X1 U19897 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16845), .ZN(n16846) );
  INV_X1 U19898 ( .A(n16846), .ZN(U277) );
  INV_X1 U19899 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16847) );
  AOI22_X1 U19900 ( .A1(n16850), .A2(n16847), .B1(n15503), .B2(U215), .ZN(U278) );
  OAI22_X1 U19901 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16850), .ZN(n16848) );
  INV_X1 U19902 ( .A(n16848), .ZN(U279) );
  OAI22_X1 U19903 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16850), .ZN(n16849) );
  INV_X1 U19904 ( .A(n16849), .ZN(U280) );
  INV_X1 U19905 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19602) );
  AOI22_X1 U19906 ( .A1(n16850), .A2(n19510), .B1(n19602), .B2(U215), .ZN(U281) );
  INV_X1 U19907 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19610) );
  AOI22_X1 U19908 ( .A1(n16850), .A2(n19505), .B1(n19610), .B2(U215), .ZN(U282) );
  INV_X1 U19909 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16851) );
  AOI222_X1 U19910 ( .A1(n19505), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16852), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16851), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16853) );
  INV_X1 U19911 ( .A(n16855), .ZN(n16854) );
  INV_X1 U19912 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19100) );
  INV_X1 U19913 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20144) );
  AOI22_X1 U19914 ( .A1(n16854), .A2(n19100), .B1(n20144), .B2(n16855), .ZN(
        U347) );
  INV_X1 U19915 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19098) );
  INV_X1 U19916 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20143) );
  AOI22_X1 U19917 ( .A1(n16854), .A2(n19098), .B1(n20143), .B2(n16855), .ZN(
        U348) );
  INV_X1 U19918 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19095) );
  INV_X1 U19919 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20142) );
  AOI22_X1 U19920 ( .A1(n16854), .A2(n19095), .B1(n20142), .B2(n16855), .ZN(
        U349) );
  INV_X1 U19921 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19094) );
  INV_X1 U19922 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20141) );
  AOI22_X1 U19923 ( .A1(n16854), .A2(n19094), .B1(n20141), .B2(n16855), .ZN(
        U350) );
  INV_X1 U19924 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19092) );
  INV_X1 U19925 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20140) );
  AOI22_X1 U19926 ( .A1(n16854), .A2(n19092), .B1(n20140), .B2(n16855), .ZN(
        U351) );
  INV_X1 U19927 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19089) );
  INV_X1 U19928 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20139) );
  AOI22_X1 U19929 ( .A1(n16854), .A2(n19089), .B1(n20139), .B2(n16855), .ZN(
        U352) );
  INV_X1 U19930 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19088) );
  INV_X1 U19931 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20138) );
  AOI22_X1 U19932 ( .A1(n16854), .A2(n19088), .B1(n20138), .B2(n16855), .ZN(
        U353) );
  INV_X1 U19933 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19086) );
  AOI22_X1 U19934 ( .A1(n16854), .A2(n19086), .B1(n20137), .B2(n16855), .ZN(
        U354) );
  INV_X1 U19935 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19139) );
  INV_X1 U19936 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20172) );
  AOI22_X1 U19937 ( .A1(n16854), .A2(n19139), .B1(n20172), .B2(n16855), .ZN(
        U356) );
  INV_X1 U19938 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19135) );
  INV_X1 U19939 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20170) );
  AOI22_X1 U19940 ( .A1(n16854), .A2(n19135), .B1(n20170), .B2(n16855), .ZN(
        U357) );
  INV_X1 U19941 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19134) );
  INV_X1 U19942 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20167) );
  AOI22_X1 U19943 ( .A1(n16854), .A2(n19134), .B1(n20167), .B2(n16855), .ZN(
        U358) );
  INV_X1 U19944 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19132) );
  INV_X1 U19945 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20166) );
  AOI22_X1 U19946 ( .A1(n16854), .A2(n19132), .B1(n20166), .B2(n16855), .ZN(
        U359) );
  INV_X1 U19947 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19130) );
  INV_X1 U19948 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20165) );
  AOI22_X1 U19949 ( .A1(n16854), .A2(n19130), .B1(n20165), .B2(n16855), .ZN(
        U360) );
  INV_X1 U19950 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19128) );
  INV_X1 U19951 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20163) );
  AOI22_X1 U19952 ( .A1(n16854), .A2(n19128), .B1(n20163), .B2(n16855), .ZN(
        U361) );
  INV_X1 U19953 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19126) );
  INV_X1 U19954 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20161) );
  AOI22_X1 U19955 ( .A1(n16854), .A2(n19126), .B1(n20161), .B2(n16855), .ZN(
        U362) );
  INV_X1 U19956 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19124) );
  INV_X1 U19957 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20159) );
  AOI22_X1 U19958 ( .A1(n16854), .A2(n19124), .B1(n20159), .B2(n16855), .ZN(
        U363) );
  INV_X1 U19959 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19122) );
  INV_X1 U19960 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20158) );
  AOI22_X1 U19961 ( .A1(n16854), .A2(n19122), .B1(n20158), .B2(n16855), .ZN(
        U364) );
  INV_X1 U19962 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19084) );
  INV_X1 U19963 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20135) );
  AOI22_X1 U19964 ( .A1(n16854), .A2(n19084), .B1(n20135), .B2(n16855), .ZN(
        U365) );
  INV_X1 U19965 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19119) );
  INV_X1 U19966 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20156) );
  AOI22_X1 U19967 ( .A1(n16854), .A2(n19119), .B1(n20156), .B2(n16855), .ZN(
        U366) );
  INV_X1 U19968 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19118) );
  INV_X1 U19969 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20155) );
  AOI22_X1 U19970 ( .A1(n16854), .A2(n19118), .B1(n20155), .B2(n16855), .ZN(
        U367) );
  INV_X1 U19971 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19116) );
  INV_X1 U19972 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20153) );
  AOI22_X1 U19973 ( .A1(n16854), .A2(n19116), .B1(n20153), .B2(n16855), .ZN(
        U368) );
  INV_X1 U19974 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19113) );
  INV_X1 U19975 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20152) );
  AOI22_X1 U19976 ( .A1(n16854), .A2(n19113), .B1(n20152), .B2(n16855), .ZN(
        U369) );
  INV_X1 U19977 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19112) );
  INV_X1 U19978 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20150) );
  AOI22_X1 U19979 ( .A1(n16854), .A2(n19112), .B1(n20150), .B2(n16855), .ZN(
        U370) );
  INV_X1 U19980 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19110) );
  INV_X1 U19981 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20149) );
  AOI22_X1 U19982 ( .A1(n16854), .A2(n19110), .B1(n20149), .B2(n16855), .ZN(
        U371) );
  INV_X1 U19983 ( .A(n16855), .ZN(n21255) );
  INV_X1 U19984 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19107) );
  INV_X1 U19985 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20148) );
  AOI22_X1 U19986 ( .A1(n21255), .A2(n19107), .B1(n20148), .B2(n16855), .ZN(
        U372) );
  INV_X1 U19987 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19106) );
  INV_X1 U19988 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20147) );
  AOI22_X1 U19989 ( .A1(n21255), .A2(n19106), .B1(n20147), .B2(n16855), .ZN(
        U373) );
  INV_X1 U19990 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19104) );
  INV_X1 U19991 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20146) );
  AOI22_X1 U19992 ( .A1(n21255), .A2(n19104), .B1(n20146), .B2(n16855), .ZN(
        U374) );
  INV_X1 U19993 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19102) );
  INV_X1 U19994 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20145) );
  AOI22_X1 U19995 ( .A1(n21255), .A2(n19102), .B1(n20145), .B2(n16855), .ZN(
        U375) );
  INV_X1 U19996 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19082) );
  INV_X1 U19997 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20134) );
  AOI22_X1 U19998 ( .A1(n21255), .A2(n19082), .B1(n20134), .B2(n16855), .ZN(
        U376) );
  INV_X1 U19999 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16857) );
  AND2_X1 U20000 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19081), .ZN(n16856) );
  MUX2_X1 U20001 ( .A(n19073), .B(n16856), .S(P3_STATE_REG_0__SCAN_IN), .Z(
        n19156) );
  OAI21_X1 U20002 ( .B1(n19079), .B2(n16857), .A(n9633), .ZN(P3_U2633) );
  NAND2_X1 U20003 ( .A1(n19206), .A2(n18986), .ZN(n17783) );
  OAI21_X1 U20004 ( .B1(n16864), .B2(n17783), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16858) );
  OAI21_X1 U20005 ( .B1(n16859), .B2(n19055), .A(n16858), .ZN(P3_U2634) );
  AOI21_X1 U20006 ( .B1(n19079), .B2(n19081), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16860) );
  AOI22_X1 U20007 ( .A1(n19151), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16860), 
        .B2(n19220), .ZN(P3_U2635) );
  INV_X1 U20008 ( .A(BS16), .ZN(n21089) );
  AOI21_X1 U20009 ( .B1(n16861), .B2(n21089), .A(n9633), .ZN(n19152) );
  INV_X1 U20010 ( .A(n19152), .ZN(n19154) );
  OAI21_X1 U20011 ( .B1(n19156), .B2(n19211), .A(n19154), .ZN(P3_U2636) );
  NOR3_X1 U20012 ( .A1(n16864), .A2(n16863), .A3(n16862), .ZN(n19040) );
  NOR2_X1 U20013 ( .A1(n19040), .A2(n19044), .ZN(n19201) );
  INV_X1 U20014 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16866) );
  OAI21_X1 U20015 ( .B1(n19201), .B2(n16866), .A(n16865), .ZN(P3_U2637) );
  NOR4_X1 U20016 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16870) );
  NOR4_X1 U20017 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16869) );
  NOR4_X1 U20018 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16868) );
  NOR4_X1 U20019 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16867) );
  NAND4_X1 U20020 ( .A1(n16870), .A2(n16869), .A3(n16868), .A4(n16867), .ZN(
        n16876) );
  NOR4_X1 U20021 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16874) );
  AOI211_X1 U20022 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16873) );
  NOR4_X1 U20023 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16872) );
  NOR4_X1 U20024 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16871) );
  NAND4_X1 U20025 ( .A1(n16874), .A2(n16873), .A3(n16872), .A4(n16871), .ZN(
        n16875) );
  NOR2_X1 U20026 ( .A1(n16876), .A2(n16875), .ZN(n19195) );
  INV_X1 U20027 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19149) );
  NOR3_X1 U20028 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16878) );
  OAI21_X1 U20029 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16878), .A(n19195), .ZN(
        n16877) );
  OAI21_X1 U20030 ( .B1(n19195), .B2(n19149), .A(n16877), .ZN(P3_U2638) );
  INV_X1 U20031 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19191) );
  INV_X1 U20032 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19155) );
  AOI21_X1 U20033 ( .B1(n19191), .B2(n19155), .A(n16878), .ZN(n16879) );
  INV_X1 U20034 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19146) );
  INV_X1 U20035 ( .A(n19195), .ZN(n19198) );
  AOI22_X1 U20036 ( .A1(n19195), .A2(n16879), .B1(n19146), .B2(n19198), .ZN(
        P3_U2639) );
  NAND3_X1 U20037 ( .A1(n19052), .A2(n19222), .A3(n19211), .ZN(n19063) );
  NOR2_X2 U20038 ( .A1(n19171), .A2(n19063), .ZN(n17210) );
  NAND2_X1 U20039 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19222), .ZN(n19056) );
  NOR2_X1 U20040 ( .A1(n19055), .A2(n19056), .ZN(n19048) );
  NOR4_X2 U20041 ( .A1(n18483), .A2(n19226), .A3(n17210), .A4(n19048), .ZN(
        n17252) );
  NOR2_X2 U20042 ( .A1(n17252), .A2(n19160), .ZN(n17242) );
  AOI211_X1 U20043 ( .C1(n19210), .C2(n19212), .A(n19208), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n19045) );
  NAND2_X1 U20044 ( .A1(n19226), .A2(n18545), .ZN(n16880) );
  AOI211_X4 U20045 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18551), .A(n19045), .B(
        n16880), .ZN(n17259) );
  AOI22_X1 U20046 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n17242), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n17259), .ZN(n16899) );
  INV_X1 U20047 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19138) );
  NAND2_X1 U20048 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16917) );
  INV_X1 U20049 ( .A(n17252), .ZN(n17257) );
  INV_X1 U20050 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19131) );
  INV_X1 U20051 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19127) );
  INV_X1 U20052 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19103) );
  INV_X1 U20053 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19096) );
  INV_X1 U20054 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19087) );
  NAND3_X1 U20055 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17213) );
  NOR2_X1 U20056 ( .A1(n19087), .A2(n17213), .ZN(n17185) );
  NAND2_X1 U20057 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17185), .ZN(n17166) );
  NAND2_X1 U20058 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n17145) );
  NOR3_X1 U20059 ( .A1(n19096), .A2(n17166), .A3(n17145), .ZN(n17084) );
  NAND4_X1 U20060 ( .A1(n17084), .A2(P3_REIP_REG_11__SCAN_IN), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n17105) );
  NOR2_X1 U20061 ( .A1(n19103), .A2(n17105), .ZN(n17074) );
  NAND3_X1 U20062 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17074), .ZN(n17019) );
  NAND3_X1 U20063 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n17011) );
  NAND2_X1 U20064 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n17012) );
  NOR2_X1 U20065 ( .A1(n17011), .A2(n17012), .ZN(n17008) );
  NAND2_X1 U20066 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17008), .ZN(n16967) );
  NOR2_X1 U20067 ( .A1(n17019), .A2(n16967), .ZN(n16980) );
  NAND4_X1 U20068 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16980), .A3(
        P3_REIP_REG_22__SCAN_IN), .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n16947) );
  NOR2_X1 U20069 ( .A1(n19127), .A2(n16947), .ZN(n16953) );
  NAND2_X1 U20070 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16953), .ZN(n16946) );
  NOR2_X1 U20071 ( .A1(n19131), .A2(n16946), .ZN(n16894) );
  OR2_X1 U20072 ( .A1(n16894), .A2(n17245), .ZN(n16945) );
  NAND2_X1 U20073 ( .A1(n17257), .A2(n16945), .ZN(n16942) );
  AOI221_X1 U20074 ( .B1(n17237), .B2(n19138), .C1(n17237), .C2(n16917), .A(
        n16942), .ZN(n16881) );
  INV_X1 U20075 ( .A(n16881), .ZN(n16913) );
  NAND2_X1 U20076 ( .A1(n19211), .A2(n19213), .ZN(n16882) );
  NOR3_X1 U20077 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17241) );
  INV_X1 U20078 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17221) );
  NAND2_X1 U20079 ( .A1(n17241), .A2(n17221), .ZN(n17219) );
  NOR2_X1 U20080 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17219), .ZN(n17203) );
  INV_X1 U20081 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17565) );
  NAND2_X1 U20082 ( .A1(n17203), .A2(n17565), .ZN(n17186) );
  NOR2_X1 U20083 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17186), .ZN(n17175) );
  INV_X1 U20084 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17165) );
  NAND2_X1 U20085 ( .A1(n17175), .A2(n17165), .ZN(n17164) );
  NOR2_X1 U20086 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17164), .ZN(n17144) );
  INV_X1 U20087 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17139) );
  NAND2_X1 U20088 ( .A1(n17144), .A2(n17139), .ZN(n17137) );
  NOR2_X1 U20089 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17137), .ZN(n17125) );
  INV_X1 U20090 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17118) );
  NAND2_X1 U20091 ( .A1(n17125), .A2(n17118), .ZN(n17117) );
  NOR2_X1 U20092 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17117), .ZN(n17099) );
  INV_X1 U20093 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17090) );
  NAND2_X1 U20094 ( .A1(n17099), .A2(n17090), .ZN(n17089) );
  NOR2_X1 U20095 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17089), .ZN(n17073) );
  INV_X1 U20096 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17068) );
  NAND2_X1 U20097 ( .A1(n17073), .A2(n17068), .ZN(n17065) );
  NOR2_X1 U20098 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17065), .ZN(n17050) );
  INV_X1 U20099 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17049) );
  NAND2_X1 U20100 ( .A1(n17050), .A2(n17049), .ZN(n17046) );
  NOR2_X1 U20101 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17046), .ZN(n17029) );
  INV_X1 U20102 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17015) );
  NAND2_X1 U20103 ( .A1(n17029), .A2(n17015), .ZN(n17013) );
  NOR2_X1 U20104 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17013), .ZN(n17004) );
  NAND2_X1 U20105 ( .A1(n17004), .A2(n17343), .ZN(n16996) );
  NOR2_X1 U20106 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16996), .ZN(n16978) );
  NAND2_X1 U20107 ( .A1(n16978), .A2(n16975), .ZN(n16974) );
  NOR2_X1 U20108 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16974), .ZN(n16960) );
  NAND2_X1 U20109 ( .A1(n16960), .A2(n17265), .ZN(n16952) );
  NOR2_X1 U20110 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16952), .ZN(n16936) );
  INV_X1 U20111 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17307) );
  NAND2_X1 U20112 ( .A1(n16936), .A2(n17307), .ZN(n16932) );
  NOR2_X1 U20113 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16932), .ZN(n16918) );
  INV_X1 U20114 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16916) );
  NAND2_X1 U20115 ( .A1(n16918), .A2(n16916), .ZN(n16900) );
  NOR2_X1 U20116 ( .A1(n17249), .A2(n16900), .ZN(n16902) );
  INV_X1 U20117 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U20118 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n16913), .B1(n16902), 
        .B2(n17270), .ZN(n16898) );
  OAI21_X1 U20119 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16892), .A(
        n16884), .ZN(n17862) );
  INV_X1 U20120 ( .A(n17862), .ZN(n16921) );
  OAI21_X1 U20121 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17853), .A(
        n16893), .ZN(n17885) );
  INV_X1 U20122 ( .A(n17885), .ZN(n16939) );
  INV_X1 U20123 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17916) );
  NOR2_X1 U20124 ( .A1(n17916), .A2(n16888), .ZN(n16891) );
  AOI21_X1 U20125 ( .B1(n17916), .B2(n16888), .A(n16891), .ZN(n17912) );
  AOI21_X1 U20126 ( .B1(n16990), .B2(n16886), .A(n17895), .ZN(n17936) );
  AOI21_X1 U20127 ( .B1(n10002), .B2(n17017), .A(n16887), .ZN(n17969) );
  INV_X1 U20128 ( .A(n17017), .ZN(n17934) );
  INV_X1 U20129 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17075) );
  INV_X1 U20130 ( .A(n18053), .ZN(n17076) );
  NOR2_X1 U20131 ( .A1(n18202), .A2(n18051), .ZN(n18050) );
  NAND2_X1 U20132 ( .A1(n17076), .A2(n18050), .ZN(n17086) );
  NOR2_X1 U20133 ( .A1(n17075), .A2(n17086), .ZN(n18013) );
  NAND2_X1 U20134 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18013), .ZN(
        n17061) );
  NOR2_X1 U20135 ( .A1(n17000), .A2(n17158), .ZN(n16992) );
  OAI21_X1 U20136 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n16887), .A(
        n16886), .ZN(n17949) );
  INV_X1 U20137 ( .A(n17949), .ZN(n16993) );
  NOR2_X1 U20138 ( .A1(n16991), .A2(n17158), .ZN(n16985) );
  NOR2_X1 U20139 ( .A1(n16984), .A2(n17158), .ZN(n16969) );
  OAI21_X1 U20140 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17895), .A(
        n16888), .ZN(n16889) );
  INV_X1 U20141 ( .A(n16889), .ZN(n17924) );
  NOR2_X1 U20142 ( .A1(n16968), .A2(n17158), .ZN(n16962) );
  NOR2_X1 U20143 ( .A1(n16961), .A2(n17158), .ZN(n16949) );
  INV_X1 U20144 ( .A(n17853), .ZN(n16890) );
  OAI21_X1 U20145 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16891), .A(
        n16890), .ZN(n17901) );
  INV_X1 U20146 ( .A(n17901), .ZN(n16950) );
  NOR2_X1 U20147 ( .A1(n16948), .A2(n17158), .ZN(n16938) );
  NOR2_X1 U20148 ( .A1(n16937), .A2(n17158), .ZN(n16928) );
  AOI21_X1 U20149 ( .B1(n17872), .B2(n16893), .A(n16892), .ZN(n17868) );
  NOR2_X1 U20150 ( .A1(n16927), .A2(n17158), .ZN(n16920) );
  NOR2_X1 U20151 ( .A1(n16921), .A2(n16920), .ZN(n16919) );
  NOR2_X1 U20152 ( .A1(n16919), .A2(n17158), .ZN(n16909) );
  NAND4_X1 U20153 ( .A1(n16885), .A2(n17210), .A3(n16908), .A4(n16901), .ZN(
        n16897) );
  INV_X1 U20154 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19143) );
  NAND2_X1 U20155 ( .A1(n17237), .A2(n16894), .ZN(n16929) );
  NOR2_X1 U20156 ( .A1(n16917), .A2(n16929), .ZN(n16905) );
  NAND2_X1 U20157 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16905), .ZN(n16904) );
  INV_X1 U20158 ( .A(n16904), .ZN(n16895) );
  OAI221_X1 U20159 ( .B1(P3_REIP_REG_31__SCAN_IN), .B2(P3_REIP_REG_30__SCAN_IN), .C1(n19141), .C2(n19143), .A(n16895), .ZN(n16896) );
  NAND4_X1 U20160 ( .A1(n16899), .A2(n16898), .A3(n16897), .A4(n16896), .ZN(
        P3_U2640) );
  AOI22_X1 U20161 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n17242), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n16913), .ZN(n16903) );
  NAND2_X1 U20162 ( .A1(n17258), .A2(n16900), .ZN(n16906) );
  INV_X1 U20163 ( .A(n17210), .ZN(n19061) );
  AOI22_X1 U20164 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17242), .B1(
        n16905), .B2(n19138), .ZN(n16915) );
  INV_X1 U20165 ( .A(n16918), .ZN(n16907) );
  AOI21_X1 U20166 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16907), .A(n16906), .ZN(
        n16912) );
  AOI211_X1 U20167 ( .C1(n16910), .C2(n16909), .A(n16908), .B(n19061), .ZN(
        n16911) );
  AOI211_X1 U20168 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16913), .A(n16912), 
        .B(n16911), .ZN(n16914) );
  OAI211_X1 U20169 ( .C1(n17244), .C2(n16916), .A(n16915), .B(n16914), .ZN(
        P3_U2642) );
  OAI21_X1 U20170 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(P3_REIP_REG_27__SCAN_IN), 
        .A(n16917), .ZN(n16926) );
  AOI22_X1 U20171 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17242), .B1(
        n17259), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16925) );
  AOI211_X1 U20172 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16932), .A(n16918), .B(
        n17249), .ZN(n16923) );
  AOI211_X1 U20173 ( .C1(n16921), .C2(n16920), .A(n16919), .B(n19061), .ZN(
        n16922) );
  AOI211_X1 U20174 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16942), .A(n16923), 
        .B(n16922), .ZN(n16924) );
  OAI211_X1 U20175 ( .C1(n16929), .C2(n16926), .A(n16925), .B(n16924), .ZN(
        P3_U2643) );
  INV_X1 U20176 ( .A(n16942), .ZN(n16935) );
  INV_X1 U20177 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19133) );
  AOI211_X1 U20178 ( .C1(n17868), .C2(n16928), .A(n16927), .B(n19061), .ZN(
        n16931) );
  OAI22_X1 U20179 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16929), .B1(n17307), 
        .B2(n17244), .ZN(n16930) );
  AOI211_X1 U20180 ( .C1(n17242), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16931), .B(n16930), .ZN(n16934) );
  OAI211_X1 U20181 ( .C1(n16936), .C2(n17307), .A(n17258), .B(n16932), .ZN(
        n16933) );
  OAI211_X1 U20182 ( .C1(n16935), .C2(n19133), .A(n16934), .B(n16933), .ZN(
        P3_U2644) );
  AOI22_X1 U20183 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17242), .B1(
        n17259), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16944) );
  AOI211_X1 U20184 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16952), .A(n16936), .B(
        n17249), .ZN(n16941) );
  AOI211_X1 U20185 ( .C1(n16939), .C2(n16938), .A(n16937), .B(n19061), .ZN(
        n16940) );
  AOI211_X1 U20186 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16942), .A(n16941), 
        .B(n16940), .ZN(n16943) );
  OAI211_X1 U20187 ( .C1(n16946), .C2(n16945), .A(n16944), .B(n16943), .ZN(
        P3_U2645) );
  AOI22_X1 U20188 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17242), .B1(
        n17259), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16957) );
  NOR2_X1 U20189 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17245), .ZN(n16958) );
  INV_X1 U20190 ( .A(n16947), .ZN(n16959) );
  OAI21_X1 U20191 ( .B1(n16959), .B2(n17245), .A(n17257), .ZN(n16973) );
  AOI211_X1 U20192 ( .C1(n16950), .C2(n16949), .A(n16948), .B(n19061), .ZN(
        n16951) );
  AOI221_X1 U20193 ( .B1(n16958), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16973), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n16951), .ZN(n16956) );
  OAI211_X1 U20194 ( .C1(n16960), .C2(n17265), .A(n17258), .B(n16952), .ZN(
        n16955) );
  INV_X1 U20195 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19129) );
  NAND3_X1 U20196 ( .A1(n17237), .A2(n16953), .A3(n19129), .ZN(n16954) );
  NAND4_X1 U20197 ( .A1(n16957), .A2(n16956), .A3(n16955), .A4(n16954), .ZN(
        P3_U2646) );
  AOI22_X1 U20198 ( .A1(n17259), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16959), 
        .B2(n16958), .ZN(n16966) );
  AOI211_X1 U20199 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16974), .A(n16960), .B(
        n17249), .ZN(n16964) );
  AOI211_X1 U20200 ( .C1(n17912), .C2(n16962), .A(n16961), .B(n19061), .ZN(
        n16963) );
  AOI211_X1 U20201 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16973), .A(n16964), 
        .B(n16963), .ZN(n16965) );
  OAI211_X1 U20202 ( .C1(n17916), .C2(n17205), .A(n16966), .B(n16965), .ZN(
        P3_U2647) );
  NAND2_X1 U20203 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16981) );
  NOR2_X1 U20204 ( .A1(n17245), .A2(n17019), .ZN(n17052) );
  INV_X1 U20205 ( .A(n17052), .ZN(n17063) );
  NOR2_X1 U20206 ( .A1(n16967), .A2(n17063), .ZN(n16995) );
  INV_X1 U20207 ( .A(n16995), .ZN(n16982) );
  INV_X1 U20208 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19125) );
  OAI21_X1 U20209 ( .B1(n16981), .B2(n16982), .A(n19125), .ZN(n16972) );
  AOI211_X1 U20210 ( .C1(n17924), .C2(n16969), .A(n16968), .B(n19061), .ZN(
        n16971) );
  OAI22_X1 U20211 ( .A1(n9999), .A2(n17205), .B1(n17244), .B2(n16975), .ZN(
        n16970) );
  AOI211_X1 U20212 ( .C1(n16973), .C2(n16972), .A(n16971), .B(n16970), .ZN(
        n16977) );
  OAI211_X1 U20213 ( .C1(n16978), .C2(n16975), .A(n17258), .B(n16974), .ZN(
        n16976) );
  NAND2_X1 U20214 ( .A1(n16977), .A2(n16976), .ZN(P3_U2648) );
  AOI211_X1 U20215 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16996), .A(n16978), .B(
        n17249), .ZN(n16979) );
  AOI21_X1 U20216 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17259), .A(n16979), .ZN(
        n16989) );
  OAI21_X1 U20217 ( .B1(n16980), .B2(n17245), .A(n17257), .ZN(n17007) );
  INV_X1 U20218 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19123) );
  INV_X1 U20219 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19121) );
  INV_X1 U20220 ( .A(n16981), .ZN(n16983) );
  AOI211_X1 U20221 ( .C1(n19123), .C2(n19121), .A(n16983), .B(n16982), .ZN(
        n16987) );
  AOI211_X1 U20222 ( .C1(n17936), .C2(n16985), .A(n16984), .B(n19061), .ZN(
        n16986) );
  AOI211_X1 U20223 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17007), .A(n16987), 
        .B(n16986), .ZN(n16988) );
  OAI211_X1 U20224 ( .C1(n16990), .C2(n17205), .A(n16989), .B(n16988), .ZN(
        P3_U2649) );
  AOI22_X1 U20225 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17242), .B1(
        n17259), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16999) );
  AOI211_X1 U20226 ( .C1(n16993), .C2(n16992), .A(n16991), .B(n19061), .ZN(
        n16994) );
  AOI221_X1 U20227 ( .B1(n16995), .B2(n19121), .C1(n17007), .C2(
        P3_REIP_REG_21__SCAN_IN), .A(n16994), .ZN(n16998) );
  OAI211_X1 U20228 ( .C1(n17004), .C2(n17343), .A(n17258), .B(n16996), .ZN(
        n16997) );
  NAND3_X1 U20229 ( .A1(n16999), .A2(n16998), .A3(n16997), .ZN(P3_U2650) );
  AOI211_X1 U20230 ( .C1(n17969), .C2(n17001), .A(n17000), .B(n19061), .ZN(
        n17006) );
  INV_X1 U20231 ( .A(n17013), .ZN(n17002) );
  OAI21_X1 U20232 ( .B1(n17002), .B2(n17357), .A(n17258), .ZN(n17003) );
  OAI22_X1 U20233 ( .A1(n17004), .A2(n17003), .B1(n17244), .B2(n17357), .ZN(
        n17005) );
  AOI211_X1 U20234 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n17007), .A(n17006), 
        .B(n17005), .ZN(n17010) );
  INV_X1 U20235 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19120) );
  NAND3_X1 U20236 ( .A1(n17008), .A2(n17052), .A3(n19120), .ZN(n17009) );
  OAI211_X1 U20237 ( .C1(n17205), .C2(n10002), .A(n17010), .B(n17009), .ZN(
        P3_U2651) );
  INV_X1 U20238 ( .A(n17011), .ZN(n17020) );
  NAND2_X1 U20239 ( .A1(n17020), .A2(n17052), .ZN(n17035) );
  OAI21_X1 U20240 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), 
        .A(n17012), .ZN(n17024) );
  OAI211_X1 U20241 ( .C1(n17029), .C2(n17015), .A(n17258), .B(n17013), .ZN(
        n17014) );
  OAI211_X1 U20242 ( .C1(n17244), .C2(n17015), .A(n18522), .B(n17014), .ZN(
        n17016) );
  AOI21_X1 U20243 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17242), .A(
        n17016), .ZN(n17023) );
  INV_X1 U20244 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17992) );
  INV_X1 U20245 ( .A(n17975), .ZN(n17038) );
  NOR2_X1 U20246 ( .A1(n17992), .A2(n17038), .ZN(n17018) );
  OAI21_X1 U20247 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17018), .A(
        n17017), .ZN(n17978) );
  INV_X1 U20248 ( .A(n17018), .ZN(n17025) );
  INV_X1 U20249 ( .A(n17058), .ZN(n17064) );
  AOI21_X1 U20250 ( .B1(n17025), .B2(n16885), .A(n17064), .ZN(n17028) );
  XOR2_X1 U20251 ( .A(n17978), .B(n17028), .Z(n17021) );
  AOI21_X1 U20252 ( .B1(n17237), .B2(n17019), .A(n17252), .ZN(n17079) );
  OAI21_X1 U20253 ( .B1(n17020), .B2(n17245), .A(n17079), .ZN(n17045) );
  AOI22_X1 U20254 ( .A1(n17210), .A2(n17021), .B1(P3_REIP_REG_19__SCAN_IN), 
        .B2(n17045), .ZN(n17022) );
  OAI211_X1 U20255 ( .C1(n17035), .C2(n17024), .A(n17023), .B(n17022), .ZN(
        P3_U2652) );
  INV_X1 U20256 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19115) );
  INV_X1 U20257 ( .A(n17045), .ZN(n17034) );
  OAI21_X1 U20258 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17975), .A(
        n17025), .ZN(n17989) );
  NAND2_X1 U20259 ( .A1(n17210), .A2(n17158), .ZN(n17232) );
  INV_X1 U20260 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17026) );
  OAI221_X1 U20261 ( .B1(n17989), .B2(n17026), .C1(n17989), .C2(n17992), .A(
        n17210), .ZN(n17027) );
  AOI22_X1 U20262 ( .A1(n17028), .A2(n17989), .B1(n17232), .B2(n17027), .ZN(
        n17032) );
  AOI211_X1 U20263 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17046), .A(n17029), .B(
        n17249), .ZN(n17031) );
  OAI22_X1 U20264 ( .A1(n17992), .A2(n17205), .B1(n17244), .B2(n17400), .ZN(
        n17030) );
  NOR4_X1 U20265 ( .A1(n18483), .A2(n17032), .A3(n17031), .A4(n17030), .ZN(
        n17033) );
  OAI221_X1 U20266 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17035), .C1(n19115), 
        .C2(n17034), .A(n17033), .ZN(P3_U2653) );
  INV_X1 U20267 ( .A(n17061), .ZN(n17036) );
  INV_X1 U20268 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20269 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17061), .B1(
        n17036), .B2(n17037), .ZN(n18018) );
  AOI21_X1 U20270 ( .B1(n17058), .B2(n18018), .A(n17158), .ZN(n17040) );
  NOR2_X1 U20271 ( .A1(n17037), .A2(n17061), .ZN(n17039) );
  OAI21_X1 U20272 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17039), .A(
        n17038), .ZN(n18000) );
  XOR2_X1 U20273 ( .A(n17040), .B(n18000), .Z(n17043) );
  NAND2_X1 U20274 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17051) );
  NOR2_X1 U20275 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17051), .ZN(n17041) );
  AOI22_X1 U20276 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17242), .B1(
        n17052), .B2(n17041), .ZN(n17042) );
  OAI211_X1 U20277 ( .C1(n19061), .C2(n17043), .A(n17042), .B(n18522), .ZN(
        n17044) );
  AOI21_X1 U20278 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n17045), .A(n17044), 
        .ZN(n17048) );
  OAI211_X1 U20279 ( .C1(n17050), .C2(n17049), .A(n17258), .B(n17046), .ZN(
        n17047) );
  OAI211_X1 U20280 ( .C1(n17049), .C2(n17244), .A(n17048), .B(n17047), .ZN(
        P3_U2654) );
  INV_X1 U20281 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19111) );
  AOI211_X1 U20282 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17065), .A(n17050), .B(
        n17249), .ZN(n17056) );
  OAI211_X1 U20283 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n17052), .B(n17051), .ZN(n17053) );
  OAI211_X1 U20284 ( .C1(n17244), .C2(n17054), .A(n18522), .B(n17053), .ZN(
        n17055) );
  AOI211_X1 U20285 ( .C1(n17242), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17056), .B(n17055), .ZN(n17060) );
  NAND2_X1 U20286 ( .A1(n17058), .A2(n18018), .ZN(n17057) );
  OAI211_X1 U20287 ( .C1(n17058), .C2(n18018), .A(n17210), .B(n17057), .ZN(
        n17059) );
  OAI211_X1 U20288 ( .C1(n17079), .C2(n19111), .A(n17060), .B(n17059), .ZN(
        P3_U2655) );
  INV_X1 U20289 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19109) );
  INV_X1 U20290 ( .A(n18013), .ZN(n17062) );
  OAI21_X1 U20291 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18013), .A(
        n17061), .ZN(n18023) );
  OAI21_X1 U20292 ( .B1(n17158), .B2(n17026), .A(n17210), .ZN(n17255) );
  AOI211_X1 U20293 ( .C1(n16885), .C2(n17062), .A(n18023), .B(n17255), .ZN(
        n17071) );
  INV_X1 U20294 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18026) );
  OAI22_X1 U20295 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n17063), .B1(n18026), 
        .B2(n17205), .ZN(n17070) );
  NAND3_X1 U20296 ( .A1(n17064), .A2(n17210), .A3(n18023), .ZN(n17067) );
  OAI211_X1 U20297 ( .C1(n17073), .C2(n17068), .A(n17258), .B(n17065), .ZN(
        n17066) );
  OAI211_X1 U20298 ( .C1(n17068), .C2(n17244), .A(n17067), .B(n17066), .ZN(
        n17069) );
  NOR4_X1 U20299 ( .A1(n18483), .A2(n17071), .A3(n17070), .A4(n17069), .ZN(
        n17072) );
  OAI21_X1 U20300 ( .B1(n17079), .B2(n19109), .A(n17072), .ZN(P3_U2656) );
  AOI211_X1 U20301 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17089), .A(n17073), .B(
        n17249), .ZN(n17081) );
  AND2_X1 U20302 ( .A1(n17237), .A2(n17074), .ZN(n17083) );
  AOI21_X1 U20303 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n17083), .A(
        P3_REIP_REG_14__SCAN_IN), .ZN(n17078) );
  AOI21_X1 U20304 ( .B1(n17075), .B2(n17086), .A(n18013), .ZN(n18038) );
  NOR2_X1 U20305 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18202), .ZN(
        n17235) );
  INV_X1 U20306 ( .A(n17235), .ZN(n17201) );
  NOR2_X1 U20307 ( .A1(n18051), .A2(n17201), .ZN(n17101) );
  AOI21_X1 U20308 ( .B1(n17076), .B2(n17101), .A(n17158), .ZN(n17088) );
  XNOR2_X1 U20309 ( .A(n18038), .B(n17088), .ZN(n17077) );
  OAI22_X1 U20310 ( .A1(n17079), .A2(n17078), .B1(n19061), .B2(n17077), .ZN(
        n17080) );
  AOI211_X1 U20311 ( .C1(n17242), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17081), .B(n17080), .ZN(n17082) );
  OAI211_X1 U20312 ( .C1(n17244), .C2(n17464), .A(n17082), .B(n18522), .ZN(
        P3_U2657) );
  INV_X1 U20313 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19105) );
  AOI22_X1 U20314 ( .A1(n17259), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n17083), 
        .B2(n19105), .ZN(n17098) );
  NAND3_X1 U20315 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_9__SCAN_IN), .ZN(n17085) );
  NAND2_X1 U20316 ( .A1(n17084), .A2(n17257), .ZN(n17124) );
  NAND2_X1 U20317 ( .A1(n17257), .A2(n17245), .ZN(n17256) );
  OAI21_X1 U20318 ( .B1(n17085), .B2(n17124), .A(n17256), .ZN(n17114) );
  OAI21_X1 U20319 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17245), .A(n17114), 
        .ZN(n17096) );
  NAND2_X1 U20320 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18050), .ZN(
        n17102) );
  INV_X1 U20321 ( .A(n17102), .ZN(n17087) );
  OAI21_X1 U20322 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17087), .A(
        n17086), .ZN(n18056) );
  AOI211_X1 U20323 ( .C1(n16885), .C2(n17102), .A(n18056), .B(n17255), .ZN(
        n17095) );
  INV_X1 U20324 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17093) );
  NAND3_X1 U20325 ( .A1(n17210), .A2(n17088), .A3(n18056), .ZN(n17092) );
  OAI211_X1 U20326 ( .C1(n17099), .C2(n17090), .A(n17258), .B(n17089), .ZN(
        n17091) );
  OAI211_X1 U20327 ( .C1(n17205), .C2(n17093), .A(n17092), .B(n17091), .ZN(
        n17094) );
  AOI211_X1 U20328 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17096), .A(n17095), 
        .B(n17094), .ZN(n17097) );
  NAND3_X1 U20329 ( .A1(n17098), .A2(n17097), .A3(n18522), .ZN(P3_U2658) );
  AOI211_X1 U20330 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17117), .A(n17099), .B(
        n17249), .ZN(n17100) );
  AOI21_X1 U20331 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17259), .A(n17100), .ZN(
        n17109) );
  NOR2_X1 U20332 ( .A1(n17101), .A2(n17158), .ZN(n17103) );
  OAI21_X1 U20333 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18050), .A(
        n17102), .ZN(n18062) );
  XNOR2_X1 U20334 ( .A(n17103), .B(n18062), .ZN(n17107) );
  INV_X1 U20335 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18066) );
  NAND2_X1 U20336 ( .A1(n17237), .A2(n19103), .ZN(n17104) );
  OAI22_X1 U20337 ( .A1(n18066), .A2(n17205), .B1(n17105), .B2(n17104), .ZN(
        n17106) );
  AOI211_X1 U20338 ( .C1(n17210), .C2(n17107), .A(n18483), .B(n17106), .ZN(
        n17108) );
  OAI211_X1 U20339 ( .C1(n19103), .C2(n17114), .A(n17109), .B(n17108), .ZN(
        P3_U2659) );
  INV_X1 U20340 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17121) );
  INV_X1 U20341 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19099) );
  INV_X1 U20342 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19097) );
  NOR2_X1 U20343 ( .A1(n19099), .A2(n19097), .ZN(n17110) );
  NOR4_X1 U20344 ( .A1(n17245), .A2(n19096), .A3(n17166), .A4(n17145), .ZN(
        n17130) );
  AOI21_X1 U20345 ( .B1(n17110), .B2(n17130), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17115) );
  NOR2_X1 U20346 ( .A1(n18202), .A2(n18112), .ZN(n17157) );
  INV_X1 U20347 ( .A(n17157), .ZN(n17172) );
  NOR2_X1 U20348 ( .A1(n18077), .A2(n17172), .ZN(n17123) );
  NAND2_X1 U20349 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17123), .ZN(
        n17122) );
  AOI21_X1 U20350 ( .B1(n17121), .B2(n17122), .A(n18050), .ZN(n18080) );
  AOI21_X1 U20351 ( .B1(n17111), .B2(n17235), .A(n17158), .ZN(n17112) );
  XNOR2_X1 U20352 ( .A(n18080), .B(n17112), .ZN(n17113) );
  OAI22_X1 U20353 ( .A1(n17115), .A2(n17114), .B1(n19061), .B2(n17113), .ZN(
        n17116) );
  AOI211_X1 U20354 ( .C1(n17259), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18483), .B(
        n17116), .ZN(n17120) );
  OAI211_X1 U20355 ( .C1(n17125), .C2(n17118), .A(n17258), .B(n17117), .ZN(
        n17119) );
  OAI211_X1 U20356 ( .C1(n17205), .C2(n17121), .A(n17120), .B(n17119), .ZN(
        P3_U2660) );
  OAI21_X1 U20357 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17123), .A(
        n17122), .ZN(n18088) );
  INV_X1 U20358 ( .A(n17123), .ZN(n17134) );
  OAI21_X1 U20359 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17134), .A(
        n16885), .ZN(n17136) );
  XNOR2_X1 U20360 ( .A(n18088), .B(n17136), .ZN(n17133) );
  NAND2_X1 U20361 ( .A1(n17256), .A2(n17124), .ZN(n17151) );
  NAND2_X1 U20362 ( .A1(n17130), .A2(n19097), .ZN(n17142) );
  AOI21_X1 U20363 ( .B1(n17151), .B2(n17142), .A(n19099), .ZN(n17129) );
  AOI211_X1 U20364 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17137), .A(n17125), .B(
        n17249), .ZN(n17128) );
  INV_X1 U20365 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17513) );
  OAI22_X1 U20366 ( .A1(n17126), .A2(n17205), .B1(n17244), .B2(n17513), .ZN(
        n17127) );
  NOR4_X1 U20367 ( .A1(n18483), .A2(n17129), .A3(n17128), .A4(n17127), .ZN(
        n17132) );
  NAND3_X1 U20368 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17130), .A3(n19099), 
        .ZN(n17131) );
  OAI211_X1 U20369 ( .C1(n19061), .C2(n17133), .A(n17132), .B(n17131), .ZN(
        P3_U2661) );
  AND2_X1 U20370 ( .A1(n18110), .A2(n17157), .ZN(n17147) );
  OAI21_X1 U20371 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17147), .A(
        n17134), .ZN(n18100) );
  OR2_X1 U20372 ( .A1(n18112), .A2(n18125), .ZN(n18111) );
  NOR2_X1 U20373 ( .A1(n18111), .A2(n17201), .ZN(n17148) );
  OAI221_X1 U20374 ( .B1(n18100), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(
        n18100), .C2(n17148), .A(n17210), .ZN(n17135) );
  AOI22_X1 U20375 ( .A1(n18100), .A2(n17136), .B1(n17232), .B2(n17135), .ZN(
        n17141) );
  OAI211_X1 U20376 ( .C1(n17144), .C2(n17139), .A(n17258), .B(n17137), .ZN(
        n17138) );
  OAI211_X1 U20377 ( .C1(n17244), .C2(n17139), .A(n18522), .B(n17138), .ZN(
        n17140) );
  AOI211_X1 U20378 ( .C1(n17242), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17141), .B(n17140), .ZN(n17143) );
  OAI211_X1 U20379 ( .C1(n17151), .C2(n19097), .A(n17143), .B(n17142), .ZN(
        P3_U2662) );
  INV_X1 U20380 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17561) );
  AOI211_X1 U20381 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17164), .A(n17144), .B(
        n17249), .ZN(n17154) );
  NOR3_X1 U20382 ( .A1(n17245), .A2(n17166), .A3(n17145), .ZN(n17146) );
  NOR2_X1 U20383 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17146), .ZN(n17152) );
  NAND2_X1 U20384 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17157), .ZN(
        n17156) );
  AOI21_X1 U20385 ( .B1(n18113), .B2(n17156), .A(n17147), .ZN(n18116) );
  NOR2_X1 U20386 ( .A1(n17148), .A2(n17158), .ZN(n17149) );
  XNOR2_X1 U20387 ( .A(n18116), .B(n17149), .ZN(n17150) );
  OAI22_X1 U20388 ( .A1(n17152), .A2(n17151), .B1(n19061), .B2(n17150), .ZN(
        n17153) );
  AOI211_X1 U20389 ( .C1(n17242), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17154), .B(n17153), .ZN(n17155) );
  OAI211_X1 U20390 ( .C1(n17244), .C2(n17561), .A(n17155), .B(n18522), .ZN(
        P3_U2663) );
  NOR3_X1 U20391 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17166), .A3(n17245), .ZN(
        n17174) );
  NAND2_X1 U20392 ( .A1(n17237), .A2(n17166), .ZN(n17188) );
  NAND2_X1 U20393 ( .A1(n17257), .A2(n17188), .ZN(n17192) );
  OAI21_X1 U20394 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17157), .A(
        n17156), .ZN(n18135) );
  INV_X1 U20395 ( .A(n18135), .ZN(n17162) );
  NAND2_X1 U20396 ( .A1(n16885), .A2(n17210), .ZN(n17216) );
  INV_X1 U20397 ( .A(n17216), .ZN(n17243) );
  OAI21_X1 U20398 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17172), .A(
        n17243), .ZN(n17182) );
  NOR2_X1 U20399 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17172), .ZN(
        n17159) );
  OAI21_X1 U20400 ( .B1(n17159), .B2(n17158), .A(n17210), .ZN(n17161) );
  AOI22_X1 U20401 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17242), .B1(
        n17259), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n17160) );
  OAI221_X1 U20402 ( .B1(n17162), .B2(n17182), .C1(n18135), .C2(n17161), .A(
        n17160), .ZN(n17163) );
  AOI221_X1 U20403 ( .B1(n17174), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n17192), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n17163), .ZN(n17170) );
  OAI211_X1 U20404 ( .C1(n17175), .C2(n17165), .A(n17258), .B(n17164), .ZN(
        n17169) );
  NOR2_X1 U20405 ( .A1(n17245), .A2(n17166), .ZN(n17167) );
  INV_X1 U20406 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19093) );
  NAND3_X1 U20407 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17167), .A3(n19093), 
        .ZN(n17168) );
  NAND4_X1 U20408 ( .A1(n17170), .A2(n18522), .A3(n17169), .A4(n17168), .ZN(
        P3_U2664) );
  NAND2_X1 U20409 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17171), .ZN(
        n17184) );
  INV_X1 U20410 ( .A(n17184), .ZN(n17173) );
  OAI21_X1 U20411 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17173), .A(
        n17172), .ZN(n18144) );
  INV_X1 U20412 ( .A(n18144), .ZN(n17183) );
  AOI211_X1 U20413 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n17242), .A(
        n18483), .B(n17174), .ZN(n17181) );
  AOI211_X1 U20414 ( .C1(n16885), .C2(n17184), .A(n18144), .B(n17255), .ZN(
        n17179) );
  AOI211_X1 U20415 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17186), .A(n17175), .B(
        n17249), .ZN(n17178) );
  AOI22_X1 U20416 ( .A1(n17192), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17259), 
        .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n17176) );
  INV_X1 U20417 ( .A(n17176), .ZN(n17177) );
  NOR3_X1 U20418 ( .A1(n17179), .A2(n17178), .A3(n17177), .ZN(n17180) );
  OAI211_X1 U20419 ( .C1(n17183), .C2(n17182), .A(n17181), .B(n17180), .ZN(
        P3_U2665) );
  NOR2_X1 U20420 ( .A1(n18202), .A2(n18153), .ZN(n17200) );
  OAI21_X1 U20421 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17200), .A(
        n17184), .ZN(n18158) );
  OAI21_X1 U20422 ( .B1(n18153), .B2(n17201), .A(n16885), .ZN(n17202) );
  XNOR2_X1 U20423 ( .A(n18158), .B(n17202), .ZN(n17194) );
  OAI22_X1 U20424 ( .A1(n18152), .A2(n17205), .B1(n17244), .B2(n17565), .ZN(
        n17191) );
  INV_X1 U20425 ( .A(n17185), .ZN(n17189) );
  OAI211_X1 U20426 ( .C1(n17203), .C2(n17565), .A(n17258), .B(n17186), .ZN(
        n17187) );
  OAI211_X1 U20427 ( .C1(n17189), .C2(n17188), .A(n18522), .B(n17187), .ZN(
        n17190) );
  AOI211_X1 U20428 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n17192), .A(n17191), .B(
        n17190), .ZN(n17193) );
  OAI21_X1 U20429 ( .B1(n19061), .B2(n17194), .A(n17193), .ZN(P3_U2666) );
  AOI21_X1 U20430 ( .B1(n17237), .B2(n17213), .A(n17252), .ZN(n17226) );
  NOR3_X1 U20431 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17245), .A3(n17213), .ZN(
        n17198) );
  NAND2_X1 U20432 ( .A1(n17195), .A2(n19226), .ZN(n17248) );
  OAI221_X1 U20433 ( .B1(n17248), .B2(n11180), .C1(n17248), .C2(n17196), .A(
        n18522), .ZN(n17197) );
  AOI211_X1 U20434 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17259), .A(n17198), .B(
        n17197), .ZN(n17212) );
  INV_X1 U20435 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17206) );
  NAND2_X1 U20436 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17199), .ZN(
        n17217) );
  AOI21_X1 U20437 ( .B1(n17206), .B2(n17217), .A(n17200), .ZN(n17204) );
  NAND2_X1 U20438 ( .A1(n17199), .A2(n17206), .ZN(n18161) );
  OAI22_X1 U20439 ( .A1(n17204), .A2(n17202), .B1(n17201), .B2(n18161), .ZN(
        n17209) );
  AOI211_X1 U20440 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17219), .A(n17203), .B(
        n17249), .ZN(n17208) );
  INV_X1 U20441 ( .A(n17204), .ZN(n18170) );
  OAI22_X1 U20442 ( .A1(n17206), .A2(n17205), .B1(n18170), .B2(n17232), .ZN(
        n17207) );
  AOI211_X1 U20443 ( .C1(n17210), .C2(n17209), .A(n17208), .B(n17207), .ZN(
        n17211) );
  OAI211_X1 U20444 ( .C1(n17226), .C2(n19087), .A(n17212), .B(n17211), .ZN(
        P3_U2667) );
  INV_X1 U20445 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19085) );
  NAND2_X1 U20446 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17236) );
  NAND2_X1 U20447 ( .A1(n17237), .A2(n17213), .ZN(n17214) );
  OAI21_X1 U20448 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18995), .A(
        n11180), .ZN(n19161) );
  OAI22_X1 U20449 ( .A1(n17236), .A2(n17214), .B1(n17248), .B2(n19161), .ZN(
        n17215) );
  AOI21_X1 U20450 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17242), .A(
        n17215), .ZN(n17225) );
  NOR2_X1 U20451 ( .A1(n18202), .A2(n18193), .ZN(n17228) );
  AOI21_X1 U20452 ( .B1(n17228), .B2(n17026), .A(n17216), .ZN(n17234) );
  OAI21_X1 U20453 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17228), .A(
        n17217), .ZN(n18183) );
  NAND2_X1 U20454 ( .A1(n17228), .A2(n17026), .ZN(n17218) );
  AOI211_X1 U20455 ( .C1(n16885), .C2(n17218), .A(n19061), .B(n18183), .ZN(
        n17223) );
  OAI211_X1 U20456 ( .C1(n17241), .C2(n17221), .A(n17258), .B(n17219), .ZN(
        n17220) );
  OAI21_X1 U20457 ( .B1(n17221), .B2(n17244), .A(n17220), .ZN(n17222) );
  AOI211_X1 U20458 ( .C1(n17234), .C2(n18183), .A(n17223), .B(n17222), .ZN(
        n17224) );
  OAI211_X1 U20459 ( .C1(n17226), .C2(n19085), .A(n17225), .B(n17224), .ZN(
        P3_U2668) );
  NOR2_X1 U20460 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17246) );
  INV_X1 U20461 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17227) );
  OAI21_X1 U20462 ( .B1(n17246), .B2(n17227), .A(n17258), .ZN(n17240) );
  INV_X1 U20463 ( .A(n17228), .ZN(n17229) );
  OAI21_X1 U20464 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17229), .ZN(n18189) );
  AOI22_X1 U20465 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17242), .B1(
        n17259), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n17231) );
  NAND2_X1 U20466 ( .A1(n19177), .A2(n19020), .ZN(n19000) );
  INV_X1 U20467 ( .A(n19000), .ZN(n19003) );
  NOR2_X1 U20468 ( .A1(n18995), .A2(n19003), .ZN(n19174) );
  INV_X1 U20469 ( .A(n17248), .ZN(n19228) );
  AOI22_X1 U20470 ( .A1(n17252), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n19174), 
        .B2(n19228), .ZN(n17230) );
  OAI211_X1 U20471 ( .C1(n18189), .C2(n17232), .A(n17231), .B(n17230), .ZN(
        n17233) );
  AOI221_X1 U20472 ( .B1(n17235), .B2(n17234), .C1(n18189), .C2(n17234), .A(
        n17233), .ZN(n17239) );
  OAI211_X1 U20473 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17237), .B(n17236), .ZN(n17238) );
  OAI211_X1 U20474 ( .C1(n17241), .C2(n17240), .A(n17239), .B(n17238), .ZN(
        P3_U2669) );
  AOI21_X1 U20475 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17243), .A(
        n17242), .ZN(n17254) );
  INV_X1 U20476 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17579) );
  OAI22_X1 U20477 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17245), .B1(n17244), 
        .B2(n17579), .ZN(n17251) );
  OR2_X1 U20478 ( .A1(n17246), .A2(n17575), .ZN(n17580) );
  NAND2_X1 U20479 ( .A1(n17247), .A2(n19020), .ZN(n19178) );
  OAI22_X1 U20480 ( .A1(n17249), .A2(n17580), .B1(n19178), .B2(n17248), .ZN(
        n17250) );
  AOI211_X1 U20481 ( .C1(n17252), .C2(P3_REIP_REG_1__SCAN_IN), .A(n17251), .B(
        n17250), .ZN(n17253) );
  OAI221_X1 U20482 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17255), .C1(
        n18202), .C2(n17254), .A(n17253), .ZN(P3_U2670) );
  NAND3_X1 U20483 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19162), .A3(
        n17257), .ZN(n17261) );
  OAI21_X1 U20484 ( .B1(n17259), .B2(n17258), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17260) );
  NAND3_X1 U20485 ( .A1(n17262), .A2(n17261), .A3(n17260), .ZN(P3_U2671) );
  INV_X1 U20486 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17264) );
  NAND4_X1 U20487 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n17372), .ZN(n17263) );
  NOR3_X1 U20488 ( .A1(n17265), .A2(n17264), .A3(n17263), .ZN(n17266) );
  NAND4_X1 U20489 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17302), .A4(n17266), .ZN(n17269) );
  NOR2_X1 U20490 ( .A1(n17270), .A2(n17269), .ZN(n17297) );
  NAND2_X1 U20491 ( .A1(n17578), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17268) );
  NAND2_X1 U20492 ( .A1(n17297), .A2(n17711), .ZN(n17267) );
  OAI22_X1 U20493 ( .A1(n17297), .A2(n17268), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17267), .ZN(P3_U2672) );
  NAND2_X1 U20494 ( .A1(n17270), .A2(n17269), .ZN(n17271) );
  NAND2_X1 U20495 ( .A1(n17271), .A2(n17578), .ZN(n17296) );
  AOI22_X1 U20496 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17272) );
  OAI21_X1 U20497 ( .B1(n11021), .B2(n17273), .A(n17272), .ZN(n17284) );
  AOI22_X1 U20498 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17281) );
  OAI22_X1 U20499 ( .A1(n17557), .A2(n17442), .B1(n17274), .B2(n18806), .ZN(
        n17279) );
  AOI22_X1 U20500 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U20501 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20502 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17275) );
  NAND3_X1 U20503 ( .A1(n17277), .A2(n17276), .A3(n17275), .ZN(n17278) );
  AOI211_X1 U20504 ( .C1(n17546), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n17279), .B(n17278), .ZN(n17280) );
  OAI211_X1 U20505 ( .C1(n10316), .C2(n17282), .A(n17281), .B(n17280), .ZN(
        n17283) );
  AOI211_X1 U20506 ( .C1(n17497), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n17284), .B(n17283), .ZN(n17295) );
  AOI22_X1 U20507 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17294) );
  INV_X1 U20508 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20509 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20510 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17285) );
  OAI211_X1 U20511 ( .C1(n10314), .C2(n17338), .A(n17286), .B(n17285), .ZN(
        n17292) );
  AOI22_X1 U20512 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17290) );
  AOI22_X1 U20513 ( .A1(n9670), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9662), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U20514 ( .A1(n9648), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17288) );
  NAND2_X1 U20515 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n17287) );
  NAND4_X1 U20516 ( .A1(n17290), .A2(n17289), .A3(n17288), .A4(n17287), .ZN(
        n17291) );
  AOI211_X1 U20517 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17292), .B(n17291), .ZN(n17293) );
  OAI211_X1 U20518 ( .C1(n17526), .C2(n17329), .A(n17294), .B(n17293), .ZN(
        n17299) );
  NAND2_X1 U20519 ( .A1(n17300), .A2(n17299), .ZN(n17298) );
  XNOR2_X1 U20520 ( .A(n17295), .B(n17298), .ZN(n17593) );
  OAI22_X1 U20521 ( .A1(n17297), .A2(n17296), .B1(n17593), .B2(n17578), .ZN(
        P3_U2673) );
  OAI21_X1 U20522 ( .B1(n17300), .B2(n17299), .A(n17298), .ZN(n17600) );
  NOR2_X1 U20523 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17308), .ZN(n17301) );
  AOI22_X1 U20524 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17303), .B1(n17302), 
        .B2(n17301), .ZN(n17304) );
  OAI21_X1 U20525 ( .B1(n17578), .B2(n17600), .A(n17304), .ZN(P3_U2674) );
  OAI211_X1 U20526 ( .C1(n17609), .C2(n17608), .A(n17583), .B(n17607), .ZN(
        n17305) );
  OAI221_X1 U20527 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17308), .C1(n17307), 
        .C2(n17306), .A(n17305), .ZN(P3_U2676) );
  AOI21_X1 U20528 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17578), .A(n17317), .ZN(
        n17310) );
  XNOR2_X1 U20529 ( .A(n17309), .B(n17313), .ZN(n17618) );
  OAI22_X1 U20530 ( .A1(n17311), .A2(n17310), .B1(n17578), .B2(n17618), .ZN(
        P3_U2677) );
  INV_X1 U20531 ( .A(n17312), .ZN(n17320) );
  AOI21_X1 U20532 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17578), .A(n17320), .ZN(
        n17316) );
  OAI21_X1 U20533 ( .B1(n17315), .B2(n17314), .A(n17313), .ZN(n17622) );
  OAI22_X1 U20534 ( .A1(n17317), .A2(n17316), .B1(n17578), .B2(n17622), .ZN(
        P3_U2678) );
  AOI21_X1 U20535 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17578), .A(n17326), .ZN(
        n17319) );
  XNOR2_X1 U20536 ( .A(n17318), .B(n17322), .ZN(n17629) );
  OAI22_X1 U20537 ( .A1(n17320), .A2(n17319), .B1(n17578), .B2(n17629), .ZN(
        P3_U2679) );
  INV_X1 U20538 ( .A(n17321), .ZN(n17342) );
  AOI21_X1 U20539 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17578), .A(n17342), .ZN(
        n17325) );
  OAI21_X1 U20540 ( .B1(n17324), .B2(n17323), .A(n17322), .ZN(n17635) );
  OAI22_X1 U20541 ( .A1(n17326), .A2(n17325), .B1(n17578), .B2(n17635), .ZN(
        P3_U2680) );
  AOI21_X1 U20542 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17578), .A(n17327), .ZN(
        n17341) );
  AOI22_X1 U20543 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17328) );
  OAI21_X1 U20544 ( .B1(n9710), .B2(n17329), .A(n17328), .ZN(n17340) );
  AOI22_X1 U20545 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17337) );
  OAI22_X1 U20546 ( .A1(n9652), .A2(n18582), .B1(n17388), .B2(n17330), .ZN(
        n17335) );
  AOI22_X1 U20547 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17333) );
  AOI22_X1 U20548 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17332) );
  AOI22_X1 U20549 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17331) );
  NAND3_X1 U20550 ( .A1(n17333), .A2(n17332), .A3(n17331), .ZN(n17334) );
  AOI211_X1 U20551 ( .C1(n9670), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17335), .B(n17334), .ZN(n17336) );
  OAI211_X1 U20552 ( .C1(n11180), .C2(n17338), .A(n17337), .B(n17336), .ZN(
        n17339) );
  AOI211_X1 U20553 ( .C1(n9655), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n17340), .B(n17339), .ZN(n17636) );
  OAI22_X1 U20554 ( .A1(n17342), .A2(n17341), .B1(n17636), .B2(n17578), .ZN(
        P3_U2681) );
  AOI22_X1 U20555 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17372), .B1(n17344), 
        .B2(n17343), .ZN(n17356) );
  AOI22_X1 U20556 ( .A1(n9670), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U20557 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U20558 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17345) );
  OAI211_X1 U20559 ( .C1(n10314), .C2(n17347), .A(n17346), .B(n17345), .ZN(
        n17353) );
  AOI22_X1 U20560 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17351) );
  AOI22_X1 U20561 ( .A1(n14248), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17350) );
  AOI22_X1 U20562 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17349) );
  NAND2_X1 U20563 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n17348) );
  NAND4_X1 U20564 ( .A1(n17351), .A2(n17350), .A3(n17349), .A4(n17348), .ZN(
        n17352) );
  AOI211_X1 U20565 ( .C1(n17547), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17353), .B(n17352), .ZN(n17354) );
  OAI211_X1 U20566 ( .C1(n9652), .C2(n18576), .A(n17355), .B(n17354), .ZN(
        n17640) );
  MUX2_X1 U20567 ( .A(n17356), .B(n17640), .S(n17583), .Z(P3_U2682) );
  AOI21_X1 U20568 ( .B1(n17357), .B2(n17384), .A(n17583), .ZN(n17358) );
  INV_X1 U20569 ( .A(n17358), .ZN(n17371) );
  AOI22_X1 U20570 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U20571 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17360) );
  AOI22_X1 U20572 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17544), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17359) );
  OAI211_X1 U20573 ( .C1(n10314), .C2(n17361), .A(n17360), .B(n17359), .ZN(
        n17367) );
  AOI22_X1 U20574 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20575 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17364) );
  AOI22_X1 U20576 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17363) );
  NAND2_X1 U20577 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n17362) );
  NAND4_X1 U20578 ( .A1(n17365), .A2(n17364), .A3(n17363), .A4(n17362), .ZN(
        n17366) );
  AOI211_X1 U20579 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17367), .B(n17366), .ZN(n17368) );
  OAI211_X1 U20580 ( .C1(n9652), .C2(n18571), .A(n17369), .B(n17368), .ZN(
        n17645) );
  INV_X1 U20581 ( .A(n17645), .ZN(n17370) );
  OAI22_X1 U20582 ( .A1(n17372), .A2(n17371), .B1(n17370), .B2(n17578), .ZN(
        P3_U2683) );
  INV_X1 U20583 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U20584 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17373) );
  OAI21_X1 U20585 ( .B1(n17522), .B2(n17374), .A(n17373), .ZN(n17383) );
  AOI22_X1 U20586 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U20587 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17375) );
  OAI21_X1 U20588 ( .B1(n9652), .B2(n18564), .A(n17375), .ZN(n17379) );
  AOI22_X1 U20589 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17377) );
  AOI22_X1 U20590 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17376) );
  OAI211_X1 U20591 ( .C1(n10314), .C2(n17484), .A(n17377), .B(n17376), .ZN(
        n17378) );
  AOI211_X1 U20592 ( .C1(n17547), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17379), .B(n17378), .ZN(n17380) );
  OAI211_X1 U20593 ( .C1(n17274), .C2(n18760), .A(n17381), .B(n17380), .ZN(
        n17382) );
  AOI211_X1 U20594 ( .C1(n17520), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17383), .B(n17382), .ZN(n17654) );
  OAI21_X1 U20595 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17385), .A(n17384), .ZN(
        n17386) );
  AOI22_X1 U20596 ( .A1(n17583), .A2(n17654), .B1(n17386), .B2(n17578), .ZN(
        P3_U2684) );
  AOI22_X1 U20597 ( .A1(n9649), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17387) );
  OAI21_X1 U20598 ( .B1(n17388), .B2(n17507), .A(n17387), .ZN(n17398) );
  AOI22_X1 U20599 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17396) );
  OAI22_X1 U20600 ( .A1(n9710), .A2(n17499), .B1(n9652), .B2(n18560), .ZN(
        n17393) );
  AOI22_X1 U20601 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20602 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20603 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17389) );
  NAND3_X1 U20604 ( .A1(n17391), .A2(n17390), .A3(n17389), .ZN(n17392) );
  AOI211_X1 U20605 ( .C1(n9641), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17393), .B(n17392), .ZN(n17395) );
  OAI211_X1 U20606 ( .C1(n17274), .C2(n11051), .A(n17396), .B(n17395), .ZN(
        n17397) );
  AOI211_X1 U20607 ( .C1(n17520), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n17398), .B(n17397), .ZN(n17659) );
  INV_X1 U20608 ( .A(n17414), .ZN(n17399) );
  OAI33_X1 U20609 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18585), .A3(n17414), 
        .B1(n17400), .B2(n17583), .B3(n17399), .ZN(n17401) );
  INV_X1 U20610 ( .A(n17401), .ZN(n17402) );
  OAI21_X1 U20611 ( .B1(n17659), .B2(n17578), .A(n17402), .ZN(P3_U2685) );
  AOI22_X1 U20612 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17501), .B1(
        n14248), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20613 ( .B1(n17500), .B2(n17532), .A(n17403), .ZN(n17413) );
  AOI22_X1 U20614 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17538), .B1(
        n17544), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17410) );
  OAI22_X1 U20615 ( .A1(n17557), .A2(n17527), .B1(n17519), .B2(n17420), .ZN(
        n17408) );
  AOI22_X1 U20616 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17546), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17541), .ZN(n17406) );
  AOI22_X1 U20617 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U20618 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17433), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9641), .ZN(n17404) );
  NAND3_X1 U20619 ( .A1(n17406), .A2(n17405), .A3(n17404), .ZN(n17407) );
  AOI211_X1 U20620 ( .C1(n9651), .C2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n17408), .B(n17407), .ZN(n17409) );
  OAI211_X1 U20621 ( .C1(n17411), .C2(n17526), .A(n17410), .B(n17409), .ZN(
        n17412) );
  AOI211_X1 U20622 ( .C1(n9655), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n17413), .B(n17412), .ZN(n17663) );
  OAI211_X1 U20623 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n17415), .A(n17414), .B(
        n17578), .ZN(n17416) );
  OAI21_X1 U20624 ( .B1(n17663), .B2(n17578), .A(n17416), .ZN(P3_U2686) );
  OR2_X1 U20625 ( .A1(n18585), .A2(n17417), .ZN(n17443) );
  AOI22_X1 U20626 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U20627 ( .B1(n10316), .B2(n18782), .A(n17418), .ZN(n17429) );
  AOI22_X1 U20628 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17427) );
  INV_X1 U20629 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18550) );
  OAI22_X1 U20630 ( .A1(n17420), .A2(n17419), .B1(n9652), .B2(n18550), .ZN(
        n17425) );
  AOI22_X1 U20631 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17423) );
  AOI22_X1 U20632 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20633 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17421) );
  NAND3_X1 U20634 ( .A1(n17423), .A2(n17422), .A3(n17421), .ZN(n17424) );
  AOI211_X1 U20635 ( .C1(n9649), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17425), .B(n17424), .ZN(n17426) );
  OAI211_X1 U20636 ( .C1(n17274), .C2(n18752), .A(n17427), .B(n17426), .ZN(
        n17428) );
  AOI211_X1 U20637 ( .C1(n9647), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17429), .B(n17428), .ZN(n17670) );
  NAND3_X1 U20638 ( .A1(n17443), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17578), 
        .ZN(n17430) );
  OAI221_X1 U20639 ( .B1(n17443), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17578), 
        .C2(n17670), .A(n17430), .ZN(P3_U2687) );
  AOI22_X1 U20640 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U20641 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20642 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17431) );
  OAI211_X1 U20643 ( .C1(n10314), .C2(n18590), .A(n17432), .B(n17431), .ZN(
        n17439) );
  AOI22_X1 U20644 ( .A1(n14248), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U20645 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20646 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17435) );
  NAND2_X1 U20647 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n17434) );
  NAND4_X1 U20648 ( .A1(n17437), .A2(n17436), .A3(n17435), .A4(n17434), .ZN(
        n17438) );
  AOI211_X1 U20649 ( .C1(n17547), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17439), .B(n17438), .ZN(n17440) );
  OAI211_X1 U20650 ( .C1(n9710), .C2(n17442), .A(n17441), .B(n17440), .ZN(
        n17671) );
  INV_X1 U20651 ( .A(n17671), .ZN(n17446) );
  OAI211_X1 U20652 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17444), .A(n17443), .B(
        n17578), .ZN(n17445) );
  OAI21_X1 U20653 ( .B1(n17446), .B2(n17578), .A(n17445), .ZN(P3_U2688) );
  NAND2_X1 U20654 ( .A1(n17578), .A2(n17460), .ZN(n17463) );
  AOI22_X1 U20655 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U20656 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U20657 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17447) );
  OAI211_X1 U20658 ( .C1(n17526), .C2(n17449), .A(n17448), .B(n17447), .ZN(
        n17456) );
  AOI22_X1 U20659 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17544), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20660 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U20661 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17452) );
  NAND2_X1 U20662 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n17451) );
  NAND4_X1 U20663 ( .A1(n17454), .A2(n17453), .A3(n17452), .A4(n17451), .ZN(
        n17455) );
  AOI211_X1 U20664 ( .C1(n9641), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n17456), .B(n17455), .ZN(n17457) );
  OAI211_X1 U20665 ( .C1(n9652), .C2(n17459), .A(n17458), .B(n17457), .ZN(
        n17676) );
  NOR3_X1 U20666 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18585), .A3(n17460), .ZN(
        n17461) );
  AOI21_X1 U20667 ( .B1(n17583), .B2(n17676), .A(n17461), .ZN(n17462) );
  OAI21_X1 U20668 ( .B1(n17464), .B2(n17463), .A(n17462), .ZN(P3_U2689) );
  OAI21_X1 U20669 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17465), .A(n17578), .ZN(
        n17481) );
  AOI22_X1 U20670 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20671 ( .B1(n17420), .B2(n17467), .A(n17466), .ZN(n17480) );
  AOI22_X1 U20672 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17477) );
  OAI22_X1 U20673 ( .A1(n17500), .A2(n17470), .B1(n11036), .B2(n17469), .ZN(
        n17475) );
  AOI22_X1 U20674 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U20675 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17544), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U20676 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17471) );
  NAND3_X1 U20677 ( .A1(n17473), .A2(n17472), .A3(n17471), .ZN(n17474) );
  AOI211_X1 U20678 ( .C1(n17538), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n17475), .B(n17474), .ZN(n17476) );
  OAI211_X1 U20679 ( .C1(n9710), .C2(n17478), .A(n17477), .B(n17476), .ZN(
        n17479) );
  AOI211_X1 U20680 ( .C1(n9647), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17480), .B(n17479), .ZN(n17686) );
  OAI22_X1 U20681 ( .A1(n17482), .A2(n17481), .B1(n17686), .B2(n17578), .ZN(
        P3_U2691) );
  AOI22_X1 U20682 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17483) );
  OAI21_X1 U20683 ( .B1(n11180), .B2(n17484), .A(n17483), .ZN(n17494) );
  AOI22_X1 U20684 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U20685 ( .A1(n9647), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17547), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17485) );
  OAI21_X1 U20686 ( .B1(n9652), .B2(n17486), .A(n17485), .ZN(n17490) );
  AOI22_X1 U20687 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U20688 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17487) );
  OAI211_X1 U20689 ( .C1(n10314), .C2(n18564), .A(n17488), .B(n17487), .ZN(
        n17489) );
  AOI211_X1 U20690 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17490), .B(n17489), .ZN(n17491) );
  OAI211_X1 U20691 ( .C1(n10316), .C2(n18760), .A(n17492), .B(n17491), .ZN(
        n17493) );
  AOI211_X1 U20692 ( .C1(n17497), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17494), .B(n17493), .ZN(n17690) );
  INV_X1 U20693 ( .A(n17564), .ZN(n17572) );
  AND3_X1 U20694 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17572), .ZN(n17567) );
  NAND2_X1 U20695 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17567), .ZN(n17558) );
  NOR2_X1 U20696 ( .A1(n17561), .A2(n17558), .ZN(n17536) );
  NAND2_X1 U20697 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17536), .ZN(n17535) );
  NOR2_X1 U20698 ( .A1(n17513), .A2(n17535), .ZN(n17516) );
  OAI21_X1 U20699 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17516), .A(n17495), .ZN(
        n17496) );
  AOI22_X1 U20700 ( .A1(n17583), .A2(n17690), .B1(n17496), .B2(n17578), .ZN(
        P3_U2692) );
  AOI22_X1 U20701 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U20702 ( .A1(n17540), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17511) );
  OAI22_X1 U20703 ( .A1(n17500), .A2(n17499), .B1(n9652), .B2(n17498), .ZN(
        n17509) );
  AOI22_X1 U20704 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17506) );
  AOI22_X1 U20705 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9649), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17503) );
  AOI22_X1 U20706 ( .A1(n9670), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17501), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17502) );
  OAI211_X1 U20707 ( .C1(n10314), .C2(n18560), .A(n17503), .B(n17502), .ZN(
        n17504) );
  AOI21_X1 U20708 ( .B1(n17547), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17504), .ZN(n17505) );
  OAI211_X1 U20709 ( .C1(n17557), .C2(n17507), .A(n17506), .B(n17505), .ZN(
        n17508) );
  AOI211_X1 U20710 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17509), .B(n17508), .ZN(n17510) );
  NAND3_X1 U20711 ( .A1(n17512), .A2(n17511), .A3(n17510), .ZN(n17696) );
  INV_X1 U20712 ( .A(n17696), .ZN(n17517) );
  AOI21_X1 U20713 ( .B1(n17513), .B2(n17535), .A(n17583), .ZN(n17514) );
  INV_X1 U20714 ( .A(n17514), .ZN(n17515) );
  OAI22_X1 U20715 ( .A1(n17517), .A2(n17578), .B1(n17516), .B2(n17515), .ZN(
        P3_U2693) );
  AOI22_X1 U20716 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14248), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17546), .ZN(n17518) );
  OAI21_X1 U20717 ( .B1(n17519), .B2(n11021), .A(n17518), .ZN(n17534) );
  AOI22_X1 U20718 ( .A1(n17538), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U20719 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U20720 ( .B1(n17523), .B2(n17522), .A(n17521), .ZN(n17529) );
  AOI22_X1 U20721 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17497), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17450), .ZN(n17525) );
  AOI22_X1 U20722 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17501), .ZN(n17524) );
  OAI211_X1 U20723 ( .C1(n17527), .C2(n17526), .A(n17525), .B(n17524), .ZN(
        n17528) );
  AOI211_X1 U20724 ( .C1(n9641), .C2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n17529), .B(n17528), .ZN(n17530) );
  OAI211_X1 U20725 ( .C1(n9709), .C2(n17532), .A(n17531), .B(n17530), .ZN(
        n17533) );
  AOI211_X1 U20726 ( .C1(n9647), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n17534), .B(n17533), .ZN(n17701) );
  OAI21_X1 U20727 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17536), .A(n17535), .ZN(
        n17537) );
  AOI22_X1 U20728 ( .A1(n17583), .A2(n17701), .B1(n17537), .B2(n17578), .ZN(
        P3_U2694) );
  NAND2_X1 U20729 ( .A1(n17578), .A2(n17558), .ZN(n17562) );
  AOI22_X1 U20730 ( .A1(n17497), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17538), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17555) );
  AOI22_X1 U20731 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9648), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U20732 ( .A1(n17501), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17541), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17542) );
  OAI211_X1 U20733 ( .C1(n10314), .C2(n18550), .A(n17543), .B(n17542), .ZN(
        n17553) );
  AOI22_X1 U20734 ( .A1(n17544), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17551) );
  AOI22_X1 U20735 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9662), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17550) );
  AOI22_X1 U20736 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17546), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17549) );
  NAND2_X1 U20737 ( .A1(n17547), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n17548) );
  NAND4_X1 U20738 ( .A1(n17551), .A2(n17550), .A3(n17549), .A4(n17548), .ZN(
        n17552) );
  AOI211_X1 U20739 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17553), .B(n17552), .ZN(n17554) );
  OAI211_X1 U20740 ( .C1(n17557), .C2(n17556), .A(n17555), .B(n17554), .ZN(
        n17706) );
  NOR3_X1 U20741 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18585), .A3(n17558), .ZN(
        n17559) );
  AOI21_X1 U20742 ( .B1(n17583), .B2(n17706), .A(n17559), .ZN(n17560) );
  OAI21_X1 U20743 ( .B1(n17561), .B2(n17562), .A(n17560), .ZN(P3_U2695) );
  NOR2_X1 U20744 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17567), .ZN(n17563) );
  OAI22_X1 U20745 ( .A1(n17563), .A2(n17562), .B1(n18590), .B2(n17578), .ZN(
        P3_U2696) );
  NOR2_X1 U20746 ( .A1(n17565), .A2(n17564), .ZN(n17569) );
  OAI21_X1 U20747 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17569), .A(n17578), .ZN(
        n17566) );
  OAI22_X1 U20748 ( .A1(n17567), .A2(n17566), .B1(n18582), .B2(n17578), .ZN(
        P3_U2697) );
  OAI21_X1 U20749 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17572), .A(n17578), .ZN(
        n17568) );
  OAI22_X1 U20750 ( .A1(n17569), .A2(n17568), .B1(n18576), .B2(n17578), .ZN(
        P3_U2698) );
  NOR2_X1 U20751 ( .A1(n17570), .A2(n17585), .ZN(n17576) );
  AND2_X1 U20752 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17576), .ZN(n17574) );
  AOI21_X1 U20753 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17578), .A(n17574), .ZN(
        n17571) );
  OAI22_X1 U20754 ( .A1(n17572), .A2(n17571), .B1(n18571), .B2(n17578), .ZN(
        P3_U2699) );
  AOI21_X1 U20755 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17578), .A(n17576), .ZN(
        n17573) );
  OAI22_X1 U20756 ( .A1(n17574), .A2(n17573), .B1(n18564), .B2(n17578), .ZN(
        P3_U2700) );
  AOI221_X1 U20757 ( .B1(n17575), .B2(n9669), .C1(n18585), .C2(n9669), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17577) );
  AOI211_X1 U20758 ( .C1(n17583), .C2(n18560), .A(n17577), .B(n17576), .ZN(
        P3_U2701) );
  INV_X1 U20759 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18555) );
  OAI222_X1 U20760 ( .A1(n17580), .A2(n17585), .B1(n17579), .B2(n9669), .C1(
        n18555), .C2(n17578), .ZN(P3_U2702) );
  INV_X1 U20761 ( .A(n9669), .ZN(n17582) );
  AOI22_X1 U20762 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17583), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17582), .ZN(n17584) );
  OAI21_X1 U20763 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17585), .A(n17584), .ZN(
        P3_U2703) );
  NAND2_X1 U20764 ( .A1(n17738), .A2(n18578), .ZN(n17649) );
  INV_X1 U20765 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17811) );
  INV_X1 U20766 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17807) );
  INV_X1 U20767 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17803) );
  INV_X1 U20768 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17801) );
  INV_X1 U20769 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17787) );
  INV_X1 U20770 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17819) );
  INV_X1 U20771 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17823) );
  INV_X1 U20772 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17821) );
  NAND4_X1 U20773 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n17587) );
  NOR3_X1 U20774 ( .A1(n17823), .A2(n17821), .A3(n17587), .ZN(n17675) );
  INV_X1 U20775 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17795) );
  INV_X1 U20776 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17793) );
  INV_X1 U20777 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17791) );
  INV_X1 U20778 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17789) );
  NOR4_X1 U20779 ( .A1(n17795), .A2(n17793), .A3(n17791), .A4(n17789), .ZN(
        n17588) );
  NAND4_X1 U20780 ( .A1(n17666), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_21__SCAN_IN), .A4(n17588), .ZN(n17631) );
  NAND2_X1 U20781 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17614), .ZN(n17610) );
  NAND2_X1 U20782 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17601), .ZN(n17597) );
  NOR2_X1 U20783 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17597), .ZN(n17591) );
  NAND2_X1 U20784 ( .A1(n17728), .A2(n17597), .ZN(n17596) );
  OAI21_X1 U20785 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17589), .A(n17596), .ZN(
        n17590) );
  AOI22_X1 U20786 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17591), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17590), .ZN(n17592) );
  OAI21_X1 U20787 ( .B1(n19610), .B2(n17649), .A(n17592), .ZN(P3_U2704) );
  INV_X1 U20788 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17815) );
  NOR2_X2 U20789 ( .A1(n18573), .A2(n17728), .ZN(n17665) );
  OAI22_X1 U20790 ( .A1(n17593), .A2(n17743), .B1(n19602), .B2(n17649), .ZN(
        n17594) );
  AOI21_X1 U20791 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17665), .A(n17594), .ZN(
        n17595) );
  OAI221_X1 U20792 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17597), .C1(n17815), 
        .C2(n17596), .A(n17595), .ZN(P3_U2705) );
  AOI22_X1 U20793 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17665), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17664), .ZN(n17599) );
  OAI211_X1 U20794 ( .C1(n17601), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17728), .B(
        n17597), .ZN(n17598) );
  OAI211_X1 U20795 ( .C1(n17600), .C2(n17743), .A(n17599), .B(n17598), .ZN(
        P3_U2706) );
  INV_X1 U20796 ( .A(n17601), .ZN(n17603) );
  OAI21_X1 U20797 ( .B1(n17738), .B2(n17811), .A(n17610), .ZN(n17602) );
  AOI22_X1 U20798 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17664), .B1(n17603), .B2(
        n17602), .ZN(n17606) );
  AOI22_X1 U20799 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17665), .B1(n17730), .B2(
        n17604), .ZN(n17605) );
  NAND2_X1 U20800 ( .A1(n17606), .A2(n17605), .ZN(P3_U2707) );
  OAI21_X1 U20801 ( .B1(n17609), .B2(n17608), .A(n17607), .ZN(n17613) );
  AOI22_X1 U20802 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17665), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17664), .ZN(n17612) );
  OAI211_X1 U20803 ( .C1(n17614), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17728), .B(
        n17610), .ZN(n17611) );
  OAI211_X1 U20804 ( .C1(n17613), .C2(n17743), .A(n17612), .B(n17611), .ZN(
        P3_U2708) );
  AOI22_X1 U20805 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17665), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17664), .ZN(n17617) );
  AOI211_X1 U20806 ( .C1(n17807), .C2(n17619), .A(n17614), .B(n17738), .ZN(
        n17615) );
  INV_X1 U20807 ( .A(n17615), .ZN(n17616) );
  OAI211_X1 U20808 ( .C1(n17618), .C2(n17743), .A(n17617), .B(n17616), .ZN(
        P3_U2709) );
  AOI22_X1 U20809 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17665), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17664), .ZN(n17621) );
  OAI211_X1 U20810 ( .C1(n17624), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17728), .B(
        n17619), .ZN(n17620) );
  OAI211_X1 U20811 ( .C1(n17622), .C2(n17743), .A(n17621), .B(n17620), .ZN(
        P3_U2710) );
  AOI22_X1 U20812 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17665), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17664), .ZN(n17628) );
  OAI21_X1 U20813 ( .B1(n17803), .B2(n17738), .A(n17623), .ZN(n17626) );
  INV_X1 U20814 ( .A(n17624), .ZN(n17625) );
  NAND2_X1 U20815 ( .A1(n17626), .A2(n17625), .ZN(n17627) );
  OAI211_X1 U20816 ( .C1(n17629), .C2(n17743), .A(n17628), .B(n17627), .ZN(
        P3_U2711) );
  AOI211_X1 U20817 ( .C1(n17801), .C2(n17631), .A(n17738), .B(n17630), .ZN(
        n17632) );
  AOI21_X1 U20818 ( .B1(n17664), .B2(BUF2_REG_23__SCAN_IN), .A(n17632), .ZN(
        n17634) );
  NAND2_X1 U20819 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17665), .ZN(n17633) );
  OAI211_X1 U20820 ( .C1(n17635), .C2(n17743), .A(n17634), .B(n17633), .ZN(
        P3_U2712) );
  NAND3_X1 U20821 ( .A1(n17711), .A2(n17666), .A3(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n17660) );
  NAND2_X1 U20822 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17650), .ZN(n17646) );
  NAND2_X1 U20823 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17642), .ZN(n17641) );
  NAND2_X1 U20824 ( .A1(n17641), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17639) );
  OAI22_X1 U20825 ( .A1(n17636), .A2(n17743), .B1(n15542), .B2(n17649), .ZN(
        n17637) );
  AOI21_X1 U20826 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17665), .A(n17637), .ZN(
        n17638) );
  OAI221_X1 U20827 ( .B1(n17641), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17639), 
        .C2(n17738), .A(n17638), .ZN(P3_U2713) );
  AOI22_X1 U20828 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17665), .B1(n17730), .B2(
        n17640), .ZN(n17644) );
  OAI211_X1 U20829 ( .C1(n17642), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17728), .B(
        n17641), .ZN(n17643) );
  OAI211_X1 U20830 ( .C1(n17649), .C2(n19594), .A(n17644), .B(n17643), .ZN(
        P3_U2714) );
  AOI22_X1 U20831 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17665), .B1(n17730), .B2(
        n17645), .ZN(n17648) );
  OAI211_X1 U20832 ( .C1(n17650), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17728), .B(
        n17646), .ZN(n17647) );
  OAI211_X1 U20833 ( .C1(n17649), .C2(n18565), .A(n17648), .B(n17647), .ZN(
        P3_U2715) );
  AOI22_X1 U20834 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17665), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17664), .ZN(n17653) );
  AOI211_X1 U20835 ( .C1(n17793), .C2(n17655), .A(n17650), .B(n17738), .ZN(
        n17651) );
  INV_X1 U20836 ( .A(n17651), .ZN(n17652) );
  OAI211_X1 U20837 ( .C1(n17654), .C2(n17743), .A(n17653), .B(n17652), .ZN(
        P3_U2716) );
  AOI22_X1 U20838 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17665), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17664), .ZN(n17658) );
  OAI211_X1 U20839 ( .C1(n17656), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17728), .B(
        n17655), .ZN(n17657) );
  OAI211_X1 U20840 ( .C1(n17659), .C2(n17743), .A(n17658), .B(n17657), .ZN(
        P3_U2717) );
  AOI22_X1 U20841 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17665), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17664), .ZN(n17662) );
  OAI211_X1 U20842 ( .C1(n17666), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17728), .B(
        n17660), .ZN(n17661) );
  OAI211_X1 U20843 ( .C1(n17663), .C2(n17743), .A(n17662), .B(n17661), .ZN(
        P3_U2718) );
  AOI22_X1 U20844 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17665), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17664), .ZN(n17669) );
  AOI211_X1 U20845 ( .C1(n17787), .C2(n17672), .A(n17738), .B(n17666), .ZN(
        n17667) );
  INV_X1 U20846 ( .A(n17667), .ZN(n17668) );
  OAI211_X1 U20847 ( .C1(n17670), .C2(n17743), .A(n17669), .B(n17668), .ZN(
        P3_U2719) );
  AOI22_X1 U20848 ( .A1(n17730), .A2(n17671), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n17741), .ZN(n17674) );
  OAI211_X1 U20849 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17677), .A(n17728), .B(
        n17672), .ZN(n17673) );
  NAND2_X1 U20850 ( .A1(n17674), .A2(n17673), .ZN(P3_U2720) );
  INV_X1 U20851 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17842) );
  INV_X1 U20852 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17837) );
  INV_X1 U20853 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17833) );
  NAND3_X1 U20854 ( .A1(n17711), .A2(n17737), .A3(n17675), .ZN(n17705) );
  NOR2_X1 U20855 ( .A1(n17833), .A2(n17705), .ZN(n17700) );
  NAND2_X1 U20856 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17700), .ZN(n17699) );
  NAND2_X1 U20857 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17694), .ZN(n17685) );
  NOR2_X1 U20858 ( .A1(n17842), .A2(n17685), .ZN(n17688) );
  NAND2_X1 U20859 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17688), .ZN(n17680) );
  AOI22_X1 U20860 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17741), .B1(n17730), .B2(
        n17676), .ZN(n17679) );
  INV_X1 U20861 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17847) );
  OR3_X1 U20862 ( .A1(n17847), .A2(n17738), .A3(n17677), .ZN(n17678) );
  OAI211_X1 U20863 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17680), .A(n17679), .B(
        n17678), .ZN(P3_U2721) );
  INV_X1 U20864 ( .A(n17680), .ZN(n17683) );
  AOI21_X1 U20865 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17728), .A(n17688), .ZN(
        n17682) );
  OAI222_X1 U20866 ( .A1(n17736), .A2(n17684), .B1(n17683), .B2(n17682), .C1(
        n17743), .C2(n17681), .ZN(P3_U2722) );
  INV_X1 U20867 ( .A(n17685), .ZN(n17692) );
  AOI21_X1 U20868 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17728), .A(n17692), .ZN(
        n17687) );
  OAI222_X1 U20869 ( .A1(n17736), .A2(n17689), .B1(n17688), .B2(n17687), .C1(
        n17743), .C2(n17686), .ZN(P3_U2723) );
  AOI21_X1 U20870 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17728), .A(n17694), .ZN(
        n17691) );
  OAI222_X1 U20871 ( .A1(n17736), .A2(n17693), .B1(n17692), .B2(n17691), .C1(
        n17743), .C2(n17690), .ZN(P3_U2724) );
  AOI211_X1 U20872 ( .C1(n17837), .C2(n17699), .A(n17738), .B(n17694), .ZN(
        n17695) );
  AOI21_X1 U20873 ( .B1(n17730), .B2(n17696), .A(n17695), .ZN(n17697) );
  OAI21_X1 U20874 ( .B1(n17698), .B2(n17736), .A(n17697), .ZN(P3_U2725) );
  INV_X1 U20875 ( .A(n17699), .ZN(n17703) );
  AOI21_X1 U20876 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17728), .A(n17700), .ZN(
        n17702) );
  OAI222_X1 U20877 ( .A1(n17736), .A2(n17704), .B1(n17703), .B2(n17702), .C1(
        n17743), .C2(n17701), .ZN(P3_U2726) );
  INV_X1 U20878 ( .A(n17705), .ZN(n17715) );
  AOI22_X1 U20879 ( .A1(n17730), .A2(n17706), .B1(n17715), .B2(n17833), .ZN(
        n17709) );
  NAND3_X1 U20880 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17728), .A3(n17707), .ZN(
        n17708) );
  OAI211_X1 U20881 ( .C1(n17736), .C2(n17710), .A(n17709), .B(n17708), .ZN(
        P3_U2727) );
  INV_X1 U20882 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17829) );
  NAND2_X1 U20883 ( .A1(n17711), .A2(n17737), .ZN(n17712) );
  NOR2_X1 U20884 ( .A1(n17823), .A2(n17732), .ZN(n17724) );
  NAND2_X1 U20885 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17727), .ZN(n17716) );
  NOR2_X1 U20886 ( .A1(n17829), .A2(n17716), .ZN(n17719) );
  AOI21_X1 U20887 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17728), .A(n17719), .ZN(
        n17714) );
  OAI222_X1 U20888 ( .A1(n18583), .A2(n17736), .B1(n17715), .B2(n17714), .C1(
        n17743), .C2(n17713), .ZN(P3_U2728) );
  INV_X1 U20889 ( .A(n17716), .ZN(n17723) );
  AOI21_X1 U20890 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17728), .A(n17723), .ZN(
        n17718) );
  OAI222_X1 U20891 ( .A1(n18577), .A2(n17736), .B1(n17719), .B2(n17718), .C1(
        n17743), .C2(n17717), .ZN(P3_U2729) );
  AOI21_X1 U20892 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17728), .A(n17727), .ZN(
        n17722) );
  INV_X1 U20893 ( .A(n17720), .ZN(n17721) );
  OAI222_X1 U20894 ( .A1(n18572), .A2(n17736), .B1(n17723), .B2(n17722), .C1(
        n17743), .C2(n17721), .ZN(P3_U2730) );
  AOI21_X1 U20895 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17728), .A(n17724), .ZN(
        n17726) );
  OAI222_X1 U20896 ( .A1(n18566), .A2(n17736), .B1(n17727), .B2(n17726), .C1(
        n17743), .C2(n17725), .ZN(P3_U2731) );
  NAND2_X1 U20897 ( .A1(n17728), .A2(n17732), .ZN(n17734) );
  AOI22_X1 U20898 ( .A1(n17741), .A2(BUF2_REG_3__SCAN_IN), .B1(n17730), .B2(
        n17729), .ZN(n17731) );
  OAI221_X1 U20899 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17732), .C1(n17823), 
        .C2(n17734), .A(n17731), .ZN(P3_U2732) );
  NOR2_X1 U20900 ( .A1(n17737), .A2(P3_EAX_REG_2__SCAN_IN), .ZN(n17733) );
  OAI222_X1 U20901 ( .A1(n17736), .A2(n18556), .B1(n17743), .B2(n17735), .C1(
        n17734), .C2(n17733), .ZN(P3_U2733) );
  AOI211_X1 U20902 ( .C1(n17819), .C2(n17739), .A(n17738), .B(n17737), .ZN(
        n17740) );
  AOI21_X1 U20903 ( .B1(n17741), .B2(BUF2_REG_1__SCAN_IN), .A(n17740), .ZN(
        n17742) );
  OAI21_X1 U20904 ( .B1(n17744), .B2(n17743), .A(n17742), .ZN(P3_U2734) );
  NAND2_X1 U20905 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17897), .ZN(n19207) );
  INV_X2 U20906 ( .A(n19207), .ZN(n17780) );
  AND2_X1 U20907 ( .A1(n17760), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20908 ( .A1(n17763), .A2(n18545), .ZN(n17762) );
  AOI22_X1 U20909 ( .A1(n17780), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17779), .ZN(n17746) );
  OAI21_X1 U20910 ( .B1(n17815), .B2(n17762), .A(n17746), .ZN(P3_U2737) );
  INV_X1 U20911 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17813) );
  AOI22_X1 U20912 ( .A1(n17780), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17747) );
  OAI21_X1 U20913 ( .B1(n17813), .B2(n17762), .A(n17747), .ZN(P3_U2738) );
  AOI22_X1 U20914 ( .A1(n17780), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17748) );
  OAI21_X1 U20915 ( .B1(n17811), .B2(n17762), .A(n17748), .ZN(P3_U2739) );
  INV_X1 U20916 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17809) );
  AOI22_X1 U20917 ( .A1(n17780), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17749) );
  OAI21_X1 U20918 ( .B1(n17809), .B2(n17762), .A(n17749), .ZN(P3_U2740) );
  AOI22_X1 U20919 ( .A1(n17780), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17750) );
  OAI21_X1 U20920 ( .B1(n17807), .B2(n17762), .A(n17750), .ZN(P3_U2741) );
  INV_X1 U20921 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17805) );
  AOI22_X1 U20922 ( .A1(n17780), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17751) );
  OAI21_X1 U20923 ( .B1(n17805), .B2(n17762), .A(n17751), .ZN(P3_U2742) );
  AOI22_X1 U20924 ( .A1(n17780), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17752) );
  OAI21_X1 U20925 ( .B1(n17803), .B2(n17762), .A(n17752), .ZN(P3_U2743) );
  AOI22_X1 U20926 ( .A1(n17780), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17753) );
  OAI21_X1 U20927 ( .B1(n17801), .B2(n17762), .A(n17753), .ZN(P3_U2744) );
  INV_X1 U20928 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U20929 ( .A1(n17780), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17754) );
  OAI21_X1 U20930 ( .B1(n17799), .B2(n17762), .A(n17754), .ZN(P3_U2745) );
  INV_X1 U20931 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17797) );
  AOI22_X1 U20932 ( .A1(n17780), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17755) );
  OAI21_X1 U20933 ( .B1(n17797), .B2(n17762), .A(n17755), .ZN(P3_U2746) );
  AOI22_X1 U20934 ( .A1(n17780), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17756) );
  OAI21_X1 U20935 ( .B1(n17795), .B2(n17762), .A(n17756), .ZN(P3_U2747) );
  AOI22_X1 U20936 ( .A1(n17780), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17757) );
  OAI21_X1 U20937 ( .B1(n17793), .B2(n17762), .A(n17757), .ZN(P3_U2748) );
  AOI22_X1 U20938 ( .A1(n17780), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17758) );
  OAI21_X1 U20939 ( .B1(n17791), .B2(n17762), .A(n17758), .ZN(P3_U2749) );
  AOI22_X1 U20940 ( .A1(n17780), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17759) );
  OAI21_X1 U20941 ( .B1(n17789), .B2(n17762), .A(n17759), .ZN(P3_U2750) );
  AOI22_X1 U20942 ( .A1(n17780), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17760), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17761) );
  OAI21_X1 U20943 ( .B1(n17787), .B2(n17762), .A(n17761), .ZN(P3_U2751) );
  AOI22_X1 U20944 ( .A1(n17780), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17764) );
  OAI21_X1 U20945 ( .B1(n9993), .B2(n17782), .A(n17764), .ZN(P3_U2752) );
  AOI22_X1 U20946 ( .A1(n17780), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17765) );
  OAI21_X1 U20947 ( .B1(n17847), .B2(n17782), .A(n17765), .ZN(P3_U2753) );
  INV_X1 U20948 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17844) );
  AOI22_X1 U20949 ( .A1(n17780), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17766) );
  OAI21_X1 U20950 ( .B1(n17844), .B2(n17782), .A(n17766), .ZN(P3_U2754) );
  AOI22_X1 U20951 ( .A1(n17780), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17767) );
  OAI21_X1 U20952 ( .B1(n17842), .B2(n17782), .A(n17767), .ZN(P3_U2755) );
  INV_X1 U20953 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17839) );
  AOI22_X1 U20954 ( .A1(n17780), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17768) );
  OAI21_X1 U20955 ( .B1(n17839), .B2(n17782), .A(n17768), .ZN(P3_U2756) );
  AOI22_X1 U20956 ( .A1(n17780), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17769) );
  OAI21_X1 U20957 ( .B1(n17837), .B2(n17782), .A(n17769), .ZN(P3_U2757) );
  INV_X1 U20958 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17835) );
  AOI22_X1 U20959 ( .A1(n17780), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17770) );
  OAI21_X1 U20960 ( .B1(n17835), .B2(n17782), .A(n17770), .ZN(P3_U2758) );
  AOI22_X1 U20961 ( .A1(n17780), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17771) );
  OAI21_X1 U20962 ( .B1(n17833), .B2(n17782), .A(n17771), .ZN(P3_U2759) );
  INV_X1 U20963 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17831) );
  AOI22_X1 U20964 ( .A1(n17780), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17772) );
  OAI21_X1 U20965 ( .B1(n17831), .B2(n17782), .A(n17772), .ZN(P3_U2760) );
  AOI22_X1 U20966 ( .A1(n17780), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17773) );
  OAI21_X1 U20967 ( .B1(n17829), .B2(n17782), .A(n17773), .ZN(P3_U2761) );
  INV_X1 U20968 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U20969 ( .A1(n17780), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17774) );
  OAI21_X1 U20970 ( .B1(n17827), .B2(n17782), .A(n17774), .ZN(P3_U2762) );
  INV_X1 U20971 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U20972 ( .A1(n17780), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17775) );
  OAI21_X1 U20973 ( .B1(n17825), .B2(n17782), .A(n17775), .ZN(P3_U2763) );
  AOI22_X1 U20974 ( .A1(n17780), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17776) );
  OAI21_X1 U20975 ( .B1(n17823), .B2(n17782), .A(n17776), .ZN(P3_U2764) );
  AOI22_X1 U20976 ( .A1(n17780), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17777) );
  OAI21_X1 U20977 ( .B1(n17821), .B2(n17782), .A(n17777), .ZN(P3_U2765) );
  AOI22_X1 U20978 ( .A1(n17780), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17778) );
  OAI21_X1 U20979 ( .B1(n17819), .B2(n17782), .A(n17778), .ZN(P3_U2766) );
  AOI22_X1 U20980 ( .A1(n17780), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17779), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17781) );
  OAI21_X1 U20981 ( .B1(n17817), .B2(n17782), .A(n17781), .ZN(P3_U2767) );
  INV_X1 U20982 ( .A(n17783), .ZN(n17784) );
  NAND2_X2 U20983 ( .A1(n17784), .A2(n19046), .ZN(n17851) );
  OAI211_X1 U20984 ( .C1(n19212), .C2(n19213), .A(n17785), .B(n17784), .ZN(
        n17845) );
  AOI22_X1 U20985 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17849), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17848), .ZN(n17786) );
  OAI21_X1 U20986 ( .B1(n17787), .B2(n17851), .A(n17786), .ZN(P3_U2768) );
  AOI22_X1 U20987 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17849), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17848), .ZN(n17788) );
  OAI21_X1 U20988 ( .B1(n17789), .B2(n17851), .A(n17788), .ZN(P3_U2769) );
  AOI22_X1 U20989 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17849), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17848), .ZN(n17790) );
  OAI21_X1 U20990 ( .B1(n17791), .B2(n17851), .A(n17790), .ZN(P3_U2770) );
  AOI22_X1 U20991 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17840), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17848), .ZN(n17792) );
  OAI21_X1 U20992 ( .B1(n17793), .B2(n17851), .A(n17792), .ZN(P3_U2771) );
  AOI22_X1 U20993 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17840), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17848), .ZN(n17794) );
  OAI21_X1 U20994 ( .B1(n17795), .B2(n17851), .A(n17794), .ZN(P3_U2772) );
  AOI22_X1 U20995 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17840), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17848), .ZN(n17796) );
  OAI21_X1 U20996 ( .B1(n17797), .B2(n17851), .A(n17796), .ZN(P3_U2773) );
  AOI22_X1 U20997 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17840), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17848), .ZN(n17798) );
  OAI21_X1 U20998 ( .B1(n17799), .B2(n17851), .A(n17798), .ZN(P3_U2774) );
  AOI22_X1 U20999 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17840), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17848), .ZN(n17800) );
  OAI21_X1 U21000 ( .B1(n17801), .B2(n17851), .A(n17800), .ZN(P3_U2775) );
  AOI22_X1 U21001 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17840), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17848), .ZN(n17802) );
  OAI21_X1 U21002 ( .B1(n17803), .B2(n17851), .A(n17802), .ZN(P3_U2776) );
  AOI22_X1 U21003 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17840), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17848), .ZN(n17804) );
  OAI21_X1 U21004 ( .B1(n17805), .B2(n17851), .A(n17804), .ZN(P3_U2777) );
  AOI22_X1 U21005 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17840), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17848), .ZN(n17806) );
  OAI21_X1 U21006 ( .B1(n17807), .B2(n17851), .A(n17806), .ZN(P3_U2778) );
  AOI22_X1 U21007 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17840), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17848), .ZN(n17808) );
  OAI21_X1 U21008 ( .B1(n17809), .B2(n17851), .A(n17808), .ZN(P3_U2779) );
  AOI22_X1 U21009 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17849), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17848), .ZN(n17810) );
  OAI21_X1 U21010 ( .B1(n17811), .B2(n17851), .A(n17810), .ZN(P3_U2780) );
  AOI22_X1 U21011 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17849), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17848), .ZN(n17812) );
  OAI21_X1 U21012 ( .B1(n17813), .B2(n17851), .A(n17812), .ZN(P3_U2781) );
  AOI22_X1 U21013 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17849), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17848), .ZN(n17814) );
  OAI21_X1 U21014 ( .B1(n17815), .B2(n17851), .A(n17814), .ZN(P3_U2782) );
  AOI22_X1 U21015 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17848), .ZN(n17816) );
  OAI21_X1 U21016 ( .B1(n17817), .B2(n17851), .A(n17816), .ZN(P3_U2783) );
  AOI22_X1 U21017 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17848), .ZN(n17818) );
  OAI21_X1 U21018 ( .B1(n17819), .B2(n17851), .A(n17818), .ZN(P3_U2784) );
  AOI22_X1 U21019 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17848), .ZN(n17820) );
  OAI21_X1 U21020 ( .B1(n17821), .B2(n17851), .A(n17820), .ZN(P3_U2785) );
  AOI22_X1 U21021 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17845), .ZN(n17822) );
  OAI21_X1 U21022 ( .B1(n17823), .B2(n17851), .A(n17822), .ZN(P3_U2786) );
  AOI22_X1 U21023 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17845), .ZN(n17824) );
  OAI21_X1 U21024 ( .B1(n17825), .B2(n17851), .A(n17824), .ZN(P3_U2787) );
  AOI22_X1 U21025 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17845), .ZN(n17826) );
  OAI21_X1 U21026 ( .B1(n17827), .B2(n17851), .A(n17826), .ZN(P3_U2788) );
  AOI22_X1 U21027 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17845), .ZN(n17828) );
  OAI21_X1 U21028 ( .B1(n17829), .B2(n17851), .A(n17828), .ZN(P3_U2789) );
  AOI22_X1 U21029 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17845), .ZN(n17830) );
  OAI21_X1 U21030 ( .B1(n17831), .B2(n17851), .A(n17830), .ZN(P3_U2790) );
  AOI22_X1 U21031 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17845), .ZN(n17832) );
  OAI21_X1 U21032 ( .B1(n17833), .B2(n17851), .A(n17832), .ZN(P3_U2791) );
  AOI22_X1 U21033 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17845), .ZN(n17834) );
  OAI21_X1 U21034 ( .B1(n17835), .B2(n17851), .A(n17834), .ZN(P3_U2792) );
  AOI22_X1 U21035 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17840), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17848), .ZN(n17836) );
  OAI21_X1 U21036 ( .B1(n17837), .B2(n17851), .A(n17836), .ZN(P3_U2793) );
  AOI22_X1 U21037 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17845), .ZN(n17838) );
  OAI21_X1 U21038 ( .B1(n17839), .B2(n17851), .A(n17838), .ZN(P3_U2794) );
  AOI22_X1 U21039 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17840), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17848), .ZN(n17841) );
  OAI21_X1 U21040 ( .B1(n17842), .B2(n17851), .A(n17841), .ZN(P3_U2795) );
  AOI22_X1 U21041 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17845), .ZN(n17843) );
  OAI21_X1 U21042 ( .B1(n17844), .B2(n17851), .A(n17843), .ZN(P3_U2796) );
  AOI22_X1 U21043 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17845), .ZN(n17846) );
  OAI21_X1 U21044 ( .B1(n17847), .B2(n17851), .A(n17846), .ZN(P3_U2797) );
  AOI22_X1 U21045 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17849), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17848), .ZN(n17850) );
  OAI21_X1 U21046 ( .B1(n9993), .B2(n17851), .A(n17850), .ZN(P3_U2798) );
  NAND2_X1 U21047 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17852), .ZN(
        n17866) );
  INV_X1 U21048 ( .A(n17897), .ZN(n18206) );
  OAI21_X1 U21049 ( .B1(n17853), .B2(n18206), .A(n18207), .ZN(n17854) );
  AOI21_X1 U21050 ( .B1(n18166), .B2(n17858), .A(n17854), .ZN(n17884) );
  OAI21_X1 U21051 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17964), .A(
        n17884), .ZN(n17867) );
  NOR2_X1 U21052 ( .A1(n18052), .A2(n17858), .ZN(n17873) );
  OAI211_X1 U21053 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17873), .B(n17859), .ZN(n17861) );
  NAND2_X1 U21054 ( .A1(n18483), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17860) );
  OAI211_X1 U21055 ( .C1(n18063), .C2(n17862), .A(n17861), .B(n17860), .ZN(
        n17863) );
  NAND2_X1 U21056 ( .A1(n18211), .A2(n18058), .ZN(n17963) );
  AOI22_X1 U21057 ( .A1(n18196), .A2(n18218), .B1(n18119), .B2(n17864), .ZN(
        n17888) );
  NAND2_X1 U21058 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17888), .ZN(
        n17875) );
  NAND3_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17963), .A3(
        n17875), .ZN(n17865) );
  AOI22_X1 U21060 ( .A1(n17970), .A2(n17868), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17867), .ZN(n17879) );
  NAND2_X1 U21061 ( .A1(n17870), .A2(n9984), .ZN(n17871) );
  XNOR2_X1 U21062 ( .A(n18109), .B(n17871), .ZN(n18224) );
  AOI22_X1 U21063 ( .A1(n18104), .A2(n18224), .B1(n17873), .B2(n17872), .ZN(
        n17878) );
  INV_X1 U21064 ( .A(n17874), .ZN(n17876) );
  OAI21_X1 U21065 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17876), .A(
        n17875), .ZN(n17877) );
  NAND2_X1 U21066 ( .A1(n18483), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18225) );
  NAND4_X1 U21067 ( .A1(n17879), .A2(n17878), .A3(n17877), .A4(n18225), .ZN(
        P3_U2803) );
  AOI21_X1 U21068 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17881), .A(
        n17880), .ZN(n18234) );
  AOI21_X1 U21069 ( .B1(n17882), .B2(n18932), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17883) );
  OAI22_X1 U21070 ( .A1(n18190), .A2(n17885), .B1(n17884), .B2(n17883), .ZN(
        n17892) );
  NOR2_X1 U21071 ( .A1(n17887), .A2(n17886), .ZN(n17890) );
  INV_X1 U21072 ( .A(n17888), .ZN(n17889) );
  MUX2_X1 U21073 ( .A(n17890), .B(n17889), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17891) );
  AOI211_X1 U21074 ( .C1(n18483), .C2(P3_REIP_REG_26__SCAN_IN), .A(n17892), 
        .B(n17891), .ZN(n17893) );
  OAI21_X1 U21075 ( .B1(n18234), .B2(n18122), .A(n17893), .ZN(P3_U2804) );
  XNOR2_X1 U21076 ( .A(n17905), .B(n17894), .ZN(n18243) );
  INV_X1 U21077 ( .A(n17895), .ZN(n17896) );
  AND2_X1 U21078 ( .A1(n17898), .A2(n18932), .ZN(n17925) );
  AOI211_X1 U21079 ( .C1(n17897), .C2(n17896), .A(n18178), .B(n17925), .ZN(
        n17928) );
  OAI21_X1 U21080 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17964), .A(
        n17928), .ZN(n17915) );
  NOR2_X1 U21081 ( .A1(n18052), .A2(n17898), .ZN(n17917) );
  OAI211_X1 U21082 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17917), .B(n17899), .ZN(n17900) );
  NAND2_X1 U21083 ( .A1(n18483), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18240) );
  OAI211_X1 U21084 ( .C1(n18063), .C2(n17901), .A(n17900), .B(n18240), .ZN(
        n17908) );
  XNOR2_X1 U21085 ( .A(n17902), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18247) );
  OAI21_X1 U21086 ( .B1(n18109), .B2(n17904), .A(n17903), .ZN(n17906) );
  XNOR2_X1 U21087 ( .A(n17906), .B(n17905), .ZN(n18242) );
  OAI22_X1 U21088 ( .A1(n18211), .A2(n18247), .B1(n18122), .B2(n18242), .ZN(
        n17907) );
  AOI211_X1 U21089 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17915), .A(
        n17908), .B(n17907), .ZN(n17909) );
  OAI21_X1 U21090 ( .B1(n18058), .B2(n18243), .A(n17909), .ZN(P3_U2805) );
  AOI21_X1 U21091 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17911), .A(
        n17910), .ZN(n18263) );
  INV_X1 U21092 ( .A(n17912), .ZN(n17913) );
  OAI22_X1 U21093 ( .A1(n18522), .A2(n19127), .B1(n18063), .B2(n17913), .ZN(
        n17914) );
  AOI221_X1 U21094 ( .B1(n17917), .B2(n17916), .C1(n17915), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17914), .ZN(n17919) );
  NOR2_X1 U21095 ( .A1(n18252), .A2(n18271), .ZN(n18249) );
  NOR2_X1 U21096 ( .A1(n18273), .A2(n18252), .ZN(n18248) );
  OAI22_X1 U21097 ( .A1(n18249), .A2(n18058), .B1(n18248), .B2(n18211), .ZN(
        n17930) );
  NOR2_X1 U21098 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18252), .ZN(
        n18258) );
  AOI22_X1 U21099 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17930), .B1(
        n18021), .B2(n18258), .ZN(n17918) );
  OAI211_X1 U21100 ( .C1(n18263), .C2(n18122), .A(n17919), .B(n17918), .ZN(
        P3_U2806) );
  AOI22_X1 U21101 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18109), .B1(
        n17920), .B2(n17938), .ZN(n17921) );
  NAND2_X1 U21102 ( .A1(n17971), .A2(n17921), .ZN(n17922) );
  XNOR2_X1 U21103 ( .A(n17922), .B(n18254), .ZN(n18269) );
  AOI22_X1 U21104 ( .A1(n17926), .A2(n17925), .B1(n17924), .B2(n17923), .ZN(
        n17927) );
  NAND2_X1 U21105 ( .A1(n18483), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18268) );
  OAI211_X1 U21106 ( .C1(n17928), .C2(n9999), .A(n17927), .B(n18268), .ZN(
        n17929) );
  AOI221_X1 U21107 ( .B1(n17931), .B2(n18254), .C1(n17930), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17929), .ZN(n17932) );
  OAI21_X1 U21108 ( .B1(n18122), .B2(n18269), .A(n17932), .ZN(P3_U2807) );
  OAI21_X1 U21109 ( .B1(n17934), .B2(n18206), .A(n18207), .ZN(n17935) );
  AOI21_X1 U21110 ( .B1(n18166), .B2(n17933), .A(n17935), .ZN(n17967) );
  OAI21_X1 U21111 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17964), .A(
        n17967), .ZN(n17951) );
  AOI22_X1 U21112 ( .A1(n17970), .A2(n17936), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17951), .ZN(n17948) );
  INV_X1 U21113 ( .A(n18011), .ZN(n17939) );
  INV_X1 U21114 ( .A(n17971), .ZN(n17937) );
  AOI221_X1 U21115 ( .B1(n17939), .B2(n17938), .C1(n18276), .C2(n17938), .A(
        n17937), .ZN(n17941) );
  XNOR2_X1 U21116 ( .A(n17941), .B(n17940), .ZN(n18283) );
  NOR2_X1 U21117 ( .A1(n18276), .A2(n18010), .ZN(n17943) );
  AOI22_X1 U21118 ( .A1(n18273), .A2(n18196), .B1(n18271), .B2(n18119), .ZN(
        n17994) );
  INV_X1 U21119 ( .A(n17994), .ZN(n18020) );
  AOI21_X1 U21120 ( .B1(n18276), .B2(n17963), .A(n18020), .ZN(n17962) );
  INV_X1 U21121 ( .A(n17962), .ZN(n17942) );
  MUX2_X1 U21122 ( .A(n17943), .B(n17942), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17944) );
  AOI21_X1 U21123 ( .B1(n18104), .B2(n18283), .A(n17944), .ZN(n17947) );
  NAND2_X1 U21124 ( .A1(n18483), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18284) );
  NOR2_X1 U21125 ( .A1(n18052), .A2(n17933), .ZN(n17953) );
  OAI211_X1 U21126 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17953), .B(n17945), .ZN(n17946) );
  NAND4_X1 U21127 ( .A1(n17948), .A2(n17947), .A3(n18284), .A4(n17946), .ZN(
        P3_U2808) );
  INV_X1 U21128 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17952) );
  OAI22_X1 U21129 ( .A1(n18522), .A2(n19121), .B1(n18063), .B2(n17949), .ZN(
        n17950) );
  AOI221_X1 U21130 ( .B1(n17953), .B2(n17952), .C1(n17951), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17950), .ZN(n17960) );
  INV_X1 U21131 ( .A(n17958), .ZN(n18290) );
  NOR3_X1 U21132 ( .A1(n17988), .A2(n18109), .A3(n17954), .ZN(n17980) );
  INV_X1 U21133 ( .A(n17955), .ZN(n17981) );
  AOI22_X1 U21134 ( .A1(n18290), .A2(n17980), .B1(n17981), .B2(n17956), .ZN(
        n17957) );
  XNOR2_X1 U21135 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17957), .ZN(
        n18295) );
  NOR2_X1 U21136 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17958), .ZN(
        n18294) );
  NAND2_X1 U21137 ( .A1(n18318), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18292) );
  NOR2_X1 U21138 ( .A1(n18010), .A2(n18292), .ZN(n17983) );
  AOI22_X1 U21139 ( .A1(n18104), .A2(n18295), .B1(n18294), .B2(n17983), .ZN(
        n17959) );
  OAI211_X1 U21140 ( .C1(n17962), .C2(n17961), .A(n17960), .B(n17959), .ZN(
        P3_U2809) );
  INV_X1 U21141 ( .A(n18292), .ZN(n18274) );
  NAND2_X1 U21142 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18274), .ZN(
        n18301) );
  AOI21_X1 U21143 ( .B1(n17963), .B2(n18301), .A(n18020), .ZN(n17987) );
  INV_X1 U21144 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18277) );
  AOI21_X1 U21145 ( .B1(n17965), .B2(n18932), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17966) );
  OAI22_X1 U21146 ( .A1(n17967), .A2(n17966), .B1(n18522), .B2(n19120), .ZN(
        n17968) );
  AOI221_X1 U21147 ( .B1(n17970), .B2(n17969), .C1(n11277), .C2(n17969), .A(
        n17968), .ZN(n17974) );
  OAI221_X1 U21148 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17995), 
        .C1(n17986), .C2(n17980), .A(n17971), .ZN(n17972) );
  XNOR2_X1 U21149 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17972), .ZN(
        n18299) );
  NOR2_X1 U21150 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17986), .ZN(
        n18298) );
  AOI22_X1 U21151 ( .A1(n18104), .A2(n18299), .B1(n17983), .B2(n18298), .ZN(
        n17973) );
  OAI211_X1 U21152 ( .C1(n17987), .C2(n18277), .A(n17974), .B(n17973), .ZN(
        P3_U2810) );
  AOI21_X1 U21153 ( .B1(n18166), .B2(n11278), .A(n18178), .ZN(n18001) );
  OAI21_X1 U21154 ( .B1(n17975), .B2(n18206), .A(n18001), .ZN(n17991) );
  NOR2_X1 U21155 ( .A1(n18052), .A2(n11278), .ZN(n17993) );
  OAI211_X1 U21156 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17993), .B(n17976), .ZN(n17977) );
  NAND2_X1 U21157 ( .A1(n18483), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18309) );
  OAI211_X1 U21158 ( .C1(n18063), .C2(n17978), .A(n17977), .B(n18309), .ZN(
        n17979) );
  AOI21_X1 U21159 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17991), .A(
        n17979), .ZN(n17985) );
  AOI21_X1 U21160 ( .B1(n17995), .B2(n17981), .A(n17980), .ZN(n17982) );
  XNOR2_X1 U21161 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n17982), .ZN(
        n18307) );
  AOI22_X1 U21162 ( .A1(n18104), .A2(n18307), .B1(n17983), .B2(n17986), .ZN(
        n17984) );
  OAI211_X1 U21163 ( .C1(n17987), .C2(n17986), .A(n17985), .B(n17984), .ZN(
        P3_U2811) );
  NAND2_X1 U21164 ( .A1(n18318), .A2(n17988), .ZN(n18326) );
  OAI22_X1 U21165 ( .A1(n18522), .A2(n19115), .B1(n18063), .B2(n17989), .ZN(
        n17990) );
  AOI221_X1 U21166 ( .B1(n17993), .B2(n17992), .C1(n17991), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17990), .ZN(n17998) );
  OAI21_X1 U21167 ( .B1(n18318), .B2(n18010), .A(n17994), .ZN(n18007) );
  AOI21_X1 U21168 ( .B1(n9883), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17995), .ZN(n17996) );
  XNOR2_X1 U21169 ( .A(n17996), .B(n17955), .ZN(n18316) );
  AOI22_X1 U21170 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18007), .B1(
        n18104), .B2(n18316), .ZN(n17997) );
  OAI211_X1 U21171 ( .C1(n18010), .C2(n18326), .A(n17998), .B(n17997), .ZN(
        P3_U2812) );
  NAND2_X1 U21172 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18005), .ZN(
        n18331) );
  AOI21_X1 U21173 ( .B1(n17999), .B2(n18932), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18002) );
  OAI22_X1 U21174 ( .A1(n18002), .A2(n18001), .B1(n18190), .B2(n18000), .ZN(
        n18003) );
  AOI21_X1 U21175 ( .B1(n18483), .B2(P3_REIP_REG_17__SCAN_IN), .A(n18003), 
        .ZN(n18009) );
  OAI21_X1 U21176 ( .B1(n18006), .B2(n18005), .A(n18004), .ZN(n18327) );
  AOI22_X1 U21177 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18007), .B1(
        n18104), .B2(n18327), .ZN(n18008) );
  OAI211_X1 U21178 ( .C1(n18010), .C2(n18331), .A(n18009), .B(n18008), .ZN(
        P3_U2813) );
  NAND2_X1 U21179 ( .A1(n9883), .A2(n11318), .ZN(n18097) );
  OAI22_X1 U21180 ( .A1(n9883), .A2(n18011), .B1(n18097), .B2(n9880), .ZN(
        n18012) );
  XNOR2_X1 U21181 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n18012), .ZN(
        n18342) );
  AOI21_X1 U21182 ( .B1(n18166), .B2(n18014), .A(n18178), .ZN(n18046) );
  OAI21_X1 U21183 ( .B1(n18013), .B2(n18206), .A(n18046), .ZN(n18025) );
  AOI22_X1 U21184 ( .A1(n18483), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18025), .ZN(n18017) );
  NOR2_X1 U21185 ( .A1(n18052), .A2(n18014), .ZN(n18027) );
  OAI211_X1 U21186 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18027), .B(n18015), .ZN(n18016) );
  OAI211_X1 U21187 ( .C1(n18063), .C2(n18018), .A(n18017), .B(n18016), .ZN(
        n18019) );
  AOI221_X1 U21188 ( .B1(n18021), .B2(n18334), .C1(n18020), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n18019), .ZN(n18022) );
  OAI21_X1 U21189 ( .B1(n18342), .B2(n18122), .A(n18022), .ZN(P3_U2814) );
  OAI21_X1 U21190 ( .B1(n18039), .B2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18273), .ZN(n18348) );
  OAI22_X1 U21191 ( .A1(n18522), .A2(n19109), .B1(n18063), .B2(n18023), .ZN(
        n18024) );
  AOI221_X1 U21192 ( .B1(n18027), .B2(n18026), .C1(n18025), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18024), .ZN(n18036) );
  AND3_X1 U21193 ( .A1(n18378), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18030) );
  AOI21_X1 U21194 ( .B1(n18028), .B2(n18030), .A(n18029), .ZN(n18031) );
  AOI221_X1 U21195 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18398), 
        .C1(n18109), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n18031), .ZN(
        n18032) );
  XNOR2_X1 U21196 ( .A(n18032), .B(n18345), .ZN(n18353) );
  NOR2_X1 U21197 ( .A1(n18343), .A2(n18058), .ZN(n18034) );
  NAND2_X1 U21198 ( .A1(n18345), .A2(n18344), .ZN(n18033) );
  AOI22_X1 U21199 ( .A1(n18104), .A2(n18353), .B1(n18034), .B2(n18033), .ZN(
        n18035) );
  OAI211_X1 U21200 ( .C1(n18211), .C2(n18348), .A(n18036), .B(n18035), .ZN(
        P3_U2815) );
  AOI21_X1 U21201 ( .B1(n18037), .B2(n18932), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18045) );
  AOI22_X1 U21202 ( .A1(n18483), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n18038), 
        .B2(n17923), .ZN(n18044) );
  AOI221_X1 U21203 ( .B1(n18404), .B2(n18361), .C1(n18347), .C2(n18361), .A(
        n18039), .ZN(n18368) );
  OAI21_X1 U21204 ( .B1(n18347), .B2(n18097), .A(n18040), .ZN(n18041) );
  XNOR2_X1 U21205 ( .A(n18041), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18366) );
  INV_X1 U21206 ( .A(n18347), .ZN(n18357) );
  OAI221_X1 U21207 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18357), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n11318), .A(n18344), .ZN(
        n18365) );
  OAI22_X1 U21208 ( .A1(n18366), .A2(n18122), .B1(n18058), .B2(n18365), .ZN(
        n18042) );
  AOI21_X1 U21209 ( .B1(n18196), .B2(n18368), .A(n18042), .ZN(n18043) );
  OAI211_X1 U21210 ( .C1(n18046), .C2(n18045), .A(n18044), .B(n18043), .ZN(
        P3_U2816) );
  INV_X1 U21211 ( .A(n18378), .ZN(n18388) );
  NOR2_X1 U21212 ( .A1(n18398), .A2(n18388), .ZN(n18389) );
  AOI22_X1 U21213 ( .A1(n18389), .A2(n18028), .B1(n18398), .B2(n18109), .ZN(
        n18047) );
  AOI21_X1 U21214 ( .B1(n18109), .B2(n18068), .A(n18047), .ZN(n18048) );
  XNOR2_X1 U21215 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18048), .ZN(
        n18387) );
  AOI21_X1 U21216 ( .B1(n18166), .B2(n18051), .A(n18178), .ZN(n18049) );
  OAI21_X1 U21217 ( .B1(n18050), .B2(n18206), .A(n18049), .ZN(n18065) );
  NOR2_X1 U21218 ( .A1(n18052), .A2(n18051), .ZN(n18067) );
  OAI211_X1 U21219 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18067), .B(n18053), .ZN(n18055) );
  NAND2_X1 U21220 ( .A1(n18483), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18054) );
  OAI211_X1 U21221 ( .C1(n18063), .C2(n18056), .A(n18055), .B(n18054), .ZN(
        n18057) );
  AOI21_X1 U21222 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18065), .A(
        n18057), .ZN(n18061) );
  INV_X1 U21223 ( .A(n18389), .ZN(n18059) );
  NOR2_X1 U21224 ( .A1(n18081), .A2(n18059), .ZN(n18380) );
  NOR2_X1 U21225 ( .A1(n18404), .A2(n18059), .ZN(n18379) );
  OAI22_X1 U21226 ( .A1(n18380), .A2(n18058), .B1(n18379), .B2(n18211), .ZN(
        n18070) );
  NOR2_X1 U21227 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18059), .ZN(
        n18374) );
  AOI22_X1 U21228 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18070), .B1(
        n18374), .B2(n18093), .ZN(n18060) );
  OAI211_X1 U21229 ( .C1(n18122), .C2(n18387), .A(n18061), .B(n18060), .ZN(
        P3_U2817) );
  NAND2_X1 U21230 ( .A1(n18483), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18396) );
  OAI21_X1 U21231 ( .B1(n18063), .B2(n18062), .A(n18396), .ZN(n18064) );
  AOI221_X1 U21232 ( .B1(n18067), .B2(n18066), .C1(n18065), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18064), .ZN(n18073) );
  OAI21_X1 U21233 ( .B1(n18388), .B2(n18097), .A(n18068), .ZN(n18069) );
  XNOR2_X1 U21234 ( .A(n18069), .B(n18398), .ZN(n18395) );
  AOI22_X1 U21235 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18070), .B1(
        n18104), .B2(n18395), .ZN(n18072) );
  NAND3_X1 U21236 ( .A1(n18378), .A2(n18398), .A3(n18093), .ZN(n18071) );
  NAND3_X1 U21237 ( .A1(n18073), .A2(n18072), .A3(n18071), .ZN(P3_U2818) );
  INV_X1 U21238 ( .A(n18097), .ZN(n18075) );
  INV_X1 U21239 ( .A(n18418), .ZN(n18082) );
  AOI21_X1 U21240 ( .B1(n18075), .B2(n18082), .A(n18074), .ZN(n18076) );
  XNOR2_X1 U21241 ( .A(n18076), .B(n18375), .ZN(n18411) );
  NOR3_X1 U21242 ( .A1(n18112), .A2(n18077), .A3(n18776), .ZN(n18102) );
  NAND2_X1 U21243 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18102), .ZN(
        n18087) );
  NAND3_X1 U21244 ( .A1(n18099), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n18087), .ZN(n18078) );
  NAND2_X1 U21245 ( .A1(n18483), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18409) );
  OAI211_X1 U21246 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18087), .A(
        n18078), .B(n18409), .ZN(n18079) );
  AOI21_X1 U21247 ( .B1(n18080), .B2(n17923), .A(n18079), .ZN(n18085) );
  INV_X1 U21248 ( .A(n18093), .ZN(n18107) );
  AOI22_X1 U21249 ( .A1(n18196), .A2(n18404), .B1(n18119), .B2(n18081), .ZN(
        n18106) );
  OAI21_X1 U21250 ( .B1(n18082), .B2(n18107), .A(n18106), .ZN(n18083) );
  NOR2_X1 U21251 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18418), .ZN(
        n18407) );
  AOI22_X1 U21252 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18083), .B1(
        n18407), .B2(n18093), .ZN(n18084) );
  OAI211_X1 U21253 ( .C1(n18411), .C2(n18122), .A(n18085), .B(n18084), .ZN(
        P3_U2819) );
  AOI22_X1 U21254 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18097), .B1(
        n18096), .B2(n11134), .ZN(n18086) );
  XOR2_X1 U21255 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18086), .Z(
        n18413) );
  NOR2_X1 U21256 ( .A1(n18522), .A2(n19099), .ZN(n18092) );
  INV_X1 U21257 ( .A(n18087), .ZN(n18090) );
  AOI21_X1 U21258 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18099), .A(
        n18102), .ZN(n18089) );
  OAI22_X1 U21259 ( .A1(n18090), .A2(n18089), .B1(n18190), .B2(n18088), .ZN(
        n18091) );
  AOI211_X1 U21260 ( .C1(n18104), .C2(n18413), .A(n18092), .B(n18091), .ZN(
        n18095) );
  OAI211_X1 U21261 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n18093), .B(n18418), .ZN(
        n18094) );
  OAI211_X1 U21262 ( .C1(n18106), .C2(n11133), .A(n18095), .B(n18094), .ZN(
        P3_U2820) );
  NAND2_X1 U21263 ( .A1(n18097), .A2(n18096), .ZN(n18098) );
  XNOR2_X1 U21264 ( .A(n18098), .B(n11134), .ZN(n18426) );
  NOR2_X1 U21265 ( .A1(n18522), .A2(n19097), .ZN(n18425) );
  NOR2_X1 U21266 ( .A1(n18112), .A2(n18776), .ZN(n18126) );
  AOI22_X1 U21267 ( .A1(n18126), .A2(n18110), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18099), .ZN(n18101) );
  OAI22_X1 U21268 ( .A1(n18102), .A2(n18101), .B1(n18190), .B2(n18100), .ZN(
        n18103) );
  AOI211_X1 U21269 ( .C1(n18104), .C2(n18426), .A(n18425), .B(n18103), .ZN(
        n18105) );
  OAI221_X1 U21270 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18107), .C1(
        n11134), .C2(n18106), .A(n18105), .ZN(P3_U2821) );
  AOI21_X1 U21271 ( .B1(n18109), .B2(n18432), .A(n18108), .ZN(n18434) );
  AOI211_X1 U21272 ( .C1(n18113), .C2(n18111), .A(n18110), .B(n18776), .ZN(
        n18115) );
  AOI21_X1 U21273 ( .B1(n18166), .B2(n18112), .A(n18178), .ZN(n18123) );
  OAI22_X1 U21274 ( .A1(n18123), .A2(n18113), .B1(n18522), .B2(n19096), .ZN(
        n18114) );
  AOI211_X1 U21275 ( .C1(n18116), .C2(n17923), .A(n18115), .B(n18114), .ZN(
        n18121) );
  AOI21_X1 U21276 ( .B1(n18118), .B2(n18442), .A(n18117), .ZN(n18436) );
  AOI22_X1 U21277 ( .A1(n18196), .A2(n18436), .B1(n18119), .B2(n9884), .ZN(
        n18120) );
  OAI211_X1 U21278 ( .C1(n18434), .C2(n18122), .A(n18121), .B(n18120), .ZN(
        P3_U2822) );
  INV_X1 U21279 ( .A(n18123), .ZN(n18124) );
  NOR2_X1 U21280 ( .A1(n18522), .A2(n19093), .ZN(n18449) );
  AOI221_X1 U21281 ( .B1(n18126), .B2(n18125), .C1(n18124), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18449), .ZN(n18134) );
  NAND2_X1 U21282 ( .A1(n18128), .A2(n18127), .ZN(n18129) );
  XNOR2_X1 U21283 ( .A(n18129), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18450) );
  AOI21_X1 U21284 ( .B1(n18132), .B2(n18131), .A(n18130), .ZN(n18451) );
  AOI22_X1 U21285 ( .A1(n18196), .A2(n18450), .B1(n18199), .B2(n18451), .ZN(
        n18133) );
  OAI211_X1 U21286 ( .C1(n18190), .C2(n18135), .A(n18134), .B(n18133), .ZN(
        P3_U2823) );
  AOI21_X1 U21287 ( .B1(n18137), .B2(n18136), .A(n9787), .ZN(n18460) );
  NAND2_X1 U21288 ( .A1(n17171), .A2(n18932), .ZN(n18138) );
  INV_X1 U21289 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19091) );
  OAI22_X1 U21290 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18138), .B1(
        n18522), .B2(n19091), .ZN(n18139) );
  AOI21_X1 U21291 ( .B1(n18199), .B2(n18460), .A(n18139), .ZN(n18143) );
  AOI21_X1 U21292 ( .B1(n18141), .B2(n18457), .A(n18140), .ZN(n18459) );
  AOI21_X1 U21293 ( .B1(n17171), .B2(n18932), .A(n18203), .ZN(n18155) );
  AOI22_X1 U21294 ( .A1(n18196), .A2(n18459), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18155), .ZN(n18142) );
  OAI211_X1 U21295 ( .C1(n18190), .C2(n18144), .A(n18143), .B(n18142), .ZN(
        P3_U2824) );
  AOI21_X1 U21296 ( .B1(n18147), .B2(n18146), .A(n18145), .ZN(n18464) );
  AOI22_X1 U21297 ( .A1(n18196), .A2(n18464), .B1(n18483), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18157) );
  AOI222_X1 U21298 ( .A1(n18467), .A2(n18151), .B1(n18467), .B2(n18150), .C1(
        n18149), .C2(n18148), .ZN(n18465) );
  OAI21_X1 U21299 ( .B1(n18178), .B2(n18153), .A(n18152), .ZN(n18154) );
  AOI22_X1 U21300 ( .A1(n18199), .A2(n18465), .B1(n18155), .B2(n18154), .ZN(
        n18156) );
  OAI211_X1 U21301 ( .C1(n18190), .C2(n18158), .A(n18157), .B(n18156), .ZN(
        P3_U2825) );
  AOI21_X1 U21302 ( .B1(n18480), .B2(n18160), .A(n18159), .ZN(n18477) );
  OAI22_X1 U21303 ( .A1(n18522), .A2(n19087), .B1(n18776), .B2(n18161), .ZN(
        n18162) );
  AOI21_X1 U21304 ( .B1(n18196), .B2(n18477), .A(n18162), .ZN(n18169) );
  AOI21_X1 U21305 ( .B1(n18165), .B2(n18164), .A(n18163), .ZN(n18475) );
  INV_X1 U21306 ( .A(n18166), .ZN(n18167) );
  OAI21_X1 U21307 ( .B1(n17199), .B2(n18167), .A(n18207), .ZN(n18180) );
  AOI22_X1 U21308 ( .A1(n18199), .A2(n18475), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18180), .ZN(n18168) );
  OAI211_X1 U21309 ( .C1(n18190), .C2(n18170), .A(n18169), .B(n18168), .ZN(
        P3_U2826) );
  AOI21_X1 U21310 ( .B1(n18173), .B2(n18172), .A(n18171), .ZN(n18482) );
  AOI22_X1 U21311 ( .A1(n18199), .A2(n18482), .B1(n18483), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n18182) );
  AOI21_X1 U21312 ( .B1(n18176), .B2(n18175), .A(n18174), .ZN(n18487) );
  OAI21_X1 U21313 ( .B1(n18178), .B2(n18193), .A(n18177), .ZN(n18179) );
  AOI22_X1 U21314 ( .A1(n18196), .A2(n18487), .B1(n18180), .B2(n18179), .ZN(
        n18181) );
  OAI211_X1 U21315 ( .C1(n18190), .C2(n18183), .A(n18182), .B(n18181), .ZN(
        P3_U2827) );
  AOI21_X1 U21316 ( .B1(n18186), .B2(n18185), .A(n18184), .ZN(n18503) );
  INV_X1 U21317 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19083) );
  NOR2_X1 U21318 ( .A1(n18522), .A2(n19083), .ZN(n18505) );
  XNOR2_X1 U21319 ( .A(n18188), .B(n18187), .ZN(n18502) );
  OAI22_X1 U21320 ( .A1(n18190), .A2(n18189), .B1(n18211), .B2(n18502), .ZN(
        n18191) );
  AOI211_X1 U21321 ( .C1(n18199), .C2(n18503), .A(n18505), .B(n18191), .ZN(
        n18192) );
  OAI221_X1 U21322 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18776), .C1(
        n18193), .C2(n18207), .A(n18192), .ZN(P3_U2828) );
  NOR2_X1 U21323 ( .A1(n18205), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18194) );
  XOR2_X1 U21324 ( .A(n18194), .B(n18198), .Z(n18519) );
  INV_X1 U21325 ( .A(n18519), .ZN(n18195) );
  AOI22_X1 U21326 ( .A1(n18196), .A2(n18195), .B1(n18483), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18201) );
  AOI21_X1 U21327 ( .B1(n18198), .B2(n18204), .A(n18197), .ZN(n18514) );
  AOI22_X1 U21328 ( .A1(n18199), .A2(n18514), .B1(n18202), .B2(n17923), .ZN(
        n18200) );
  OAI211_X1 U21329 ( .C1(n18203), .C2(n18202), .A(n18201), .B(n18200), .ZN(
        P3_U2829) );
  OAI21_X1 U21330 ( .B1(n18205), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18204), .ZN(n18526) );
  INV_X1 U21331 ( .A(n18526), .ZN(n18524) );
  NAND3_X1 U21332 ( .A1(n19171), .A2(n18207), .A3(n18206), .ZN(n18208) );
  AOI22_X1 U21333 ( .A1(n18483), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18208), .ZN(n18209) );
  OAI221_X1 U21334 ( .B1(n18524), .B2(n18211), .C1(n18526), .C2(n18210), .A(
        n18209), .ZN(P3_U2830) );
  NAND2_X1 U21335 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18214) );
  NOR2_X1 U21336 ( .A1(n19188), .A2(n18414), .ZN(n18399) );
  NAND2_X1 U21337 ( .A1(n18315), .A2(n18399), .ZN(n18337) );
  OAI21_X1 U21338 ( .B1(n18276), .B2(n18337), .A(n19015), .ZN(n18278) );
  OAI221_X1 U21339 ( .B1(n18493), .B2(n18213), .C1(n18493), .C2(n18212), .A(
        n18278), .ZN(n18251) );
  AOI21_X1 U21340 ( .B1(n18472), .B2(n18214), .A(n18251), .ZN(n18235) );
  INV_X1 U21341 ( .A(n18501), .ZN(n18990) );
  OAI22_X1 U21342 ( .A1(n19007), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18400), .B2(n18215), .ZN(n18216) );
  AOI211_X1 U21343 ( .C1(n18990), .C2(n18218), .A(n18217), .B(n18216), .ZN(
        n18219) );
  OAI211_X1 U21344 ( .C1(n18220), .C2(n18401), .A(n18235), .B(n18219), .ZN(
        n18227) );
  AOI21_X1 U21345 ( .B1(n19002), .B2(n18228), .A(n18227), .ZN(n18222) );
  AOI221_X1 U21346 ( .B1(n18222), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n18221), .C2(n11149), .A(n18510), .ZN(n18223) );
  AOI21_X1 U21347 ( .B1(n9631), .B2(n18224), .A(n18223), .ZN(n18226) );
  OAI211_X1 U21348 ( .C1(n18511), .C2(n11149), .A(n18226), .B(n18225), .ZN(
        P3_U2835) );
  NAND2_X1 U21349 ( .A1(n18483), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18233) );
  NOR2_X1 U21350 ( .A1(n18227), .A2(n18228), .ZN(n18229) );
  OAI22_X1 U21351 ( .A1(n18510), .A2(n18229), .B1(n18511), .B2(n18228), .ZN(
        n18230) );
  OAI21_X1 U21352 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18231), .A(
        n18230), .ZN(n18232) );
  OAI211_X1 U21353 ( .C1(n18234), .C2(n21258), .A(n18233), .B(n18232), .ZN(
        P3_U2836) );
  OAI211_X1 U21354 ( .C1(n18236), .C2(n19023), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18235), .ZN(n18237) );
  OAI221_X1 U21355 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18239), 
        .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18238), .A(n18237), .ZN(
        n18241) );
  OAI21_X1 U21356 ( .B1(n18466), .B2(n18241), .A(n18240), .ZN(n18245) );
  OAI22_X1 U21357 ( .A1(n18431), .A2(n18243), .B1(n21258), .B2(n18242), .ZN(
        n18244) );
  AOI211_X1 U21358 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18520), .A(
        n18245), .B(n18244), .ZN(n18246) );
  OAI21_X1 U21359 ( .B1(n18518), .B2(n18247), .A(n18246), .ZN(P3_U2837) );
  OAI22_X1 U21360 ( .A1(n18249), .A2(n18401), .B1(n18248), .B2(n18501), .ZN(
        n18250) );
  NOR3_X1 U21361 ( .A1(n18520), .A2(n18251), .A3(n18250), .ZN(n18257) );
  OAI22_X1 U21362 ( .A1(n18992), .A2(n18254), .B1(n18253), .B2(n18252), .ZN(
        n18255) );
  AOI21_X1 U21363 ( .B1(n18257), .B2(n18255), .A(n18483), .ZN(n18265) );
  AOI21_X1 U21364 ( .B1(n18440), .B2(n18257), .A(n18256), .ZN(n18260) );
  NOR2_X1 U21365 ( .A1(n18293), .A2(n18510), .ZN(n18259) );
  AOI22_X1 U21366 ( .A1(n18265), .A2(n18260), .B1(n18259), .B2(n18258), .ZN(
        n18262) );
  NAND2_X1 U21367 ( .A1(n18483), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18261) );
  OAI211_X1 U21368 ( .C1(n18263), .C2(n21258), .A(n18262), .B(n18261), .ZN(
        P3_U2838) );
  NOR2_X1 U21369 ( .A1(n18520), .A2(n18264), .ZN(n18266) );
  OAI21_X1 U21370 ( .B1(n18266), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n18265), .ZN(n18267) );
  OAI211_X1 U21371 ( .C1(n18269), .C2(n21258), .A(n18268), .B(n18267), .ZN(
        P3_U2839) );
  INV_X1 U21372 ( .A(n18270), .ZN(n18282) );
  AOI22_X1 U21373 ( .A1(n18990), .A2(n18273), .B1(n18272), .B2(n18271), .ZN(
        n18338) );
  OAI221_X1 U21374 ( .B1(n19023), .B2(n18319), .C1(n19023), .C2(n18274), .A(
        n18338), .ZN(n18275) );
  AOI221_X1 U21375 ( .B1(n18317), .B2(n19002), .C1(n18301), .C2(n19002), .A(
        n18275), .ZN(n18288) );
  NAND2_X1 U21376 ( .A1(n18501), .A2(n18401), .ZN(n18417) );
  AOI22_X1 U21377 ( .A1(n19002), .A2(n18277), .B1(n18276), .B2(n18417), .ZN(
        n18289) );
  NAND3_X1 U21378 ( .A1(n18288), .A2(n18289), .A3(n18278), .ZN(n18280) );
  OAI22_X1 U21379 ( .A1(n18382), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n18290), .B2(n19023), .ZN(n18279) );
  NOR2_X1 U21380 ( .A1(n18280), .A2(n18279), .ZN(n18281) );
  MUX2_X1 U21381 ( .A(n18282), .B(n18281), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n18286) );
  AOI22_X1 U21382 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18520), .B1(
        n9631), .B2(n18283), .ZN(n18285) );
  OAI211_X1 U21383 ( .C1(n18510), .C2(n18286), .A(n18285), .B(n18284), .ZN(
        P3_U2840) );
  OAI21_X1 U21384 ( .B1(n18337), .B2(n18292), .A(n19015), .ZN(n18287) );
  NAND3_X1 U21385 ( .A1(n18288), .A2(n18521), .A3(n18287), .ZN(n18300) );
  NOR2_X1 U21386 ( .A1(n18992), .A2(n19015), .ZN(n18509) );
  OAI21_X1 U21387 ( .B1(n18290), .B2(n18509), .A(n18289), .ZN(n18291) );
  OAI21_X1 U21388 ( .B1(n18300), .B2(n18291), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18297) );
  NOR3_X1 U21389 ( .A1(n18293), .A2(n18466), .A3(n18292), .ZN(n18306) );
  AOI22_X1 U21390 ( .A1(n9631), .A2(n18295), .B1(n18294), .B2(n18306), .ZN(
        n18296) );
  OAI221_X1 U21391 ( .B1(n18483), .B2(n18297), .C1(n18522), .C2(n19121), .A(
        n18296), .ZN(P3_U2841) );
  AOI22_X1 U21392 ( .A1(n9631), .A2(n18299), .B1(n18298), .B2(n18306), .ZN(
        n18305) );
  AOI21_X1 U21393 ( .B1(n18417), .B2(n18301), .A(n18300), .ZN(n18302) );
  NOR2_X1 U21394 ( .A1(n18483), .A2(n18302), .ZN(n18308) );
  NOR3_X1 U21395 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18509), .A3(
        n19222), .ZN(n18303) );
  OAI21_X1 U21396 ( .B1(n18308), .B2(n18303), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18304) );
  OAI211_X1 U21397 ( .C1(n19120), .C2(n18522), .A(n18305), .B(n18304), .ZN(
        P3_U2842) );
  INV_X1 U21398 ( .A(n18306), .ZN(n18311) );
  AOI22_X1 U21399 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18308), .B1(
        n9631), .B2(n18307), .ZN(n18310) );
  OAI211_X1 U21400 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18311), .A(
        n18310), .B(n18309), .ZN(P3_U2843) );
  OAI22_X1 U21401 ( .A1(n19023), .A2(n18498), .B1(n18471), .B2(n18491), .ZN(
        n18312) );
  INV_X1 U21402 ( .A(n18312), .ZN(n18484) );
  NOR2_X1 U21403 ( .A1(n18484), .A2(n18441), .ZN(n18448) );
  NAND2_X1 U21404 ( .A1(n18313), .A2(n18448), .ZN(n18346) );
  NOR2_X1 U21405 ( .A1(n18510), .A2(n18346), .ZN(n18371) );
  AOI22_X1 U21406 ( .A1(n18315), .A2(n18371), .B1(n18521), .B2(n18314), .ZN(
        n18332) );
  AOI22_X1 U21407 ( .A1(n18483), .A2(P3_REIP_REG_18__SCAN_IN), .B1(n9631), 
        .B2(n18316), .ZN(n18325) );
  NOR2_X1 U21408 ( .A1(n18400), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18495) );
  NOR3_X1 U21409 ( .A1(n18495), .A2(n18334), .A3(n18317), .ZN(n18322) );
  OAI21_X1 U21410 ( .B1(n18319), .B2(n19023), .A(n18318), .ZN(n18320) );
  OAI21_X1 U21411 ( .B1(n18992), .B2(n18417), .A(n18320), .ZN(n18321) );
  OAI211_X1 U21412 ( .C1(n18493), .C2(n18322), .A(n18338), .B(n18321), .ZN(
        n18328) );
  OAI21_X1 U21413 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18493), .A(
        n18521), .ZN(n18323) );
  OAI211_X1 U21414 ( .C1(n18328), .C2(n18323), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n18522), .ZN(n18324) );
  OAI211_X1 U21415 ( .C1(n18332), .C2(n18326), .A(n18325), .B(n18324), .ZN(
        P3_U2844) );
  AOI22_X1 U21416 ( .A1(n18483), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n9631), 
        .B2(n18327), .ZN(n18330) );
  OAI221_X1 U21417 ( .B1(n18520), .B2(n18521), .C1(n18520), .C2(n18328), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18329) );
  OAI211_X1 U21418 ( .C1(n18332), .C2(n18331), .A(n18330), .B(n18329), .ZN(
        P3_U2845) );
  INV_X1 U21419 ( .A(n18332), .ZN(n18333) );
  AOI22_X1 U21420 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18483), .B1(n18334), 
        .B2(n18333), .ZN(n18341) );
  AOI22_X1 U21421 ( .A1(n18992), .A2(n18376), .B1(n19002), .B2(n18414), .ZN(
        n18358) );
  AOI21_X1 U21422 ( .B1(n18335), .B2(n18358), .A(n18382), .ZN(n18336) );
  AOI211_X1 U21423 ( .C1(n18337), .C2(n19015), .A(n18345), .B(n18336), .ZN(
        n18350) );
  OAI211_X1 U21424 ( .C1(n18440), .C2(n18350), .A(n18521), .B(n18338), .ZN(
        n18339) );
  NAND3_X1 U21425 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18522), .A3(
        n18339), .ZN(n18340) );
  OAI211_X1 U21426 ( .C1(n18342), .C2(n21258), .A(n18341), .B(n18340), .ZN(
        P3_U2846) );
  AOI211_X1 U21427 ( .C1(n18345), .C2(n18344), .A(n18343), .B(n18401), .ZN(
        n18352) );
  NOR2_X1 U21428 ( .A1(n18347), .A2(n18346), .ZN(n18363) );
  AOI21_X1 U21429 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18363), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18349) );
  OAI22_X1 U21430 ( .A1(n18350), .A2(n18349), .B1(n18501), .B2(n18348), .ZN(
        n18351) );
  AOI211_X1 U21431 ( .C1(n18354), .C2(n18353), .A(n18352), .B(n18351), .ZN(
        n18356) );
  AOI22_X1 U21432 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18520), .B1(
        n18483), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18355) );
  OAI21_X1 U21433 ( .B1(n18356), .B2(n18466), .A(n18355), .ZN(P3_U2847) );
  INV_X1 U21434 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19108) );
  AOI21_X1 U21435 ( .B1(n18399), .B2(n18389), .A(n18400), .ZN(n18384) );
  OAI22_X1 U21436 ( .A1(n19007), .A2(n18357), .B1(n18389), .B2(n19023), .ZN(
        n18360) );
  OAI21_X1 U21437 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18509), .A(
        n18358), .ZN(n18359) );
  NOR4_X1 U21438 ( .A1(n18384), .A2(n18361), .A3(n18360), .A4(n18359), .ZN(
        n18362) );
  NOR2_X1 U21439 ( .A1(n18362), .A2(n18510), .ZN(n18364) );
  AOI222_X1 U21440 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18364), 
        .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18520), .C1(n18364), 
        .C2(n18363), .ZN(n18370) );
  OAI22_X1 U21441 ( .A1(n18366), .A2(n21258), .B1(n18431), .B2(n18365), .ZN(
        n18367) );
  AOI21_X1 U21442 ( .B1(n18527), .B2(n18368), .A(n18367), .ZN(n18369) );
  OAI211_X1 U21443 ( .C1(n18522), .C2(n19108), .A(n18370), .B(n18369), .ZN(
        P3_U2848) );
  AOI21_X1 U21444 ( .B1(n18372), .B2(n11318), .A(n18371), .ZN(n18373) );
  OAI21_X1 U21445 ( .B1(n18404), .B2(n18518), .A(n18373), .ZN(n18412) );
  AOI22_X1 U21446 ( .A1(n18483), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18374), 
        .B2(n18412), .ZN(n18386) );
  AOI21_X1 U21447 ( .B1(n19002), .B2(n18375), .A(n18398), .ZN(n18391) );
  AND2_X1 U21448 ( .A1(n18992), .A2(n18376), .ZN(n18403) );
  OAI21_X1 U21449 ( .B1(n18418), .B2(n18414), .A(n19002), .ZN(n18377) );
  OAI21_X1 U21450 ( .B1(n18378), .B2(n19023), .A(n18377), .ZN(n18405) );
  OAI22_X1 U21451 ( .A1(n18380), .A2(n18401), .B1(n18379), .B2(n18501), .ZN(
        n18381) );
  NOR3_X1 U21452 ( .A1(n18403), .A2(n18405), .A3(n18381), .ZN(n18390) );
  OAI211_X1 U21453 ( .C1(n18382), .C2(n18391), .A(n18521), .B(n18390), .ZN(
        n18383) );
  OAI211_X1 U21454 ( .C1(n18384), .C2(n18383), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18522), .ZN(n18385) );
  OAI211_X1 U21455 ( .C1(n18387), .C2(n21258), .A(n18386), .B(n18385), .ZN(
        P3_U2849) );
  INV_X1 U21456 ( .A(n18412), .ZN(n18430) );
  OAI22_X1 U21457 ( .A1(n18430), .A2(n18388), .B1(n18398), .B2(n18510), .ZN(
        n18394) );
  AND2_X1 U21458 ( .A1(n18399), .A2(n18389), .ZN(n18392) );
  OAI211_X1 U21459 ( .C1(n18392), .C2(n18400), .A(n18391), .B(n18390), .ZN(
        n18393) );
  AOI22_X1 U21460 ( .A1(n9631), .A2(n18395), .B1(n18394), .B2(n18393), .ZN(
        n18397) );
  OAI211_X1 U21461 ( .C1(n18511), .C2(n18398), .A(n18397), .B(n18396), .ZN(
        P3_U2850) );
  OAI22_X1 U21462 ( .A1(n11318), .A2(n18401), .B1(n18400), .B2(n18399), .ZN(
        n18402) );
  AOI211_X1 U21463 ( .C1(n18404), .C2(n18990), .A(n18403), .B(n18402), .ZN(
        n18416) );
  AOI221_X1 U21464 ( .B1(n19015), .B2(n18418), .C1(n18417), .C2(n18418), .A(
        n18405), .ZN(n18406) );
  OAI221_X1 U21465 ( .B1(n18466), .B2(n18416), .C1(n18466), .C2(n18406), .A(
        n18511), .ZN(n18408) );
  AOI22_X1 U21466 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18408), .B1(
        n18407), .B2(n18412), .ZN(n18410) );
  OAI211_X1 U21467 ( .C1(n18411), .C2(n21258), .A(n18410), .B(n18409), .ZN(
        P3_U2851) );
  NAND2_X1 U21468 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18412), .ZN(
        n18423) );
  AOI22_X1 U21469 ( .A1(n18483), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n9631), 
        .B2(n18413), .ZN(n18422) );
  NAND2_X1 U21470 ( .A1(n19002), .A2(n18414), .ZN(n18415) );
  NAND3_X1 U21471 ( .A1(n18521), .A2(n18416), .A3(n18415), .ZN(n18424) );
  NAND2_X1 U21472 ( .A1(n18418), .A2(n18417), .ZN(n18419) );
  OAI21_X1 U21473 ( .B1(n18440), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18419), .ZN(n18420) );
  OAI211_X1 U21474 ( .C1(n18424), .C2(n18420), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18522), .ZN(n18421) );
  OAI211_X1 U21475 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n18423), .A(
        n18422), .B(n18421), .ZN(P3_U2852) );
  NAND2_X1 U21476 ( .A1(n18522), .A2(n18424), .ZN(n18429) );
  AOI21_X1 U21477 ( .B1(n9631), .B2(n18426), .A(n18425), .ZN(n18428) );
  OAI221_X1 U21478 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18430), .C1(
        n11134), .C2(n18429), .A(n18428), .ZN(P3_U2853) );
  OAI22_X1 U21479 ( .A1(n18434), .A2(n21258), .B1(n18432), .B2(n18431), .ZN(
        n18435) );
  AOI21_X1 U21480 ( .B1(n18527), .B2(n18436), .A(n18435), .ZN(n18446) );
  NAND2_X1 U21481 ( .A1(n18483), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18445) );
  OAI22_X1 U21482 ( .A1(n18438), .A2(n19023), .B1(n18493), .B2(n18437), .ZN(
        n18439) );
  NOR2_X1 U21483 ( .A1(n18495), .A2(n18439), .ZN(n18455) );
  OAI211_X1 U21484 ( .C1(n18440), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18455), .ZN(n18447) );
  OAI221_X1 U21485 ( .B1(n18520), .B2(n18515), .C1(n18520), .C2(n18447), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18444) );
  NOR3_X1 U21486 ( .A1(n18484), .A2(n18441), .A3(n18510), .ZN(n18458) );
  NAND4_X1 U21487 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n18458), .A4(n18442), .ZN(
        n18443) );
  NAND4_X1 U21488 ( .A1(n18446), .A2(n18445), .A3(n18444), .A4(n18443), .ZN(
        P3_U2854) );
  OAI221_X1 U21489 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18448), .A(n18447), .ZN(
        n18454) );
  AOI21_X1 U21490 ( .B1(n18520), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18449), .ZN(n18453) );
  AOI22_X1 U21491 ( .A1(n18525), .A2(n18451), .B1(n18527), .B2(n18450), .ZN(
        n18452) );
  OAI211_X1 U21492 ( .C1(n18466), .C2(n18454), .A(n18453), .B(n18452), .ZN(
        P3_U2855) );
  OAI21_X1 U21493 ( .B1(n18455), .B2(n18466), .A(n18511), .ZN(n18463) );
  NOR2_X1 U21494 ( .A1(n18522), .A2(n19091), .ZN(n18456) );
  AOI221_X1 U21495 ( .B1(n18458), .B2(n18457), .C1(n18463), .C2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n18456), .ZN(n18462) );
  AOI22_X1 U21496 ( .A1(n18525), .A2(n18460), .B1(n18527), .B2(n18459), .ZN(
        n18461) );
  NAND2_X1 U21497 ( .A1(n18462), .A2(n18461), .ZN(P3_U2856) );
  AOI22_X1 U21498 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18463), .B1(
        n18483), .B2(P3_REIP_REG_5__SCAN_IN), .ZN(n18470) );
  AOI22_X1 U21499 ( .A1(n18525), .A2(n18465), .B1(n18527), .B2(n18464), .ZN(
        n18469) );
  NOR3_X1 U21500 ( .A1(n18484), .A2(n18466), .A3(n18490), .ZN(n18476) );
  NAND3_X1 U21501 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18476), .A3(
        n18467), .ZN(n18468) );
  NAND3_X1 U21502 ( .A1(n18470), .A2(n18469), .A3(n18468), .ZN(P3_U2857) );
  INV_X1 U21503 ( .A(n18498), .ZN(n18474) );
  AOI211_X1 U21504 ( .C1(n18472), .C2(n18471), .A(n18495), .B(n18490), .ZN(
        n18473) );
  OAI21_X1 U21505 ( .B1(n19023), .B2(n18474), .A(n18473), .ZN(n18485) );
  AOI21_X1 U21506 ( .B1(n18515), .B2(n18485), .A(n18520), .ZN(n18481) );
  AOI22_X1 U21507 ( .A1(n18483), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18525), 
        .B2(n18475), .ZN(n18479) );
  AOI22_X1 U21508 ( .A1(n18477), .A2(n18527), .B1(n18476), .B2(n18480), .ZN(
        n18478) );
  OAI211_X1 U21509 ( .C1(n18481), .C2(n18480), .A(n18479), .B(n18478), .ZN(
        P3_U2858) );
  AOI22_X1 U21510 ( .A1(n18483), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18525), 
        .B2(n18482), .ZN(n18489) );
  AOI21_X1 U21511 ( .B1(n18484), .B2(n18490), .A(n18510), .ZN(n18486) );
  AOI22_X1 U21512 ( .A1(n18527), .A2(n18487), .B1(n18486), .B2(n18485), .ZN(
        n18488) );
  OAI211_X1 U21513 ( .C1(n18490), .C2(n18511), .A(n18489), .B(n18488), .ZN(
        P3_U2859) );
  OR2_X1 U21514 ( .A1(n19173), .A2(n18491), .ZN(n18497) );
  NAND2_X1 U21515 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18492) );
  OAI22_X1 U21516 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18493), .B1(
        n19023), .B2(n18492), .ZN(n18494) );
  NOR2_X1 U21517 ( .A1(n18495), .A2(n18494), .ZN(n18496) );
  MUX2_X1 U21518 ( .A(n18497), .B(n18496), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18500) );
  NAND2_X1 U21519 ( .A1(n18992), .A2(n18498), .ZN(n18499) );
  OAI211_X1 U21520 ( .C1(n18502), .C2(n18501), .A(n18500), .B(n18499), .ZN(
        n18504) );
  AOI22_X1 U21521 ( .A1(n18521), .A2(n18504), .B1(n18525), .B2(n18503), .ZN(
        n18507) );
  INV_X1 U21522 ( .A(n18505), .ZN(n18506) );
  OAI211_X1 U21523 ( .C1(n18511), .C2(n18508), .A(n18507), .B(n18506), .ZN(
        P3_U2860) );
  NOR2_X1 U21524 ( .A1(n18522), .A2(n19191), .ZN(n18513) );
  OR3_X1 U21525 ( .A1(n18510), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18509), .ZN(n18528) );
  AOI21_X1 U21526 ( .B1(n18511), .B2(n18528), .A(n19173), .ZN(n18512) );
  AOI211_X1 U21527 ( .C1(n18514), .C2(n18525), .A(n18513), .B(n18512), .ZN(
        n18517) );
  OAI211_X1 U21528 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19002), .A(
        n18515), .B(n19173), .ZN(n18516) );
  OAI211_X1 U21529 ( .C1(n18519), .C2(n18518), .A(n18517), .B(n18516), .ZN(
        P3_U2861) );
  AOI21_X1 U21530 ( .B1(n18521), .B2(n19002), .A(n18520), .ZN(n18530) );
  INV_X1 U21531 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19197) );
  NOR2_X1 U21532 ( .A1(n18522), .A2(n19197), .ZN(n18523) );
  AOI221_X1 U21533 ( .B1(n18527), .B2(n18526), .C1(n18525), .C2(n18524), .A(
        n18523), .ZN(n18529) );
  OAI211_X1 U21534 ( .C1(n18530), .C2(n19188), .A(n18529), .B(n18528), .ZN(
        P3_U2862) );
  OAI211_X1 U21535 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18531), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n19051)
         );
  INV_X1 U21536 ( .A(n18532), .ZN(n18591) );
  OAI21_X1 U21537 ( .B1(n18535), .B2(n18533), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18534) );
  OAI221_X1 U21538 ( .B1(n18535), .B2(n19051), .C1(n18535), .C2(n18591), .A(
        n18534), .ZN(P3_U2863) );
  INV_X1 U21539 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18541) );
  NOR2_X1 U21540 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18541), .ZN(
        n18852) );
  NOR2_X1 U21541 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19030), .ZN(
        n18726) );
  NOR2_X1 U21542 ( .A1(n18852), .A2(n18726), .ZN(n18537) );
  OAI22_X1 U21543 ( .A1(n18538), .A2(n18541), .B1(n18537), .B2(n18536), .ZN(
        P3_U2866) );
  NOR2_X1 U21544 ( .A1(n18540), .A2(n18539), .ZN(P3_U2867) );
  NOR2_X1 U21545 ( .A1(n18541), .A2(n18724), .ZN(n18930) );
  NAND2_X1 U21546 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18930), .ZN(
        n18983) );
  INV_X1 U21547 ( .A(n18983), .ZN(n18627) );
  NOR2_X1 U21548 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19032) );
  INV_X1 U21549 ( .A(n19032), .ZN(n18747) );
  NOR2_X1 U21550 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18633) );
  INV_X1 U21551 ( .A(n18633), .ZN(n18632) );
  NOR2_X1 U21552 ( .A1(n18747), .A2(n18632), .ZN(n18647) );
  CLKBUF_X1 U21553 ( .A(n18647), .Z(n18651) );
  NOR2_X1 U21554 ( .A1(n18627), .A2(n18651), .ZN(n18610) );
  OAI21_X1 U21555 ( .B1(n19010), .B2(n19160), .A(n18905), .ZN(n18748) );
  NAND2_X1 U21556 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18547) );
  NOR2_X1 U21557 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19012), .ZN(
        n18807) );
  NOR2_X1 U21558 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19010), .ZN(
        n18778) );
  NOR2_X1 U21559 ( .A1(n18807), .A2(n18778), .ZN(n18856) );
  OR2_X1 U21560 ( .A1(n18547), .A2(n18856), .ZN(n18901) );
  OAI22_X1 U21561 ( .A1(n18610), .A2(n18748), .B1(n18776), .B2(n18901), .ZN(
        n18589) );
  AND2_X1 U21562 ( .A1(n18932), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18928) );
  INV_X1 U21563 ( .A(n18807), .ZN(n18542) );
  NOR2_X2 U21564 ( .A1(n18542), .A2(n18547), .ZN(n18906) );
  AND2_X1 U21565 ( .A1(n18905), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18927) );
  INV_X1 U21566 ( .A(n19056), .ZN(n18900) );
  NOR2_X1 U21567 ( .A1(n18900), .A2(n18610), .ZN(n18584) );
  AOI22_X1 U21568 ( .A1(n18928), .A2(n18906), .B1(n18927), .B2(n18584), .ZN(
        n18549) );
  NOR2_X1 U21569 ( .A1(n18544), .A2(n18543), .ZN(n18586) );
  NAND2_X1 U21570 ( .A1(n18586), .A2(n18545), .ZN(n18936) );
  INV_X1 U21571 ( .A(n18936), .ZN(n18779) );
  NOR2_X2 U21572 ( .A1(n18546), .A2(n18776), .ZN(n18933) );
  NOR2_X1 U21573 ( .A1(n18547), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18931) );
  INV_X1 U21574 ( .A(n18931), .ZN(n18878) );
  NOR2_X2 U21575 ( .A1(n19010), .A2(n18878), .ZN(n18975) );
  AOI22_X1 U21576 ( .A1(n18651), .A2(n18779), .B1(n18933), .B2(n18975), .ZN(
        n18548) );
  OAI211_X1 U21577 ( .C1(n18550), .C2(n18589), .A(n18549), .B(n18548), .ZN(
        P3_U2868) );
  AND2_X1 U21578 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18932), .ZN(n18938) );
  AND2_X1 U21579 ( .A1(n18905), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18937) );
  AOI22_X1 U21580 ( .A1(n18938), .A2(n18975), .B1(n18937), .B2(n18584), .ZN(
        n18554) );
  NAND2_X1 U21581 ( .A1(n18586), .A2(n18551), .ZN(n18942) );
  INV_X1 U21582 ( .A(n18942), .ZN(n18552) );
  NOR2_X2 U21583 ( .A1(n18776), .A2(n14163), .ZN(n18939) );
  AOI22_X1 U21584 ( .A1(n18647), .A2(n18552), .B1(n18939), .B2(n18906), .ZN(
        n18553) );
  OAI211_X1 U21585 ( .C1(n18555), .C2(n18589), .A(n18554), .B(n18553), .ZN(
        P3_U2869) );
  AND2_X1 U21586 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18932), .ZN(n18944) );
  NOR2_X2 U21587 ( .A1(n18656), .A2(n18556), .ZN(n18943) );
  AOI22_X1 U21588 ( .A1(n18944), .A2(n18975), .B1(n18943), .B2(n18584), .ZN(
        n18559) );
  NAND2_X1 U21589 ( .A1(n18586), .A2(n18557), .ZN(n18948) );
  INV_X1 U21590 ( .A(n18948), .ZN(n18755) );
  NOR2_X2 U21591 ( .A1(n18776), .A2(n19581), .ZN(n18945) );
  AOI22_X1 U21592 ( .A1(n18647), .A2(n18755), .B1(n18945), .B2(n18906), .ZN(
        n18558) );
  OAI211_X1 U21593 ( .C1(n18560), .C2(n18589), .A(n18559), .B(n18558), .ZN(
        P3_U2870) );
  AND2_X1 U21594 ( .A1(n18932), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18950) );
  AND2_X1 U21595 ( .A1(n18905), .A2(BUF2_REG_3__SCAN_IN), .ZN(n18949) );
  AOI22_X1 U21596 ( .A1(n18950), .A2(n18906), .B1(n18949), .B2(n18584), .ZN(
        n18563) );
  NAND2_X1 U21597 ( .A1(n18586), .A2(n18561), .ZN(n18954) );
  INV_X1 U21598 ( .A(n18954), .ZN(n18787) );
  NOR2_X2 U21599 ( .A1(n15503), .A2(n18776), .ZN(n18951) );
  AOI22_X1 U21600 ( .A1(n18647), .A2(n18787), .B1(n18951), .B2(n18975), .ZN(
        n18562) );
  OAI211_X1 U21601 ( .C1(n18564), .C2(n18589), .A(n18563), .B(n18562), .ZN(
        P3_U2871) );
  NOR2_X2 U21602 ( .A1(n18776), .A2(n18565), .ZN(n18956) );
  NOR2_X2 U21603 ( .A1(n18656), .A2(n18566), .ZN(n18955) );
  AOI22_X1 U21604 ( .A1(n18956), .A2(n18906), .B1(n18955), .B2(n18584), .ZN(
        n18570) );
  NAND2_X1 U21605 ( .A1(n18586), .A2(n18567), .ZN(n18960) );
  INV_X1 U21606 ( .A(n18960), .ZN(n18568) );
  AND2_X1 U21607 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18932), .ZN(n18957) );
  AOI22_X1 U21608 ( .A1(n18651), .A2(n18568), .B1(n18957), .B2(n18975), .ZN(
        n18569) );
  OAI211_X1 U21609 ( .C1(n18571), .C2(n18589), .A(n18570), .B(n18569), .ZN(
        P3_U2872) );
  NOR2_X2 U21610 ( .A1(n18776), .A2(n19594), .ZN(n18962) );
  NOR2_X2 U21611 ( .A1(n18656), .A2(n18572), .ZN(n18961) );
  AOI22_X1 U21612 ( .A1(n18962), .A2(n18906), .B1(n18961), .B2(n18584), .ZN(
        n18575) );
  NAND2_X1 U21613 ( .A1(n18586), .A2(n18573), .ZN(n18966) );
  INV_X1 U21614 ( .A(n18966), .ZN(n18793) );
  AND2_X1 U21615 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18932), .ZN(n18963) );
  AOI22_X1 U21616 ( .A1(n18651), .A2(n18793), .B1(n18963), .B2(n18975), .ZN(
        n18574) );
  OAI211_X1 U21617 ( .C1(n18576), .C2(n18589), .A(n18575), .B(n18574), .ZN(
        P3_U2873) );
  NOR2_X2 U21618 ( .A1(n19602), .A2(n18776), .ZN(n18969) );
  NOR2_X2 U21619 ( .A1(n18656), .A2(n18577), .ZN(n18967) );
  AOI22_X1 U21620 ( .A1(n18969), .A2(n18975), .B1(n18967), .B2(n18584), .ZN(
        n18581) );
  NAND2_X1 U21621 ( .A1(n18586), .A2(n18578), .ZN(n18972) );
  INV_X1 U21622 ( .A(n18972), .ZN(n18579) );
  NOR2_X2 U21623 ( .A1(n18776), .A2(n15542), .ZN(n18968) );
  AOI22_X1 U21624 ( .A1(n18651), .A2(n18579), .B1(n18968), .B2(n18906), .ZN(
        n18580) );
  OAI211_X1 U21625 ( .C1(n18582), .C2(n18589), .A(n18581), .B(n18580), .ZN(
        P3_U2874) );
  NOR2_X2 U21626 ( .A1(n18656), .A2(n18583), .ZN(n18974) );
  NOR2_X2 U21627 ( .A1(n18776), .A2(n19610), .ZN(n18978) );
  AOI22_X1 U21628 ( .A1(n18974), .A2(n18584), .B1(n18978), .B2(n18975), .ZN(
        n18588) );
  NAND2_X1 U21629 ( .A1(n18586), .A2(n18585), .ZN(n18982) );
  INV_X1 U21630 ( .A(n18982), .ZN(n18802) );
  AND2_X1 U21631 ( .A1(n18932), .A2(BUF2_REG_23__SCAN_IN), .ZN(n18976) );
  AOI22_X1 U21632 ( .A1(n18651), .A2(n18802), .B1(n18976), .B2(n18906), .ZN(
        n18587) );
  OAI211_X1 U21633 ( .C1(n18590), .C2(n18589), .A(n18588), .B(n18587), .ZN(
        P3_U2875) );
  NAND2_X1 U21634 ( .A1(n18633), .A2(n18778), .ZN(n18634) );
  NAND2_X1 U21635 ( .A1(n19012), .A2(n19056), .ZN(n18777) );
  NOR2_X1 U21636 ( .A1(n18632), .A2(n18777), .ZN(n18606) );
  AOI22_X1 U21637 ( .A1(n18627), .A2(n18928), .B1(n18927), .B2(n18606), .ZN(
        n18593) );
  NAND2_X1 U21638 ( .A1(n18905), .A2(n18591), .ZN(n18832) );
  NOR2_X1 U21639 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18832), .ZN(
        n18680) );
  AOI22_X1 U21640 ( .A1(n18932), .A2(n18930), .B1(n18633), .B2(n18680), .ZN(
        n18607) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18607), .B1(
        n18933), .B2(n18906), .ZN(n18592) );
  OAI211_X1 U21642 ( .C1(n18634), .C2(n18936), .A(n18593), .B(n18592), .ZN(
        P3_U2876) );
  AOI22_X1 U21643 ( .A1(n18938), .A2(n18906), .B1(n18937), .B2(n18606), .ZN(
        n18595) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18607), .B1(
        n18627), .B2(n18939), .ZN(n18594) );
  OAI211_X1 U21645 ( .C1(n18634), .C2(n18942), .A(n18595), .B(n18594), .ZN(
        P3_U2877) );
  AOI22_X1 U21646 ( .A1(n18944), .A2(n18906), .B1(n18943), .B2(n18606), .ZN(
        n18597) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18607), .B1(
        n18627), .B2(n18945), .ZN(n18596) );
  OAI211_X1 U21648 ( .C1(n18634), .C2(n18948), .A(n18597), .B(n18596), .ZN(
        P3_U2878) );
  AOI22_X1 U21649 ( .A1(n18951), .A2(n18906), .B1(n18949), .B2(n18606), .ZN(
        n18599) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18607), .B1(
        n18627), .B2(n18950), .ZN(n18598) );
  OAI211_X1 U21651 ( .C1(n18634), .C2(n18954), .A(n18599), .B(n18598), .ZN(
        P3_U2879) );
  AOI22_X1 U21652 ( .A1(n18957), .A2(n18906), .B1(n18955), .B2(n18606), .ZN(
        n18601) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18607), .B1(
        n18627), .B2(n18956), .ZN(n18600) );
  OAI211_X1 U21654 ( .C1(n18634), .C2(n18960), .A(n18601), .B(n18600), .ZN(
        P3_U2880) );
  AOI22_X1 U21655 ( .A1(n18963), .A2(n18906), .B1(n18961), .B2(n18606), .ZN(
        n18603) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18607), .B1(
        n18627), .B2(n18962), .ZN(n18602) );
  OAI211_X1 U21657 ( .C1(n18634), .C2(n18966), .A(n18603), .B(n18602), .ZN(
        P3_U2881) );
  AOI22_X1 U21658 ( .A1(n18627), .A2(n18968), .B1(n18967), .B2(n18606), .ZN(
        n18605) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18607), .B1(
        n18969), .B2(n18906), .ZN(n18604) );
  OAI211_X1 U21660 ( .C1(n18634), .C2(n18972), .A(n18605), .B(n18604), .ZN(
        P3_U2882) );
  AOI22_X1 U21661 ( .A1(n18627), .A2(n18976), .B1(n18974), .B2(n18606), .ZN(
        n18609) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18607), .B1(
        n18978), .B2(n18906), .ZN(n18608) );
  OAI211_X1 U21663 ( .C1(n18634), .C2(n18982), .A(n18609), .B(n18608), .ZN(
        P3_U2883) );
  NAND2_X1 U21664 ( .A1(n18807), .A2(n18633), .ZN(n18631) );
  AOI21_X1 U21665 ( .B1(n18631), .B2(n18634), .A(n18900), .ZN(n18626) );
  AOI22_X1 U21666 ( .A1(n18651), .A2(n18928), .B1(n18927), .B2(n18626), .ZN(
        n18613) );
  INV_X1 U21667 ( .A(n18631), .ZN(n18697) );
  AOI221_X1 U21668 ( .B1(n18610), .B2(n18634), .C1(n18902), .C2(n18634), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18611) );
  OAI21_X1 U21669 ( .B1(n18697), .B2(n18611), .A(n18905), .ZN(n18628) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18628), .B1(
        n18627), .B2(n18933), .ZN(n18612) );
  OAI211_X1 U21671 ( .C1(n18631), .C2(n18936), .A(n18613), .B(n18612), .ZN(
        P3_U2884) );
  AOI22_X1 U21672 ( .A1(n18651), .A2(n18939), .B1(n18626), .B2(n18937), .ZN(
        n18615) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18628), .B1(
        n18627), .B2(n18938), .ZN(n18614) );
  OAI211_X1 U21674 ( .C1(n18631), .C2(n18942), .A(n18615), .B(n18614), .ZN(
        P3_U2885) );
  AOI22_X1 U21675 ( .A1(n18651), .A2(n18945), .B1(n18626), .B2(n18943), .ZN(
        n18617) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18628), .B1(
        n18627), .B2(n18944), .ZN(n18616) );
  OAI211_X1 U21677 ( .C1(n18631), .C2(n18948), .A(n18617), .B(n18616), .ZN(
        P3_U2886) );
  AOI22_X1 U21678 ( .A1(n18651), .A2(n18950), .B1(n18626), .B2(n18949), .ZN(
        n18619) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18628), .B1(
        n18627), .B2(n18951), .ZN(n18618) );
  OAI211_X1 U21680 ( .C1(n18631), .C2(n18954), .A(n18619), .B(n18618), .ZN(
        P3_U2887) );
  AOI22_X1 U21681 ( .A1(n18651), .A2(n18956), .B1(n18626), .B2(n18955), .ZN(
        n18621) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18628), .B1(
        n18627), .B2(n18957), .ZN(n18620) );
  OAI211_X1 U21683 ( .C1(n18631), .C2(n18960), .A(n18621), .B(n18620), .ZN(
        P3_U2888) );
  AOI22_X1 U21684 ( .A1(n18627), .A2(n18963), .B1(n18626), .B2(n18961), .ZN(
        n18623) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18628), .B1(
        n18647), .B2(n18962), .ZN(n18622) );
  OAI211_X1 U21686 ( .C1(n18631), .C2(n18966), .A(n18623), .B(n18622), .ZN(
        P3_U2889) );
  AOI22_X1 U21687 ( .A1(n18651), .A2(n18968), .B1(n18626), .B2(n18967), .ZN(
        n18625) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18628), .B1(
        n18627), .B2(n18969), .ZN(n18624) );
  OAI211_X1 U21689 ( .C1(n18631), .C2(n18972), .A(n18625), .B(n18624), .ZN(
        P3_U2890) );
  AOI22_X1 U21690 ( .A1(n18627), .A2(n18978), .B1(n18626), .B2(n18974), .ZN(
        n18630) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18628), .B1(
        n18651), .B2(n18976), .ZN(n18629) );
  OAI211_X1 U21692 ( .C1(n18631), .C2(n18982), .A(n18630), .B(n18629), .ZN(
        P3_U2891) );
  NOR2_X1 U21693 ( .A1(n19012), .A2(n18632), .ZN(n18681) );
  NAND2_X1 U21694 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18681), .ZN(
        n18655) );
  INV_X1 U21695 ( .A(n18655), .ZN(n18718) );
  AOI21_X1 U21696 ( .B1(n19012), .B2(n18902), .A(n18656), .ZN(n18725) );
  OAI211_X1 U21697 ( .C1(n18718), .C2(n19160), .A(n18633), .B(n18725), .ZN(
        n18652) );
  AND2_X1 U21698 ( .A1(n19056), .A2(n18681), .ZN(n18650) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18652), .B1(
        n18927), .B2(n18650), .ZN(n18636) );
  INV_X1 U21700 ( .A(n18634), .ZN(n18674) );
  AOI22_X1 U21701 ( .A1(n18674), .A2(n18928), .B1(n18651), .B2(n18933), .ZN(
        n18635) );
  OAI211_X1 U21702 ( .C1(n18936), .C2(n18655), .A(n18636), .B(n18635), .ZN(
        P3_U2892) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18652), .B1(
        n18937), .B2(n18650), .ZN(n18638) );
  AOI22_X1 U21704 ( .A1(n18674), .A2(n18939), .B1(n18647), .B2(n18938), .ZN(
        n18637) );
  OAI211_X1 U21705 ( .C1(n18942), .C2(n18655), .A(n18638), .B(n18637), .ZN(
        P3_U2893) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18652), .B1(
        n18943), .B2(n18650), .ZN(n18640) );
  AOI22_X1 U21707 ( .A1(n18674), .A2(n18945), .B1(n18647), .B2(n18944), .ZN(
        n18639) );
  OAI211_X1 U21708 ( .C1(n18948), .C2(n18655), .A(n18640), .B(n18639), .ZN(
        P3_U2894) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18652), .B1(
        n18949), .B2(n18650), .ZN(n18642) );
  AOI22_X1 U21710 ( .A1(n18674), .A2(n18950), .B1(n18647), .B2(n18951), .ZN(
        n18641) );
  OAI211_X1 U21711 ( .C1(n18954), .C2(n18655), .A(n18642), .B(n18641), .ZN(
        P3_U2895) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18652), .B1(
        n18955), .B2(n18650), .ZN(n18644) );
  AOI22_X1 U21713 ( .A1(n18674), .A2(n18956), .B1(n18647), .B2(n18957), .ZN(
        n18643) );
  OAI211_X1 U21714 ( .C1(n18960), .C2(n18655), .A(n18644), .B(n18643), .ZN(
        P3_U2896) );
  AOI22_X1 U21715 ( .A1(n18674), .A2(n18962), .B1(n18961), .B2(n18650), .ZN(
        n18646) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18652), .B1(
        n18651), .B2(n18963), .ZN(n18645) );
  OAI211_X1 U21717 ( .C1(n18966), .C2(n18655), .A(n18646), .B(n18645), .ZN(
        P3_U2897) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18652), .B1(
        n18967), .B2(n18650), .ZN(n18649) );
  AOI22_X1 U21719 ( .A1(n18674), .A2(n18968), .B1(n18647), .B2(n18969), .ZN(
        n18648) );
  OAI211_X1 U21720 ( .C1(n18972), .C2(n18655), .A(n18649), .B(n18648), .ZN(
        P3_U2898) );
  AOI22_X1 U21721 ( .A1(n18674), .A2(n18976), .B1(n18974), .B2(n18650), .ZN(
        n18654) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18652), .B1(
        n18651), .B2(n18978), .ZN(n18653) );
  OAI211_X1 U21723 ( .C1(n18982), .C2(n18655), .A(n18654), .B(n18653), .ZN(
        P3_U2899) );
  NAND2_X1 U21724 ( .A1(n19032), .A2(n18726), .ZN(n18678) );
  INV_X1 U21725 ( .A(n18678), .ZN(n18742) );
  NOR2_X1 U21726 ( .A1(n18718), .A2(n18742), .ZN(n18702) );
  NOR2_X1 U21727 ( .A1(n18900), .A2(n18702), .ZN(n18673) );
  AOI22_X1 U21728 ( .A1(n18697), .A2(n18928), .B1(n18927), .B2(n18673), .ZN(
        n18660) );
  NOR2_X1 U21729 ( .A1(n18697), .A2(n18674), .ZN(n18657) );
  OAI22_X1 U21730 ( .A1(n18657), .A2(n18776), .B1(n18702), .B2(n18656), .ZN(
        n18658) );
  OAI21_X1 U21731 ( .B1(n18742), .B2(n19160), .A(n18658), .ZN(n18675) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18675), .B1(
        n18674), .B2(n18933), .ZN(n18659) );
  OAI211_X1 U21733 ( .C1(n18936), .C2(n18678), .A(n18660), .B(n18659), .ZN(
        P3_U2900) );
  AOI22_X1 U21734 ( .A1(n18697), .A2(n18939), .B1(n18937), .B2(n18673), .ZN(
        n18662) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18675), .B1(
        n18674), .B2(n18938), .ZN(n18661) );
  OAI211_X1 U21736 ( .C1(n18942), .C2(n18678), .A(n18662), .B(n18661), .ZN(
        P3_U2901) );
  AOI22_X1 U21737 ( .A1(n18674), .A2(n18944), .B1(n18943), .B2(n18673), .ZN(
        n18664) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18675), .B1(
        n18697), .B2(n18945), .ZN(n18663) );
  OAI211_X1 U21739 ( .C1(n18948), .C2(n18678), .A(n18664), .B(n18663), .ZN(
        P3_U2902) );
  AOI22_X1 U21740 ( .A1(n18697), .A2(n18950), .B1(n18949), .B2(n18673), .ZN(
        n18666) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18675), .B1(
        n18674), .B2(n18951), .ZN(n18665) );
  OAI211_X1 U21742 ( .C1(n18954), .C2(n18678), .A(n18666), .B(n18665), .ZN(
        P3_U2903) );
  AOI22_X1 U21743 ( .A1(n18697), .A2(n18956), .B1(n18955), .B2(n18673), .ZN(
        n18668) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18675), .B1(
        n18674), .B2(n18957), .ZN(n18667) );
  OAI211_X1 U21745 ( .C1(n18960), .C2(n18678), .A(n18668), .B(n18667), .ZN(
        P3_U2904) );
  AOI22_X1 U21746 ( .A1(n18697), .A2(n18962), .B1(n18961), .B2(n18673), .ZN(
        n18670) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18675), .B1(
        n18674), .B2(n18963), .ZN(n18669) );
  OAI211_X1 U21748 ( .C1(n18966), .C2(n18678), .A(n18670), .B(n18669), .ZN(
        P3_U2905) );
  AOI22_X1 U21749 ( .A1(n18697), .A2(n18968), .B1(n18967), .B2(n18673), .ZN(
        n18672) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18675), .B1(
        n18674), .B2(n18969), .ZN(n18671) );
  OAI211_X1 U21751 ( .C1(n18972), .C2(n18678), .A(n18672), .B(n18671), .ZN(
        P3_U2906) );
  AOI22_X1 U21752 ( .A1(n18674), .A2(n18978), .B1(n18974), .B2(n18673), .ZN(
        n18677) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18675), .B1(
        n18697), .B2(n18976), .ZN(n18676) );
  OAI211_X1 U21754 ( .C1(n18982), .C2(n18678), .A(n18677), .B(n18676), .ZN(
        P3_U2907) );
  NAND2_X1 U21755 ( .A1(n18778), .A2(n18726), .ZN(n18701) );
  INV_X1 U21756 ( .A(n18726), .ZN(n18679) );
  NOR2_X1 U21757 ( .A1(n18679), .A2(n18777), .ZN(n18696) );
  AOI22_X1 U21758 ( .A1(n18697), .A2(n18933), .B1(n18927), .B2(n18696), .ZN(
        n18683) );
  AOI22_X1 U21759 ( .A1(n18932), .A2(n18681), .B1(n18726), .B2(n18680), .ZN(
        n18698) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18698), .B1(
        n18928), .B2(n18718), .ZN(n18682) );
  OAI211_X1 U21761 ( .C1(n18936), .C2(n18701), .A(n18683), .B(n18682), .ZN(
        P3_U2908) );
  AOI22_X1 U21762 ( .A1(n18937), .A2(n18696), .B1(n18939), .B2(n18718), .ZN(
        n18685) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18698), .B1(
        n18697), .B2(n18938), .ZN(n18684) );
  OAI211_X1 U21764 ( .C1(n18942), .C2(n18701), .A(n18685), .B(n18684), .ZN(
        P3_U2909) );
  AOI22_X1 U21765 ( .A1(n18945), .A2(n18718), .B1(n18943), .B2(n18696), .ZN(
        n18687) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18698), .B1(
        n18697), .B2(n18944), .ZN(n18686) );
  OAI211_X1 U21767 ( .C1(n18948), .C2(n18701), .A(n18687), .B(n18686), .ZN(
        P3_U2910) );
  AOI22_X1 U21768 ( .A1(n18697), .A2(n18951), .B1(n18949), .B2(n18696), .ZN(
        n18689) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18698), .B1(
        n18950), .B2(n18718), .ZN(n18688) );
  OAI211_X1 U21770 ( .C1(n18954), .C2(n18701), .A(n18689), .B(n18688), .ZN(
        P3_U2911) );
  AOI22_X1 U21771 ( .A1(n18956), .A2(n18718), .B1(n18955), .B2(n18696), .ZN(
        n18691) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18698), .B1(
        n18697), .B2(n18957), .ZN(n18690) );
  OAI211_X1 U21773 ( .C1(n18960), .C2(n18701), .A(n18691), .B(n18690), .ZN(
        P3_U2912) );
  AOI22_X1 U21774 ( .A1(n18962), .A2(n18718), .B1(n18961), .B2(n18696), .ZN(
        n18693) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18698), .B1(
        n18697), .B2(n18963), .ZN(n18692) );
  OAI211_X1 U21776 ( .C1(n18966), .C2(n18701), .A(n18693), .B(n18692), .ZN(
        P3_U2913) );
  AOI22_X1 U21777 ( .A1(n18697), .A2(n18969), .B1(n18967), .B2(n18696), .ZN(
        n18695) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18698), .B1(
        n18968), .B2(n18718), .ZN(n18694) );
  OAI211_X1 U21779 ( .C1(n18972), .C2(n18701), .A(n18695), .B(n18694), .ZN(
        P3_U2914) );
  AOI22_X1 U21780 ( .A1(n18976), .A2(n18718), .B1(n18974), .B2(n18696), .ZN(
        n18700) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18698), .B1(
        n18697), .B2(n18978), .ZN(n18699) );
  OAI211_X1 U21782 ( .C1(n18982), .C2(n18701), .A(n18700), .B(n18699), .ZN(
        P3_U2915) );
  NAND2_X1 U21783 ( .A1(n18807), .A2(n18726), .ZN(n18723) );
  INV_X1 U21784 ( .A(n18701), .ZN(n18770) );
  INV_X1 U21785 ( .A(n18723), .ZN(n18800) );
  NOR2_X1 U21786 ( .A1(n18770), .A2(n18800), .ZN(n18749) );
  NOR2_X1 U21787 ( .A1(n18900), .A2(n18749), .ZN(n18719) );
  AOI22_X1 U21788 ( .A1(n18928), .A2(n18742), .B1(n18927), .B2(n18719), .ZN(
        n18705) );
  OAI21_X1 U21789 ( .B1(n18702), .B2(n18902), .A(n18749), .ZN(n18703) );
  OAI211_X1 U21790 ( .C1(n18800), .C2(n19160), .A(n18905), .B(n18703), .ZN(
        n18720) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18720), .B1(
        n18933), .B2(n18718), .ZN(n18704) );
  OAI211_X1 U21792 ( .C1(n18936), .C2(n18723), .A(n18705), .B(n18704), .ZN(
        P3_U2916) );
  AOI22_X1 U21793 ( .A1(n18938), .A2(n18718), .B1(n18937), .B2(n18719), .ZN(
        n18707) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18720), .B1(
        n18939), .B2(n18742), .ZN(n18706) );
  OAI211_X1 U21795 ( .C1(n18942), .C2(n18723), .A(n18707), .B(n18706), .ZN(
        P3_U2917) );
  AOI22_X1 U21796 ( .A1(n18944), .A2(n18718), .B1(n18943), .B2(n18719), .ZN(
        n18709) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18720), .B1(
        n18945), .B2(n18742), .ZN(n18708) );
  OAI211_X1 U21798 ( .C1(n18948), .C2(n18723), .A(n18709), .B(n18708), .ZN(
        P3_U2918) );
  AOI22_X1 U21799 ( .A1(n18950), .A2(n18742), .B1(n18949), .B2(n18719), .ZN(
        n18711) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18720), .B1(
        n18951), .B2(n18718), .ZN(n18710) );
  OAI211_X1 U21801 ( .C1(n18954), .C2(n18723), .A(n18711), .B(n18710), .ZN(
        P3_U2919) );
  AOI22_X1 U21802 ( .A1(n18956), .A2(n18742), .B1(n18955), .B2(n18719), .ZN(
        n18713) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18720), .B1(
        n18957), .B2(n18718), .ZN(n18712) );
  OAI211_X1 U21804 ( .C1(n18960), .C2(n18723), .A(n18713), .B(n18712), .ZN(
        P3_U2920) );
  AOI22_X1 U21805 ( .A1(n18963), .A2(n18718), .B1(n18961), .B2(n18719), .ZN(
        n18715) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18720), .B1(
        n18962), .B2(n18742), .ZN(n18714) );
  OAI211_X1 U21807 ( .C1(n18966), .C2(n18723), .A(n18715), .B(n18714), .ZN(
        P3_U2921) );
  AOI22_X1 U21808 ( .A1(n18968), .A2(n18742), .B1(n18967), .B2(n18719), .ZN(
        n18717) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18720), .B1(
        n18969), .B2(n18718), .ZN(n18716) );
  OAI211_X1 U21810 ( .C1(n18972), .C2(n18723), .A(n18717), .B(n18716), .ZN(
        P3_U2922) );
  AOI22_X1 U21811 ( .A1(n18974), .A2(n18719), .B1(n18978), .B2(n18718), .ZN(
        n18722) );
  AOI22_X1 U21812 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18720), .B1(
        n18976), .B2(n18742), .ZN(n18721) );
  OAI211_X1 U21813 ( .C1(n18982), .C2(n18723), .A(n18722), .B(n18721), .ZN(
        P3_U2923) );
  OR2_X1 U21814 ( .A1(n18724), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18775) );
  NOR2_X2 U21815 ( .A1(n19010), .A2(n18775), .ZN(n18826) );
  INV_X1 U21816 ( .A(n18826), .ZN(n18746) );
  NOR2_X1 U21817 ( .A1(n18900), .A2(n18775), .ZN(n18741) );
  AOI22_X1 U21818 ( .A1(n18933), .A2(n18742), .B1(n18927), .B2(n18741), .ZN(
        n18728) );
  OAI211_X1 U21819 ( .C1(n18826), .C2(n19160), .A(n18726), .B(n18725), .ZN(
        n18743) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18743), .B1(
        n18928), .B2(n18770), .ZN(n18727) );
  OAI211_X1 U21821 ( .C1(n18936), .C2(n18746), .A(n18728), .B(n18727), .ZN(
        P3_U2924) );
  AOI22_X1 U21822 ( .A1(n18937), .A2(n18741), .B1(n18939), .B2(n18770), .ZN(
        n18730) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18743), .B1(
        n18938), .B2(n18742), .ZN(n18729) );
  OAI211_X1 U21824 ( .C1(n18942), .C2(n18746), .A(n18730), .B(n18729), .ZN(
        P3_U2925) );
  AOI22_X1 U21825 ( .A1(n18944), .A2(n18742), .B1(n18943), .B2(n18741), .ZN(
        n18732) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18743), .B1(
        n18945), .B2(n18770), .ZN(n18731) );
  OAI211_X1 U21827 ( .C1(n18948), .C2(n18746), .A(n18732), .B(n18731), .ZN(
        P3_U2926) );
  AOI22_X1 U21828 ( .A1(n18950), .A2(n18770), .B1(n18949), .B2(n18741), .ZN(
        n18734) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18743), .B1(
        n18951), .B2(n18742), .ZN(n18733) );
  OAI211_X1 U21830 ( .C1(n18954), .C2(n18746), .A(n18734), .B(n18733), .ZN(
        P3_U2927) );
  AOI22_X1 U21831 ( .A1(n18956), .A2(n18770), .B1(n18955), .B2(n18741), .ZN(
        n18736) );
  AOI22_X1 U21832 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18743), .B1(
        n18957), .B2(n18742), .ZN(n18735) );
  OAI211_X1 U21833 ( .C1(n18960), .C2(n18746), .A(n18736), .B(n18735), .ZN(
        P3_U2928) );
  AOI22_X1 U21834 ( .A1(n18962), .A2(n18770), .B1(n18961), .B2(n18741), .ZN(
        n18738) );
  AOI22_X1 U21835 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18743), .B1(
        n18963), .B2(n18742), .ZN(n18737) );
  OAI211_X1 U21836 ( .C1(n18966), .C2(n18746), .A(n18738), .B(n18737), .ZN(
        P3_U2929) );
  AOI22_X1 U21837 ( .A1(n18968), .A2(n18770), .B1(n18967), .B2(n18741), .ZN(
        n18740) );
  AOI22_X1 U21838 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18743), .B1(
        n18969), .B2(n18742), .ZN(n18739) );
  OAI211_X1 U21839 ( .C1(n18972), .C2(n18746), .A(n18740), .B(n18739), .ZN(
        P3_U2930) );
  AOI22_X1 U21840 ( .A1(n18976), .A2(n18770), .B1(n18974), .B2(n18741), .ZN(
        n18745) );
  AOI22_X1 U21841 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18743), .B1(
        n18978), .B2(n18742), .ZN(n18744) );
  OAI211_X1 U21842 ( .C1(n18982), .C2(n18746), .A(n18745), .B(n18744), .ZN(
        P3_U2931) );
  INV_X1 U21843 ( .A(n18852), .ZN(n18831) );
  NOR2_X2 U21844 ( .A1(n18747), .A2(n18831), .ZN(n18848) );
  NOR2_X1 U21845 ( .A1(n18848), .A2(n18826), .ZN(n18809) );
  AOI221_X1 U21846 ( .B1(n18749), .B2(n18809), .C1(n18902), .C2(n18809), .A(
        n18748), .ZN(n18761) );
  NOR2_X1 U21847 ( .A1(n18900), .A2(n18809), .ZN(n18768) );
  AOI22_X1 U21848 ( .A1(n18933), .A2(n18770), .B1(n18927), .B2(n18768), .ZN(
        n18751) );
  AOI22_X1 U21849 ( .A1(n18779), .A2(n18848), .B1(n18928), .B2(n18800), .ZN(
        n18750) );
  OAI211_X1 U21850 ( .C1(n18761), .C2(n18752), .A(n18751), .B(n18750), .ZN(
        P3_U2932) );
  INV_X1 U21851 ( .A(n18848), .ZN(n18773) );
  AOI22_X1 U21852 ( .A1(n18938), .A2(n18770), .B1(n18937), .B2(n18768), .ZN(
        n18754) );
  INV_X1 U21853 ( .A(n18761), .ZN(n18769) );
  AOI22_X1 U21854 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18769), .B1(
        n18939), .B2(n18800), .ZN(n18753) );
  OAI211_X1 U21855 ( .C1(n18942), .C2(n18773), .A(n18754), .B(n18753), .ZN(
        P3_U2933) );
  AOI22_X1 U21856 ( .A1(n18944), .A2(n18770), .B1(n18943), .B2(n18768), .ZN(
        n18757) );
  AOI22_X1 U21857 ( .A1(n18755), .A2(n18848), .B1(n18945), .B2(n18800), .ZN(
        n18756) );
  OAI211_X1 U21858 ( .C1(n18761), .C2(n11051), .A(n18757), .B(n18756), .ZN(
        P3_U2934) );
  AOI22_X1 U21859 ( .A1(n18950), .A2(n18800), .B1(n18949), .B2(n18768), .ZN(
        n18759) );
  AOI22_X1 U21860 ( .A1(n18951), .A2(n18770), .B1(n18787), .B2(n18848), .ZN(
        n18758) );
  OAI211_X1 U21861 ( .C1(n18761), .C2(n18760), .A(n18759), .B(n18758), .ZN(
        P3_U2935) );
  AOI22_X1 U21862 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18769), .B1(
        n18955), .B2(n18768), .ZN(n18763) );
  AOI22_X1 U21863 ( .A1(n18957), .A2(n18770), .B1(n18956), .B2(n18800), .ZN(
        n18762) );
  OAI211_X1 U21864 ( .C1(n18960), .C2(n18773), .A(n18763), .B(n18762), .ZN(
        P3_U2936) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18769), .B1(
        n18961), .B2(n18768), .ZN(n18765) );
  AOI22_X1 U21866 ( .A1(n18962), .A2(n18800), .B1(n18963), .B2(n18770), .ZN(
        n18764) );
  OAI211_X1 U21867 ( .C1(n18966), .C2(n18773), .A(n18765), .B(n18764), .ZN(
        P3_U2937) );
  AOI22_X1 U21868 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18769), .B1(
        n18967), .B2(n18768), .ZN(n18767) );
  AOI22_X1 U21869 ( .A1(n18969), .A2(n18770), .B1(n18968), .B2(n18800), .ZN(
        n18766) );
  OAI211_X1 U21870 ( .C1(n18972), .C2(n18773), .A(n18767), .B(n18766), .ZN(
        P3_U2938) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18769), .B1(
        n18974), .B2(n18768), .ZN(n18772) );
  AOI22_X1 U21872 ( .A1(n18976), .A2(n18800), .B1(n18978), .B2(n18770), .ZN(
        n18771) );
  OAI211_X1 U21873 ( .C1(n18982), .C2(n18773), .A(n18772), .B(n18771), .ZN(
        P3_U2939) );
  NAND2_X1 U21874 ( .A1(n18852), .A2(n19012), .ZN(n18774) );
  OAI22_X1 U21875 ( .A1(n18776), .A2(n18775), .B1(n18832), .B2(n18774), .ZN(
        n18805) );
  NOR2_X1 U21876 ( .A1(n18831), .A2(n18777), .ZN(n18801) );
  AOI22_X1 U21877 ( .A1(n18933), .A2(n18800), .B1(n18927), .B2(n18801), .ZN(
        n18781) );
  NAND2_X1 U21878 ( .A1(n18778), .A2(n18852), .ZN(n18808) );
  INV_X1 U21879 ( .A(n18808), .ZN(n18874) );
  AOI22_X1 U21880 ( .A1(n18779), .A2(n18874), .B1(n18928), .B2(n18826), .ZN(
        n18780) );
  OAI211_X1 U21881 ( .C1(n18782), .C2(n18805), .A(n18781), .B(n18780), .ZN(
        P3_U2940) );
  AOI22_X1 U21882 ( .A1(n18938), .A2(n18800), .B1(n18937), .B2(n18801), .ZN(
        n18784) );
  INV_X1 U21883 ( .A(n18805), .ZN(n18797) );
  AOI22_X1 U21884 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18797), .B1(
        n18939), .B2(n18826), .ZN(n18783) );
  OAI211_X1 U21885 ( .C1(n18942), .C2(n18808), .A(n18784), .B(n18783), .ZN(
        P3_U2941) );
  AOI22_X1 U21886 ( .A1(n18945), .A2(n18826), .B1(n18943), .B2(n18801), .ZN(
        n18786) );
  AOI22_X1 U21887 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18797), .B1(
        n18944), .B2(n18800), .ZN(n18785) );
  OAI211_X1 U21888 ( .C1(n18948), .C2(n18808), .A(n18786), .B(n18785), .ZN(
        P3_U2942) );
  AOI22_X1 U21889 ( .A1(n18951), .A2(n18800), .B1(n18949), .B2(n18801), .ZN(
        n18789) );
  AOI22_X1 U21890 ( .A1(n18787), .A2(n18874), .B1(n18950), .B2(n18826), .ZN(
        n18788) );
  OAI211_X1 U21891 ( .C1(n18790), .C2(n18805), .A(n18789), .B(n18788), .ZN(
        P3_U2943) );
  AOI22_X1 U21892 ( .A1(n18957), .A2(n18800), .B1(n18955), .B2(n18801), .ZN(
        n18792) );
  AOI22_X1 U21893 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18797), .B1(
        n18956), .B2(n18826), .ZN(n18791) );
  OAI211_X1 U21894 ( .C1(n18960), .C2(n18808), .A(n18792), .B(n18791), .ZN(
        P3_U2944) );
  AOI22_X1 U21895 ( .A1(n18963), .A2(n18800), .B1(n18961), .B2(n18801), .ZN(
        n18795) );
  AOI22_X1 U21896 ( .A1(n18962), .A2(n18826), .B1(n18793), .B2(n18874), .ZN(
        n18794) );
  OAI211_X1 U21897 ( .C1(n18796), .C2(n18805), .A(n18795), .B(n18794), .ZN(
        P3_U2945) );
  AOI22_X1 U21898 ( .A1(n18968), .A2(n18826), .B1(n18967), .B2(n18801), .ZN(
        n18799) );
  AOI22_X1 U21899 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18797), .B1(
        n18969), .B2(n18800), .ZN(n18798) );
  OAI211_X1 U21900 ( .C1(n18972), .C2(n18808), .A(n18799), .B(n18798), .ZN(
        P3_U2946) );
  AOI22_X1 U21901 ( .A1(n18974), .A2(n18801), .B1(n18978), .B2(n18800), .ZN(
        n18804) );
  AOI22_X1 U21902 ( .A1(n18976), .A2(n18826), .B1(n18802), .B2(n18874), .ZN(
        n18803) );
  OAI211_X1 U21903 ( .C1(n18806), .C2(n18805), .A(n18804), .B(n18803), .ZN(
        P3_U2947) );
  NAND2_X1 U21904 ( .A1(n18807), .A2(n18852), .ZN(n18830) );
  AOI22_X1 U21905 ( .A1(n18933), .A2(n18826), .B1(n18927), .B2(n18825), .ZN(
        n18812) );
  INV_X1 U21906 ( .A(n18830), .ZN(n18895) );
  AOI221_X1 U21907 ( .B1(n18809), .B2(n18808), .C1(n18902), .C2(n18808), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18810) );
  OAI21_X1 U21908 ( .B1(n18895), .B2(n18810), .A(n18905), .ZN(n18827) );
  AOI22_X1 U21909 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18827), .B1(
        n18928), .B2(n18848), .ZN(n18811) );
  OAI211_X1 U21910 ( .C1(n18936), .C2(n18830), .A(n18812), .B(n18811), .ZN(
        P3_U2948) );
  AOI22_X1 U21911 ( .A1(n18938), .A2(n18826), .B1(n18937), .B2(n18825), .ZN(
        n18814) );
  AOI22_X1 U21912 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18827), .B1(
        n18939), .B2(n18848), .ZN(n18813) );
  OAI211_X1 U21913 ( .C1(n18942), .C2(n18830), .A(n18814), .B(n18813), .ZN(
        P3_U2949) );
  AOI22_X1 U21914 ( .A1(n18945), .A2(n18848), .B1(n18943), .B2(n18825), .ZN(
        n18816) );
  AOI22_X1 U21915 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18827), .B1(
        n18944), .B2(n18826), .ZN(n18815) );
  OAI211_X1 U21916 ( .C1(n18948), .C2(n18830), .A(n18816), .B(n18815), .ZN(
        P3_U2950) );
  AOI22_X1 U21917 ( .A1(n18951), .A2(n18826), .B1(n18949), .B2(n18825), .ZN(
        n18818) );
  AOI22_X1 U21918 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18827), .B1(
        n18950), .B2(n18848), .ZN(n18817) );
  OAI211_X1 U21919 ( .C1(n18954), .C2(n18830), .A(n18818), .B(n18817), .ZN(
        P3_U2951) );
  AOI22_X1 U21920 ( .A1(n18957), .A2(n18826), .B1(n18955), .B2(n18825), .ZN(
        n18820) );
  AOI22_X1 U21921 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18827), .B1(
        n18956), .B2(n18848), .ZN(n18819) );
  OAI211_X1 U21922 ( .C1(n18960), .C2(n18830), .A(n18820), .B(n18819), .ZN(
        P3_U2952) );
  AOI22_X1 U21923 ( .A1(n18962), .A2(n18848), .B1(n18961), .B2(n18825), .ZN(
        n18822) );
  AOI22_X1 U21924 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18827), .B1(
        n18963), .B2(n18826), .ZN(n18821) );
  OAI211_X1 U21925 ( .C1(n18966), .C2(n18830), .A(n18822), .B(n18821), .ZN(
        P3_U2953) );
  AOI22_X1 U21926 ( .A1(n18968), .A2(n18848), .B1(n18967), .B2(n18825), .ZN(
        n18824) );
  AOI22_X1 U21927 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18827), .B1(
        n18969), .B2(n18826), .ZN(n18823) );
  OAI211_X1 U21928 ( .C1(n18972), .C2(n18830), .A(n18824), .B(n18823), .ZN(
        P3_U2954) );
  AOI22_X1 U21929 ( .A1(n18976), .A2(n18848), .B1(n18974), .B2(n18825), .ZN(
        n18829) );
  AOI22_X1 U21930 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18827), .B1(
        n18978), .B2(n18826), .ZN(n18828) );
  OAI211_X1 U21931 ( .C1(n18982), .C2(n18830), .A(n18829), .B(n18828), .ZN(
        P3_U2955) );
  NOR2_X1 U21932 ( .A1(n19012), .A2(n18831), .ZN(n18879) );
  NAND2_X1 U21933 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18879), .ZN(
        n18854) );
  AND2_X1 U21934 ( .A1(n19056), .A2(n18879), .ZN(n18847) );
  AOI22_X1 U21935 ( .A1(n18933), .A2(n18848), .B1(n18927), .B2(n18847), .ZN(
        n18834) );
  INV_X1 U21936 ( .A(n18832), .ZN(n18929) );
  OAI211_X1 U21937 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18932), .A(
        n18929), .B(n18852), .ZN(n18849) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18849), .B1(
        n18928), .B2(n18874), .ZN(n18833) );
  OAI211_X1 U21939 ( .C1(n18936), .C2(n18854), .A(n18834), .B(n18833), .ZN(
        P3_U2956) );
  AOI22_X1 U21940 ( .A1(n18937), .A2(n18847), .B1(n18939), .B2(n18874), .ZN(
        n18836) );
  AOI22_X1 U21941 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18849), .B1(
        n18938), .B2(n18848), .ZN(n18835) );
  OAI211_X1 U21942 ( .C1(n18942), .C2(n18854), .A(n18836), .B(n18835), .ZN(
        P3_U2957) );
  AOI22_X1 U21943 ( .A1(n18945), .A2(n18874), .B1(n18943), .B2(n18847), .ZN(
        n18838) );
  AOI22_X1 U21944 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18849), .B1(
        n18944), .B2(n18848), .ZN(n18837) );
  OAI211_X1 U21945 ( .C1(n18948), .C2(n18854), .A(n18838), .B(n18837), .ZN(
        P3_U2958) );
  AOI22_X1 U21946 ( .A1(n18950), .A2(n18874), .B1(n18949), .B2(n18847), .ZN(
        n18840) );
  AOI22_X1 U21947 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18849), .B1(
        n18951), .B2(n18848), .ZN(n18839) );
  OAI211_X1 U21948 ( .C1(n18954), .C2(n18854), .A(n18840), .B(n18839), .ZN(
        P3_U2959) );
  AOI22_X1 U21949 ( .A1(n18956), .A2(n18874), .B1(n18955), .B2(n18847), .ZN(
        n18842) );
  AOI22_X1 U21950 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18849), .B1(
        n18957), .B2(n18848), .ZN(n18841) );
  OAI211_X1 U21951 ( .C1(n18960), .C2(n18854), .A(n18842), .B(n18841), .ZN(
        P3_U2960) );
  AOI22_X1 U21952 ( .A1(n18963), .A2(n18848), .B1(n18961), .B2(n18847), .ZN(
        n18844) );
  AOI22_X1 U21953 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18849), .B1(
        n18962), .B2(n18874), .ZN(n18843) );
  OAI211_X1 U21954 ( .C1(n18966), .C2(n18854), .A(n18844), .B(n18843), .ZN(
        P3_U2961) );
  AOI22_X1 U21955 ( .A1(n18969), .A2(n18848), .B1(n18967), .B2(n18847), .ZN(
        n18846) );
  AOI22_X1 U21956 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18849), .B1(
        n18968), .B2(n18874), .ZN(n18845) );
  OAI211_X1 U21957 ( .C1(n18972), .C2(n18854), .A(n18846), .B(n18845), .ZN(
        P3_U2962) );
  AOI22_X1 U21958 ( .A1(n18976), .A2(n18874), .B1(n18974), .B2(n18847), .ZN(
        n18851) );
  AOI22_X1 U21959 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18849), .B1(
        n18978), .B2(n18848), .ZN(n18850) );
  OAI211_X1 U21960 ( .C1(n18982), .C2(n18854), .A(n18851), .B(n18850), .ZN(
        P3_U2963) );
  NAND2_X1 U21961 ( .A1(n18931), .A2(n19010), .ZN(n18877) );
  INV_X1 U21962 ( .A(n18877), .ZN(n18977) );
  NAND2_X1 U21963 ( .A1(n18853), .A2(n18852), .ZN(n18855) );
  INV_X1 U21964 ( .A(n18854), .ZN(n18922) );
  NOR2_X1 U21965 ( .A1(n18922), .A2(n18977), .ZN(n18903) );
  OAI21_X1 U21966 ( .B1(n18856), .B2(n18855), .A(n18903), .ZN(n18857) );
  OAI211_X1 U21967 ( .C1(n18977), .C2(n19160), .A(n18905), .B(n18857), .ZN(
        n18873) );
  NOR2_X1 U21968 ( .A1(n18900), .A2(n18903), .ZN(n18872) );
  AOI22_X1 U21969 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18873), .B1(
        n18927), .B2(n18872), .ZN(n18859) );
  AOI22_X1 U21970 ( .A1(n18933), .A2(n18874), .B1(n18928), .B2(n18895), .ZN(
        n18858) );
  OAI211_X1 U21971 ( .C1(n18936), .C2(n18877), .A(n18859), .B(n18858), .ZN(
        P3_U2964) );
  AOI22_X1 U21972 ( .A1(n18937), .A2(n18872), .B1(n18939), .B2(n18895), .ZN(
        n18861) );
  AOI22_X1 U21973 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18873), .B1(
        n18938), .B2(n18874), .ZN(n18860) );
  OAI211_X1 U21974 ( .C1(n18942), .C2(n18877), .A(n18861), .B(n18860), .ZN(
        P3_U2965) );
  AOI22_X1 U21975 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18873), .B1(
        n18943), .B2(n18872), .ZN(n18863) );
  AOI22_X1 U21976 ( .A1(n18944), .A2(n18874), .B1(n18945), .B2(n18895), .ZN(
        n18862) );
  OAI211_X1 U21977 ( .C1(n18948), .C2(n18877), .A(n18863), .B(n18862), .ZN(
        P3_U2966) );
  AOI22_X1 U21978 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18873), .B1(
        n18949), .B2(n18872), .ZN(n18865) );
  AOI22_X1 U21979 ( .A1(n18951), .A2(n18874), .B1(n18950), .B2(n18895), .ZN(
        n18864) );
  OAI211_X1 U21980 ( .C1(n18954), .C2(n18877), .A(n18865), .B(n18864), .ZN(
        P3_U2967) );
  AOI22_X1 U21981 ( .A1(n18956), .A2(n18895), .B1(n18955), .B2(n18872), .ZN(
        n18867) );
  AOI22_X1 U21982 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18873), .B1(
        n18957), .B2(n18874), .ZN(n18866) );
  OAI211_X1 U21983 ( .C1(n18960), .C2(n18877), .A(n18867), .B(n18866), .ZN(
        P3_U2968) );
  AOI22_X1 U21984 ( .A1(n18962), .A2(n18895), .B1(n18961), .B2(n18872), .ZN(
        n18869) );
  AOI22_X1 U21985 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18873), .B1(
        n18963), .B2(n18874), .ZN(n18868) );
  OAI211_X1 U21986 ( .C1(n18966), .C2(n18877), .A(n18869), .B(n18868), .ZN(
        P3_U2969) );
  AOI22_X1 U21987 ( .A1(n18968), .A2(n18895), .B1(n18967), .B2(n18872), .ZN(
        n18871) );
  AOI22_X1 U21988 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18873), .B1(
        n18969), .B2(n18874), .ZN(n18870) );
  OAI211_X1 U21989 ( .C1(n18972), .C2(n18877), .A(n18871), .B(n18870), .ZN(
        P3_U2970) );
  AOI22_X1 U21990 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18873), .B1(
        n18974), .B2(n18872), .ZN(n18876) );
  AOI22_X1 U21991 ( .A1(n18976), .A2(n18895), .B1(n18978), .B2(n18874), .ZN(
        n18875) );
  OAI211_X1 U21992 ( .C1(n18982), .C2(n18877), .A(n18876), .B(n18875), .ZN(
        P3_U2971) );
  INV_X1 U21993 ( .A(n18975), .ZN(n18899) );
  NOR2_X1 U21994 ( .A1(n18900), .A2(n18878), .ZN(n18894) );
  AOI22_X1 U21995 ( .A1(n18928), .A2(n18922), .B1(n18927), .B2(n18894), .ZN(
        n18881) );
  AOI22_X1 U21996 ( .A1(n18932), .A2(n18879), .B1(n18931), .B2(n18929), .ZN(
        n18896) );
  AOI22_X1 U21997 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18896), .B1(
        n18933), .B2(n18895), .ZN(n18880) );
  OAI211_X1 U21998 ( .C1(n18936), .C2(n18899), .A(n18881), .B(n18880), .ZN(
        P3_U2972) );
  AOI22_X1 U21999 ( .A1(n18938), .A2(n18895), .B1(n18937), .B2(n18894), .ZN(
        n18883) );
  AOI22_X1 U22000 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18896), .B1(
        n18939), .B2(n18922), .ZN(n18882) );
  OAI211_X1 U22001 ( .C1(n18942), .C2(n18899), .A(n18883), .B(n18882), .ZN(
        P3_U2973) );
  AOI22_X1 U22002 ( .A1(n18944), .A2(n18895), .B1(n18943), .B2(n18894), .ZN(
        n18885) );
  AOI22_X1 U22003 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18896), .B1(
        n18945), .B2(n18922), .ZN(n18884) );
  OAI211_X1 U22004 ( .C1(n18948), .C2(n18899), .A(n18885), .B(n18884), .ZN(
        P3_U2974) );
  AOI22_X1 U22005 ( .A1(n18951), .A2(n18895), .B1(n18949), .B2(n18894), .ZN(
        n18887) );
  AOI22_X1 U22006 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18896), .B1(
        n18950), .B2(n18922), .ZN(n18886) );
  OAI211_X1 U22007 ( .C1(n18954), .C2(n18899), .A(n18887), .B(n18886), .ZN(
        P3_U2975) );
  AOI22_X1 U22008 ( .A1(n18957), .A2(n18895), .B1(n18955), .B2(n18894), .ZN(
        n18889) );
  AOI22_X1 U22009 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18896), .B1(
        n18956), .B2(n18922), .ZN(n18888) );
  OAI211_X1 U22010 ( .C1(n18960), .C2(n18899), .A(n18889), .B(n18888), .ZN(
        P3_U2976) );
  AOI22_X1 U22011 ( .A1(n18962), .A2(n18922), .B1(n18961), .B2(n18894), .ZN(
        n18891) );
  AOI22_X1 U22012 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18896), .B1(
        n18963), .B2(n18895), .ZN(n18890) );
  OAI211_X1 U22013 ( .C1(n18966), .C2(n18899), .A(n18891), .B(n18890), .ZN(
        P3_U2977) );
  AOI22_X1 U22014 ( .A1(n18969), .A2(n18895), .B1(n18967), .B2(n18894), .ZN(
        n18893) );
  AOI22_X1 U22015 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18896), .B1(
        n18968), .B2(n18922), .ZN(n18892) );
  OAI211_X1 U22016 ( .C1(n18972), .C2(n18899), .A(n18893), .B(n18892), .ZN(
        P3_U2978) );
  AOI22_X1 U22017 ( .A1(n18976), .A2(n18922), .B1(n18974), .B2(n18894), .ZN(
        n18898) );
  AOI22_X1 U22018 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18896), .B1(
        n18978), .B2(n18895), .ZN(n18897) );
  OAI211_X1 U22019 ( .C1(n18982), .C2(n18899), .A(n18898), .B(n18897), .ZN(
        P3_U2979) );
  INV_X1 U22020 ( .A(n18906), .ZN(n18926) );
  NOR2_X1 U22021 ( .A1(n18900), .A2(n18901), .ZN(n18921) );
  AOI22_X1 U22022 ( .A1(n18928), .A2(n18977), .B1(n18927), .B2(n18921), .ZN(
        n18908) );
  OAI21_X1 U22023 ( .B1(n18903), .B2(n18902), .A(n18901), .ZN(n18904) );
  OAI211_X1 U22024 ( .C1(n18906), .C2(n19160), .A(n18905), .B(n18904), .ZN(
        n18923) );
  AOI22_X1 U22025 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18923), .B1(
        n18933), .B2(n18922), .ZN(n18907) );
  OAI211_X1 U22026 ( .C1(n18936), .C2(n18926), .A(n18908), .B(n18907), .ZN(
        P3_U2980) );
  AOI22_X1 U22027 ( .A1(n18938), .A2(n18922), .B1(n18937), .B2(n18921), .ZN(
        n18910) );
  AOI22_X1 U22028 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18923), .B1(
        n18939), .B2(n18977), .ZN(n18909) );
  OAI211_X1 U22029 ( .C1(n18942), .C2(n18926), .A(n18910), .B(n18909), .ZN(
        P3_U2981) );
  AOI22_X1 U22030 ( .A1(n18945), .A2(n18977), .B1(n18943), .B2(n18921), .ZN(
        n18912) );
  AOI22_X1 U22031 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18923), .B1(
        n18944), .B2(n18922), .ZN(n18911) );
  OAI211_X1 U22032 ( .C1(n18948), .C2(n18926), .A(n18912), .B(n18911), .ZN(
        P3_U2982) );
  AOI22_X1 U22033 ( .A1(n18951), .A2(n18922), .B1(n18949), .B2(n18921), .ZN(
        n18914) );
  AOI22_X1 U22034 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18923), .B1(
        n18950), .B2(n18977), .ZN(n18913) );
  OAI211_X1 U22035 ( .C1(n18954), .C2(n18926), .A(n18914), .B(n18913), .ZN(
        P3_U2983) );
  AOI22_X1 U22036 ( .A1(n18957), .A2(n18922), .B1(n18955), .B2(n18921), .ZN(
        n18916) );
  AOI22_X1 U22037 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18923), .B1(
        n18956), .B2(n18977), .ZN(n18915) );
  OAI211_X1 U22038 ( .C1(n18960), .C2(n18926), .A(n18916), .B(n18915), .ZN(
        P3_U2984) );
  AOI22_X1 U22039 ( .A1(n18962), .A2(n18977), .B1(n18961), .B2(n18921), .ZN(
        n18918) );
  AOI22_X1 U22040 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18923), .B1(
        n18963), .B2(n18922), .ZN(n18917) );
  OAI211_X1 U22041 ( .C1(n18966), .C2(n18926), .A(n18918), .B(n18917), .ZN(
        P3_U2985) );
  AOI22_X1 U22042 ( .A1(n18969), .A2(n18922), .B1(n18967), .B2(n18921), .ZN(
        n18920) );
  AOI22_X1 U22043 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18923), .B1(
        n18968), .B2(n18977), .ZN(n18919) );
  OAI211_X1 U22044 ( .C1(n18972), .C2(n18926), .A(n18920), .B(n18919), .ZN(
        P3_U2986) );
  AOI22_X1 U22045 ( .A1(n18976), .A2(n18977), .B1(n18974), .B2(n18921), .ZN(
        n18925) );
  AOI22_X1 U22046 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18923), .B1(
        n18978), .B2(n18922), .ZN(n18924) );
  OAI211_X1 U22047 ( .C1(n18982), .C2(n18926), .A(n18925), .B(n18924), .ZN(
        P3_U2987) );
  AND2_X1 U22048 ( .A1(n19056), .A2(n18930), .ZN(n18973) );
  AOI22_X1 U22049 ( .A1(n18928), .A2(n18975), .B1(n18927), .B2(n18973), .ZN(
        n18935) );
  AOI22_X1 U22050 ( .A1(n18932), .A2(n18931), .B1(n18930), .B2(n18929), .ZN(
        n18979) );
  AOI22_X1 U22051 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18979), .B1(
        n18933), .B2(n18977), .ZN(n18934) );
  OAI211_X1 U22052 ( .C1(n18983), .C2(n18936), .A(n18935), .B(n18934), .ZN(
        P3_U2988) );
  AOI22_X1 U22053 ( .A1(n18938), .A2(n18977), .B1(n18937), .B2(n18973), .ZN(
        n18941) );
  AOI22_X1 U22054 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18979), .B1(
        n18939), .B2(n18975), .ZN(n18940) );
  OAI211_X1 U22055 ( .C1(n18983), .C2(n18942), .A(n18941), .B(n18940), .ZN(
        P3_U2989) );
  AOI22_X1 U22056 ( .A1(n18944), .A2(n18977), .B1(n18943), .B2(n18973), .ZN(
        n18947) );
  AOI22_X1 U22057 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18979), .B1(
        n18945), .B2(n18975), .ZN(n18946) );
  OAI211_X1 U22058 ( .C1(n18983), .C2(n18948), .A(n18947), .B(n18946), .ZN(
        P3_U2990) );
  AOI22_X1 U22059 ( .A1(n18950), .A2(n18975), .B1(n18949), .B2(n18973), .ZN(
        n18953) );
  AOI22_X1 U22060 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18979), .B1(
        n18951), .B2(n18977), .ZN(n18952) );
  OAI211_X1 U22061 ( .C1(n18983), .C2(n18954), .A(n18953), .B(n18952), .ZN(
        P3_U2991) );
  AOI22_X1 U22062 ( .A1(n18956), .A2(n18975), .B1(n18955), .B2(n18973), .ZN(
        n18959) );
  AOI22_X1 U22063 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18979), .B1(
        n18957), .B2(n18977), .ZN(n18958) );
  OAI211_X1 U22064 ( .C1(n18983), .C2(n18960), .A(n18959), .B(n18958), .ZN(
        P3_U2992) );
  AOI22_X1 U22065 ( .A1(n18962), .A2(n18975), .B1(n18961), .B2(n18973), .ZN(
        n18965) );
  AOI22_X1 U22066 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18979), .B1(
        n18963), .B2(n18977), .ZN(n18964) );
  OAI211_X1 U22067 ( .C1(n18983), .C2(n18966), .A(n18965), .B(n18964), .ZN(
        P3_U2993) );
  AOI22_X1 U22068 ( .A1(n18968), .A2(n18975), .B1(n18967), .B2(n18973), .ZN(
        n18971) );
  AOI22_X1 U22069 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18979), .B1(
        n18969), .B2(n18977), .ZN(n18970) );
  OAI211_X1 U22070 ( .C1(n18983), .C2(n18972), .A(n18971), .B(n18970), .ZN(
        P3_U2994) );
  AOI22_X1 U22071 ( .A1(n18976), .A2(n18975), .B1(n18974), .B2(n18973), .ZN(
        n18981) );
  AOI22_X1 U22072 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18979), .B1(
        n18978), .B2(n18977), .ZN(n18980) );
  OAI211_X1 U22073 ( .C1(n18983), .C2(n18982), .A(n18981), .B(n18980), .ZN(
        P3_U2995) );
  AND2_X1 U22074 ( .A1(n19014), .A2(n18984), .ZN(n18985) );
  OAI22_X1 U22075 ( .A1(n18988), .A2(n18987), .B1(n18986), .B2(n18985), .ZN(
        n18989) );
  AOI221_X1 U22076 ( .B1(n18992), .B2(n18991), .C1(n18990), .C2(n18991), .A(
        n18989), .ZN(n19203) );
  AOI211_X1 U22077 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19029), .A(
        n18994), .B(n18993), .ZN(n19043) );
  INV_X1 U22078 ( .A(n18995), .ZN(n18999) );
  OAI21_X1 U22079 ( .B1(n18998), .B2(n18997), .A(n18996), .ZN(n19018) );
  AOI22_X1 U22080 ( .A1(n19026), .A2(n19002), .B1(n18999), .B2(n19018), .ZN(
        n19001) );
  NAND2_X1 U22081 ( .A1(n19001), .A2(n19000), .ZN(n19166) );
  NOR2_X1 U22082 ( .A1(n19029), .A2(n19166), .ZN(n19005) );
  NOR2_X1 U22083 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19002), .ZN(
        n19008) );
  OAI22_X1 U22084 ( .A1(n19003), .A2(n19023), .B1(n19008), .B2(n19026), .ZN(
        n19163) );
  NAND2_X1 U22085 ( .A1(n19167), .A2(n19163), .ZN(n19004) );
  OAI22_X1 U22086 ( .A1(n19005), .A2(n19167), .B1(n19029), .B2(n19004), .ZN(
        n19039) );
  NOR2_X1 U22087 ( .A1(n19006), .A2(n19015), .ZN(n19009) );
  OAI22_X1 U22088 ( .A1(n19009), .A2(n19178), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19008), .ZN(n19183) );
  OR3_X1 U22089 ( .A1(n19187), .A2(n19012), .A3(n19010), .ZN(n19011) );
  AOI22_X1 U22090 ( .A1(n19187), .A2(n19012), .B1(n19183), .B2(n19011), .ZN(
        n19013) );
  NOR2_X1 U22091 ( .A1(n19029), .A2(n19013), .ZN(n19031) );
  AOI21_X1 U22092 ( .B1(n19185), .B2(n19177), .A(n19014), .ZN(n19027) );
  NAND2_X1 U22093 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19015), .ZN(
        n19016) );
  AOI211_X1 U22094 ( .C1(n19017), .C2(n19016), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n19185), .ZN(n19025) );
  AOI21_X1 U22095 ( .B1(n19185), .B2(n19019), .A(n19018), .ZN(n19022) );
  NAND2_X1 U22096 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19020), .ZN(
        n19021) );
  OAI22_X1 U22097 ( .A1(n19174), .A2(n19023), .B1(n19022), .B2(n19021), .ZN(
        n19024) );
  AOI211_X1 U22098 ( .C1(n19027), .C2(n19026), .A(n19025), .B(n19024), .ZN(
        n19170) );
  INV_X1 U22099 ( .A(n19029), .ZN(n19028) );
  AOI22_X1 U22100 ( .A1(n19029), .A2(n19177), .B1(n19170), .B2(n19028), .ZN(
        n19033) );
  OAI22_X1 U22101 ( .A1(n19032), .A2(n19031), .B1(n19030), .B2(n19033), .ZN(
        n19034) );
  INV_X1 U22102 ( .A(n19033), .ZN(n19035) );
  OAI221_X1 U22103 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n19034), .A(n19035), .ZN(
        n19038) );
  NOR2_X1 U22104 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19037) );
  OAI21_X1 U22105 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19035), .A(
        n19034), .ZN(n19036) );
  AOI22_X1 U22106 ( .A1(n19039), .A2(n19038), .B1(n19037), .B2(n19036), .ZN(
        n19042) );
  OAI21_X1 U22107 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19040), .ZN(n19041) );
  NAND4_X1 U22108 ( .A1(n19203), .A2(n19043), .A3(n19042), .A4(n19041), .ZN(
        n19049) );
  AOI211_X1 U22109 ( .C1(n19046), .C2(n19045), .A(n19044), .B(n19049), .ZN(
        n19157) );
  NOR2_X1 U22110 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19213), .ZN(n19054) );
  NOR2_X1 U22111 ( .A1(n19157), .A2(n19054), .ZN(n19057) );
  NOR2_X1 U22112 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19215) );
  NOR2_X1 U22113 ( .A1(n19213), .A2(n19207), .ZN(n19053) );
  AOI211_X1 U22114 ( .C1(n19186), .C2(n19215), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n19053), .ZN(n19047) );
  AOI211_X1 U22115 ( .C1(n19206), .C2(n19049), .A(n19048), .B(n19047), .ZN(
        n19050) );
  OAI221_X1 U22116 ( .B1(n19052), .B2(n19057), .C1(n19052), .C2(n19051), .A(
        n19050), .ZN(P3_U2996) );
  INV_X1 U22117 ( .A(n19053), .ZN(n19060) );
  NAND3_X1 U22118 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n19054), .ZN(n19062) );
  INV_X1 U22119 ( .A(n19055), .ZN(n19058) );
  NAND3_X1 U22120 ( .A1(n19058), .A2(n19057), .A3(n19056), .ZN(n19059) );
  NAND4_X1 U22121 ( .A1(n19061), .A2(n19060), .A3(n19062), .A4(n19059), .ZN(
        P3_U2997) );
  INV_X1 U22122 ( .A(n19215), .ZN(n19064) );
  AND4_X1 U22123 ( .A1(n19064), .A2(n19063), .A3(n19062), .A4(n19158), .ZN(
        P3_U2998) );
  AND2_X1 U22124 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n9634), .ZN(P3_U2999) );
  AND2_X1 U22125 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n9633), .ZN(P3_U3000) );
  AND2_X1 U22126 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n9634), .ZN(P3_U3001) );
  AND2_X1 U22127 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n9633), .ZN(P3_U3002) );
  AND2_X1 U22128 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n9634), .ZN(P3_U3003) );
  AND2_X1 U22129 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n9633), .ZN(P3_U3004) );
  AND2_X1 U22130 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n9633), .ZN(P3_U3005) );
  AND2_X1 U22131 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n9634), .ZN(P3_U3006) );
  AND2_X1 U22132 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n9633), .ZN(P3_U3007) );
  AND2_X1 U22133 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n9634), .ZN(P3_U3008) );
  AND2_X1 U22134 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n9633), .ZN(P3_U3009) );
  AND2_X1 U22135 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n9634), .ZN(P3_U3010) );
  AND2_X1 U22136 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n9633), .ZN(P3_U3011) );
  AND2_X1 U22137 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n9634), .ZN(P3_U3012) );
  AND2_X1 U22138 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n9633), .ZN(P3_U3013) );
  AND2_X1 U22139 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n9634), .ZN(P3_U3014) );
  AND2_X1 U22140 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n9633), .ZN(P3_U3015) );
  AND2_X1 U22141 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n9634), .ZN(P3_U3016) );
  AND2_X1 U22142 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n9634), .ZN(P3_U3017) );
  AND2_X1 U22143 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n9633), .ZN(P3_U3018) );
  AND2_X1 U22144 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n9634), .ZN(P3_U3019) );
  AND2_X1 U22145 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n9633), .ZN(P3_U3020) );
  AND2_X1 U22146 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n9633), .ZN(P3_U3021)
         );
  AND2_X1 U22147 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n9634), .ZN(P3_U3022)
         );
  AND2_X1 U22148 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n9633), .ZN(P3_U3023)
         );
  AND2_X1 U22149 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n9634), .ZN(P3_U3024)
         );
  AND2_X1 U22150 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n9633), .ZN(P3_U3025)
         );
  AND2_X1 U22151 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n9634), .ZN(P3_U3026)
         );
  AND2_X1 U22152 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n9633), .ZN(P3_U3027)
         );
  AND2_X1 U22153 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n9634), .ZN(P3_U3028)
         );
  NOR2_X1 U22154 ( .A1(n19081), .A2(n21190), .ZN(n19077) );
  INV_X1 U22155 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19072) );
  AOI211_X1 U22156 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n19077), .B(
        n19072), .ZN(n19068) );
  NOR2_X1 U22157 ( .A1(n19213), .A2(n19073), .ZN(n19074) );
  OAI21_X1 U22158 ( .B1(n19074), .B2(n19079), .A(n19081), .ZN(n19067) );
  NAND3_X1 U22159 ( .A1(NA), .A2(n19079), .A3(n19073), .ZN(n19066) );
  OAI211_X1 U22160 ( .C1(n19151), .C2(n19068), .A(n19067), .B(n19066), .ZN(
        P3_U3029) );
  NAND2_X1 U22161 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n19071) );
  NOR2_X1 U22162 ( .A1(n19077), .A2(n19072), .ZN(n19069) );
  AOI22_X1 U22163 ( .A1(n19208), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n19069), .ZN(n19070) );
  OAI211_X1 U22164 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(n19071), .A(n19070), 
        .B(n19210), .ZN(P3_U3030) );
  INV_X1 U22165 ( .A(NA), .ZN(n21230) );
  AOI221_X1 U22166 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n19079), .C1(n21230), 
        .C2(n19079), .A(n19074), .ZN(n19080) );
  AOI22_X1 U22167 ( .A1(n21230), .A2(n19074), .B1(n19073), .B2(n19072), .ZN(
        n19075) );
  INV_X1 U22168 ( .A(n19075), .ZN(n19076) );
  OAI22_X1 U22169 ( .A1(n19077), .A2(n19076), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19078) );
  OAI22_X1 U22170 ( .A1(n19080), .A2(n19081), .B1(n19079), .B2(n19078), .ZN(
        P3_U3031) );
  OAI222_X1 U22171 ( .A1(n19191), .A2(n19137), .B1(n19082), .B2(n19151), .C1(
        n19083), .C2(n19140), .ZN(P3_U3032) );
  OAI222_X1 U22172 ( .A1(n19140), .A2(n19085), .B1(n19084), .B2(n19151), .C1(
        n19083), .C2(n19144), .ZN(P3_U3033) );
  OAI222_X1 U22173 ( .A1(n19140), .A2(n19087), .B1(n19086), .B2(n19151), .C1(
        n19085), .C2(n19137), .ZN(P3_U3034) );
  INV_X1 U22174 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19090) );
  OAI222_X1 U22175 ( .A1(n19140), .A2(n19090), .B1(n19088), .B2(n19151), .C1(
        n19087), .C2(n19137), .ZN(P3_U3035) );
  OAI222_X1 U22176 ( .A1(n19090), .A2(n19137), .B1(n19089), .B2(n19151), .C1(
        n19091), .C2(n19140), .ZN(P3_U3036) );
  OAI222_X1 U22177 ( .A1(n19140), .A2(n19093), .B1(n19092), .B2(n19151), .C1(
        n19091), .C2(n19137), .ZN(P3_U3037) );
  OAI222_X1 U22178 ( .A1(n19140), .A2(n19096), .B1(n19094), .B2(n19151), .C1(
        n19093), .C2(n19137), .ZN(P3_U3038) );
  OAI222_X1 U22179 ( .A1(n19096), .A2(n19137), .B1(n19095), .B2(n19151), .C1(
        n19097), .C2(n19140), .ZN(P3_U3039) );
  OAI222_X1 U22180 ( .A1(n19140), .A2(n19099), .B1(n19098), .B2(n19151), .C1(
        n19097), .C2(n19137), .ZN(P3_U3040) );
  INV_X1 U22181 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19101) );
  OAI222_X1 U22182 ( .A1(n19140), .A2(n19101), .B1(n19100), .B2(n19151), .C1(
        n19099), .C2(n19137), .ZN(P3_U3041) );
  OAI222_X1 U22183 ( .A1(n19140), .A2(n19103), .B1(n19102), .B2(n19151), .C1(
        n19101), .C2(n19137), .ZN(P3_U3042) );
  OAI222_X1 U22184 ( .A1(n19140), .A2(n19105), .B1(n19104), .B2(n19151), .C1(
        n19103), .C2(n19137), .ZN(P3_U3043) );
  OAI222_X1 U22185 ( .A1(n19140), .A2(n19108), .B1(n19106), .B2(n19151), .C1(
        n19105), .C2(n19137), .ZN(P3_U3044) );
  OAI222_X1 U22186 ( .A1(n19108), .A2(n19137), .B1(n19107), .B2(n19151), .C1(
        n19109), .C2(n19140), .ZN(P3_U3045) );
  OAI222_X1 U22187 ( .A1(n19140), .A2(n19111), .B1(n19110), .B2(n19151), .C1(
        n19109), .C2(n19137), .ZN(P3_U3046) );
  INV_X1 U22188 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19114) );
  OAI222_X1 U22189 ( .A1(n19140), .A2(n19114), .B1(n19112), .B2(n19151), .C1(
        n19111), .C2(n19144), .ZN(P3_U3047) );
  OAI222_X1 U22190 ( .A1(n19114), .A2(n19137), .B1(n19113), .B2(n19151), .C1(
        n19115), .C2(n19140), .ZN(P3_U3048) );
  INV_X1 U22191 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19117) );
  OAI222_X1 U22192 ( .A1(n19140), .A2(n19117), .B1(n19116), .B2(n19151), .C1(
        n19115), .C2(n19144), .ZN(P3_U3049) );
  OAI222_X1 U22193 ( .A1(n19140), .A2(n19120), .B1(n19118), .B2(n19151), .C1(
        n19117), .C2(n19144), .ZN(P3_U3050) );
  OAI222_X1 U22194 ( .A1(n19120), .A2(n19137), .B1(n19119), .B2(n19151), .C1(
        n19121), .C2(n19140), .ZN(P3_U3051) );
  OAI222_X1 U22195 ( .A1(n19140), .A2(n19123), .B1(n19122), .B2(n19151), .C1(
        n19121), .C2(n19144), .ZN(P3_U3052) );
  OAI222_X1 U22196 ( .A1(n19140), .A2(n19125), .B1(n19124), .B2(n19151), .C1(
        n19123), .C2(n19144), .ZN(P3_U3053) );
  OAI222_X1 U22197 ( .A1(n19140), .A2(n19127), .B1(n19126), .B2(n19151), .C1(
        n19125), .C2(n19144), .ZN(P3_U3054) );
  OAI222_X1 U22198 ( .A1(n19140), .A2(n19129), .B1(n19128), .B2(n19151), .C1(
        n19127), .C2(n19144), .ZN(P3_U3055) );
  OAI222_X1 U22199 ( .A1(n19140), .A2(n19131), .B1(n19130), .B2(n19151), .C1(
        n19129), .C2(n19137), .ZN(P3_U3056) );
  OAI222_X1 U22200 ( .A1(n19140), .A2(n19133), .B1(n19132), .B2(n19151), .C1(
        n19131), .C2(n19137), .ZN(P3_U3057) );
  INV_X1 U22201 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19136) );
  OAI222_X1 U22202 ( .A1(n19140), .A2(n19136), .B1(n19134), .B2(n19151), .C1(
        n19133), .C2(n19137), .ZN(P3_U3058) );
  OAI222_X1 U22203 ( .A1(n19136), .A2(n19137), .B1(n19135), .B2(n19151), .C1(
        n19138), .C2(n19140), .ZN(P3_U3059) );
  OAI222_X1 U22204 ( .A1(n19140), .A2(n19143), .B1(n19139), .B2(n19151), .C1(
        n19138), .C2(n19137), .ZN(P3_U3060) );
  INV_X1 U22205 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19142) );
  OAI222_X1 U22206 ( .A1(n19144), .A2(n19143), .B1(n19142), .B2(n19151), .C1(
        n19141), .C2(n19140), .ZN(P3_U3061) );
  INV_X1 U22207 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19145) );
  AOI22_X1 U22208 ( .A1(n19151), .A2(n19146), .B1(n19145), .B2(n19220), .ZN(
        P3_U3274) );
  INV_X1 U22209 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19193) );
  INV_X1 U22210 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19147) );
  AOI22_X1 U22211 ( .A1(n19151), .A2(n19193), .B1(n19147), .B2(n19220), .ZN(
        P3_U3275) );
  INV_X1 U22212 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19148) );
  AOI22_X1 U22213 ( .A1(n19151), .A2(n19149), .B1(n19148), .B2(n19220), .ZN(
        P3_U3276) );
  INV_X1 U22214 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19199) );
  INV_X1 U22215 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19150) );
  AOI22_X1 U22216 ( .A1(n19151), .A2(n19199), .B1(n19150), .B2(n19220), .ZN(
        P3_U3277) );
  INV_X1 U22217 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19153) );
  AOI21_X1 U22218 ( .B1(n9634), .B2(n19153), .A(n19152), .ZN(P3_U3280) );
  OAI21_X1 U22219 ( .B1(n19156), .B2(n19155), .A(n19154), .ZN(P3_U3281) );
  INV_X1 U22220 ( .A(n19157), .ZN(n19159) );
  OAI221_X1 U22221 ( .B1(n19160), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19160), 
        .C2(n19159), .A(n19158), .ZN(P3_U3282) );
  INV_X1 U22222 ( .A(n19189), .ZN(n19190) );
  INV_X1 U22223 ( .A(n19161), .ZN(n19165) );
  NOR2_X1 U22224 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19162), .ZN(
        n19164) );
  AOI22_X1 U22225 ( .A1(n19186), .A2(n19165), .B1(n19164), .B2(n19163), .ZN(
        n19169) );
  AOI21_X1 U22226 ( .B1(n19223), .B2(n19166), .A(n19190), .ZN(n19168) );
  OAI22_X1 U22227 ( .A1(n19190), .A2(n19169), .B1(n19168), .B2(n19167), .ZN(
        P3_U3285) );
  INV_X1 U22228 ( .A(n19170), .ZN(n19175) );
  NOR2_X1 U22229 ( .A1(n19171), .A2(n19188), .ZN(n19180) );
  AOI22_X1 U22230 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19173), .B2(n19172), .ZN(
        n19179) );
  AOI222_X1 U22231 ( .A1(n19175), .A2(n19223), .B1(n19180), .B2(n19179), .C1(
        n19186), .C2(n19174), .ZN(n19176) );
  AOI22_X1 U22232 ( .A1(n19190), .A2(n19177), .B1(n19176), .B2(n19189), .ZN(
        P3_U3288) );
  INV_X1 U22233 ( .A(n19178), .ZN(n19182) );
  INV_X1 U22234 ( .A(n19179), .ZN(n19181) );
  AOI222_X1 U22235 ( .A1(n19183), .A2(n19223), .B1(n19186), .B2(n19182), .C1(
        n19181), .C2(n19180), .ZN(n19184) );
  AOI22_X1 U22236 ( .A1(n19190), .A2(n19185), .B1(n19184), .B2(n19189), .ZN(
        P3_U3289) );
  AOI21_X1 U22237 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19192) );
  AOI22_X1 U22238 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19192), .B2(n19191), .ZN(n19194) );
  AOI22_X1 U22239 ( .A1(n19195), .A2(n19194), .B1(n19193), .B2(n19198), .ZN(
        P3_U3292) );
  NOR2_X1 U22240 ( .A1(n19198), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19196) );
  AOI22_X1 U22241 ( .A1(n19199), .A2(n19198), .B1(n19197), .B2(n19196), .ZN(
        P3_U3293) );
  INV_X1 U22242 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19200) );
  AOI22_X1 U22243 ( .A1(n19151), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19200), 
        .B2(n19220), .ZN(P3_U3294) );
  INV_X1 U22244 ( .A(n19201), .ZN(n19204) );
  NAND2_X1 U22245 ( .A1(n19204), .A2(P3_MORE_REG_SCAN_IN), .ZN(n19202) );
  OAI21_X1 U22246 ( .B1(n19204), .B2(n19203), .A(n19202), .ZN(P3_U3295) );
  OAI22_X1 U22247 ( .A1(n19208), .A2(n19207), .B1(n19206), .B2(n19205), .ZN(
        n19209) );
  NOR2_X1 U22248 ( .A1(n19226), .A2(n19209), .ZN(n19219) );
  AOI21_X1 U22249 ( .B1(n19212), .B2(n19211), .A(n19210), .ZN(n19214) );
  OAI211_X1 U22250 ( .C1(n19224), .C2(n19214), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19213), .ZN(n19216) );
  AOI21_X1 U22251 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19216), .A(n19215), 
        .ZN(n19218) );
  NAND2_X1 U22252 ( .A1(n19219), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19217) );
  OAI21_X1 U22253 ( .B1(n19219), .B2(n19218), .A(n19217), .ZN(P3_U3296) );
  INV_X1 U22254 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19229) );
  INV_X1 U22255 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19221) );
  AOI22_X1 U22256 ( .A1(n19151), .A2(n19229), .B1(n19221), .B2(n19220), .ZN(
        P3_U3297) );
  AOI21_X1 U22257 ( .B1(n19223), .B2(n19222), .A(n19226), .ZN(n19230) );
  INV_X1 U22258 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19227) );
  INV_X1 U22259 ( .A(n19224), .ZN(n19225) );
  AOI22_X1 U22260 ( .A1(n19230), .A2(n19227), .B1(n19226), .B2(n19225), .ZN(
        P3_U3298) );
  AOI21_X1 U22261 ( .B1(n19230), .B2(n19229), .A(n19228), .ZN(P3_U3299) );
  INV_X1 U22262 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19235) );
  INV_X1 U22263 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19231) );
  INV_X1 U22264 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20133) );
  NAND2_X1 U22265 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20133), .ZN(n20121) );
  AOI22_X1 U22266 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20121), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19235), .ZN(n20186) );
  INV_X1 U22267 ( .A(n20186), .ZN(n20115) );
  OAI21_X1 U22268 ( .B1(n19235), .B2(n19231), .A(n20115), .ZN(P2_U2815) );
  INV_X1 U22269 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19234) );
  NAND2_X1 U22270 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19761), .ZN(n19232) );
  OAI22_X1 U22271 ( .A1(n20253), .A2(n19234), .B1(n19233), .B2(n19232), .ZN(
        P2_U2816) );
  INV_X1 U22272 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20125) );
  OR2_X1 U22273 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20125), .ZN(n20271) );
  INV_X2 U22274 ( .A(n20271), .ZN(n20274) );
  OR2_X1 U22275 ( .A1(n20124), .A2(n20274), .ZN(n20118) );
  AOI21_X1 U22276 ( .B1(n19235), .B2(n20118), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19236) );
  AOI21_X1 U22277 ( .B1(n20274), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n19236), 
        .ZN(P2_U2817) );
  OAI21_X1 U22278 ( .B1(n20124), .B2(BS16), .A(n20186), .ZN(n20184) );
  OAI21_X1 U22279 ( .B1(n20186), .B2(n19820), .A(n20184), .ZN(P2_U2818) );
  NOR2_X1 U22280 ( .A1(n19238), .A2(n19237), .ZN(n20250) );
  OAI21_X1 U22281 ( .B1(n20250), .B2(n11632), .A(n19239), .ZN(P2_U2819) );
  NOR4_X1 U22282 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19243) );
  NOR4_X1 U22283 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19242) );
  NOR4_X1 U22284 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19241) );
  NOR4_X1 U22285 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19240) );
  NAND4_X1 U22286 ( .A1(n19243), .A2(n19242), .A3(n19241), .A4(n19240), .ZN(
        n19249) );
  NOR4_X1 U22287 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19247) );
  AOI211_X1 U22288 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19246) );
  NOR4_X1 U22289 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19245) );
  NOR4_X1 U22290 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19244) );
  NAND4_X1 U22291 ( .A1(n19247), .A2(n19246), .A3(n19245), .A4(n19244), .ZN(
        n19248) );
  NOR2_X1 U22292 ( .A1(n19249), .A2(n19248), .ZN(n19257) );
  INV_X1 U22293 ( .A(n19257), .ZN(n19256) );
  NOR2_X1 U22294 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19256), .ZN(n19250) );
  INV_X1 U22295 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20182) );
  AOI22_X1 U22296 ( .A1(n19250), .A2(n19251), .B1(n19256), .B2(n20182), .ZN(
        P2_U2820) );
  OR3_X1 U22297 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19255) );
  INV_X1 U22298 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20180) );
  AOI22_X1 U22299 ( .A1(n19250), .A2(n19255), .B1(n19256), .B2(n20180), .ZN(
        P2_U2821) );
  INV_X1 U22300 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20185) );
  NAND2_X1 U22301 ( .A1(n19250), .A2(n20185), .ZN(n19254) );
  OAI21_X1 U22302 ( .B1(n10459), .B2(n19251), .A(n19257), .ZN(n19252) );
  OAI21_X1 U22303 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19257), .A(n19252), 
        .ZN(n19253) );
  OAI221_X1 U22304 ( .B1(n19254), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19254), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19253), .ZN(P2_U2822) );
  INV_X1 U22305 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20178) );
  OAI221_X1 U22306 ( .B1(n19257), .B2(n20178), .C1(n19256), .C2(n19255), .A(
        n19254), .ZN(P2_U2823) );
  AOI22_X1 U22307 ( .A1(n19259), .A2(n19425), .B1(n19258), .B2(n19420), .ZN(
        n19268) );
  AOI211_X1 U22308 ( .C1(n19262), .C2(n19261), .A(n19260), .B(n19394), .ZN(
        n19266) );
  AOI22_X1 U22309 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19431), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19402), .ZN(n19263) );
  OAI21_X1 U22310 ( .B1(n19264), .B2(n19423), .A(n19263), .ZN(n19265) );
  AOI211_X1 U22311 ( .C1(P2_EBX_REG_20__SCAN_IN), .C2(n19406), .A(n19266), .B(
        n19265), .ZN(n19267) );
  NAND2_X1 U22312 ( .A1(n19268), .A2(n19267), .ZN(P2_U2835) );
  AOI211_X1 U22313 ( .C1(n19271), .C2(n19270), .A(n19394), .B(n19269), .ZN(
        n19278) );
  NOR2_X1 U22314 ( .A1(n19272), .A2(n19423), .ZN(n19277) );
  NOR2_X1 U22315 ( .A1(n19273), .A2(n19389), .ZN(n19276) );
  AOI22_X1 U22316 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n19406), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19431), .ZN(n19274) );
  OAI211_X1 U22317 ( .C1(n19416), .C2(n20154), .A(n19274), .B(n19364), .ZN(
        n19275) );
  NOR4_X1 U22318 ( .A1(n19278), .A2(n19277), .A3(n19276), .A4(n19275), .ZN(
        n19279) );
  OAI21_X1 U22319 ( .B1(n19280), .B2(n19408), .A(n19279), .ZN(P2_U2836) );
  INV_X1 U22320 ( .A(n19281), .ZN(n19288) );
  NAND2_X1 U22321 ( .A1(n19393), .A2(n19411), .ZN(n19429) );
  AOI22_X1 U22322 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19431), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19402), .ZN(n19282) );
  OAI211_X1 U22323 ( .C1(n19429), .C2(n19283), .A(n19333), .B(n19282), .ZN(
        n19284) );
  AOI21_X1 U22324 ( .B1(n19406), .B2(P2_EBX_REG_17__SCAN_IN), .A(n19284), .ZN(
        n19285) );
  OAI21_X1 U22325 ( .B1(n19286), .B2(n19389), .A(n19285), .ZN(n19287) );
  AOI21_X1 U22326 ( .B1(n19288), .B2(n12839), .A(n19287), .ZN(n19295) );
  AOI21_X1 U22327 ( .B1(n19291), .B2(n19290), .A(n19289), .ZN(n19292) );
  AOI22_X1 U22328 ( .A1(n19293), .A2(n19420), .B1(n19427), .B2(n19292), .ZN(
        n19294) );
  NAND2_X1 U22329 ( .A1(n19295), .A2(n19294), .ZN(P2_U2838) );
  OAI22_X1 U22330 ( .A1(n19296), .A2(n19423), .B1(n10321), .B2(n19386), .ZN(
        n19297) );
  AOI211_X1 U22331 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19402), .A(n16616), 
        .B(n19297), .ZN(n19307) );
  NOR2_X1 U22332 ( .A1(n19393), .A2(n19298), .ZN(n19299) );
  XNOR2_X1 U22333 ( .A(n19300), .B(n19299), .ZN(n19305) );
  INV_X1 U22334 ( .A(n19301), .ZN(n19303) );
  OAI22_X1 U22335 ( .A1(n19303), .A2(n19389), .B1(n19408), .B2(n19302), .ZN(
        n19304) );
  AOI21_X1 U22336 ( .B1(n19305), .B2(n19411), .A(n19304), .ZN(n19306) );
  OAI211_X1 U22337 ( .C1(n19418), .C2(n14071), .A(n19307), .B(n19306), .ZN(
        P2_U2839) );
  OAI21_X1 U22338 ( .B1(n10948), .B2(n19416), .A(n19364), .ZN(n19310) );
  OAI22_X1 U22339 ( .A1(n19308), .A2(n19423), .B1(n10599), .B2(n19418), .ZN(
        n19309) );
  AOI211_X1 U22340 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19431), .A(
        n19310), .B(n19309), .ZN(n19317) );
  NAND2_X1 U22341 ( .A1(n9658), .A2(n19311), .ZN(n19312) );
  XNOR2_X1 U22342 ( .A(n19313), .B(n19312), .ZN(n19315) );
  AOI22_X1 U22343 ( .A1(n19315), .A2(n19411), .B1(n19425), .B2(n19314), .ZN(
        n19316) );
  OAI211_X1 U22344 ( .C1(n19442), .C2(n19408), .A(n19317), .B(n19316), .ZN(
        P2_U2840) );
  INV_X1 U22345 ( .A(n19427), .ZN(n19318) );
  AOI211_X1 U22346 ( .C1(n19327), .C2(n19320), .A(n19319), .B(n19318), .ZN(
        n19326) );
  NAND2_X1 U22347 ( .A1(n19321), .A2(n12839), .ZN(n19324) );
  AOI22_X1 U22348 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19431), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19402), .ZN(n19323) );
  NAND2_X1 U22349 ( .A1(n19406), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n19322) );
  NAND4_X1 U22350 ( .A1(n19324), .A2(n19323), .A3(n19333), .A4(n19322), .ZN(
        n19325) );
  NOR2_X1 U22351 ( .A1(n19326), .A2(n19325), .ZN(n19332) );
  INV_X1 U22352 ( .A(n19327), .ZN(n19328) );
  OAI22_X1 U22353 ( .A1(n19329), .A2(n19389), .B1(n19429), .B2(n19328), .ZN(
        n19330) );
  INV_X1 U22354 ( .A(n19330), .ZN(n19331) );
  OAI211_X1 U22355 ( .C1(n19447), .C2(n19408), .A(n19332), .B(n19331), .ZN(
        P2_U2842) );
  OAI21_X1 U22356 ( .B1(n10888), .B2(n19416), .A(n19333), .ZN(n19336) );
  OAI22_X1 U22357 ( .A1(n19334), .A2(n19423), .B1(n19418), .B2(n10578), .ZN(
        n19335) );
  AOI211_X1 U22358 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n19431), .A(
        n19336), .B(n19335), .ZN(n19343) );
  NAND2_X1 U22359 ( .A1(n9658), .A2(n19337), .ZN(n19338) );
  XNOR2_X1 U22360 ( .A(n19339), .B(n19338), .ZN(n19341) );
  AOI22_X1 U22361 ( .A1(n19341), .A2(n19411), .B1(n19425), .B2(n19340), .ZN(
        n19342) );
  OAI211_X1 U22362 ( .C1(n19452), .C2(n19408), .A(n19343), .B(n19342), .ZN(
        P2_U2844) );
  AOI22_X1 U22363 ( .A1(P2_EBX_REG_10__SCAN_IN), .A2(n19406), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19431), .ZN(n19344) );
  OAI21_X1 U22364 ( .B1(n19345), .B2(n19423), .A(n19344), .ZN(n19346) );
  AOI211_X1 U22365 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19402), .A(n16616), 
        .B(n19346), .ZN(n19353) );
  NOR2_X1 U22366 ( .A1(n19393), .A2(n19347), .ZN(n19349) );
  XNOR2_X1 U22367 ( .A(n19349), .B(n19348), .ZN(n19351) );
  AOI22_X1 U22368 ( .A1(n19351), .A2(n19411), .B1(n19425), .B2(n19350), .ZN(
        n19352) );
  OAI211_X1 U22369 ( .C1(n19455), .C2(n19408), .A(n19353), .B(n19352), .ZN(
        P2_U2845) );
  OAI21_X1 U22370 ( .B1(n10855), .B2(n19416), .A(n19364), .ZN(n19356) );
  OAI22_X1 U22371 ( .A1(n19354), .A2(n19423), .B1(n10570), .B2(n19418), .ZN(
        n19355) );
  AOI211_X1 U22372 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19431), .A(
        n19356), .B(n19355), .ZN(n19363) );
  NAND2_X1 U22373 ( .A1(n9658), .A2(n19357), .ZN(n19358) );
  XNOR2_X1 U22374 ( .A(n19359), .B(n19358), .ZN(n19361) );
  AOI22_X1 U22375 ( .A1(n19361), .A2(n19411), .B1(n19425), .B2(n19360), .ZN(
        n19362) );
  OAI211_X1 U22376 ( .C1(n19457), .C2(n19408), .A(n19363), .B(n19362), .ZN(
        P2_U2846) );
  OAI21_X1 U22377 ( .B1(n16058), .B2(n19416), .A(n19364), .ZN(n19367) );
  OAI22_X1 U22378 ( .A1(n19365), .A2(n19423), .B1(n19418), .B2(n10560), .ZN(
        n19366) );
  AOI211_X1 U22379 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19431), .A(
        n19367), .B(n19366), .ZN(n19374) );
  NOR2_X1 U22380 ( .A1(n19393), .A2(n19368), .ZN(n19370) );
  XNOR2_X1 U22381 ( .A(n19370), .B(n19369), .ZN(n19372) );
  AOI22_X1 U22382 ( .A1(n19372), .A2(n19411), .B1(n19425), .B2(n19371), .ZN(
        n19373) );
  OAI211_X1 U22383 ( .C1(n19408), .C2(n19465), .A(n19374), .B(n19373), .ZN(
        P2_U2849) );
  AOI22_X1 U22384 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(n19406), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19431), .ZN(n19375) );
  OAI21_X1 U22385 ( .B1(n19376), .B2(n19423), .A(n19375), .ZN(n19377) );
  AOI211_X1 U22386 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19402), .A(n16616), .B(
        n19377), .ZN(n19385) );
  NAND2_X1 U22387 ( .A1(n9658), .A2(n19378), .ZN(n19380) );
  XNOR2_X1 U22388 ( .A(n19381), .B(n19380), .ZN(n19383) );
  AOI22_X1 U22389 ( .A1(n19383), .A2(n19411), .B1(n19425), .B2(n19382), .ZN(
        n19384) );
  OAI211_X1 U22390 ( .C1(n19408), .C2(n19472), .A(n19385), .B(n19384), .ZN(
        P2_U2850) );
  OAI22_X1 U22391 ( .A1(n19387), .A2(n19423), .B1(n10070), .B2(n19386), .ZN(
        n19388) );
  AOI211_X1 U22392 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19402), .A(n16616), .B(
        n19388), .ZN(n19401) );
  AOI22_X1 U22393 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19406), .B1(n19420), .B2(
        n19474), .ZN(n19400) );
  OAI22_X1 U22394 ( .A1(n19476), .A2(n19390), .B1(n19389), .B2(n19558), .ZN(
        n19391) );
  INV_X1 U22395 ( .A(n19391), .ZN(n19399) );
  INV_X1 U22396 ( .A(n19563), .ZN(n19397) );
  NOR2_X1 U22397 ( .A1(n19393), .A2(n19392), .ZN(n19396) );
  AOI21_X1 U22398 ( .B1(n19397), .B2(n19396), .A(n19394), .ZN(n19395) );
  OAI21_X1 U22399 ( .B1(n19397), .B2(n19396), .A(n19395), .ZN(n19398) );
  NAND4_X1 U22400 ( .A1(n19401), .A2(n19400), .A3(n19399), .A4(n19398), .ZN(
        P2_U2851) );
  AOI22_X1 U22401 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19431), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19402), .ZN(n19403) );
  OAI21_X1 U22402 ( .B1(n19423), .B2(n19404), .A(n19403), .ZN(n19405) );
  AOI21_X1 U22403 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n19406), .A(n19405), .ZN(
        n19407) );
  OAI21_X1 U22404 ( .B1(n19409), .B2(n19408), .A(n19407), .ZN(n19410) );
  AOI21_X1 U22405 ( .B1(n9644), .B2(n19425), .A(n19410), .ZN(n19414) );
  AOI22_X1 U22406 ( .A1(n19412), .A2(n19411), .B1(n19428), .B2(n20224), .ZN(
        n19413) );
  OAI211_X1 U22407 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19429), .A(
        n19414), .B(n19413), .ZN(P2_U2854) );
  INV_X1 U22408 ( .A(n19415), .ZN(n19499) );
  OAI22_X1 U22409 ( .A1(n19418), .A2(n19417), .B1(n19416), .B2(n19251), .ZN(
        n19419) );
  AOI21_X1 U22410 ( .B1(n19420), .B2(n19499), .A(n19419), .ZN(n19421) );
  OAI21_X1 U22411 ( .B1(n19423), .B2(n19422), .A(n19421), .ZN(n19424) );
  AOI21_X1 U22412 ( .B1(n13050), .B2(n19425), .A(n19424), .ZN(n19434) );
  AOI22_X1 U22413 ( .A1(n19500), .A2(n19428), .B1(n19427), .B2(n19426), .ZN(
        n19433) );
  INV_X1 U22414 ( .A(n19429), .ZN(n19430) );
  OAI21_X1 U22415 ( .B1(n19431), .B2(n19430), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19432) );
  NAND3_X1 U22416 ( .A1(n19434), .A2(n19433), .A3(n19432), .ZN(P2_U2855) );
  INV_X1 U22417 ( .A(n19435), .ZN(n19437) );
  AOI22_X1 U22418 ( .A1(n19437), .A2(n19495), .B1(n19436), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19440) );
  AOI22_X1 U22419 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19494), .B1(n19438), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19439) );
  NAND2_X1 U22420 ( .A1(n19440), .A2(n19439), .ZN(P2_U2888) );
  OAI222_X1 U22421 ( .A1(n19442), .A2(n19473), .B1(n13022), .B2(n19466), .C1(
        n19441), .C2(n19503), .ZN(P2_U2904) );
  INV_X1 U22422 ( .A(n19443), .ZN(n19445) );
  AOI22_X1 U22423 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19494), .B1(n19546), 
        .B2(n19459), .ZN(n19444) );
  OAI21_X1 U22424 ( .B1(n19473), .B2(n19445), .A(n19444), .ZN(P2_U2905) );
  INV_X1 U22425 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19515) );
  OAI222_X1 U22426 ( .A1(n19447), .A2(n19473), .B1(n19515), .B2(n19466), .C1(
        n19503), .C2(n19446), .ZN(P2_U2906) );
  INV_X1 U22427 ( .A(n19448), .ZN(n19450) );
  INV_X1 U22428 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19517) );
  OAI222_X1 U22429 ( .A1(n19450), .A2(n19473), .B1(n19517), .B2(n19466), .C1(
        n19503), .C2(n19449), .ZN(P2_U2907) );
  INV_X1 U22430 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19519) );
  OAI222_X1 U22431 ( .A1(n19452), .A2(n19473), .B1(n19519), .B2(n19466), .C1(
        n19503), .C2(n19451), .ZN(P2_U2908) );
  AOI22_X1 U22432 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19494), .B1(n19453), 
        .B2(n19459), .ZN(n19454) );
  OAI21_X1 U22433 ( .B1(n19473), .B2(n19455), .A(n19454), .ZN(P2_U2909) );
  INV_X1 U22434 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19523) );
  OAI222_X1 U22435 ( .A1(n19457), .A2(n19473), .B1(n19523), .B2(n19466), .C1(
        n19503), .C2(n19456), .ZN(P2_U2910) );
  INV_X1 U22436 ( .A(n19458), .ZN(n19462) );
  AOI22_X1 U22437 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19494), .B1(n19460), .B2(
        n19459), .ZN(n19461) );
  OAI21_X1 U22438 ( .B1(n19473), .B2(n19462), .A(n19461), .ZN(P2_U2911) );
  INV_X1 U22439 ( .A(n19463), .ZN(n19464) );
  INV_X1 U22440 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19527) );
  OAI222_X1 U22441 ( .A1(n19464), .A2(n19473), .B1(n19527), .B2(n19466), .C1(
        n19503), .C2(n19616), .ZN(P2_U2912) );
  INV_X1 U22442 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19529) );
  OAI222_X1 U22443 ( .A1(n19465), .A2(n19473), .B1(n19529), .B2(n19466), .C1(
        n19503), .C2(n19604), .ZN(P2_U2913) );
  INV_X1 U22444 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19531) );
  OAI22_X1 U22445 ( .A1(n19531), .A2(n19466), .B1(n19598), .B2(n19503), .ZN(
        n19467) );
  INV_X1 U22446 ( .A(n19467), .ZN(n19471) );
  AOI21_X1 U22447 ( .B1(n20213), .B2(n20210), .A(n19468), .ZN(n19484) );
  XNOR2_X1 U22448 ( .A(n20204), .B(n20206), .ZN(n19483) );
  NOR2_X1 U22449 ( .A1(n19484), .A2(n19483), .ZN(n19482) );
  AOI21_X1 U22450 ( .B1(n20206), .B2(n20204), .A(n19482), .ZN(n19469) );
  NOR2_X1 U22451 ( .A1(n19469), .A2(n19474), .ZN(n19475) );
  OR3_X1 U22452 ( .A1(n19475), .A2(n19476), .A3(n19490), .ZN(n19470) );
  OAI211_X1 U22453 ( .C1(n19473), .C2(n19472), .A(n19471), .B(n19470), .ZN(
        P2_U2914) );
  AOI22_X1 U22454 ( .A1(n19495), .A2(n19474), .B1(n19494), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19479) );
  XOR2_X1 U22455 ( .A(n19476), .B(n19475), .Z(n19477) );
  NAND2_X1 U22456 ( .A1(n19477), .A2(n19497), .ZN(n19478) );
  OAI211_X1 U22457 ( .C1(n19480), .C2(n19503), .A(n19479), .B(n19478), .ZN(
        P2_U2915) );
  INV_X1 U22458 ( .A(n20206), .ZN(n19481) );
  AOI22_X1 U22459 ( .A1(n19481), .A2(n19495), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19494), .ZN(n19487) );
  AOI21_X1 U22460 ( .B1(n19484), .B2(n19483), .A(n19482), .ZN(n19485) );
  OR2_X1 U22461 ( .A1(n19485), .A2(n19490), .ZN(n19486) );
  OAI211_X1 U22462 ( .C1(n19587), .C2(n19503), .A(n19487), .B(n19486), .ZN(
        P2_U2916) );
  AOI22_X1 U22463 ( .A1(n19495), .A2(n20227), .B1(n19494), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19493) );
  AOI21_X1 U22464 ( .B1(n19496), .B2(n19489), .A(n19488), .ZN(n19491) );
  OR2_X1 U22465 ( .A1(n19491), .A2(n19490), .ZN(n19492) );
  OAI211_X1 U22466 ( .C1(n19578), .C2(n19503), .A(n19493), .B(n19492), .ZN(
        P2_U2918) );
  AOI22_X1 U22467 ( .A1(n19495), .A2(n19499), .B1(n19494), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19502) );
  INV_X1 U22468 ( .A(n19496), .ZN(n19498) );
  OAI211_X1 U22469 ( .C1(n19500), .C2(n19499), .A(n19498), .B(n19497), .ZN(
        n19501) );
  OAI211_X1 U22470 ( .C1(n19504), .C2(n19503), .A(n19502), .B(n19501), .ZN(
        P2_U2919) );
  NOR2_X1 U22471 ( .A1(n19509), .A2(n19505), .ZN(P2_U2920) );
  INV_X1 U22472 ( .A(n19506), .ZN(n19507) );
  AOI22_X1 U22473 ( .A1(n19507), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n20255), .ZN(n19508) );
  OAI21_X1 U22474 ( .B1(n19510), .B2(n19509), .A(n19508), .ZN(P2_U2921) );
  AOI22_X1 U22475 ( .A1(n20255), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19511) );
  OAI21_X1 U22476 ( .B1(n13022), .B2(n19542), .A(n19511), .ZN(P2_U2936) );
  INV_X1 U22477 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19513) );
  AOI22_X1 U22478 ( .A1(n20255), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19512) );
  OAI21_X1 U22479 ( .B1(n19513), .B2(n19542), .A(n19512), .ZN(P2_U2937) );
  AOI22_X1 U22480 ( .A1(n20255), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19514) );
  OAI21_X1 U22481 ( .B1(n19515), .B2(n19542), .A(n19514), .ZN(P2_U2938) );
  AOI22_X1 U22482 ( .A1(n20255), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19516) );
  OAI21_X1 U22483 ( .B1(n19517), .B2(n19542), .A(n19516), .ZN(P2_U2939) );
  AOI22_X1 U22484 ( .A1(n20255), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19518) );
  OAI21_X1 U22485 ( .B1(n19519), .B2(n19542), .A(n19518), .ZN(P2_U2940) );
  AOI22_X1 U22486 ( .A1(n20255), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19520) );
  OAI21_X1 U22487 ( .B1(n19521), .B2(n19542), .A(n19520), .ZN(P2_U2941) );
  AOI22_X1 U22488 ( .A1(n20255), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19522) );
  OAI21_X1 U22489 ( .B1(n19523), .B2(n19542), .A(n19522), .ZN(P2_U2942) );
  AOI22_X1 U22490 ( .A1(n20255), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19524) );
  OAI21_X1 U22491 ( .B1(n19525), .B2(n19542), .A(n19524), .ZN(P2_U2943) );
  AOI22_X1 U22492 ( .A1(n20255), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19526) );
  OAI21_X1 U22493 ( .B1(n19527), .B2(n19542), .A(n19526), .ZN(P2_U2944) );
  AOI22_X1 U22494 ( .A1(n20255), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19528) );
  OAI21_X1 U22495 ( .B1(n19529), .B2(n19542), .A(n19528), .ZN(P2_U2945) );
  AOI22_X1 U22496 ( .A1(n20255), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19530) );
  OAI21_X1 U22497 ( .B1(n19531), .B2(n19542), .A(n19530), .ZN(P2_U2946) );
  INV_X1 U22498 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19533) );
  AOI22_X1 U22499 ( .A1(n20255), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19532) );
  OAI21_X1 U22500 ( .B1(n19533), .B2(n19542), .A(n19532), .ZN(P2_U2947) );
  INV_X1 U22501 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19535) );
  AOI22_X1 U22502 ( .A1(n20255), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19534) );
  OAI21_X1 U22503 ( .B1(n19535), .B2(n19542), .A(n19534), .ZN(P2_U2948) );
  INV_X1 U22504 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19537) );
  AOI22_X1 U22505 ( .A1(n20255), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19536) );
  OAI21_X1 U22506 ( .B1(n19537), .B2(n19542), .A(n19536), .ZN(P2_U2949) );
  INV_X1 U22507 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19539) );
  AOI22_X1 U22508 ( .A1(n20255), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19538) );
  OAI21_X1 U22509 ( .B1(n19539), .B2(n19542), .A(n19538), .ZN(P2_U2950) );
  INV_X1 U22510 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19543) );
  AOI22_X1 U22511 ( .A1(n20255), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19540), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19541) );
  OAI21_X1 U22512 ( .B1(n19543), .B2(n19542), .A(n19541), .ZN(P2_U2951) );
  AOI22_X1 U22513 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19545), .B1(n19544), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19548) );
  NAND2_X1 U22514 ( .A1(n19547), .A2(n19546), .ZN(n19549) );
  NAND2_X1 U22515 ( .A1(n19548), .A2(n19549), .ZN(P2_U2966) );
  AOI22_X1 U22516 ( .A1(n19545), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13113), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19550) );
  NAND2_X1 U22517 ( .A1(n19550), .A2(n19549), .ZN(P2_U2981) );
  AOI22_X1 U22518 ( .A1(n19551), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n16616), .ZN(n19562) );
  NAND2_X1 U22519 ( .A1(n19553), .A2(n19552), .ZN(n19557) );
  NAND2_X1 U22520 ( .A1(n19555), .A2(n19554), .ZN(n19556) );
  OAI211_X1 U22521 ( .C1(n19559), .C2(n19558), .A(n19557), .B(n19556), .ZN(
        n19560) );
  INV_X1 U22522 ( .A(n19560), .ZN(n19561) );
  OAI211_X1 U22523 ( .C1(n19564), .C2(n19563), .A(n19562), .B(n19561), .ZN(
        P2_U3010) );
  NOR2_X1 U22524 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19565), .ZN(
        n19615) );
  AOI22_X1 U22525 ( .A1(n20092), .A2(n20055), .B1(n20046), .B2(n19615), .ZN(
        n19575) );
  NOR2_X1 U22526 ( .A1(n20092), .A2(n19639), .ZN(n19566) );
  OAI21_X1 U22527 ( .B1(n19566), .B2(n19820), .A(n20196), .ZN(n19573) );
  INV_X1 U22528 ( .A(n20051), .ZN(n20098) );
  NOR2_X1 U22529 ( .A1(n19573), .A2(n20098), .ZN(n19567) );
  AOI211_X1 U22530 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19569), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19567), .ZN(n19568) );
  NOR2_X1 U22531 ( .A1(n20098), .A2(n19615), .ZN(n19572) );
  INV_X1 U22532 ( .A(n19569), .ZN(n19570) );
  OAI21_X1 U22533 ( .B1(n19570), .B2(n19615), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19571) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19618), .B1(
        n20047), .B2(n19617), .ZN(n19574) );
  OAI211_X1 U22535 ( .C1(n20058), .C2(n19636), .A(n19575), .B(n19574), .ZN(
        P2_U3048) );
  OAI22_X1 U22536 ( .A1(n19576), .A2(n19611), .B1(n14163), .B2(n19609), .ZN(
        n20061) );
  AOI22_X1 U22537 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19608), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19607), .ZN(n20064) );
  NOR2_X2 U22538 ( .A1(n10493), .A2(n19596), .ZN(n20059) );
  INV_X1 U22539 ( .A(n20059), .ZN(n19864) );
  INV_X1 U22540 ( .A(n19615), .ZN(n19590) );
  OAI22_X1 U22541 ( .A1(n20106), .A2(n20064), .B1(n19864), .B2(n19590), .ZN(
        n19577) );
  INV_X1 U22542 ( .A(n19577), .ZN(n19580) );
  NOR2_X2 U22543 ( .A1(n19578), .A2(n19764), .ZN(n20060) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19618), .B1(
        n20060), .B2(n19617), .ZN(n19579) );
  OAI211_X1 U22545 ( .C1(n20018), .C2(n19636), .A(n19580), .B(n19579), .ZN(
        P2_U3049) );
  OAI22_X1 U22546 ( .A1(n19582), .A2(n19611), .B1(n19581), .B2(n19609), .ZN(
        n20067) );
  AOI22_X1 U22547 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19608), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19607), .ZN(n20070) );
  NOR2_X2 U22548 ( .A1(n10499), .A2(n19596), .ZN(n20065) );
  AOI22_X1 U22549 ( .A1(n20092), .A2(n19982), .B1(n20065), .B2(n19615), .ZN(
        n19585) );
  NOR2_X2 U22550 ( .A1(n19583), .A2(n19764), .ZN(n20066) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19618), .B1(
        n20066), .B2(n19617), .ZN(n19584) );
  OAI211_X1 U22552 ( .C1(n19985), .C2(n19636), .A(n19585), .B(n19584), .ZN(
        P2_U3050) );
  AOI22_X1 U22553 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19608), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19607), .ZN(n20076) );
  AOI22_X1 U22554 ( .A1(n20092), .A2(n20073), .B1(n20071), .B2(n19615), .ZN(
        n19589) );
  NOR2_X2 U22555 ( .A1(n19587), .A2(n19764), .ZN(n20072) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19618), .B1(
        n20072), .B2(n19617), .ZN(n19588) );
  OAI211_X1 U22557 ( .C1(n20076), .C2(n19636), .A(n19589), .B(n19588), .ZN(
        P2_U3051) );
  INV_X1 U22558 ( .A(n20079), .ZN(n20029) );
  OAI22_X1 U22559 ( .A1(n20106), .A2(n20082), .B1(n19873), .B2(n19590), .ZN(
        n19591) );
  INV_X1 U22560 ( .A(n19591), .ZN(n19593) );
  AOI22_X1 U22561 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19618), .B1(
        n20078), .B2(n19617), .ZN(n19592) );
  OAI211_X1 U22562 ( .C1(n20029), .C2(n19636), .A(n19593), .B(n19592), .ZN(
        P2_U3052) );
  AOI22_X1 U22563 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19608), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19607), .ZN(n20088) );
  INV_X1 U22564 ( .A(n20088), .ZN(n19990) );
  NOR2_X2 U22565 ( .A1(n19597), .A2(n19596), .ZN(n20083) );
  AOI22_X1 U22566 ( .A1(n20092), .A2(n19990), .B1(n20083), .B2(n19615), .ZN(
        n19600) );
  NOR2_X2 U22567 ( .A1(n19598), .A2(n19764), .ZN(n20084) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19618), .B1(
        n20084), .B2(n19617), .ZN(n19599) );
  OAI211_X1 U22569 ( .C1(n19993), .C2(n19636), .A(n19600), .B(n19599), .ZN(
        P2_U3053) );
  AOI22_X1 U22570 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19608), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19607), .ZN(n19997) );
  OAI22_X2 U22571 ( .A1(n19602), .A2(n19609), .B1(n19601), .B2(n19611), .ZN(
        n19994) );
  AND2_X1 U22572 ( .A1(n19603), .A2(n19613), .ZN(n20089) );
  AOI22_X1 U22573 ( .A1(n20092), .A2(n19994), .B1(n20089), .B2(n19615), .ZN(
        n19606) );
  NOR2_X2 U22574 ( .A1(n19604), .A2(n19764), .ZN(n20090) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19618), .B1(
        n20090), .B2(n19617), .ZN(n19605) );
  OAI211_X1 U22576 ( .C1(n19997), .C2(n19636), .A(n19606), .B(n19605), .ZN(
        P2_U3054) );
  OAI22_X2 U22577 ( .A1(n19612), .A2(n19611), .B1(n19610), .B2(n19609), .ZN(
        n20101) );
  AOI22_X1 U22578 ( .A1(n20092), .A2(n20101), .B1(n20097), .B2(n19615), .ZN(
        n19620) );
  NOR2_X2 U22579 ( .A1(n19616), .A2(n19764), .ZN(n20099) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19618), .B1(
        n20099), .B2(n19617), .ZN(n19619) );
  OAI211_X1 U22581 ( .C1(n20107), .C2(n19636), .A(n19620), .B(n19619), .ZN(
        P2_U3055) );
  AOI22_X1 U22582 ( .A1(n19638), .A2(n20047), .B1(n20046), .B2(n19637), .ZN(
        n19623) );
  AOI22_X1 U22583 ( .A1(n19639), .A2(n20055), .B1(n19669), .B2(n19621), .ZN(
        n19622) );
  OAI211_X1 U22584 ( .C1(n19625), .C2(n19624), .A(n19623), .B(n19622), .ZN(
        P2_U3056) );
  AOI22_X1 U22585 ( .A1(n19638), .A2(n20060), .B1(n20059), .B2(n19637), .ZN(
        n19627) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19640), .B1(
        n19669), .B2(n20061), .ZN(n19626) );
  OAI211_X1 U22587 ( .C1(n20064), .C2(n19636), .A(n19627), .B(n19626), .ZN(
        P2_U3057) );
  AOI22_X1 U22588 ( .A1(n19638), .A2(n20066), .B1(n20065), .B2(n19637), .ZN(
        n19629) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n19982), .ZN(n19628) );
  OAI211_X1 U22590 ( .C1(n19985), .C2(n19643), .A(n19629), .B(n19628), .ZN(
        P2_U3058) );
  AOI22_X1 U22591 ( .A1(n19638), .A2(n20072), .B1(n20071), .B2(n19637), .ZN(
        n19631) );
  INV_X1 U22592 ( .A(n20076), .ZN(n20021) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19640), .B1(
        n19669), .B2(n20021), .ZN(n19630) );
  OAI211_X1 U22594 ( .C1(n20024), .C2(n19636), .A(n19631), .B(n19630), .ZN(
        P2_U3059) );
  AOI22_X1 U22595 ( .A1(n19638), .A2(n20084), .B1(n20083), .B2(n19637), .ZN(
        n19633) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19640), .B1(
        n19669), .B2(n20085), .ZN(n19632) );
  OAI211_X1 U22597 ( .C1(n20088), .C2(n19636), .A(n19633), .B(n19632), .ZN(
        P2_U3061) );
  INV_X1 U22598 ( .A(n19994), .ZN(n20096) );
  AOI22_X1 U22599 ( .A1(n19638), .A2(n20090), .B1(n20089), .B2(n19637), .ZN(
        n19635) );
  INV_X1 U22600 ( .A(n19997), .ZN(n20091) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19640), .B1(
        n19669), .B2(n20091), .ZN(n19634) );
  OAI211_X1 U22602 ( .C1(n20096), .C2(n19636), .A(n19635), .B(n19634), .ZN(
        P2_U3062) );
  AOI22_X1 U22603 ( .A1(n19638), .A2(n20099), .B1(n20097), .B2(n19637), .ZN(
        n19642) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n20101), .ZN(n19641) );
  OAI211_X1 U22605 ( .C1(n20107), .C2(n19643), .A(n19642), .B(n19641), .ZN(
        P2_U3063) );
  INV_X1 U22606 ( .A(n19647), .ZN(n19644) );
  NOR2_X1 U22607 ( .A1(n20229), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19887) );
  AND2_X1 U22608 ( .A1(n19887), .A2(n19675), .ZN(n19667) );
  OAI21_X1 U22609 ( .B1(n19644), .B2(n19667), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19645) );
  OR2_X1 U22610 ( .A1(n19673), .A2(n19890), .ZN(n19648) );
  NAND2_X1 U22611 ( .A1(n19645), .A2(n19648), .ZN(n19668) );
  AOI22_X1 U22612 ( .A1(n19668), .A2(n20047), .B1(n20046), .B2(n19667), .ZN(
        n19654) );
  INV_X1 U22613 ( .A(n19667), .ZN(n19646) );
  OAI21_X1 U22614 ( .B1(n19647), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19646), 
        .ZN(n19651) );
  OAI21_X1 U22615 ( .B1(n19702), .B2(n19669), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19649) );
  NAND2_X1 U22616 ( .A1(n19649), .A2(n19648), .ZN(n19650) );
  MUX2_X1 U22617 ( .A(n19651), .B(n19650), .S(n20196), .Z(n19652) );
  NAND2_X1 U22618 ( .A1(n19652), .A2(n20053), .ZN(n19670) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n20055), .ZN(n19653) );
  OAI211_X1 U22620 ( .C1(n20058), .C2(n19698), .A(n19654), .B(n19653), .ZN(
        P2_U3064) );
  AOI22_X1 U22621 ( .A1(n19668), .A2(n20060), .B1(n20059), .B2(n19667), .ZN(
        n19656) );
  INV_X1 U22622 ( .A(n20064), .ZN(n20015) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n20015), .ZN(n19655) );
  OAI211_X1 U22624 ( .C1(n20018), .C2(n19698), .A(n19656), .B(n19655), .ZN(
        P2_U3065) );
  AOI22_X1 U22625 ( .A1(n19668), .A2(n20066), .B1(n20065), .B2(n19667), .ZN(
        n19658) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n19982), .ZN(n19657) );
  OAI211_X1 U22627 ( .C1(n19985), .C2(n19698), .A(n19658), .B(n19657), .ZN(
        P2_U3066) );
  AOI22_X1 U22628 ( .A1(n19668), .A2(n20072), .B1(n20071), .B2(n19667), .ZN(
        n19660) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n20073), .ZN(n19659) );
  OAI211_X1 U22630 ( .C1(n20076), .C2(n19698), .A(n19660), .B(n19659), .ZN(
        P2_U3067) );
  AOI22_X1 U22631 ( .A1(n19668), .A2(n20078), .B1(n20077), .B2(n19667), .ZN(
        n19662) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n20025), .ZN(n19661) );
  OAI211_X1 U22633 ( .C1(n20029), .C2(n19698), .A(n19662), .B(n19661), .ZN(
        P2_U3068) );
  AOI22_X1 U22634 ( .A1(n19668), .A2(n20084), .B1(n20083), .B2(n19667), .ZN(
        n19664) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n19990), .ZN(n19663) );
  OAI211_X1 U22636 ( .C1(n19993), .C2(n19698), .A(n19664), .B(n19663), .ZN(
        P2_U3069) );
  AOI22_X1 U22637 ( .A1(n19668), .A2(n20090), .B1(n20089), .B2(n19667), .ZN(
        n19666) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n19994), .ZN(n19665) );
  OAI211_X1 U22639 ( .C1(n19997), .C2(n19698), .A(n19666), .B(n19665), .ZN(
        P2_U3070) );
  AOI22_X1 U22640 ( .A1(n19668), .A2(n20099), .B1(n20097), .B2(n19667), .ZN(
        n19672) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19670), .B1(
        n19669), .B2(n20101), .ZN(n19671) );
  OAI211_X1 U22642 ( .C1(n20107), .C2(n19698), .A(n19672), .B(n19671), .ZN(
        P2_U3071) );
  NOR2_X1 U22643 ( .A1(n19673), .A2(n19917), .ZN(n19701) );
  AOI22_X1 U22644 ( .A1(n19702), .A2(n20055), .B1(n20046), .B2(n19701), .ZN(
        n19685) );
  AOI21_X1 U22645 ( .B1(n19794), .B2(n19674), .A(n20202), .ZN(n19679) );
  NAND2_X1 U22646 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19675), .ZN(
        n19682) );
  INV_X1 U22647 ( .A(n19701), .ZN(n19686) );
  NAND2_X1 U22648 ( .A1(n19676), .A2(n19686), .ZN(n19680) );
  NOR2_X1 U22649 ( .A1(n19680), .A2(n19761), .ZN(n19677) );
  AOI21_X1 U22650 ( .B1(n19679), .B2(n19682), .A(n19677), .ZN(n19678) );
  OAI211_X1 U22651 ( .C1(n19701), .C2(n20205), .A(n19678), .B(n20053), .ZN(
        n19704) );
  INV_X1 U22652 ( .A(n19679), .ZN(n19683) );
  INV_X1 U22653 ( .A(n19680), .ZN(n19681) );
  OAI22_X1 U22654 ( .A1(n19683), .A2(n19682), .B1(n19681), .B2(n19761), .ZN(
        n19703) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19704), .B1(
        n20047), .B2(n19703), .ZN(n19684) );
  OAI211_X1 U22656 ( .C1(n20058), .C2(n19707), .A(n19685), .B(n19684), .ZN(
        P2_U3072) );
  OAI22_X1 U22657 ( .A1(n19698), .A2(n20064), .B1(n19686), .B2(n19864), .ZN(
        n19687) );
  INV_X1 U22658 ( .A(n19687), .ZN(n19689) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19704), .B1(
        n20060), .B2(n19703), .ZN(n19688) );
  OAI211_X1 U22660 ( .C1(n20018), .C2(n19707), .A(n19689), .B(n19688), .ZN(
        P2_U3073) );
  AOI22_X1 U22661 ( .A1(n19702), .A2(n19982), .B1(n19701), .B2(n20065), .ZN(
        n19691) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19704), .B1(
        n20066), .B2(n19703), .ZN(n19690) );
  OAI211_X1 U22663 ( .C1(n19985), .C2(n19707), .A(n19691), .B(n19690), .ZN(
        P2_U3074) );
  AOI22_X1 U22664 ( .A1(n19733), .A2(n20021), .B1(n19701), .B2(n20071), .ZN(
        n19693) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19704), .B1(
        n20072), .B2(n19703), .ZN(n19692) );
  OAI211_X1 U22666 ( .C1(n20024), .C2(n19698), .A(n19693), .B(n19692), .ZN(
        P2_U3075) );
  AOI22_X1 U22667 ( .A1(n19733), .A2(n20079), .B1(n20077), .B2(n19701), .ZN(
        n19695) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19704), .B1(
        n20078), .B2(n19703), .ZN(n19694) );
  OAI211_X1 U22669 ( .C1(n20082), .C2(n19698), .A(n19695), .B(n19694), .ZN(
        P2_U3076) );
  AOI22_X1 U22670 ( .A1(n19733), .A2(n20085), .B1(n19701), .B2(n20083), .ZN(
        n19697) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19704), .B1(
        n20084), .B2(n19703), .ZN(n19696) );
  OAI211_X1 U22672 ( .C1(n20088), .C2(n19698), .A(n19697), .B(n19696), .ZN(
        P2_U3077) );
  AOI22_X1 U22673 ( .A1(n19702), .A2(n19994), .B1(n19701), .B2(n20089), .ZN(
        n19700) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19704), .B1(
        n20090), .B2(n19703), .ZN(n19699) );
  OAI211_X1 U22675 ( .C1(n19997), .C2(n19707), .A(n19700), .B(n19699), .ZN(
        P2_U3078) );
  AOI22_X1 U22676 ( .A1(n19702), .A2(n20101), .B1(n19701), .B2(n20097), .ZN(
        n19706) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19704), .B1(
        n20099), .B2(n19703), .ZN(n19705) );
  OAI211_X1 U22678 ( .C1(n20107), .C2(n19707), .A(n19706), .B(n19705), .ZN(
        P2_U3079) );
  NAND2_X1 U22679 ( .A1(n19708), .A2(n20209), .ZN(n19715) );
  INV_X1 U22680 ( .A(n19709), .ZN(n19712) );
  NOR2_X1 U22681 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19710), .ZN(
        n19731) );
  OAI21_X1 U22682 ( .B1(n19712), .B2(n19731), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19711) );
  OAI21_X1 U22683 ( .B1(n19715), .B2(n20202), .A(n19711), .ZN(n19732) );
  AOI22_X1 U22684 ( .A1(n19732), .A2(n20047), .B1(n20046), .B2(n19731), .ZN(
        n19718) );
  OAI21_X1 U22685 ( .B1(n19733), .B2(n19751), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19714) );
  AOI211_X1 U22686 ( .C1(n19712), .C2(n20205), .A(n20196), .B(n19731), .ZN(
        n19713) );
  AOI211_X1 U22687 ( .C1(n19715), .C2(n19714), .A(n19764), .B(n19713), .ZN(
        n19716) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n20055), .ZN(n19717) );
  OAI211_X1 U22689 ( .C1(n20058), .C2(n19748), .A(n19718), .B(n19717), .ZN(
        P2_U3080) );
  AOI22_X1 U22690 ( .A1(n19732), .A2(n20060), .B1(n20059), .B2(n19731), .ZN(
        n19720) );
  AOI22_X1 U22691 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n20015), .ZN(n19719) );
  OAI211_X1 U22692 ( .C1(n20018), .C2(n19748), .A(n19720), .B(n19719), .ZN(
        P2_U3081) );
  AOI22_X1 U22693 ( .A1(n19732), .A2(n20066), .B1(n20065), .B2(n19731), .ZN(
        n19722) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n19982), .ZN(n19721) );
  OAI211_X1 U22695 ( .C1(n19985), .C2(n19748), .A(n19722), .B(n19721), .ZN(
        P2_U3082) );
  AOI22_X1 U22696 ( .A1(n19732), .A2(n20072), .B1(n20071), .B2(n19731), .ZN(
        n19724) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n20073), .ZN(n19723) );
  OAI211_X1 U22698 ( .C1(n20076), .C2(n19748), .A(n19724), .B(n19723), .ZN(
        P2_U3083) );
  AOI22_X1 U22699 ( .A1(n19732), .A2(n20078), .B1(n20077), .B2(n19731), .ZN(
        n19726) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n20025), .ZN(n19725) );
  OAI211_X1 U22701 ( .C1(n20029), .C2(n19748), .A(n19726), .B(n19725), .ZN(
        P2_U3084) );
  AOI22_X1 U22702 ( .A1(n19732), .A2(n20084), .B1(n20083), .B2(n19731), .ZN(
        n19728) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n19990), .ZN(n19727) );
  OAI211_X1 U22704 ( .C1(n19993), .C2(n19748), .A(n19728), .B(n19727), .ZN(
        P2_U3085) );
  AOI22_X1 U22705 ( .A1(n19732), .A2(n20090), .B1(n20089), .B2(n19731), .ZN(
        n19730) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n19994), .ZN(n19729) );
  OAI211_X1 U22707 ( .C1(n19997), .C2(n19748), .A(n19730), .B(n19729), .ZN(
        P2_U3086) );
  AOI22_X1 U22708 ( .A1(n19732), .A2(n20099), .B1(n20097), .B2(n19731), .ZN(
        n19736) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n20101), .ZN(n19735) );
  OAI211_X1 U22710 ( .C1(n20107), .C2(n19748), .A(n19736), .B(n19735), .ZN(
        P2_U3087) );
  AOI22_X1 U22711 ( .A1(n19751), .A2(n20015), .B1(n9804), .B2(n20059), .ZN(
        n19738) );
  AOI22_X1 U22712 ( .A1(n20060), .A2(n19752), .B1(n19771), .B2(n20061), .ZN(
        n19737) );
  OAI211_X1 U22713 ( .C1(n19739), .C2(n11401), .A(n19738), .B(n19737), .ZN(
        P2_U3089) );
  AOI22_X1 U22714 ( .A1(n19771), .A2(n20067), .B1(n9804), .B2(n20065), .ZN(
        n19741) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19753), .B1(
        n20066), .B2(n19752), .ZN(n19740) );
  OAI211_X1 U22716 ( .C1(n20070), .C2(n19748), .A(n19741), .B(n19740), .ZN(
        P2_U3090) );
  AOI22_X1 U22717 ( .A1(n19771), .A2(n20021), .B1(n9804), .B2(n20071), .ZN(
        n19743) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19753), .B1(
        n20072), .B2(n19752), .ZN(n19742) );
  OAI211_X1 U22719 ( .C1(n20024), .C2(n19748), .A(n19743), .B(n19742), .ZN(
        P2_U3091) );
  AOI22_X1 U22720 ( .A1(n19771), .A2(n20079), .B1(n9804), .B2(n20077), .ZN(
        n19745) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19753), .B1(
        n20078), .B2(n19752), .ZN(n19744) );
  OAI211_X1 U22722 ( .C1(n20082), .C2(n19748), .A(n19745), .B(n19744), .ZN(
        P2_U3092) );
  AOI22_X1 U22723 ( .A1(n19771), .A2(n20085), .B1(n9804), .B2(n20083), .ZN(
        n19747) );
  AOI22_X1 U22724 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19753), .B1(
        n20084), .B2(n19752), .ZN(n19746) );
  OAI211_X1 U22725 ( .C1(n20088), .C2(n19748), .A(n19747), .B(n19746), .ZN(
        P2_U3093) );
  AOI22_X1 U22726 ( .A1(n19751), .A2(n19994), .B1(n9804), .B2(n20089), .ZN(
        n19750) );
  AOI22_X1 U22727 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19753), .B1(
        n20090), .B2(n19752), .ZN(n19749) );
  OAI211_X1 U22728 ( .C1(n19997), .C2(n19787), .A(n19750), .B(n19749), .ZN(
        P2_U3094) );
  AOI22_X1 U22729 ( .A1(n19751), .A2(n20101), .B1(n9804), .B2(n20097), .ZN(
        n19755) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19753), .B1(
        n20099), .B2(n19752), .ZN(n19754) );
  OAI211_X1 U22731 ( .C1(n20107), .C2(n19787), .A(n19755), .B(n19754), .ZN(
        P2_U3095) );
  INV_X1 U22732 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19761) );
  NAND2_X1 U22733 ( .A1(n20209), .A2(n20042), .ZN(n19796) );
  NOR2_X1 U22734 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19796), .ZN(
        n19782) );
  NOR2_X1 U22735 ( .A1(n19763), .A2(n19782), .ZN(n19757) );
  OR2_X1 U22736 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19757), .ZN(n19760) );
  INV_X1 U22737 ( .A(n19758), .ZN(n19759) );
  NOR3_X1 U22738 ( .A1(n19759), .A2(n19782), .A3(n19761), .ZN(n19765) );
  AOI21_X1 U22739 ( .B1(n19761), .B2(n19760), .A(n19765), .ZN(n19783) );
  AOI22_X1 U22740 ( .A1(n19783), .A2(n20047), .B1(n20046), .B2(n19782), .ZN(
        n19768) );
  AOI21_X1 U22741 ( .B1(n19787), .B2(n19813), .A(n19820), .ZN(n19762) );
  AOI221_X1 U22742 ( .B1(n20205), .B2(n19763), .C1(n20205), .C2(n19762), .A(
        n19782), .ZN(n19766) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19784), .B1(
        n19771), .B2(n20055), .ZN(n19767) );
  OAI211_X1 U22744 ( .C1(n20058), .C2(n19813), .A(n19768), .B(n19767), .ZN(
        P2_U3096) );
  AOI22_X1 U22745 ( .A1(n19783), .A2(n20060), .B1(n20059), .B2(n19782), .ZN(
        n19770) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19784), .B1(
        n19815), .B2(n20061), .ZN(n19769) );
  OAI211_X1 U22747 ( .C1(n20064), .C2(n19787), .A(n19770), .B(n19769), .ZN(
        P2_U3097) );
  AOI22_X1 U22748 ( .A1(n19783), .A2(n20066), .B1(n20065), .B2(n19782), .ZN(
        n19773) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19784), .B1(
        n19771), .B2(n19982), .ZN(n19772) );
  OAI211_X1 U22750 ( .C1(n19985), .C2(n19813), .A(n19773), .B(n19772), .ZN(
        P2_U3098) );
  AOI22_X1 U22751 ( .A1(n19783), .A2(n20072), .B1(n20071), .B2(n19782), .ZN(
        n19775) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19784), .B1(
        n19815), .B2(n20021), .ZN(n19774) );
  OAI211_X1 U22753 ( .C1(n20024), .C2(n19787), .A(n19775), .B(n19774), .ZN(
        P2_U3099) );
  AOI22_X1 U22754 ( .A1(n19783), .A2(n20078), .B1(n20077), .B2(n19782), .ZN(
        n19777) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19784), .B1(
        n19815), .B2(n20079), .ZN(n19776) );
  OAI211_X1 U22756 ( .C1(n20082), .C2(n19787), .A(n19777), .B(n19776), .ZN(
        P2_U3100) );
  AOI22_X1 U22757 ( .A1(n19783), .A2(n20084), .B1(n20083), .B2(n19782), .ZN(
        n19779) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19784), .B1(
        n19815), .B2(n20085), .ZN(n19778) );
  OAI211_X1 U22759 ( .C1(n20088), .C2(n19787), .A(n19779), .B(n19778), .ZN(
        P2_U3101) );
  AOI22_X1 U22760 ( .A1(n19783), .A2(n20090), .B1(n20089), .B2(n19782), .ZN(
        n19781) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19784), .B1(
        n19815), .B2(n20091), .ZN(n19780) );
  OAI211_X1 U22762 ( .C1(n20096), .C2(n19787), .A(n19781), .B(n19780), .ZN(
        P2_U3102) );
  INV_X1 U22763 ( .A(n20101), .ZN(n20041) );
  AOI22_X1 U22764 ( .A1(n19783), .A2(n20099), .B1(n20097), .B2(n19782), .ZN(
        n19786) );
  INV_X1 U22765 ( .A(n20107), .ZN(n20035) );
  AOI22_X1 U22766 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19784), .B1(
        n19815), .B2(n20035), .ZN(n19785) );
  OAI211_X1 U22767 ( .C1(n20041), .C2(n19787), .A(n19786), .B(n19785), .ZN(
        P2_U3103) );
  INV_X1 U22768 ( .A(n19789), .ZN(n19790) );
  NOR2_X1 U22769 ( .A1(n20239), .A2(n19796), .ZN(n19828) );
  NOR3_X1 U22770 ( .A1(n19790), .A2(n19828), .A3(n19761), .ZN(n19793) );
  INV_X1 U22771 ( .A(n19796), .ZN(n19791) );
  AOI21_X1 U22772 ( .B1(n19791), .B2(n20205), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19792) );
  NOR2_X1 U22773 ( .A1(n19793), .A2(n19792), .ZN(n19814) );
  AOI22_X1 U22774 ( .A1(n19814), .A2(n20047), .B1(n20046), .B2(n19828), .ZN(
        n19800) );
  INV_X1 U22775 ( .A(n19793), .ZN(n19798) );
  INV_X1 U22776 ( .A(n19828), .ZN(n19825) );
  NAND2_X1 U22777 ( .A1(n19795), .A2(n19794), .ZN(n20201) );
  AOI22_X1 U22778 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19825), .B1(n19796), 
        .B2(n20201), .ZN(n19797) );
  NAND3_X1 U22779 ( .A1(n19798), .A2(n20053), .A3(n19797), .ZN(n19816) );
  AOI22_X1 U22780 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n20055), .ZN(n19799) );
  OAI211_X1 U22781 ( .C1(n20058), .C2(n19844), .A(n19800), .B(n19799), .ZN(
        P2_U3104) );
  AOI22_X1 U22782 ( .A1(n19814), .A2(n20060), .B1(n20059), .B2(n19828), .ZN(
        n19802) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n20015), .ZN(n19801) );
  OAI211_X1 U22784 ( .C1(n20018), .C2(n19844), .A(n19802), .B(n19801), .ZN(
        P2_U3105) );
  AOI22_X1 U22785 ( .A1(n19814), .A2(n20066), .B1(n20065), .B2(n19828), .ZN(
        n19804) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19982), .ZN(n19803) );
  OAI211_X1 U22787 ( .C1(n19985), .C2(n19844), .A(n19804), .B(n19803), .ZN(
        P2_U3106) );
  AOI22_X1 U22788 ( .A1(n19814), .A2(n20072), .B1(n20071), .B2(n19828), .ZN(
        n19806) );
  INV_X1 U22789 ( .A(n19844), .ZN(n19848) );
  AOI22_X1 U22790 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19816), .B1(
        n19848), .B2(n20021), .ZN(n19805) );
  OAI211_X1 U22791 ( .C1(n20024), .C2(n19813), .A(n19806), .B(n19805), .ZN(
        P2_U3107) );
  AOI22_X1 U22792 ( .A1(n19814), .A2(n20078), .B1(n20077), .B2(n19828), .ZN(
        n19808) );
  AOI22_X1 U22793 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19816), .B1(
        n19848), .B2(n20079), .ZN(n19807) );
  OAI211_X1 U22794 ( .C1(n20082), .C2(n19813), .A(n19808), .B(n19807), .ZN(
        P2_U3108) );
  AOI22_X1 U22795 ( .A1(n19814), .A2(n20084), .B1(n20083), .B2(n19828), .ZN(
        n19810) );
  AOI22_X1 U22796 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n19990), .ZN(n19809) );
  OAI211_X1 U22797 ( .C1(n19993), .C2(n19844), .A(n19810), .B(n19809), .ZN(
        P2_U3109) );
  AOI22_X1 U22798 ( .A1(n19814), .A2(n20090), .B1(n20089), .B2(n19828), .ZN(
        n19812) );
  AOI22_X1 U22799 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19816), .B1(
        n19848), .B2(n20091), .ZN(n19811) );
  OAI211_X1 U22800 ( .C1(n20096), .C2(n19813), .A(n19812), .B(n19811), .ZN(
        P2_U3110) );
  AOI22_X1 U22801 ( .A1(n19814), .A2(n20099), .B1(n20097), .B2(n19828), .ZN(
        n19818) );
  AOI22_X1 U22802 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19816), .B1(
        n19815), .B2(n20101), .ZN(n19817) );
  OAI211_X1 U22803 ( .C1(n20107), .C2(n19844), .A(n19818), .B(n19817), .ZN(
        P2_U3111) );
  NOR2_X1 U22804 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20209), .ZN(
        n19921) );
  NAND2_X1 U22805 ( .A1(n19921), .A2(n20229), .ZN(n19860) );
  NOR2_X1 U22806 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19860), .ZN(
        n19847) );
  AOI22_X1 U22807 ( .A1(n19848), .A2(n20055), .B1(n20046), .B2(n19847), .ZN(
        n19833) );
  NAND3_X1 U22808 ( .A1(n19886), .A2(n20196), .A3(n19844), .ZN(n19822) );
  AND2_X1 U22809 ( .A1(n20196), .A2(n19820), .ZN(n20199) );
  INV_X1 U22810 ( .A(n20199), .ZN(n19821) );
  NAND2_X1 U22811 ( .A1(n19822), .A2(n19821), .ZN(n19827) );
  INV_X1 U22812 ( .A(n19823), .ZN(n19829) );
  AOI21_X1 U22813 ( .B1(n19829), .B2(n20205), .A(n20196), .ZN(n19824) );
  AOI21_X1 U22814 ( .B1(n19827), .B2(n19825), .A(n19824), .ZN(n19826) );
  OAI21_X1 U22815 ( .B1(n19847), .B2(n19828), .A(n19827), .ZN(n19831) );
  OAI21_X1 U22816 ( .B1(n19829), .B2(n19847), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19830) );
  NAND2_X1 U22817 ( .A1(n19831), .A2(n19830), .ZN(n19849) );
  AOI22_X1 U22818 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19850), .B1(
        n20047), .B2(n19849), .ZN(n19832) );
  OAI211_X1 U22819 ( .C1(n20058), .C2(n19886), .A(n19833), .B(n19832), .ZN(
        P2_U3112) );
  INV_X1 U22820 ( .A(n19886), .ZN(n19879) );
  AOI22_X1 U22821 ( .A1(n19879), .A2(n20061), .B1(n20059), .B2(n19847), .ZN(
        n19835) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20060), .ZN(n19834) );
  OAI211_X1 U22823 ( .C1(n20064), .C2(n19844), .A(n19835), .B(n19834), .ZN(
        P2_U3113) );
  AOI22_X1 U22824 ( .A1(n19879), .A2(n20067), .B1(n20065), .B2(n19847), .ZN(
        n19837) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20066), .ZN(n19836) );
  OAI211_X1 U22826 ( .C1(n20070), .C2(n19844), .A(n19837), .B(n19836), .ZN(
        P2_U3114) );
  AOI22_X1 U22827 ( .A1(n19848), .A2(n20073), .B1(n20071), .B2(n19847), .ZN(
        n19839) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20072), .ZN(n19838) );
  OAI211_X1 U22829 ( .C1(n20076), .C2(n19886), .A(n19839), .B(n19838), .ZN(
        P2_U3115) );
  AOI22_X1 U22830 ( .A1(n19879), .A2(n20079), .B1(n20077), .B2(n19847), .ZN(
        n19841) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20078), .ZN(n19840) );
  OAI211_X1 U22832 ( .C1(n20082), .C2(n19844), .A(n19841), .B(n19840), .ZN(
        P2_U3116) );
  AOI22_X1 U22833 ( .A1(n19879), .A2(n20085), .B1(n20083), .B2(n19847), .ZN(
        n19843) );
  AOI22_X1 U22834 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20084), .ZN(n19842) );
  OAI211_X1 U22835 ( .C1(n20088), .C2(n19844), .A(n19843), .B(n19842), .ZN(
        P2_U3117) );
  AOI22_X1 U22836 ( .A1(n19848), .A2(n19994), .B1(n20089), .B2(n19847), .ZN(
        n19846) );
  AOI22_X1 U22837 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20090), .ZN(n19845) );
  OAI211_X1 U22838 ( .C1(n19997), .C2(n19886), .A(n19846), .B(n19845), .ZN(
        P2_U3118) );
  AOI22_X1 U22839 ( .A1(n19848), .A2(n20101), .B1(n20097), .B2(n19847), .ZN(
        n19852) );
  AOI22_X1 U22840 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19850), .B1(
        n19849), .B2(n20099), .ZN(n19851) );
  OAI211_X1 U22841 ( .C1(n20107), .C2(n19886), .A(n19852), .B(n19851), .ZN(
        P2_U3119) );
  INV_X1 U22842 ( .A(n19921), .ZN(n19918) );
  NOR2_X1 U22843 ( .A1(n19853), .A2(n19918), .ZN(n19893) );
  AOI22_X1 U22844 ( .A1(n19879), .A2(n20055), .B1(n20046), .B2(n19893), .ZN(
        n19863) );
  NAND2_X1 U22845 ( .A1(n19854), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20050) );
  OAI21_X1 U22846 ( .B1(n20050), .B2(n19855), .A(n20196), .ZN(n19861) );
  INV_X1 U22847 ( .A(n19860), .ZN(n19857) );
  INV_X1 U22848 ( .A(n19893), .ZN(n19872) );
  OAI211_X1 U22849 ( .C1(n11446), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20202), 
        .B(n19872), .ZN(n19856) );
  OAI211_X1 U22850 ( .C1(n19861), .C2(n19857), .A(n20053), .B(n19856), .ZN(
        n19883) );
  INV_X1 U22851 ( .A(n11446), .ZN(n19858) );
  OAI21_X1 U22852 ( .B1(n19858), .B2(n19893), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19859) );
  OAI21_X1 U22853 ( .B1(n19861), .B2(n19860), .A(n19859), .ZN(n19882) );
  AOI22_X1 U22854 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19883), .B1(
        n20047), .B2(n19882), .ZN(n19862) );
  OAI211_X1 U22855 ( .C1(n20058), .C2(n19891), .A(n19863), .B(n19862), .ZN(
        P2_U3120) );
  OAI22_X1 U22856 ( .A1(n19886), .A2(n20064), .B1(n19864), .B2(n19872), .ZN(
        n19865) );
  INV_X1 U22857 ( .A(n19865), .ZN(n19867) );
  AOI22_X1 U22858 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19883), .B1(
        n20060), .B2(n19882), .ZN(n19866) );
  OAI211_X1 U22859 ( .C1(n20018), .C2(n19891), .A(n19867), .B(n19866), .ZN(
        P2_U3121) );
  AOI22_X1 U22860 ( .A1(n19913), .A2(n20067), .B1(n20065), .B2(n19893), .ZN(
        n19869) );
  AOI22_X1 U22861 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19883), .B1(
        n20066), .B2(n19882), .ZN(n19868) );
  OAI211_X1 U22862 ( .C1(n20070), .C2(n19886), .A(n19869), .B(n19868), .ZN(
        P2_U3122) );
  AOI22_X1 U22863 ( .A1(n19879), .A2(n20073), .B1(n20071), .B2(n19893), .ZN(
        n19871) );
  AOI22_X1 U22864 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19883), .B1(
        n20072), .B2(n19882), .ZN(n19870) );
  OAI211_X1 U22865 ( .C1(n20076), .C2(n19891), .A(n19871), .B(n19870), .ZN(
        P2_U3123) );
  OAI22_X1 U22866 ( .A1(n19886), .A2(n20082), .B1(n19873), .B2(n19872), .ZN(
        n19874) );
  INV_X1 U22867 ( .A(n19874), .ZN(n19876) );
  AOI22_X1 U22868 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19883), .B1(
        n20078), .B2(n19882), .ZN(n19875) );
  OAI211_X1 U22869 ( .C1(n20029), .C2(n19891), .A(n19876), .B(n19875), .ZN(
        P2_U3124) );
  AOI22_X1 U22870 ( .A1(n19879), .A2(n19990), .B1(n20083), .B2(n19893), .ZN(
        n19878) );
  AOI22_X1 U22871 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19883), .B1(
        n20084), .B2(n19882), .ZN(n19877) );
  OAI211_X1 U22872 ( .C1(n19993), .C2(n19891), .A(n19878), .B(n19877), .ZN(
        P2_U3125) );
  AOI22_X1 U22873 ( .A1(n19879), .A2(n19994), .B1(n20089), .B2(n19893), .ZN(
        n19881) );
  AOI22_X1 U22874 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19883), .B1(
        n20090), .B2(n19882), .ZN(n19880) );
  OAI211_X1 U22875 ( .C1(n19997), .C2(n19891), .A(n19881), .B(n19880), .ZN(
        P2_U3126) );
  AOI22_X1 U22876 ( .A1(n19913), .A2(n20035), .B1(n20097), .B2(n19893), .ZN(
        n19885) );
  AOI22_X1 U22877 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19883), .B1(
        n20099), .B2(n19882), .ZN(n19884) );
  OAI211_X1 U22878 ( .C1(n20041), .C2(n19886), .A(n19885), .B(n19884), .ZN(
        P2_U3127) );
  AND2_X1 U22879 ( .A1(n19887), .A2(n19921), .ZN(n19911) );
  OAI21_X1 U22880 ( .B1(n19888), .B2(n19911), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19889) );
  OAI21_X1 U22881 ( .B1(n19918), .B2(n19890), .A(n19889), .ZN(n19912) );
  AOI22_X1 U22882 ( .A1(n19912), .A2(n20047), .B1(n20046), .B2(n19911), .ZN(
        n19898) );
  AOI21_X1 U22883 ( .B1(n19948), .B2(n19891), .A(n19820), .ZN(n19892) );
  OAI21_X1 U22884 ( .B1(n19893), .B2(n19892), .A(n20205), .ZN(n19894) );
  AOI21_X1 U22885 ( .B1(n19895), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19894), 
        .ZN(n19896) );
  AOI22_X1 U22886 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19914), .B1(
        n19913), .B2(n20055), .ZN(n19897) );
  OAI211_X1 U22887 ( .C1(n20058), .C2(n19948), .A(n19898), .B(n19897), .ZN(
        P2_U3128) );
  AOI22_X1 U22888 ( .A1(n19912), .A2(n20060), .B1(n20059), .B2(n19911), .ZN(
        n19900) );
  AOI22_X1 U22889 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19914), .B1(
        n19913), .B2(n20015), .ZN(n19899) );
  OAI211_X1 U22890 ( .C1(n20018), .C2(n19948), .A(n19900), .B(n19899), .ZN(
        P2_U3129) );
  AOI22_X1 U22891 ( .A1(n19912), .A2(n20066), .B1(n20065), .B2(n19911), .ZN(
        n19902) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19914), .B1(
        n19913), .B2(n19982), .ZN(n19901) );
  OAI211_X1 U22893 ( .C1(n19985), .C2(n19948), .A(n19902), .B(n19901), .ZN(
        P2_U3130) );
  AOI22_X1 U22894 ( .A1(n19912), .A2(n20072), .B1(n20071), .B2(n19911), .ZN(
        n19904) );
  AOI22_X1 U22895 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19914), .B1(
        n19913), .B2(n20073), .ZN(n19903) );
  OAI211_X1 U22896 ( .C1(n20076), .C2(n19948), .A(n19904), .B(n19903), .ZN(
        P2_U3131) );
  AOI22_X1 U22897 ( .A1(n19912), .A2(n20078), .B1(n20077), .B2(n19911), .ZN(
        n19906) );
  AOI22_X1 U22898 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19914), .B1(
        n19913), .B2(n20025), .ZN(n19905) );
  OAI211_X1 U22899 ( .C1(n20029), .C2(n19948), .A(n19906), .B(n19905), .ZN(
        P2_U3132) );
  AOI22_X1 U22900 ( .A1(n19912), .A2(n20084), .B1(n20083), .B2(n19911), .ZN(
        n19908) );
  AOI22_X1 U22901 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19914), .B1(
        n19913), .B2(n19990), .ZN(n19907) );
  OAI211_X1 U22902 ( .C1(n19993), .C2(n19948), .A(n19908), .B(n19907), .ZN(
        P2_U3133) );
  AOI22_X1 U22903 ( .A1(n19912), .A2(n20090), .B1(n20089), .B2(n19911), .ZN(
        n19910) );
  AOI22_X1 U22904 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19914), .B1(
        n19913), .B2(n19994), .ZN(n19909) );
  OAI211_X1 U22905 ( .C1(n19997), .C2(n19948), .A(n19910), .B(n19909), .ZN(
        P2_U3134) );
  AOI22_X1 U22906 ( .A1(n19912), .A2(n20099), .B1(n20097), .B2(n19911), .ZN(
        n19916) );
  AOI22_X1 U22907 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19914), .B1(
        n19913), .B2(n20101), .ZN(n19915) );
  OAI211_X1 U22908 ( .C1(n20107), .C2(n19948), .A(n19916), .B(n19915), .ZN(
        P2_U3135) );
  INV_X1 U22909 ( .A(n19965), .ZN(n19942) );
  NOR2_X1 U22910 ( .A1(n19918), .A2(n19917), .ZN(n19943) );
  NOR2_X1 U22911 ( .A1(n19943), .A2(n19761), .ZN(n19919) );
  NAND2_X1 U22912 ( .A1(n19920), .A2(n19919), .ZN(n19924) );
  NAND2_X1 U22913 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19921), .ZN(
        n19923) );
  OAI21_X1 U22914 ( .B1(n19923), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19761), 
        .ZN(n19922) );
  AOI22_X1 U22915 ( .A1(n19944), .A2(n20047), .B1(n20046), .B2(n19943), .ZN(
        n19928) );
  OAI21_X1 U22916 ( .B1(n20050), .B2(n20197), .A(n19923), .ZN(n19925) );
  AND2_X1 U22917 ( .A1(n19925), .A2(n19924), .ZN(n19926) );
  OAI211_X1 U22918 ( .C1(n19943), .C2(n20205), .A(n19926), .B(n20053), .ZN(
        n19945) );
  AOI22_X1 U22919 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19945), .B1(
        n19939), .B2(n20055), .ZN(n19927) );
  OAI211_X1 U22920 ( .C1(n20058), .C2(n19942), .A(n19928), .B(n19927), .ZN(
        P2_U3136) );
  AOI22_X1 U22921 ( .A1(n19944), .A2(n20060), .B1(n20059), .B2(n19943), .ZN(
        n19930) );
  AOI22_X1 U22922 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19945), .B1(
        n19965), .B2(n20061), .ZN(n19929) );
  OAI211_X1 U22923 ( .C1(n20064), .C2(n19948), .A(n19930), .B(n19929), .ZN(
        P2_U3137) );
  AOI22_X1 U22924 ( .A1(n19944), .A2(n20066), .B1(n20065), .B2(n19943), .ZN(
        n19932) );
  AOI22_X1 U22925 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19945), .B1(
        n19939), .B2(n19982), .ZN(n19931) );
  OAI211_X1 U22926 ( .C1(n19985), .C2(n19942), .A(n19932), .B(n19931), .ZN(
        P2_U3138) );
  AOI22_X1 U22927 ( .A1(n19944), .A2(n20072), .B1(n20071), .B2(n19943), .ZN(
        n19934) );
  AOI22_X1 U22928 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19945), .B1(
        n19965), .B2(n20021), .ZN(n19933) );
  OAI211_X1 U22929 ( .C1(n20024), .C2(n19948), .A(n19934), .B(n19933), .ZN(
        P2_U3139) );
  AOI22_X1 U22930 ( .A1(n19944), .A2(n20078), .B1(n20077), .B2(n19943), .ZN(
        n19936) );
  AOI22_X1 U22931 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19945), .B1(
        n19965), .B2(n20079), .ZN(n19935) );
  OAI211_X1 U22932 ( .C1(n20082), .C2(n19948), .A(n19936), .B(n19935), .ZN(
        P2_U3140) );
  AOI22_X1 U22933 ( .A1(n19944), .A2(n20084), .B1(n20083), .B2(n19943), .ZN(
        n19938) );
  AOI22_X1 U22934 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19945), .B1(
        n19965), .B2(n20085), .ZN(n19937) );
  OAI211_X1 U22935 ( .C1(n20088), .C2(n19948), .A(n19938), .B(n19937), .ZN(
        P2_U3141) );
  AOI22_X1 U22936 ( .A1(n19944), .A2(n20090), .B1(n20089), .B2(n19943), .ZN(
        n19941) );
  AOI22_X1 U22937 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19945), .B1(
        n19939), .B2(n19994), .ZN(n19940) );
  OAI211_X1 U22938 ( .C1(n19997), .C2(n19942), .A(n19941), .B(n19940), .ZN(
        P2_U3142) );
  AOI22_X1 U22939 ( .A1(n19944), .A2(n20099), .B1(n20097), .B2(n19943), .ZN(
        n19947) );
  AOI22_X1 U22940 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19945), .B1(
        n19965), .B2(n20035), .ZN(n19946) );
  OAI211_X1 U22941 ( .C1(n20041), .C2(n19948), .A(n19947), .B(n19946), .ZN(
        P2_U3143) );
  AOI22_X1 U22942 ( .A1(n19964), .A2(n20060), .B1(n19963), .B2(n20059), .ZN(
        n19950) );
  AOI22_X1 U22943 ( .A1(n19999), .A2(n20061), .B1(n19965), .B2(n20015), .ZN(
        n19949) );
  OAI211_X1 U22944 ( .C1(n19969), .C2(n11402), .A(n19950), .B(n19949), .ZN(
        P2_U3145) );
  INV_X1 U22945 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n19953) );
  AOI22_X1 U22946 ( .A1(n19964), .A2(n20066), .B1(n19963), .B2(n20065), .ZN(
        n19952) );
  AOI22_X1 U22947 ( .A1(n19999), .A2(n20067), .B1(n19965), .B2(n19982), .ZN(
        n19951) );
  OAI211_X1 U22948 ( .C1(n19969), .C2(n19953), .A(n19952), .B(n19951), .ZN(
        P2_U3146) );
  AOI22_X1 U22949 ( .A1(n19964), .A2(n20072), .B1(n19963), .B2(n20071), .ZN(
        n19955) );
  AOI22_X1 U22950 ( .A1(n19965), .A2(n20073), .B1(n19999), .B2(n20021), .ZN(
        n19954) );
  OAI211_X1 U22951 ( .C1(n19969), .C2(n11345), .A(n19955), .B(n19954), .ZN(
        P2_U3147) );
  INV_X1 U22952 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n19958) );
  AOI22_X1 U22953 ( .A1(n19964), .A2(n20078), .B1(n19963), .B2(n20077), .ZN(
        n19957) );
  AOI22_X1 U22954 ( .A1(n19999), .A2(n20079), .B1(n19965), .B2(n20025), .ZN(
        n19956) );
  OAI211_X1 U22955 ( .C1(n19969), .C2(n19958), .A(n19957), .B(n19956), .ZN(
        P2_U3148) );
  AOI22_X1 U22956 ( .A1(n19964), .A2(n20084), .B1(n19963), .B2(n20083), .ZN(
        n19960) );
  AOI22_X1 U22957 ( .A1(n19999), .A2(n20085), .B1(n19965), .B2(n19990), .ZN(
        n19959) );
  OAI211_X1 U22958 ( .C1(n19969), .C2(n11445), .A(n19960), .B(n19959), .ZN(
        P2_U3149) );
  AOI22_X1 U22959 ( .A1(n19964), .A2(n20090), .B1(n19963), .B2(n20089), .ZN(
        n19962) );
  AOI22_X1 U22960 ( .A1(n19965), .A2(n19994), .B1(n19999), .B2(n20091), .ZN(
        n19961) );
  OAI211_X1 U22961 ( .C1(n19969), .C2(n11486), .A(n19962), .B(n19961), .ZN(
        P2_U3150) );
  INV_X1 U22962 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n19968) );
  AOI22_X1 U22963 ( .A1(n19964), .A2(n20099), .B1(n19963), .B2(n20097), .ZN(
        n19967) );
  AOI22_X1 U22964 ( .A1(n19965), .A2(n20101), .B1(n19999), .B2(n20035), .ZN(
        n19966) );
  OAI211_X1 U22965 ( .C1(n19969), .C2(n19968), .A(n19967), .B(n19966), .ZN(
        P2_U3151) );
  INV_X1 U22966 ( .A(n11450), .ZN(n19971) );
  NOR2_X1 U22967 ( .A1(n20239), .A2(n19973), .ZN(n20005) );
  OAI21_X1 U22968 ( .B1(n19971), .B2(n20005), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19972) );
  OAI21_X1 U22969 ( .B1(n19973), .B2(n20202), .A(n19972), .ZN(n19998) );
  AOI22_X1 U22970 ( .A1(n19998), .A2(n20047), .B1(n20046), .B2(n20005), .ZN(
        n19979) );
  OAI21_X1 U22971 ( .B1(n20050), .B2(n19974), .A(n19973), .ZN(n19977) );
  INV_X1 U22972 ( .A(n20005), .ZN(n19975) );
  OAI211_X1 U22973 ( .C1(n11450), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20202), 
        .B(n19975), .ZN(n19976) );
  NAND3_X1 U22974 ( .A1(n19977), .A2(n20053), .A3(n19976), .ZN(n20000) );
  AOI22_X1 U22975 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n20055), .ZN(n19978) );
  OAI211_X1 U22976 ( .C1(n20058), .C2(n20040), .A(n19979), .B(n19978), .ZN(
        P2_U3152) );
  AOI22_X1 U22977 ( .A1(n19998), .A2(n20060), .B1(n20059), .B2(n20005), .ZN(
        n19981) );
  AOI22_X1 U22978 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n20015), .ZN(n19980) );
  OAI211_X1 U22979 ( .C1(n20018), .C2(n20040), .A(n19981), .B(n19980), .ZN(
        P2_U3153) );
  AOI22_X1 U22980 ( .A1(n19998), .A2(n20066), .B1(n20065), .B2(n20005), .ZN(
        n19984) );
  AOI22_X1 U22981 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n19982), .ZN(n19983) );
  OAI211_X1 U22982 ( .C1(n19985), .C2(n20040), .A(n19984), .B(n19983), .ZN(
        P2_U3154) );
  AOI22_X1 U22983 ( .A1(n19998), .A2(n20072), .B1(n20071), .B2(n20005), .ZN(
        n19987) );
  AOI22_X1 U22984 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n20073), .ZN(n19986) );
  OAI211_X1 U22985 ( .C1(n20076), .C2(n20040), .A(n19987), .B(n19986), .ZN(
        P2_U3155) );
  AOI22_X1 U22986 ( .A1(n19998), .A2(n20078), .B1(n20077), .B2(n20005), .ZN(
        n19989) );
  AOI22_X1 U22987 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n20025), .ZN(n19988) );
  OAI211_X1 U22988 ( .C1(n20029), .C2(n20040), .A(n19989), .B(n19988), .ZN(
        P2_U3156) );
  AOI22_X1 U22989 ( .A1(n19998), .A2(n20084), .B1(n20083), .B2(n20005), .ZN(
        n19992) );
  AOI22_X1 U22990 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n19990), .ZN(n19991) );
  OAI211_X1 U22991 ( .C1(n19993), .C2(n20040), .A(n19992), .B(n19991), .ZN(
        P2_U3157) );
  AOI22_X1 U22992 ( .A1(n19998), .A2(n20090), .B1(n20089), .B2(n20005), .ZN(
        n19996) );
  AOI22_X1 U22993 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n19994), .ZN(n19995) );
  OAI211_X1 U22994 ( .C1(n19997), .C2(n20040), .A(n19996), .B(n19995), .ZN(
        P2_U3158) );
  AOI22_X1 U22995 ( .A1(n19998), .A2(n20099), .B1(n20097), .B2(n20005), .ZN(
        n20002) );
  AOI22_X1 U22996 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20000), .B1(
        n19999), .B2(n20101), .ZN(n20001) );
  OAI211_X1 U22997 ( .C1(n20107), .C2(n20040), .A(n20002), .B(n20001), .ZN(
        P2_U3159) );
  NOR3_X2 U22998 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20209), .A3(
        n20048), .ZN(n20034) );
  AOI22_X1 U22999 ( .A1(n20026), .A2(n20055), .B1(n20046), .B2(n20034), .ZN(
        n20014) );
  NOR3_X1 U23000 ( .A1(n20026), .A2(n20102), .A3(n20202), .ZN(n20004) );
  NOR2_X1 U23001 ( .A1(n20004), .A2(n20199), .ZN(n20012) );
  NOR2_X1 U23002 ( .A1(n20034), .A2(n20005), .ZN(n20011) );
  INV_X1 U23003 ( .A(n20011), .ZN(n20008) );
  INV_X1 U23004 ( .A(n20034), .ZN(n20006) );
  OAI211_X1 U23005 ( .C1(n20009), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20202), 
        .B(n20006), .ZN(n20007) );
  OAI211_X1 U23006 ( .C1(n20012), .C2(n20008), .A(n20053), .B(n20007), .ZN(
        n20037) );
  OAI21_X1 U23007 ( .B1(n11373), .B2(n20034), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20010) );
  AOI22_X1 U23008 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20037), .B1(
        n20047), .B2(n20036), .ZN(n20013) );
  OAI211_X1 U23009 ( .C1(n20058), .C2(n20095), .A(n20014), .B(n20013), .ZN(
        P2_U3160) );
  AOI22_X1 U23010 ( .A1(n20026), .A2(n20015), .B1(n20059), .B2(n20034), .ZN(
        n20017) );
  AOI22_X1 U23011 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20037), .B1(
        n20060), .B2(n20036), .ZN(n20016) );
  OAI211_X1 U23012 ( .C1(n20018), .C2(n20095), .A(n20017), .B(n20016), .ZN(
        P2_U3161) );
  AOI22_X1 U23013 ( .A1(n20102), .A2(n20067), .B1(n20065), .B2(n20034), .ZN(
        n20020) );
  AOI22_X1 U23014 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20037), .B1(
        n20066), .B2(n20036), .ZN(n20019) );
  OAI211_X1 U23015 ( .C1(n20070), .C2(n20040), .A(n20020), .B(n20019), .ZN(
        P2_U3162) );
  AOI22_X1 U23016 ( .A1(n20102), .A2(n20021), .B1(n20071), .B2(n20034), .ZN(
        n20023) );
  AOI22_X1 U23017 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20037), .B1(
        n20072), .B2(n20036), .ZN(n20022) );
  OAI211_X1 U23018 ( .C1(n20024), .C2(n20040), .A(n20023), .B(n20022), .ZN(
        P2_U3163) );
  AOI22_X1 U23019 ( .A1(n20026), .A2(n20025), .B1(n20077), .B2(n20034), .ZN(
        n20028) );
  AOI22_X1 U23020 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20037), .B1(
        n20078), .B2(n20036), .ZN(n20027) );
  OAI211_X1 U23021 ( .C1(n20029), .C2(n20095), .A(n20028), .B(n20027), .ZN(
        P2_U3164) );
  AOI22_X1 U23022 ( .A1(n20102), .A2(n20085), .B1(n20083), .B2(n20034), .ZN(
        n20031) );
  AOI22_X1 U23023 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20037), .B1(
        n20084), .B2(n20036), .ZN(n20030) );
  OAI211_X1 U23024 ( .C1(n20088), .C2(n20040), .A(n20031), .B(n20030), .ZN(
        P2_U3165) );
  AOI22_X1 U23025 ( .A1(n20102), .A2(n20091), .B1(n20089), .B2(n20034), .ZN(
        n20033) );
  AOI22_X1 U23026 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20037), .B1(
        n20090), .B2(n20036), .ZN(n20032) );
  OAI211_X1 U23027 ( .C1(n20096), .C2(n20040), .A(n20033), .B(n20032), .ZN(
        P2_U3166) );
  AOI22_X1 U23028 ( .A1(n20102), .A2(n20035), .B1(n20097), .B2(n20034), .ZN(
        n20039) );
  AOI22_X1 U23029 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20037), .B1(
        n20099), .B2(n20036), .ZN(n20038) );
  OAI211_X1 U23030 ( .C1(n20041), .C2(n20040), .A(n20039), .B(n20038), .ZN(
        P2_U3167) );
  NAND2_X1 U23031 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20042), .ZN(
        n20045) );
  INV_X1 U23032 ( .A(n11447), .ZN(n20043) );
  OAI21_X1 U23033 ( .B1(n20043), .B2(n20098), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20044) );
  OAI21_X1 U23034 ( .B1(n20045), .B2(n20202), .A(n20044), .ZN(n20100) );
  AOI22_X1 U23035 ( .A1(n20100), .A2(n20047), .B1(n20098), .B2(n20046), .ZN(
        n20057) );
  OAI22_X1 U23036 ( .A1(n20050), .A2(n20049), .B1(n20048), .B2(n20209), .ZN(
        n20054) );
  OAI211_X1 U23037 ( .C1(n11447), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20202), 
        .B(n20051), .ZN(n20052) );
  NAND3_X1 U23038 ( .A1(n20054), .A2(n20053), .A3(n20052), .ZN(n20103) );
  AOI22_X1 U23039 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20103), .B1(
        n20102), .B2(n20055), .ZN(n20056) );
  OAI211_X1 U23040 ( .C1(n20058), .C2(n20106), .A(n20057), .B(n20056), .ZN(
        P2_U3168) );
  AOI22_X1 U23041 ( .A1(n20100), .A2(n20060), .B1(n20098), .B2(n20059), .ZN(
        n20063) );
  AOI22_X1 U23042 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20103), .B1(
        n20092), .B2(n20061), .ZN(n20062) );
  OAI211_X1 U23043 ( .C1(n20064), .C2(n20095), .A(n20063), .B(n20062), .ZN(
        P2_U3169) );
  AOI22_X1 U23044 ( .A1(n20100), .A2(n20066), .B1(n20098), .B2(n20065), .ZN(
        n20069) );
  AOI22_X1 U23045 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20103), .B1(
        n20092), .B2(n20067), .ZN(n20068) );
  OAI211_X1 U23046 ( .C1(n20070), .C2(n20095), .A(n20069), .B(n20068), .ZN(
        P2_U3170) );
  AOI22_X1 U23047 ( .A1(n20100), .A2(n20072), .B1(n20098), .B2(n20071), .ZN(
        n20075) );
  AOI22_X1 U23048 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20103), .B1(
        n20102), .B2(n20073), .ZN(n20074) );
  OAI211_X1 U23049 ( .C1(n20076), .C2(n20106), .A(n20075), .B(n20074), .ZN(
        P2_U3171) );
  AOI22_X1 U23050 ( .A1(n20100), .A2(n20078), .B1(n20098), .B2(n20077), .ZN(
        n20081) );
  AOI22_X1 U23051 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20103), .B1(
        n20092), .B2(n20079), .ZN(n20080) );
  OAI211_X1 U23052 ( .C1(n20082), .C2(n20095), .A(n20081), .B(n20080), .ZN(
        P2_U3172) );
  AOI22_X1 U23053 ( .A1(n20100), .A2(n20084), .B1(n20098), .B2(n20083), .ZN(
        n20087) );
  AOI22_X1 U23054 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20103), .B1(
        n20092), .B2(n20085), .ZN(n20086) );
  OAI211_X1 U23055 ( .C1(n20088), .C2(n20095), .A(n20087), .B(n20086), .ZN(
        P2_U3173) );
  AOI22_X1 U23056 ( .A1(n20100), .A2(n20090), .B1(n20098), .B2(n20089), .ZN(
        n20094) );
  AOI22_X1 U23057 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20103), .B1(
        n20092), .B2(n20091), .ZN(n20093) );
  OAI211_X1 U23058 ( .C1(n20096), .C2(n20095), .A(n20094), .B(n20093), .ZN(
        P2_U3174) );
  AOI22_X1 U23059 ( .A1(n20100), .A2(n20099), .B1(n20098), .B2(n20097), .ZN(
        n20105) );
  AOI22_X1 U23060 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20103), .B1(
        n20102), .B2(n20101), .ZN(n20104) );
  OAI211_X1 U23061 ( .C1(n20107), .C2(n20106), .A(n20105), .B(n20104), .ZN(
        P2_U3175) );
  AOI21_X1 U23062 ( .B1(n20110), .B2(n20109), .A(n20108), .ZN(n20114) );
  OAI221_X1 U23063 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20205), .C1(
        P2_STATE2_REG_2__SCAN_IN), .C2(n20257), .A(n20111), .ZN(n20112) );
  OAI22_X1 U23064 ( .A1(n20114), .A2(n10598), .B1(n20113), .B2(n20112), .ZN(
        P2_U3177) );
  AND2_X1 U23065 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20115), .ZN(
        P2_U3179) );
  AND2_X1 U23066 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20115), .ZN(
        P2_U3180) );
  AND2_X1 U23067 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20115), .ZN(
        P2_U3181) );
  AND2_X1 U23068 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20115), .ZN(
        P2_U3182) );
  AND2_X1 U23069 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20115), .ZN(
        P2_U3183) );
  AND2_X1 U23070 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20115), .ZN(
        P2_U3184) );
  AND2_X1 U23071 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20115), .ZN(
        P2_U3185) );
  AND2_X1 U23072 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20115), .ZN(
        P2_U3186) );
  AND2_X1 U23073 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20115), .ZN(
        P2_U3187) );
  AND2_X1 U23074 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20115), .ZN(
        P2_U3188) );
  AND2_X1 U23075 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20115), .ZN(
        P2_U3189) );
  AND2_X1 U23076 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20115), .ZN(
        P2_U3190) );
  AND2_X1 U23077 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20115), .ZN(
        P2_U3191) );
  AND2_X1 U23078 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20115), .ZN(
        P2_U3192) );
  AND2_X1 U23079 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20115), .ZN(
        P2_U3193) );
  AND2_X1 U23080 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20115), .ZN(
        P2_U3194) );
  AND2_X1 U23081 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20115), .ZN(
        P2_U3195) );
  AND2_X1 U23082 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20115), .ZN(
        P2_U3196) );
  AND2_X1 U23083 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20115), .ZN(
        P2_U3197) );
  AND2_X1 U23084 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20115), .ZN(
        P2_U3198) );
  AND2_X1 U23085 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20115), .ZN(
        P2_U3199) );
  AND2_X1 U23086 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20115), .ZN(
        P2_U3200) );
  AND2_X1 U23087 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20115), .ZN(P2_U3201) );
  AND2_X1 U23088 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20115), .ZN(P2_U3202) );
  AND2_X1 U23089 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20115), .ZN(P2_U3203) );
  AND2_X1 U23090 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20115), .ZN(P2_U3204) );
  AND2_X1 U23091 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20115), .ZN(P2_U3205) );
  AND2_X1 U23092 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20115), .ZN(P2_U3206) );
  AND2_X1 U23093 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20115), .ZN(P2_U3207) );
  AND2_X1 U23094 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20115), .ZN(P2_U3208) );
  NAND2_X1 U23095 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20128), .ZN(n20122) );
  NAND3_X1 U23096 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20122), .ZN(n20116) );
  NOR3_X1 U23097 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21230), .ZN(n20130) );
  AOI21_X1 U23098 ( .B1(n20133), .B2(n20116), .A(n20130), .ZN(n20117) );
  OAI221_X1 U23099 ( .B1(n20118), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20118), .C2(n21190), .A(n20117), .ZN(P2_U3209) );
  AOI21_X1 U23100 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21190), .A(n20133), 
        .ZN(n20126) );
  INV_X1 U23101 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20270) );
  NOR3_X1 U23102 ( .A1(n20126), .A2(n20270), .A3(n19235), .ZN(n20119) );
  NOR2_X1 U23103 ( .A1(n20119), .A2(n20262), .ZN(n20120) );
  OAI211_X1 U23104 ( .C1(n21190), .C2(n20121), .A(n20120), .B(n20122), .ZN(
        P2_U3210) );
  INV_X1 U23105 ( .A(n20122), .ZN(n20123) );
  AOI22_X1 U23106 ( .A1(n20124), .A2(n20270), .B1(n20123), .B2(n21230), .ZN(
        n20132) );
  OAI21_X1 U23107 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20131) );
  NOR2_X1 U23108 ( .A1(n20125), .A2(n20133), .ZN(n20127) );
  AOI21_X1 U23109 ( .B1(n20128), .B2(n20127), .A(n20126), .ZN(n20129) );
  OAI22_X1 U23110 ( .A1(n20132), .A2(n20131), .B1(n20130), .B2(n20129), .ZN(
        P2_U3211) );
  OAI222_X1 U23111 ( .A1(n20176), .A2(n10535), .B1(n20134), .B2(n20274), .C1(
        n10459), .C2(n20173), .ZN(P2_U3212) );
  OAI222_X1 U23112 ( .A1(n20176), .A2(n20136), .B1(n20135), .B2(n20274), .C1(
        n10535), .C2(n20173), .ZN(P2_U3213) );
  OAI222_X1 U23113 ( .A1(n20176), .A2(n10760), .B1(n20137), .B2(n20274), .C1(
        n20136), .C2(n20173), .ZN(P2_U3214) );
  OAI222_X1 U23114 ( .A1(n20176), .A2(n10794), .B1(n20138), .B2(n20274), .C1(
        n10760), .C2(n20173), .ZN(P2_U3215) );
  OAI222_X1 U23115 ( .A1(n20176), .A2(n16058), .B1(n20139), .B2(n20274), .C1(
        n10794), .C2(n20173), .ZN(P2_U3216) );
  OAI222_X1 U23116 ( .A1(n20176), .A2(n10567), .B1(n20140), .B2(n20274), .C1(
        n16058), .C2(n20173), .ZN(P2_U3217) );
  OAI222_X1 U23117 ( .A1(n20176), .A2(n13912), .B1(n20141), .B2(n20274), .C1(
        n10567), .C2(n20173), .ZN(P2_U3218) );
  OAI222_X1 U23118 ( .A1(n20176), .A2(n10855), .B1(n20142), .B2(n20274), .C1(
        n13912), .C2(n20173), .ZN(P2_U3219) );
  OAI222_X1 U23119 ( .A1(n20176), .A2(n10577), .B1(n20143), .B2(n20274), .C1(
        n10855), .C2(n20173), .ZN(P2_U3220) );
  OAI222_X1 U23120 ( .A1(n20176), .A2(n10888), .B1(n20144), .B2(n20274), .C1(
        n10577), .C2(n20173), .ZN(P2_U3221) );
  OAI222_X1 U23121 ( .A1(n20176), .A2(n10585), .B1(n20145), .B2(n20274), .C1(
        n10888), .C2(n20173), .ZN(P2_U3222) );
  OAI222_X1 U23122 ( .A1(n20176), .A2(n10591), .B1(n20146), .B2(n20274), .C1(
        n10585), .C2(n20173), .ZN(P2_U3223) );
  OAI222_X1 U23123 ( .A1(n20176), .A2(n14045), .B1(n20147), .B2(n20274), .C1(
        n10591), .C2(n20173), .ZN(P2_U3224) );
  OAI222_X1 U23124 ( .A1(n20176), .A2(n10948), .B1(n20148), .B2(n20274), .C1(
        n14045), .C2(n20173), .ZN(P2_U3225) );
  OAI222_X1 U23125 ( .A1(n20176), .A2(n10952), .B1(n20149), .B2(n20274), .C1(
        n10948), .C2(n20173), .ZN(P2_U3226) );
  OAI222_X1 U23126 ( .A1(n20176), .A2(n20151), .B1(n20150), .B2(n20274), .C1(
        n10952), .C2(n20173), .ZN(P2_U3227) );
  OAI222_X1 U23127 ( .A1(n20176), .A2(n15696), .B1(n20152), .B2(n20274), .C1(
        n20151), .C2(n20173), .ZN(P2_U3228) );
  OAI222_X1 U23128 ( .A1(n20176), .A2(n20154), .B1(n20153), .B2(n20274), .C1(
        n15696), .C2(n20173), .ZN(P2_U3229) );
  OAI222_X1 U23129 ( .A1(n20176), .A2(n15674), .B1(n20155), .B2(n20274), .C1(
        n20154), .C2(n20173), .ZN(P2_U3230) );
  OAI222_X1 U23130 ( .A1(n20176), .A2(n20157), .B1(n20156), .B2(n20274), .C1(
        n15674), .C2(n20173), .ZN(P2_U3231) );
  OAI222_X1 U23131 ( .A1(n20176), .A2(n10965), .B1(n20158), .B2(n20274), .C1(
        n20157), .C2(n20173), .ZN(P2_U3232) );
  OAI222_X1 U23132 ( .A1(n20176), .A2(n20160), .B1(n20159), .B2(n20274), .C1(
        n10965), .C2(n20173), .ZN(P2_U3233) );
  OAI222_X1 U23133 ( .A1(n20176), .A2(n20162), .B1(n20161), .B2(n20274), .C1(
        n20160), .C2(n20173), .ZN(P2_U3234) );
  OAI222_X1 U23134 ( .A1(n20176), .A2(n20164), .B1(n20163), .B2(n20274), .C1(
        n20162), .C2(n20173), .ZN(P2_U3235) );
  OAI222_X1 U23135 ( .A1(n20176), .A2(n15615), .B1(n20165), .B2(n20274), .C1(
        n20164), .C2(n20173), .ZN(P2_U3236) );
  OAI222_X1 U23136 ( .A1(n20176), .A2(n20168), .B1(n20166), .B2(n20274), .C1(
        n15615), .C2(n20173), .ZN(P2_U3237) );
  OAI222_X1 U23137 ( .A1(n20173), .A2(n20168), .B1(n20167), .B2(n20274), .C1(
        n20169), .C2(n20176), .ZN(P2_U3238) );
  OAI222_X1 U23138 ( .A1(n20176), .A2(n20171), .B1(n20170), .B2(n20274), .C1(
        n20169), .C2(n20173), .ZN(P2_U3239) );
  OAI222_X1 U23139 ( .A1(n20176), .A2(n20174), .B1(n20172), .B2(n20274), .C1(
        n20171), .C2(n20173), .ZN(P2_U3240) );
  INV_X1 U23140 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20175) );
  OAI222_X1 U23141 ( .A1(n20176), .A2(n11698), .B1(n20175), .B2(n20274), .C1(
        n20174), .C2(n20173), .ZN(P2_U3241) );
  INV_X1 U23142 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20177) );
  AOI22_X1 U23143 ( .A1(n20274), .A2(n20178), .B1(n20177), .B2(n20271), .ZN(
        P2_U3585) );
  MUX2_X1 U23144 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20274), .Z(P2_U3586) );
  INV_X1 U23145 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20179) );
  AOI22_X1 U23146 ( .A1(n20274), .A2(n20180), .B1(n20179), .B2(n20271), .ZN(
        P2_U3587) );
  INV_X1 U23147 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20181) );
  AOI22_X1 U23148 ( .A1(n20274), .A2(n20182), .B1(n20181), .B2(n20271), .ZN(
        P2_U3588) );
  OAI21_X1 U23149 ( .B1(n20186), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20184), 
        .ZN(n20183) );
  INV_X1 U23150 ( .A(n20183), .ZN(P2_U3591) );
  OAI21_X1 U23151 ( .B1(n20186), .B2(n20185), .A(n20184), .ZN(P2_U3592) );
  INV_X1 U23152 ( .A(n20187), .ZN(n20189) );
  AOI222_X1 U23153 ( .A1(n20191), .A2(n20198), .B1(n20224), .B2(n20190), .C1(
        n20189), .C2(n20188), .ZN(n20193) );
  AOI22_X1 U23154 ( .A1(n20195), .A2(n20194), .B1(n20193), .B2(n20192), .ZN(
        P2_U3600) );
  INV_X1 U23155 ( .A(n20238), .ZN(n20237) );
  NAND2_X1 U23156 ( .A1(n20196), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20225) );
  NOR2_X1 U23157 ( .A1(n20197), .A2(n20225), .ZN(n20217) );
  NOR2_X1 U23158 ( .A1(n20199), .A2(n20198), .ZN(n20200) );
  OAI21_X1 U23159 ( .B1(n20224), .B2(n20202), .A(n20200), .ZN(n20211) );
  NOR2_X1 U23160 ( .A1(n20217), .A2(n20211), .ZN(n20203) );
  OAI222_X1 U23161 ( .A1(n20206), .A2(n20205), .B1(n20204), .B2(n20203), .C1(
        n20202), .C2(n20201), .ZN(n20207) );
  INV_X1 U23162 ( .A(n20207), .ZN(n20208) );
  AOI22_X1 U23163 ( .A1(n20237), .A2(n20209), .B1(n20208), .B2(n20238), .ZN(
        P2_U3602) );
  INV_X1 U23164 ( .A(n20210), .ZN(n20212) );
  NAND2_X1 U23165 ( .A1(n20212), .A2(n20211), .ZN(n20215) );
  OR2_X1 U23166 ( .A1(n20213), .A2(n20205), .ZN(n20214) );
  NAND2_X1 U23167 ( .A1(n20215), .A2(n20214), .ZN(n20216) );
  NOR2_X1 U23168 ( .A1(n20217), .A2(n20216), .ZN(n20218) );
  AOI22_X1 U23169 ( .A1(n20237), .A2(n20219), .B1(n20218), .B2(n20238), .ZN(
        P2_U3603) );
  INV_X1 U23170 ( .A(n20220), .ZN(n20233) );
  AND2_X1 U23171 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20221) );
  OR3_X1 U23172 ( .A1(n20222), .A2(n20233), .A3(n20221), .ZN(n20223) );
  OAI21_X1 U23173 ( .B1(n20225), .B2(n20224), .A(n20223), .ZN(n20226) );
  AOI21_X1 U23174 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20227), .A(n20226), 
        .ZN(n20228) );
  AOI22_X1 U23175 ( .A1(n20237), .A2(n20229), .B1(n20228), .B2(n20238), .ZN(
        P2_U3604) );
  INV_X1 U23176 ( .A(n20230), .ZN(n20232) );
  OAI22_X1 U23177 ( .A1(n20234), .A2(n20233), .B1(n20232), .B2(n20231), .ZN(
        n20235) );
  AOI21_X1 U23178 ( .B1(n20239), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20235), 
        .ZN(n20236) );
  OAI22_X1 U23179 ( .A1(n20239), .A2(n20238), .B1(n20237), .B2(n20236), .ZN(
        P2_U3605) );
  INV_X1 U23180 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20240) );
  AOI22_X1 U23181 ( .A1(n20274), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20240), 
        .B2(n20271), .ZN(P2_U3608) );
  INV_X1 U23182 ( .A(n20241), .ZN(n20248) );
  INV_X1 U23183 ( .A(n20242), .ZN(n20247) );
  INV_X1 U23184 ( .A(n20243), .ZN(n20244) );
  NAND2_X1 U23185 ( .A1(n20245), .A2(n20244), .ZN(n20246) );
  OAI211_X1 U23186 ( .C1(n20249), .C2(n20248), .A(n20247), .B(n20246), .ZN(
        n20251) );
  MUX2_X1 U23187 ( .A(P2_MORE_REG_SCAN_IN), .B(n20251), .S(n20250), .Z(
        P2_U3609) );
  AOI21_X1 U23188 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20252), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20254) );
  AOI211_X1 U23189 ( .C1(n20255), .C2(n20257), .A(n20254), .B(n20253), .ZN(
        n20269) );
  OAI21_X1 U23190 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n20256), .ZN(n20261) );
  NAND2_X1 U23191 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20257), .ZN(n20260) );
  NOR3_X1 U23192 ( .A1(n20262), .A2(n20258), .A3(n10468), .ZN(n20259) );
  AOI21_X1 U23193 ( .B1(n20261), .B2(n20260), .A(n20259), .ZN(n20268) );
  NAND2_X1 U23194 ( .A1(n20262), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20265) );
  INV_X1 U23195 ( .A(n20263), .ZN(n20264) );
  AND3_X1 U23196 ( .A1(n20265), .A2(n20264), .A3(n10493), .ZN(n20266) );
  NOR2_X1 U23197 ( .A1(n20269), .A2(n20266), .ZN(n20267) );
  AOI22_X1 U23198 ( .A1(n20270), .A2(n20269), .B1(n20268), .B2(n20267), .ZN(
        P2_U3610) );
  INV_X1 U23199 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20272) );
  AOI22_X1 U23200 ( .A1(n20274), .A2(n20273), .B1(n20272), .B2(n20271), .ZN(
        P2_U3611) );
  NAND2_X1 U23201 ( .A1(n13206), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21053) );
  INV_X1 U23202 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21123) );
  AOI21_X1 U23203 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20952), .A(n21013), 
        .ZN(n21019) );
  OAI21_X1 U23204 ( .B1(n21013), .B2(n21123), .A(n21015), .ZN(P1_U2802) );
  INV_X1 U23205 ( .A(n20275), .ZN(n20277) );
  OAI21_X1 U23206 ( .B1(n20277), .B2(n20276), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20278) );
  OAI21_X1 U23207 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20279), .A(n20278), 
        .ZN(P1_U2803) );
  NOR2_X1 U23208 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20281) );
  OAI21_X1 U23209 ( .B1(n20281), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21053), .ZN(
        n20280) );
  OAI21_X1 U23210 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21053), .A(n20280), 
        .ZN(P1_U2804) );
  OAI21_X1 U23211 ( .B1(BS16), .B2(n20281), .A(n21019), .ZN(n21017) );
  OAI21_X1 U23212 ( .B1(n21019), .B2(n21172), .A(n21017), .ZN(P1_U2805) );
  INV_X1 U23213 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20283) );
  OAI21_X1 U23214 ( .B1(n20284), .B2(n20283), .A(n20282), .ZN(P1_U2806) );
  NOR4_X1 U23215 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20288) );
  NOR4_X1 U23216 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20287) );
  NOR4_X1 U23217 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20286) );
  NOR4_X1 U23218 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20285) );
  NAND4_X1 U23219 ( .A1(n20288), .A2(n20287), .A3(n20286), .A4(n20285), .ZN(
        n20294) );
  NOR4_X1 U23220 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20292) );
  AOI211_X1 U23221 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20291) );
  NOR4_X1 U23222 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20290) );
  NOR4_X1 U23223 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20289) );
  NAND4_X1 U23224 ( .A1(n20292), .A2(n20291), .A3(n20290), .A4(n20289), .ZN(
        n20293) );
  NOR2_X1 U23225 ( .A1(n20294), .A2(n20293), .ZN(n21040) );
  INV_X1 U23226 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21058) );
  NOR3_X1 U23227 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20296) );
  OAI21_X1 U23228 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20296), .A(n21040), .ZN(
        n20295) );
  OAI21_X1 U23229 ( .B1(n21040), .B2(n21058), .A(n20295), .ZN(P1_U2807) );
  INV_X1 U23230 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21018) );
  AOI21_X1 U23231 ( .B1(n13461), .B2(n21018), .A(n20296), .ZN(n20297) );
  INV_X1 U23232 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21211) );
  INV_X1 U23233 ( .A(n21040), .ZN(n21037) );
  AOI22_X1 U23234 ( .A1(n21040), .A2(n20297), .B1(n21211), .B2(n21037), .ZN(
        P1_U2808) );
  NAND4_X1 U23235 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .A4(n15127), .ZN(n20304) );
  AOI22_X1 U23236 ( .A1(n20362), .A2(n20376), .B1(n20360), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n20298) );
  OAI21_X1 U23237 ( .B1(n15127), .B2(n20299), .A(n20298), .ZN(n20300) );
  AOI211_X1 U23238 ( .C1(n20348), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20346), .B(n20300), .ZN(n20303) );
  AOI22_X1 U23239 ( .A1(n20377), .A2(n20328), .B1(n20349), .B2(n20301), .ZN(
        n20302) );
  OAI211_X1 U23240 ( .C1(n20343), .C2(n20304), .A(n20303), .B(n20302), .ZN(
        P1_U2832) );
  NAND2_X1 U23241 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20313) );
  INV_X1 U23242 ( .A(n20313), .ZN(n20306) );
  OR2_X1 U23243 ( .A1(n20307), .A2(n20305), .ZN(n20357) );
  OAI21_X1 U23244 ( .B1(n20307), .B2(n20306), .A(n20357), .ZN(n20322) );
  OAI21_X1 U23245 ( .B1(n20365), .B2(n20309), .A(n20308), .ZN(n20310) );
  AOI21_X1 U23246 ( .B1(n20360), .B2(P1_EBX_REG_7__SCAN_IN), .A(n20310), .ZN(
        n20311) );
  OAI21_X1 U23247 ( .B1(n20312), .B2(n20320), .A(n20311), .ZN(n20315) );
  NOR3_X1 U23248 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20343), .A3(n20313), .ZN(
        n20314) );
  AOI211_X1 U23249 ( .C1(P1_REIP_REG_7__SCAN_IN), .C2(n20322), .A(n20315), .B(
        n20314), .ZN(n20318) );
  NAND2_X1 U23250 ( .A1(n20316), .A2(n20328), .ZN(n20317) );
  OAI211_X1 U23251 ( .C1(n20375), .C2(n20319), .A(n20318), .B(n20317), .ZN(
        P1_U2833) );
  NOR2_X1 U23252 ( .A1(n20320), .A2(n20380), .ZN(n20321) );
  AOI211_X1 U23253 ( .C1(n20348), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20346), .B(n20321), .ZN(n20324) );
  NAND2_X1 U23254 ( .A1(n20322), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n20323) );
  OAI211_X1 U23255 ( .C1(n20386), .C2(n20325), .A(n20324), .B(n20323), .ZN(
        n20327) );
  NOR3_X1 U23256 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20343), .A3(n20966), .ZN(
        n20326) );
  AOI211_X1 U23257 ( .C1(n20384), .C2(n20328), .A(n20327), .B(n20326), .ZN(
        n20329) );
  OAI21_X1 U23258 ( .B1(n20330), .B2(n20375), .A(n20329), .ZN(P1_U2834) );
  NAND2_X1 U23259 ( .A1(n20360), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n20337) );
  NAND2_X1 U23260 ( .A1(n20362), .A2(n20331), .ZN(n20336) );
  INV_X1 U23261 ( .A(n20332), .ZN(n20333) );
  AOI21_X1 U23262 ( .B1(n20349), .B2(n20333), .A(n20346), .ZN(n20335) );
  NAND2_X1 U23263 ( .A1(n20348), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n20334) );
  AND4_X1 U23264 ( .A1(n20337), .A2(n20336), .A3(n20335), .A4(n20334), .ZN(
        n20340) );
  NAND2_X1 U23265 ( .A1(n20338), .A2(n20371), .ZN(n20339) );
  OAI211_X1 U23266 ( .C1(n20357), .C2(n20966), .A(n20340), .B(n20339), .ZN(
        n20341) );
  INV_X1 U23267 ( .A(n20341), .ZN(n20342) );
  OAI21_X1 U23268 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20343), .A(n20342), .ZN(
        P1_U2835) );
  NAND2_X1 U23269 ( .A1(n20344), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20358) );
  AOI22_X1 U23270 ( .A1(n20362), .A2(n20345), .B1(n20360), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n20353) );
  AOI21_X1 U23271 ( .B1(n20363), .B2(n20347), .A(n20346), .ZN(n20352) );
  AOI22_X1 U23272 ( .A1(n20350), .A2(n20349), .B1(n20348), .B2(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20351) );
  NAND3_X1 U23273 ( .A1(n20353), .A2(n20352), .A3(n20351), .ZN(n20354) );
  AOI21_X1 U23274 ( .B1(n20355), .B2(n20371), .A(n20354), .ZN(n20356) );
  OAI221_X1 U23275 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(n20358), .C1(n13706), 
        .C2(n20357), .A(n20356), .ZN(P1_U2836) );
  INV_X1 U23276 ( .A(n20359), .ZN(n20361) );
  AOI22_X1 U23277 ( .A1(n20362), .A2(n20361), .B1(n20360), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n20374) );
  INV_X1 U23278 ( .A(n20363), .ZN(n20364) );
  OAI22_X1 U23279 ( .A1(n13462), .A2(n20365), .B1(n20364), .B2(n20693), .ZN(
        n20370) );
  INV_X1 U23280 ( .A(n20366), .ZN(n20368) );
  AOI21_X1 U23281 ( .B1(n20368), .B2(n13461), .A(n20367), .ZN(n20369) );
  AOI211_X1 U23282 ( .C1(n20372), .C2(n20371), .A(n20370), .B(n20369), .ZN(
        n20373) );
  OAI211_X1 U23283 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20375), .A(
        n20374), .B(n20373), .ZN(P1_U2839) );
  AOI22_X1 U23284 ( .A1(n20377), .A2(n20383), .B1(n20382), .B2(n20376), .ZN(
        n20378) );
  OAI21_X1 U23285 ( .B1(n20387), .B2(n20379), .A(n20378), .ZN(P1_U2864) );
  INV_X1 U23286 ( .A(n20380), .ZN(n20381) );
  AOI22_X1 U23287 ( .A1(n20384), .A2(n20383), .B1(n20382), .B2(n20381), .ZN(
        n20385) );
  OAI21_X1 U23288 ( .B1(n20387), .B2(n20386), .A(n20385), .ZN(P1_U2866) );
  AOI22_X1 U23289 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20388), .B1(n20409), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20389) );
  OAI21_X1 U23290 ( .B1(n20390), .B2(n21049), .A(n20389), .ZN(P1_U2921) );
  INV_X1 U23291 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20392) );
  AOI22_X1 U23292 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20391) );
  OAI21_X1 U23293 ( .B1(n20392), .B2(n20416), .A(n20391), .ZN(P1_U2922) );
  INV_X1 U23294 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20394) );
  AOI22_X1 U23295 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20393) );
  OAI21_X1 U23296 ( .B1(n20394), .B2(n20416), .A(n20393), .ZN(P1_U2923) );
  AOI22_X1 U23297 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20395) );
  OAI21_X1 U23298 ( .B1(n14984), .B2(n20416), .A(n20395), .ZN(P1_U2924) );
  AOI22_X1 U23299 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20396) );
  OAI21_X1 U23300 ( .B1(n20397), .B2(n20416), .A(n20396), .ZN(P1_U2925) );
  INV_X1 U23301 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20399) );
  AOI22_X1 U23302 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20398) );
  OAI21_X1 U23303 ( .B1(n20399), .B2(n20416), .A(n20398), .ZN(P1_U2926) );
  AOI22_X1 U23304 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20400), .B1(n20409), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20401) );
  OAI21_X1 U23305 ( .B1(n14111), .B2(n20416), .A(n20401), .ZN(P1_U2927) );
  INV_X1 U23306 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20403) );
  AOI22_X1 U23307 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20402) );
  OAI21_X1 U23308 ( .B1(n20403), .B2(n20416), .A(n20402), .ZN(P1_U2928) );
  AOI22_X1 U23309 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20404) );
  OAI21_X1 U23310 ( .B1(n12077), .B2(n20416), .A(n20404), .ZN(P1_U2929) );
  AOI22_X1 U23311 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20405) );
  OAI21_X1 U23312 ( .B1(n12153), .B2(n20416), .A(n20405), .ZN(P1_U2930) );
  AOI22_X1 U23313 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20406) );
  OAI21_X1 U23314 ( .B1(n12144), .B2(n20416), .A(n20406), .ZN(P1_U2931) );
  INV_X1 U23315 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20408) );
  AOI22_X1 U23316 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20407) );
  OAI21_X1 U23317 ( .B1(n20408), .B2(n20416), .A(n20407), .ZN(P1_U2932) );
  AOI22_X1 U23318 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20410) );
  OAI21_X1 U23319 ( .B1(n12125), .B2(n20416), .A(n20410), .ZN(P1_U2933) );
  AOI22_X1 U23320 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20411) );
  OAI21_X1 U23321 ( .B1(n20412), .B2(n20416), .A(n20411), .ZN(P1_U2934) );
  AOI22_X1 U23322 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20413) );
  OAI21_X1 U23323 ( .B1(n12108), .B2(n20416), .A(n20413), .ZN(P1_U2935) );
  AOI22_X1 U23324 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20414), .B1(n20409), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20415) );
  OAI21_X1 U23325 ( .B1(n12116), .B2(n20416), .A(n20415), .ZN(P1_U2936) );
  AOI22_X1 U23326 ( .A1(n20439), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20438), .ZN(n20418) );
  NAND2_X1 U23327 ( .A1(n20426), .A2(n20417), .ZN(n20428) );
  NAND2_X1 U23328 ( .A1(n20418), .A2(n20428), .ZN(P1_U2945) );
  AOI22_X1 U23329 ( .A1(n20439), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20420) );
  NAND2_X1 U23330 ( .A1(n20426), .A2(n20419), .ZN(n20432) );
  NAND2_X1 U23331 ( .A1(n20420), .A2(n20432), .ZN(P1_U2947) );
  AOI22_X1 U23332 ( .A1(n20439), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20422) );
  NAND2_X1 U23333 ( .A1(n20426), .A2(n20421), .ZN(n20434) );
  NAND2_X1 U23334 ( .A1(n20422), .A2(n20434), .ZN(P1_U2949) );
  AOI22_X1 U23335 ( .A1(n20439), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20424) );
  NAND2_X1 U23336 ( .A1(n20426), .A2(n20423), .ZN(n20436) );
  NAND2_X1 U23337 ( .A1(n20424), .A2(n20436), .ZN(P1_U2950) );
  AOI22_X1 U23338 ( .A1(n20439), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20438), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20427) );
  NAND2_X1 U23339 ( .A1(n20426), .A2(n20425), .ZN(n20440) );
  NAND2_X1 U23340 ( .A1(n20427), .A2(n20440), .ZN(P1_U2951) );
  AOI22_X1 U23341 ( .A1(n20439), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20429) );
  NAND2_X1 U23342 ( .A1(n20429), .A2(n20428), .ZN(P1_U2960) );
  AOI22_X1 U23343 ( .A1(n20439), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20438), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20431) );
  NAND2_X1 U23344 ( .A1(n20431), .A2(n20430), .ZN(P1_U2961) );
  AOI22_X1 U23345 ( .A1(n20439), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20438), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20433) );
  NAND2_X1 U23346 ( .A1(n20433), .A2(n20432), .ZN(P1_U2962) );
  AOI22_X1 U23347 ( .A1(n20439), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20438), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20435) );
  NAND2_X1 U23348 ( .A1(n20435), .A2(n20434), .ZN(P1_U2964) );
  AOI22_X1 U23349 ( .A1(n20439), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20438), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20437) );
  NAND2_X1 U23350 ( .A1(n20437), .A2(n20436), .ZN(P1_U2965) );
  AOI22_X1 U23351 ( .A1(n20439), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20438), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20441) );
  NAND2_X1 U23352 ( .A1(n20441), .A2(n20440), .ZN(P1_U2966) );
  INV_X1 U23353 ( .A(n20442), .ZN(n20444) );
  OAI211_X1 U23354 ( .C1(n20446), .C2(n20445), .A(n20444), .B(n20443), .ZN(
        n20449) );
  INV_X1 U23355 ( .A(n20447), .ZN(n20448) );
  AOI211_X1 U23356 ( .C1(n20451), .C2(n20450), .A(n20449), .B(n20448), .ZN(
        n20452) );
  OAI221_X1 U23357 ( .B1(n20455), .B2(n20454), .C1(n20455), .C2(n20453), .A(
        n20452), .ZN(P1_U3031) );
  NOR2_X1 U23358 ( .A1(n20456), .A2(n21032), .ZN(P1_U3032) );
  INV_X1 U23359 ( .A(n20757), .ZN(n20894) );
  NAND3_X1 U23360 ( .A1(n21034), .A2(n12762), .A3(n20692), .ZN(n20493) );
  NOR2_X1 U23361 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20493), .ZN(
        n20487) );
  AOI22_X1 U23362 ( .A1(n20881), .A2(n20487), .B1(n9807), .B2(n20938), .ZN(
        n20470) );
  INV_X1 U23363 ( .A(n20517), .ZN(n20458) );
  OAI21_X1 U23364 ( .B1(n20458), .B2(n20938), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20459) );
  NAND2_X1 U23365 ( .A1(n20459), .A2(n20889), .ZN(n20468) );
  OR2_X1 U23366 ( .A1(n13342), .A2(n20460), .ZN(n20548) );
  NOR2_X1 U23367 ( .A1(n20548), .A2(n11995), .ZN(n20466) );
  INV_X1 U23368 ( .A(n20461), .ZN(n20462) );
  NAND2_X1 U23369 ( .A1(n20462), .A2(n20753), .ZN(n20584) );
  INV_X1 U23370 ( .A(n20487), .ZN(n20463) );
  AOI22_X1 U23371 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20584), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20463), .ZN(n20465) );
  NAND2_X1 U23372 ( .A1(n20464), .A2(n20845), .ZN(n20521) );
  OAI211_X1 U23373 ( .C1(n20468), .C2(n20466), .A(n20465), .B(n20759), .ZN(
        n20489) );
  INV_X1 U23374 ( .A(n20466), .ZN(n20467) );
  INV_X1 U23375 ( .A(n20755), .ZN(n20695) );
  OAI22_X1 U23376 ( .A1(n20468), .A2(n20467), .B1(n20695), .B2(n20584), .ZN(
        n20488) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20489), .B1(
        n20880), .B2(n20488), .ZN(n20469) );
  OAI211_X1 U23378 ( .C1(n20894), .C2(n20517), .A(n20470), .B(n20469), .ZN(
        P1_U3033) );
  INV_X1 U23379 ( .A(n20823), .ZN(n20900) );
  AOI22_X1 U23380 ( .A1(n20896), .A2(n20487), .B1(n9811), .B2(n20938), .ZN(
        n20473) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20489), .B1(
        n20895), .B2(n20488), .ZN(n20472) );
  OAI211_X1 U23382 ( .C1(n20900), .C2(n20517), .A(n20473), .B(n20472), .ZN(
        P1_U3034) );
  INV_X1 U23383 ( .A(n20771), .ZN(n20906) );
  AOI22_X1 U23384 ( .A1(n20902), .A2(n20487), .B1(n9813), .B2(n20938), .ZN(
        n20475) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20489), .B1(
        n20901), .B2(n20488), .ZN(n20474) );
  OAI211_X1 U23386 ( .C1(n20906), .C2(n20517), .A(n20475), .B(n20474), .ZN(
        P1_U3035) );
  INV_X1 U23387 ( .A(n20909), .ZN(n20860) );
  AOI22_X1 U23388 ( .A1(n20908), .A2(n20487), .B1(n20857), .B2(n20938), .ZN(
        n20478) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20489), .B1(
        n20907), .B2(n20488), .ZN(n20477) );
  OAI211_X1 U23390 ( .C1(n20860), .C2(n20517), .A(n20478), .B(n20477), .ZN(
        P1_U3036) );
  INV_X1 U23391 ( .A(n20778), .ZN(n20918) );
  AOI22_X1 U23392 ( .A1(n20914), .A2(n20487), .B1(n20915), .B2(n20938), .ZN(
        n20480) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20489), .B1(
        n20913), .B2(n20488), .ZN(n20479) );
  OAI211_X1 U23394 ( .C1(n20918), .C2(n20517), .A(n20480), .B(n20479), .ZN(
        P1_U3037) );
  INV_X1 U23395 ( .A(n20828), .ZN(n20924) );
  AOI22_X1 U23396 ( .A1(n20920), .A2(n20487), .B1(n20921), .B2(n20938), .ZN(
        n20483) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20489), .B1(
        n20919), .B2(n20488), .ZN(n20482) );
  OAI211_X1 U23398 ( .C1(n20924), .C2(n20517), .A(n20483), .B(n20482), .ZN(
        P1_U3038) );
  INV_X1 U23399 ( .A(n20832), .ZN(n20932) );
  AOI22_X1 U23400 ( .A1(n20926), .A2(n20487), .B1(n9809), .B2(n20938), .ZN(
        n20486) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20489), .B1(
        n20925), .B2(n20488), .ZN(n20485) );
  OAI211_X1 U23402 ( .C1(n20932), .C2(n20517), .A(n20486), .B(n20485), .ZN(
        P1_U3039) );
  INV_X1 U23403 ( .A(n9805), .ZN(n20874) );
  AOI22_X1 U23404 ( .A1(n20933), .A2(n20487), .B1(n20869), .B2(n20938), .ZN(
        n20491) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20489), .B1(
        n20936), .B2(n20488), .ZN(n20490) );
  OAI211_X1 U23406 ( .C1(n20874), .C2(n20517), .A(n20491), .B(n20490), .ZN(
        P1_U3040) );
  NOR2_X1 U23407 ( .A1(n20721), .A2(n20493), .ZN(n20512) );
  INV_X1 U23408 ( .A(n20548), .ZN(n20492) );
  INV_X1 U23409 ( .A(n13944), .ZN(n20722) );
  AOI21_X1 U23410 ( .B1(n20492), .B2(n20722), .A(n20512), .ZN(n20494) );
  OAI22_X1 U23411 ( .A1(n20494), .A2(n20883), .B1(n20493), .B2(n21042), .ZN(
        n20513) );
  AOI22_X1 U23412 ( .A1(n20881), .A2(n20512), .B1(n20880), .B2(n20513), .ZN(
        n20499) );
  INV_X1 U23413 ( .A(n20493), .ZN(n20496) );
  INV_X1 U23414 ( .A(n20552), .ZN(n20560) );
  OAI211_X1 U23415 ( .C1(n20560), .C2(n21172), .A(n20889), .B(n20494), .ZN(
        n20495) );
  OAI211_X1 U23416 ( .C1(n20889), .C2(n20496), .A(n20888), .B(n20495), .ZN(
        n20514) );
  INV_X1 U23417 ( .A(n20728), .ZN(n20497) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20514), .B1(
        n20541), .B2(n20757), .ZN(n20498) );
  OAI211_X1 U23419 ( .C1(n9806), .C2(n20517), .A(n20499), .B(n20498), .ZN(
        P1_U3041) );
  AOI22_X1 U23420 ( .A1(n20896), .A2(n20512), .B1(n20895), .B2(n20513), .ZN(
        n20501) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20514), .B1(
        n20541), .B2(n20823), .ZN(n20500) );
  OAI211_X1 U23422 ( .C1(n9810), .C2(n20517), .A(n20501), .B(n20500), .ZN(
        P1_U3042) );
  AOI22_X1 U23423 ( .A1(n20902), .A2(n20512), .B1(n20901), .B2(n20513), .ZN(
        n20503) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20514), .B1(
        n20541), .B2(n20771), .ZN(n20502) );
  OAI211_X1 U23425 ( .C1(n9812), .C2(n20517), .A(n20503), .B(n20502), .ZN(
        P1_U3043) );
  AOI22_X1 U23426 ( .A1(n20908), .A2(n20512), .B1(n20907), .B2(n20513), .ZN(
        n20505) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20514), .B1(
        n20541), .B2(n20909), .ZN(n20504) );
  OAI211_X1 U23428 ( .C1(n20912), .C2(n20517), .A(n20505), .B(n20504), .ZN(
        P1_U3044) );
  AOI22_X1 U23429 ( .A1(n20914), .A2(n20512), .B1(n20913), .B2(n20513), .ZN(
        n20507) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20514), .B1(
        n20541), .B2(n20778), .ZN(n20506) );
  OAI211_X1 U23431 ( .C1(n20739), .C2(n20517), .A(n20507), .B(n20506), .ZN(
        P1_U3045) );
  AOI22_X1 U23432 ( .A1(n20920), .A2(n20512), .B1(n20919), .B2(n20513), .ZN(
        n20509) );
  AOI22_X1 U23433 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20514), .B1(
        n20541), .B2(n20828), .ZN(n20508) );
  OAI211_X1 U23434 ( .C1(n20831), .C2(n20517), .A(n20509), .B(n20508), .ZN(
        P1_U3046) );
  AOI22_X1 U23435 ( .A1(n20926), .A2(n20512), .B1(n20925), .B2(n20513), .ZN(
        n20511) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20514), .B1(
        n20541), .B2(n20832), .ZN(n20510) );
  OAI211_X1 U23437 ( .C1(n9808), .C2(n20517), .A(n20511), .B(n20510), .ZN(
        P1_U3047) );
  INV_X1 U23438 ( .A(n20869), .ZN(n20943) );
  AOI22_X1 U23439 ( .A1(n20936), .A2(n20513), .B1(n20933), .B2(n20512), .ZN(
        n20516) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20514), .B1(
        n20541), .B2(n20937), .ZN(n20515) );
  OAI211_X1 U23441 ( .C1(n20943), .C2(n20517), .A(n20516), .B(n20515), .ZN(
        P1_U3048) );
  NOR3_X1 U23442 ( .A1(n20575), .A2(n20541), .A3(n20883), .ZN(n20519) );
  NOR2_X1 U23443 ( .A1(n20519), .A2(n20725), .ZN(n20525) );
  INV_X1 U23444 ( .A(n20525), .ZN(n20520) );
  NOR2_X1 U23445 ( .A1(n20548), .A2(n20693), .ZN(n20524) );
  NOR3_X1 U23446 ( .A1(n20692), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20554) );
  NAND2_X1 U23447 ( .A1(n20721), .A2(n20554), .ZN(n20522) );
  INV_X1 U23448 ( .A(n20522), .ZN(n20540) );
  AOI22_X1 U23449 ( .A1(n20881), .A2(n20540), .B1(n20757), .B2(n20575), .ZN(
        n20527) );
  NOR2_X1 U23450 ( .A1(n10294), .A2(n21042), .ZN(n20637) );
  AOI211_X1 U23451 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20522), .A(n20637), 
        .B(n20521), .ZN(n20523) );
  OAI21_X1 U23452 ( .B1(n20525), .B2(n20524), .A(n20523), .ZN(n20542) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n9807), .ZN(n20526) );
  OAI211_X1 U23454 ( .C1(n20545), .C2(n20767), .A(n20527), .B(n20526), .ZN(
        P1_U3049) );
  AOI22_X1 U23455 ( .A1(n20896), .A2(n20540), .B1(n20823), .B2(n20575), .ZN(
        n20529) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n9811), .ZN(n20528) );
  OAI211_X1 U23457 ( .C1(n20545), .C2(n20770), .A(n20529), .B(n20528), .ZN(
        P1_U3050) );
  AOI22_X1 U23458 ( .A1(n20902), .A2(n20540), .B1(n20771), .B2(n20575), .ZN(
        n20531) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n9813), .ZN(n20530) );
  OAI211_X1 U23460 ( .C1(n20545), .C2(n20774), .A(n20531), .B(n20530), .ZN(
        P1_U3051) );
  AOI22_X1 U23461 ( .A1(n20908), .A2(n20540), .B1(n20909), .B2(n20575), .ZN(
        n20533) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20857), .ZN(n20532) );
  OAI211_X1 U23463 ( .C1(n20545), .C2(n20777), .A(n20533), .B(n20532), .ZN(
        P1_U3052) );
  AOI22_X1 U23464 ( .A1(n20914), .A2(n20540), .B1(n20915), .B2(n20541), .ZN(
        n20535) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20542), .B1(
        n20575), .B2(n20778), .ZN(n20534) );
  OAI211_X1 U23466 ( .C1(n20545), .C2(n20781), .A(n20535), .B(n20534), .ZN(
        P1_U3053) );
  AOI22_X1 U23467 ( .A1(n20920), .A2(n20540), .B1(n20828), .B2(n20575), .ZN(
        n20537) );
  AOI22_X1 U23468 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20921), .ZN(n20536) );
  OAI211_X1 U23469 ( .C1(n20545), .C2(n20784), .A(n20537), .B(n20536), .ZN(
        P1_U3054) );
  AOI22_X1 U23470 ( .A1(n20926), .A2(n20540), .B1(n9809), .B2(n20541), .ZN(
        n20539) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20542), .B1(
        n20575), .B2(n20832), .ZN(n20538) );
  OAI211_X1 U23472 ( .C1(n20545), .C2(n20787), .A(n20539), .B(n20538), .ZN(
        P1_U3055) );
  AOI22_X1 U23473 ( .A1(n20933), .A2(n20540), .B1(n9805), .B2(n20575), .ZN(
        n20544) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20542), .B1(
        n20541), .B2(n20869), .ZN(n20543) );
  OAI211_X1 U23475 ( .C1(n20545), .C2(n20793), .A(n20544), .B(n20543), .ZN(
        P1_U3056) );
  AND2_X1 U23476 ( .A1(n20547), .A2(n20546), .ZN(n20796) );
  INV_X1 U23477 ( .A(n20796), .ZN(n20875) );
  OR2_X1 U23478 ( .A1(n20548), .A2(n20875), .ZN(n20550) );
  NOR2_X1 U23479 ( .A1(n20795), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20576) );
  INV_X1 U23480 ( .A(n20576), .ZN(n20549) );
  AND2_X1 U23481 ( .A1(n20550), .A2(n20549), .ZN(n20556) );
  INV_X1 U23482 ( .A(n20556), .ZN(n20553) );
  INV_X1 U23483 ( .A(n20551), .ZN(n20882) );
  OAI21_X1 U23484 ( .B1(n20552), .B2(n20883), .A(n20882), .ZN(n20557) );
  AOI22_X1 U23485 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20554), .B1(n20553), 
        .B2(n20557), .ZN(n20580) );
  AOI22_X1 U23486 ( .A1(n20881), .A2(n20576), .B1(n9807), .B2(n20575), .ZN(
        n20562) );
  OAI21_X1 U23487 ( .B1(n20889), .B2(n20554), .A(n20888), .ZN(n20555) );
  AOI21_X1 U23488 ( .B1(n20557), .B2(n20556), .A(n20555), .ZN(n20558) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20577), .B1(
        n20605), .B2(n20757), .ZN(n20561) );
  OAI211_X1 U23490 ( .C1(n20580), .C2(n20767), .A(n20562), .B(n20561), .ZN(
        P1_U3057) );
  AOI22_X1 U23491 ( .A1(n20896), .A2(n20576), .B1(n20605), .B2(n20823), .ZN(
        n20564) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20577), .B1(
        n20575), .B2(n9811), .ZN(n20563) );
  OAI211_X1 U23493 ( .C1(n20580), .C2(n20770), .A(n20564), .B(n20563), .ZN(
        P1_U3058) );
  AOI22_X1 U23494 ( .A1(n20902), .A2(n20576), .B1(n9813), .B2(n20575), .ZN(
        n20566) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20577), .B1(
        n20605), .B2(n20771), .ZN(n20565) );
  OAI211_X1 U23496 ( .C1(n20580), .C2(n20774), .A(n20566), .B(n20565), .ZN(
        P1_U3059) );
  AOI22_X1 U23497 ( .A1(n20908), .A2(n20576), .B1(n20857), .B2(n20575), .ZN(
        n20568) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20577), .B1(
        n20605), .B2(n20909), .ZN(n20567) );
  OAI211_X1 U23499 ( .C1(n20580), .C2(n20777), .A(n20568), .B(n20567), .ZN(
        P1_U3060) );
  AOI22_X1 U23500 ( .A1(n20914), .A2(n20576), .B1(n20915), .B2(n20575), .ZN(
        n20570) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20577), .B1(
        n20605), .B2(n20778), .ZN(n20569) );
  OAI211_X1 U23502 ( .C1(n20580), .C2(n20781), .A(n20570), .B(n20569), .ZN(
        P1_U3061) );
  AOI22_X1 U23503 ( .A1(n20920), .A2(n20576), .B1(n20921), .B2(n20575), .ZN(
        n20572) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20577), .B1(
        n20605), .B2(n20828), .ZN(n20571) );
  OAI211_X1 U23505 ( .C1(n20580), .C2(n20784), .A(n20572), .B(n20571), .ZN(
        P1_U3062) );
  AOI22_X1 U23506 ( .A1(n20926), .A2(n20576), .B1(n20605), .B2(n20832), .ZN(
        n20574) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20577), .B1(
        n20575), .B2(n9809), .ZN(n20573) );
  OAI211_X1 U23508 ( .C1(n20580), .C2(n20787), .A(n20574), .B(n20573), .ZN(
        P1_U3063) );
  AOI22_X1 U23509 ( .A1(n20933), .A2(n20576), .B1(n20869), .B2(n20575), .ZN(
        n20579) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20577), .B1(
        n20605), .B2(n9805), .ZN(n20578) );
  OAI211_X1 U23511 ( .C1(n20580), .C2(n20793), .A(n20579), .B(n20578), .ZN(
        P1_U3064) );
  NAND3_X1 U23512 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21034), .A3(
        n20692), .ZN(n20609) );
  NOR2_X1 U23513 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20609), .ZN(
        n20603) );
  NOR2_X1 U23514 ( .A1(n13570), .A2(n20583), .ZN(n20663) );
  NAND2_X1 U23515 ( .A1(n20663), .A2(n20693), .ZN(n20586) );
  OAI22_X1 U23516 ( .A1(n20586), .A2(n20883), .B1(n20584), .B2(n20845), .ZN(
        n20604) );
  AOI22_X1 U23517 ( .A1(n20881), .A2(n20603), .B1(n20880), .B2(n20604), .ZN(
        n20590) );
  INV_X1 U23518 ( .A(n20632), .ZN(n20585) );
  OAI21_X1 U23519 ( .B1(n20605), .B2(n20585), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20587) );
  AOI21_X1 U23520 ( .B1(n20587), .B2(n20586), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20588) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20606), .B1(
        n20605), .B2(n9807), .ZN(n20589) );
  OAI211_X1 U23522 ( .C1(n20894), .C2(n20632), .A(n20590), .B(n20589), .ZN(
        P1_U3065) );
  AOI22_X1 U23523 ( .A1(n20896), .A2(n20603), .B1(n20895), .B2(n20604), .ZN(
        n20592) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20606), .B1(
        n20605), .B2(n9811), .ZN(n20591) );
  OAI211_X1 U23525 ( .C1(n20900), .C2(n20632), .A(n20592), .B(n20591), .ZN(
        P1_U3066) );
  AOI22_X1 U23526 ( .A1(n20902), .A2(n20603), .B1(n20901), .B2(n20604), .ZN(
        n20594) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20606), .B1(
        n20605), .B2(n9813), .ZN(n20593) );
  OAI211_X1 U23528 ( .C1(n20906), .C2(n20632), .A(n20594), .B(n20593), .ZN(
        P1_U3067) );
  AOI22_X1 U23529 ( .A1(n20908), .A2(n20603), .B1(n20907), .B2(n20604), .ZN(
        n20596) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20606), .B1(
        n20605), .B2(n20857), .ZN(n20595) );
  OAI211_X1 U23531 ( .C1(n20860), .C2(n20632), .A(n20596), .B(n20595), .ZN(
        P1_U3068) );
  AOI22_X1 U23532 ( .A1(n20914), .A2(n20603), .B1(n20913), .B2(n20604), .ZN(
        n20598) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20606), .B1(
        n20605), .B2(n20915), .ZN(n20597) );
  OAI211_X1 U23534 ( .C1(n20918), .C2(n20632), .A(n20598), .B(n20597), .ZN(
        P1_U3069) );
  AOI22_X1 U23535 ( .A1(n20920), .A2(n20603), .B1(n20919), .B2(n20604), .ZN(
        n20600) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20606), .B1(
        n20605), .B2(n20921), .ZN(n20599) );
  OAI211_X1 U23537 ( .C1(n20924), .C2(n20632), .A(n20600), .B(n20599), .ZN(
        P1_U3070) );
  AOI22_X1 U23538 ( .A1(n20926), .A2(n20603), .B1(n20925), .B2(n20604), .ZN(
        n20602) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20606), .B1(
        n20605), .B2(n9809), .ZN(n20601) );
  OAI211_X1 U23540 ( .C1(n20932), .C2(n20632), .A(n20602), .B(n20601), .ZN(
        P1_U3071) );
  AOI22_X1 U23541 ( .A1(n20936), .A2(n20604), .B1(n20933), .B2(n20603), .ZN(
        n20608) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20606), .B1(
        n20605), .B2(n20869), .ZN(n20607) );
  OAI211_X1 U23543 ( .C1(n20874), .C2(n20632), .A(n20608), .B(n20607), .ZN(
        P1_U3072) );
  NOR2_X1 U23544 ( .A1(n20721), .A2(n20609), .ZN(n20627) );
  AOI21_X1 U23545 ( .B1(n20663), .B2(n20722), .A(n20627), .ZN(n20610) );
  OAI22_X1 U23546 ( .A1(n20610), .A2(n20883), .B1(n20609), .B2(n21042), .ZN(
        n20628) );
  AOI22_X1 U23547 ( .A1(n20881), .A2(n20627), .B1(n20880), .B2(n20628), .ZN(
        n20614) );
  INV_X1 U23548 ( .A(n20609), .ZN(n20612) );
  OAI211_X1 U23549 ( .C1(n21024), .C2(n21172), .A(n20889), .B(n20610), .ZN(
        n20611) );
  OAI211_X1 U23550 ( .C1(n20889), .C2(n20612), .A(n20888), .B(n20611), .ZN(
        n20629) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20629), .B1(
        n20656), .B2(n20757), .ZN(n20613) );
  OAI211_X1 U23552 ( .C1(n9806), .C2(n20632), .A(n20614), .B(n20613), .ZN(
        P1_U3073) );
  AOI22_X1 U23553 ( .A1(n20896), .A2(n20627), .B1(n20895), .B2(n20628), .ZN(
        n20616) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20629), .B1(
        n20656), .B2(n20823), .ZN(n20615) );
  OAI211_X1 U23555 ( .C1(n9810), .C2(n20632), .A(n20616), .B(n20615), .ZN(
        P1_U3074) );
  AOI22_X1 U23556 ( .A1(n20902), .A2(n20627), .B1(n20901), .B2(n20628), .ZN(
        n20618) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20629), .B1(
        n20656), .B2(n20771), .ZN(n20617) );
  OAI211_X1 U23558 ( .C1(n9812), .C2(n20632), .A(n20618), .B(n20617), .ZN(
        P1_U3075) );
  AOI22_X1 U23559 ( .A1(n20908), .A2(n20627), .B1(n20907), .B2(n20628), .ZN(
        n20620) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20629), .B1(
        n20656), .B2(n20909), .ZN(n20619) );
  OAI211_X1 U23561 ( .C1(n20912), .C2(n20632), .A(n20620), .B(n20619), .ZN(
        P1_U3076) );
  AOI22_X1 U23562 ( .A1(n20914), .A2(n20627), .B1(n20913), .B2(n20628), .ZN(
        n20622) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20629), .B1(
        n20656), .B2(n20778), .ZN(n20621) );
  OAI211_X1 U23564 ( .C1(n20739), .C2(n20632), .A(n20622), .B(n20621), .ZN(
        P1_U3077) );
  AOI22_X1 U23565 ( .A1(n20920), .A2(n20627), .B1(n20919), .B2(n20628), .ZN(
        n20624) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20629), .B1(
        n20656), .B2(n20828), .ZN(n20623) );
  OAI211_X1 U23567 ( .C1(n20831), .C2(n20632), .A(n20624), .B(n20623), .ZN(
        P1_U3078) );
  AOI22_X1 U23568 ( .A1(n20926), .A2(n20627), .B1(n20925), .B2(n20628), .ZN(
        n20626) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20629), .B1(
        n20656), .B2(n20832), .ZN(n20625) );
  OAI211_X1 U23570 ( .C1(n9808), .C2(n20632), .A(n20626), .B(n20625), .ZN(
        P1_U3079) );
  AOI22_X1 U23571 ( .A1(n20936), .A2(n20628), .B1(n20933), .B2(n20627), .ZN(
        n20631) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20629), .B1(
        n20656), .B2(n20937), .ZN(n20630) );
  OAI211_X1 U23573 ( .C1(n20943), .C2(n20632), .A(n20631), .B(n20630), .ZN(
        P1_U3080) );
  INV_X1 U23574 ( .A(n20656), .ZN(n20633) );
  NAND2_X1 U23575 ( .A1(n20633), .A2(n20889), .ZN(n20634) );
  INV_X1 U23576 ( .A(n20725), .ZN(n21027) );
  OAI21_X1 U23577 ( .B1(n20634), .B2(n20686), .A(n21027), .ZN(n20639) );
  AND2_X1 U23578 ( .A1(n20663), .A2(n11995), .ZN(n20636) );
  INV_X1 U23579 ( .A(n20845), .ZN(n20635) );
  AOI22_X1 U23580 ( .A1(n20639), .A2(n20636), .B1(n20635), .B2(n10294), .ZN(
        n20660) );
  INV_X1 U23581 ( .A(n20669), .ZN(n20664) );
  NOR2_X1 U23582 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20664), .ZN(
        n20655) );
  AOI22_X1 U23583 ( .A1(n20881), .A2(n20655), .B1(n9807), .B2(n20656), .ZN(
        n20642) );
  INV_X1 U23584 ( .A(n20636), .ZN(n20638) );
  AOI21_X1 U23585 ( .B1(n20639), .B2(n20638), .A(n20637), .ZN(n20640) );
  OAI211_X1 U23586 ( .C1(n20655), .C2(n20760), .A(n20849), .B(n20640), .ZN(
        n20657) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20657), .B1(
        n20686), .B2(n20757), .ZN(n20641) );
  OAI211_X1 U23588 ( .C1(n20660), .C2(n20767), .A(n20642), .B(n20641), .ZN(
        P1_U3081) );
  AOI22_X1 U23589 ( .A1(n20896), .A2(n20655), .B1(n9811), .B2(n20656), .ZN(
        n20644) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20657), .B1(
        n20686), .B2(n20823), .ZN(n20643) );
  OAI211_X1 U23591 ( .C1(n20660), .C2(n20770), .A(n20644), .B(n20643), .ZN(
        P1_U3082) );
  AOI22_X1 U23592 ( .A1(n20902), .A2(n20655), .B1(n9813), .B2(n20656), .ZN(
        n20646) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20657), .B1(
        n20686), .B2(n20771), .ZN(n20645) );
  OAI211_X1 U23594 ( .C1(n20660), .C2(n20774), .A(n20646), .B(n20645), .ZN(
        P1_U3083) );
  AOI22_X1 U23595 ( .A1(n20908), .A2(n20655), .B1(n20909), .B2(n20686), .ZN(
        n20648) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20857), .ZN(n20647) );
  OAI211_X1 U23597 ( .C1(n20660), .C2(n20777), .A(n20648), .B(n20647), .ZN(
        P1_U3084) );
  AOI22_X1 U23598 ( .A1(n20914), .A2(n20655), .B1(n20778), .B2(n20686), .ZN(
        n20650) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20915), .ZN(n20649) );
  OAI211_X1 U23600 ( .C1(n20660), .C2(n20781), .A(n20650), .B(n20649), .ZN(
        P1_U3085) );
  AOI22_X1 U23601 ( .A1(n20920), .A2(n20655), .B1(n20921), .B2(n20656), .ZN(
        n20652) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20657), .B1(
        n20686), .B2(n20828), .ZN(n20651) );
  OAI211_X1 U23603 ( .C1(n20660), .C2(n20784), .A(n20652), .B(n20651), .ZN(
        P1_U3086) );
  AOI22_X1 U23604 ( .A1(n20926), .A2(n20655), .B1(n20832), .B2(n20686), .ZN(
        n20654) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n9809), .ZN(n20653) );
  OAI211_X1 U23606 ( .C1(n20660), .C2(n20787), .A(n20654), .B(n20653), .ZN(
        P1_U3087) );
  AOI22_X1 U23607 ( .A1(n20933), .A2(n20655), .B1(n9805), .B2(n20686), .ZN(
        n20659) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20657), .B1(
        n20656), .B2(n20869), .ZN(n20658) );
  OAI211_X1 U23609 ( .C1(n20660), .C2(n20793), .A(n20659), .B(n20658), .ZN(
        P1_U3088) );
  INV_X1 U23610 ( .A(n20662), .ZN(n20684) );
  AOI21_X1 U23611 ( .B1(n20663), .B2(n20796), .A(n20684), .ZN(n20666) );
  OAI22_X1 U23612 ( .A1(n20666), .A2(n20883), .B1(n20664), .B2(n21042), .ZN(
        n20685) );
  AOI22_X1 U23613 ( .A1(n20881), .A2(n20684), .B1(n20880), .B2(n20685), .ZN(
        n20671) );
  OAI21_X1 U23614 ( .B1(n20665), .B2(n20883), .A(n20882), .ZN(n20667) );
  NAND2_X1 U23615 ( .A1(n20667), .A2(n20666), .ZN(n20668) );
  OAI211_X1 U23616 ( .C1(n20669), .C2(n20889), .A(n20888), .B(n20668), .ZN(
        n20687) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n9807), .ZN(n20670) );
  OAI211_X1 U23618 ( .C1(n20894), .C2(n20696), .A(n20671), .B(n20670), .ZN(
        P1_U3089) );
  AOI22_X1 U23619 ( .A1(n20896), .A2(n20684), .B1(n20895), .B2(n20685), .ZN(
        n20673) );
  AOI22_X1 U23620 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n9811), .ZN(n20672) );
  OAI211_X1 U23621 ( .C1(n20900), .C2(n20696), .A(n20673), .B(n20672), .ZN(
        P1_U3090) );
  AOI22_X1 U23622 ( .A1(n20902), .A2(n20684), .B1(n20901), .B2(n20685), .ZN(
        n20675) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n9813), .ZN(n20674) );
  OAI211_X1 U23624 ( .C1(n20906), .C2(n20696), .A(n20675), .B(n20674), .ZN(
        P1_U3091) );
  AOI22_X1 U23625 ( .A1(n20908), .A2(n20684), .B1(n20907), .B2(n20685), .ZN(
        n20677) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20857), .ZN(n20676) );
  OAI211_X1 U23627 ( .C1(n20860), .C2(n20696), .A(n20677), .B(n20676), .ZN(
        P1_U3092) );
  AOI22_X1 U23628 ( .A1(n20914), .A2(n20684), .B1(n20913), .B2(n20685), .ZN(
        n20679) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20915), .ZN(n20678) );
  OAI211_X1 U23630 ( .C1(n20918), .C2(n20696), .A(n20679), .B(n20678), .ZN(
        P1_U3093) );
  AOI22_X1 U23631 ( .A1(n20920), .A2(n20684), .B1(n20919), .B2(n20685), .ZN(
        n20681) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20921), .ZN(n20680) );
  OAI211_X1 U23633 ( .C1(n20924), .C2(n20696), .A(n20681), .B(n20680), .ZN(
        P1_U3094) );
  AOI22_X1 U23634 ( .A1(n20926), .A2(n20684), .B1(n20925), .B2(n20685), .ZN(
        n20683) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n9809), .ZN(n20682) );
  OAI211_X1 U23636 ( .C1(n20932), .C2(n20696), .A(n20683), .B(n20682), .ZN(
        P1_U3095) );
  AOI22_X1 U23637 ( .A1(n20936), .A2(n20685), .B1(n20684), .B2(n20933), .ZN(
        n20689) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20687), .B1(
        n20686), .B2(n20869), .ZN(n20688) );
  OAI211_X1 U23639 ( .C1(n20874), .C2(n20696), .A(n20689), .B(n20688), .ZN(
        P1_U3096) );
  INV_X1 U23640 ( .A(n21020), .ZN(n20691) );
  NAND3_X1 U23641 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12762), .A3(
        n20692), .ZN(n20723) );
  NOR2_X1 U23642 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20723), .ZN(
        n20715) );
  AND2_X1 U23643 ( .A1(n13342), .A2(n13570), .ZN(n20797) );
  AOI21_X1 U23644 ( .B1(n20797), .B2(n20693), .A(n20715), .ZN(n20698) );
  OAI22_X1 U23645 ( .A1(n20698), .A2(n20883), .B1(n20695), .B2(n20694), .ZN(
        n20716) );
  AOI22_X1 U23646 ( .A1(n20881), .A2(n20715), .B1(n20880), .B2(n20716), .ZN(
        n20702) );
  INV_X1 U23647 ( .A(n20749), .ZN(n20697) );
  OAI21_X1 U23648 ( .B1(n20697), .B2(n20717), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20699) );
  NAND2_X1 U23649 ( .A1(n20699), .A2(n20698), .ZN(n20700) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20718), .B1(
        n20717), .B2(n9807), .ZN(n20701) );
  OAI211_X1 U23651 ( .C1(n20894), .C2(n20749), .A(n20702), .B(n20701), .ZN(
        P1_U3097) );
  AOI22_X1 U23652 ( .A1(n20896), .A2(n20715), .B1(n20895), .B2(n20716), .ZN(
        n20704) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20718), .B1(
        n20717), .B2(n9811), .ZN(n20703) );
  OAI211_X1 U23654 ( .C1(n20900), .C2(n20749), .A(n20704), .B(n20703), .ZN(
        P1_U3098) );
  AOI22_X1 U23655 ( .A1(n20902), .A2(n20715), .B1(n20901), .B2(n20716), .ZN(
        n20706) );
  AOI22_X1 U23656 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20718), .B1(
        n20717), .B2(n9813), .ZN(n20705) );
  OAI211_X1 U23657 ( .C1(n20906), .C2(n20749), .A(n20706), .B(n20705), .ZN(
        P1_U3099) );
  AOI22_X1 U23658 ( .A1(n20908), .A2(n20715), .B1(n20907), .B2(n20716), .ZN(
        n20708) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20718), .B1(
        n20717), .B2(n20857), .ZN(n20707) );
  OAI211_X1 U23660 ( .C1(n20860), .C2(n20749), .A(n20708), .B(n20707), .ZN(
        P1_U3100) );
  AOI22_X1 U23661 ( .A1(n20914), .A2(n20715), .B1(n20913), .B2(n20716), .ZN(
        n20710) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20718), .B1(
        n20717), .B2(n20915), .ZN(n20709) );
  OAI211_X1 U23663 ( .C1(n20918), .C2(n20749), .A(n20710), .B(n20709), .ZN(
        P1_U3101) );
  AOI22_X1 U23664 ( .A1(n20920), .A2(n20715), .B1(n20919), .B2(n20716), .ZN(
        n20712) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20718), .B1(
        n20717), .B2(n20921), .ZN(n20711) );
  OAI211_X1 U23666 ( .C1(n20924), .C2(n20749), .A(n20712), .B(n20711), .ZN(
        P1_U3102) );
  AOI22_X1 U23667 ( .A1(n20926), .A2(n20715), .B1(n20925), .B2(n20716), .ZN(
        n20714) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20718), .B1(
        n20717), .B2(n9809), .ZN(n20713) );
  OAI211_X1 U23669 ( .C1(n20932), .C2(n20749), .A(n20714), .B(n20713), .ZN(
        P1_U3103) );
  AOI22_X1 U23670 ( .A1(n20936), .A2(n20716), .B1(n20933), .B2(n20715), .ZN(
        n20720) );
  AOI22_X1 U23671 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20718), .B1(
        n20717), .B2(n20869), .ZN(n20719) );
  OAI211_X1 U23672 ( .C1(n20874), .C2(n20749), .A(n20720), .B(n20719), .ZN(
        P1_U3104) );
  NOR2_X1 U23673 ( .A1(n20721), .A2(n20723), .ZN(n20744) );
  AOI21_X1 U23674 ( .B1(n20797), .B2(n20722), .A(n20744), .ZN(n20724) );
  OAI22_X1 U23675 ( .A1(n20724), .A2(n20883), .B1(n20723), .B2(n21042), .ZN(
        n20745) );
  AOI22_X1 U23676 ( .A1(n20881), .A2(n20744), .B1(n20880), .B2(n20745), .ZN(
        n20730) );
  INV_X1 U23677 ( .A(n20723), .ZN(n20727) );
  OAI21_X1 U23678 ( .B1(n21020), .B2(n20725), .A(n20724), .ZN(n20726) );
  OAI211_X1 U23679 ( .C1(n20889), .C2(n20727), .A(n20888), .B(n20726), .ZN(
        n20746) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20746), .B1(
        n20789), .B2(n20757), .ZN(n20729) );
  OAI211_X1 U23681 ( .C1(n9806), .C2(n20749), .A(n20730), .B(n20729), .ZN(
        P1_U3105) );
  AOI22_X1 U23682 ( .A1(n20896), .A2(n20744), .B1(n20895), .B2(n20745), .ZN(
        n20732) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20746), .B1(
        n20789), .B2(n20823), .ZN(n20731) );
  OAI211_X1 U23684 ( .C1(n9810), .C2(n20749), .A(n20732), .B(n20731), .ZN(
        P1_U3106) );
  AOI22_X1 U23685 ( .A1(n20902), .A2(n20744), .B1(n20901), .B2(n20745), .ZN(
        n20734) );
  AOI22_X1 U23686 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20746), .B1(
        n20789), .B2(n20771), .ZN(n20733) );
  OAI211_X1 U23687 ( .C1(n9812), .C2(n20749), .A(n20734), .B(n20733), .ZN(
        P1_U3107) );
  AOI22_X1 U23688 ( .A1(n20908), .A2(n20744), .B1(n20907), .B2(n20745), .ZN(
        n20736) );
  AOI22_X1 U23689 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20746), .B1(
        n20789), .B2(n20909), .ZN(n20735) );
  OAI211_X1 U23690 ( .C1(n20912), .C2(n20749), .A(n20736), .B(n20735), .ZN(
        P1_U3108) );
  AOI22_X1 U23691 ( .A1(n20914), .A2(n20744), .B1(n20913), .B2(n20745), .ZN(
        n20738) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20746), .B1(
        n20789), .B2(n20778), .ZN(n20737) );
  OAI211_X1 U23693 ( .C1(n20739), .C2(n20749), .A(n20738), .B(n20737), .ZN(
        P1_U3109) );
  AOI22_X1 U23694 ( .A1(n20920), .A2(n20744), .B1(n20919), .B2(n20745), .ZN(
        n20741) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20746), .B1(
        n20789), .B2(n20828), .ZN(n20740) );
  OAI211_X1 U23696 ( .C1(n20831), .C2(n20749), .A(n20741), .B(n20740), .ZN(
        P1_U3110) );
  AOI22_X1 U23697 ( .A1(n20926), .A2(n20744), .B1(n20925), .B2(n20745), .ZN(
        n20743) );
  AOI22_X1 U23698 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20746), .B1(
        n20789), .B2(n20832), .ZN(n20742) );
  OAI211_X1 U23699 ( .C1(n9808), .C2(n20749), .A(n20743), .B(n20742), .ZN(
        P1_U3111) );
  AOI22_X1 U23700 ( .A1(n20936), .A2(n20745), .B1(n20933), .B2(n20744), .ZN(
        n20748) );
  AOI22_X1 U23701 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20746), .B1(
        n20789), .B2(n9805), .ZN(n20747) );
  OAI211_X1 U23702 ( .C1(n20943), .C2(n20749), .A(n20748), .B(n20747), .ZN(
        P1_U3112) );
  NAND3_X1 U23703 ( .A1(n20756), .A2(n20751), .A3(n20889), .ZN(n20752) );
  NAND2_X1 U23704 ( .A1(n20752), .A2(n21027), .ZN(n20763) );
  AND2_X1 U23705 ( .A1(n20797), .A2(n11995), .ZN(n20758) );
  OR2_X1 U23706 ( .A1(n20753), .A2(n21034), .ZN(n20844) );
  INV_X1 U23707 ( .A(n20844), .ZN(n20754) );
  AOI22_X1 U23708 ( .A1(n20763), .A2(n20758), .B1(n20755), .B2(n20754), .ZN(
        n20794) );
  NAND3_X1 U23709 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n12762), .ZN(n20799) );
  NOR2_X1 U23710 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20799), .ZN(
        n20788) );
  AOI22_X1 U23711 ( .A1(n20757), .A2(n20819), .B1(n20881), .B2(n20788), .ZN(
        n20766) );
  INV_X1 U23712 ( .A(n20758), .ZN(n20762) );
  NAND2_X1 U23713 ( .A1(n20844), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20848) );
  OAI211_X1 U23714 ( .C1(n20760), .C2(n20788), .A(n20848), .B(n20759), .ZN(
        n20761) );
  AOI21_X1 U23715 ( .B1(n20763), .B2(n20762), .A(n20761), .ZN(n20764) );
  AOI22_X1 U23716 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20790), .B1(
        n20789), .B2(n9807), .ZN(n20765) );
  OAI211_X1 U23717 ( .C1(n20794), .C2(n20767), .A(n20766), .B(n20765), .ZN(
        P1_U3113) );
  AOI22_X1 U23718 ( .A1(n20896), .A2(n20788), .B1(n20823), .B2(n20819), .ZN(
        n20769) );
  AOI22_X1 U23719 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20790), .B1(
        n20789), .B2(n9811), .ZN(n20768) );
  OAI211_X1 U23720 ( .C1(n20794), .C2(n20770), .A(n20769), .B(n20768), .ZN(
        P1_U3114) );
  AOI22_X1 U23721 ( .A1(n9813), .A2(n20789), .B1(n20902), .B2(n20788), .ZN(
        n20773) );
  AOI22_X1 U23722 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20790), .B1(
        n20819), .B2(n20771), .ZN(n20772) );
  OAI211_X1 U23723 ( .C1(n20794), .C2(n20774), .A(n20773), .B(n20772), .ZN(
        P1_U3115) );
  AOI22_X1 U23724 ( .A1(n20908), .A2(n20788), .B1(n20909), .B2(n20819), .ZN(
        n20776) );
  AOI22_X1 U23725 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20790), .B1(
        n20789), .B2(n20857), .ZN(n20775) );
  OAI211_X1 U23726 ( .C1(n20794), .C2(n20777), .A(n20776), .B(n20775), .ZN(
        P1_U3116) );
  AOI22_X1 U23727 ( .A1(n20915), .A2(n20789), .B1(n20914), .B2(n20788), .ZN(
        n20780) );
  AOI22_X1 U23728 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20790), .B1(
        n20819), .B2(n20778), .ZN(n20779) );
  OAI211_X1 U23729 ( .C1(n20794), .C2(n20781), .A(n20780), .B(n20779), .ZN(
        P1_U3117) );
  AOI22_X1 U23730 ( .A1(n20920), .A2(n20788), .B1(n20921), .B2(n20789), .ZN(
        n20783) );
  AOI22_X1 U23731 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20790), .B1(
        n20819), .B2(n20828), .ZN(n20782) );
  OAI211_X1 U23732 ( .C1(n20794), .C2(n20784), .A(n20783), .B(n20782), .ZN(
        P1_U3118) );
  AOI22_X1 U23733 ( .A1(n20926), .A2(n20788), .B1(n9809), .B2(n20789), .ZN(
        n20786) );
  AOI22_X1 U23734 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20790), .B1(
        n20819), .B2(n20832), .ZN(n20785) );
  OAI211_X1 U23735 ( .C1(n20794), .C2(n20787), .A(n20786), .B(n20785), .ZN(
        P1_U3119) );
  AOI22_X1 U23736 ( .A1(n20869), .A2(n20789), .B1(n20933), .B2(n20788), .ZN(
        n20792) );
  AOI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20790), .B1(
        n20819), .B2(n9805), .ZN(n20791) );
  OAI211_X1 U23738 ( .C1(n20794), .C2(n20793), .A(n20792), .B(n20791), .ZN(
        P1_U3120) );
  NOR2_X1 U23739 ( .A1(n20795), .A2(n21034), .ZN(n20817) );
  AOI21_X1 U23740 ( .B1(n20797), .B2(n20796), .A(n20817), .ZN(n20798) );
  OAI22_X1 U23741 ( .A1(n20798), .A2(n20883), .B1(n20799), .B2(n21042), .ZN(
        n20818) );
  AOI22_X1 U23742 ( .A1(n20881), .A2(n20817), .B1(n20880), .B2(n20818), .ZN(
        n20804) );
  INV_X1 U23743 ( .A(n20799), .ZN(n20802) );
  INV_X1 U23744 ( .A(n20800), .ZN(n21023) );
  NOR2_X1 U23745 ( .A1(n21020), .A2(n21023), .ZN(n20801) );
  OAI21_X1 U23746 ( .B1(n20802), .B2(n20801), .A(n20888), .ZN(n20820) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20820), .B1(
        n20819), .B2(n9807), .ZN(n20803) );
  OAI211_X1 U23748 ( .C1(n20894), .C2(n20841), .A(n20804), .B(n20803), .ZN(
        P1_U3121) );
  AOI22_X1 U23749 ( .A1(n20896), .A2(n20817), .B1(n20895), .B2(n20818), .ZN(
        n20806) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20820), .B1(
        n20819), .B2(n9811), .ZN(n20805) );
  OAI211_X1 U23751 ( .C1(n20900), .C2(n20841), .A(n20806), .B(n20805), .ZN(
        P1_U3122) );
  AOI22_X1 U23752 ( .A1(n20902), .A2(n20817), .B1(n20901), .B2(n20818), .ZN(
        n20808) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20820), .B1(
        n20819), .B2(n9813), .ZN(n20807) );
  OAI211_X1 U23754 ( .C1(n20906), .C2(n20841), .A(n20808), .B(n20807), .ZN(
        P1_U3123) );
  AOI22_X1 U23755 ( .A1(n20908), .A2(n20817), .B1(n20907), .B2(n20818), .ZN(
        n20810) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20820), .B1(
        n20819), .B2(n20857), .ZN(n20809) );
  OAI211_X1 U23757 ( .C1(n20860), .C2(n20841), .A(n20810), .B(n20809), .ZN(
        P1_U3124) );
  AOI22_X1 U23758 ( .A1(n20914), .A2(n20817), .B1(n20913), .B2(n20818), .ZN(
        n20812) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20820), .B1(
        n20819), .B2(n20915), .ZN(n20811) );
  OAI211_X1 U23760 ( .C1(n20918), .C2(n20841), .A(n20812), .B(n20811), .ZN(
        P1_U3125) );
  AOI22_X1 U23761 ( .A1(n20920), .A2(n20817), .B1(n20919), .B2(n20818), .ZN(
        n20814) );
  AOI22_X1 U23762 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20820), .B1(
        n20819), .B2(n20921), .ZN(n20813) );
  OAI211_X1 U23763 ( .C1(n20924), .C2(n20841), .A(n20814), .B(n20813), .ZN(
        P1_U3126) );
  AOI22_X1 U23764 ( .A1(n20926), .A2(n20817), .B1(n20925), .B2(n20818), .ZN(
        n20816) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20820), .B1(
        n20819), .B2(n9809), .ZN(n20815) );
  OAI211_X1 U23766 ( .C1(n20932), .C2(n20841), .A(n20816), .B(n20815), .ZN(
        P1_U3127) );
  AOI22_X1 U23767 ( .A1(n20936), .A2(n20818), .B1(n20933), .B2(n20817), .ZN(
        n20822) );
  AOI22_X1 U23768 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20820), .B1(
        n20819), .B2(n20869), .ZN(n20821) );
  OAI211_X1 U23769 ( .C1(n20874), .C2(n20841), .A(n20822), .B(n20821), .ZN(
        P1_U3128) );
  AOI22_X1 U23770 ( .A1(n20896), .A2(n20836), .B1(n20835), .B2(n20823), .ZN(
        n20825) );
  AOI22_X1 U23771 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20838), .B1(
        n20895), .B2(n20837), .ZN(n20824) );
  OAI211_X1 U23772 ( .C1(n9810), .C2(n20841), .A(n20825), .B(n20824), .ZN(
        P1_U3130) );
  AOI22_X1 U23773 ( .A1(n20908), .A2(n20836), .B1(n20835), .B2(n20909), .ZN(
        n20827) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20838), .B1(
        n20907), .B2(n20837), .ZN(n20826) );
  OAI211_X1 U23775 ( .C1(n20912), .C2(n20841), .A(n20827), .B(n20826), .ZN(
        P1_U3132) );
  AOI22_X1 U23776 ( .A1(n20920), .A2(n20836), .B1(n20835), .B2(n20828), .ZN(
        n20830) );
  AOI22_X1 U23777 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20838), .B1(
        n20919), .B2(n20837), .ZN(n20829) );
  OAI211_X1 U23778 ( .C1(n20831), .C2(n20841), .A(n20830), .B(n20829), .ZN(
        P1_U3134) );
  AOI22_X1 U23779 ( .A1(n20926), .A2(n20836), .B1(n20835), .B2(n20832), .ZN(
        n20834) );
  AOI22_X1 U23780 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20838), .B1(
        n20925), .B2(n20837), .ZN(n20833) );
  OAI211_X1 U23781 ( .C1(n9808), .C2(n20841), .A(n20834), .B(n20833), .ZN(
        P1_U3135) );
  AOI22_X1 U23782 ( .A1(n20933), .A2(n20836), .B1(n20835), .B2(n20937), .ZN(
        n20840) );
  AOI22_X1 U23783 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20838), .B1(
        n20936), .B2(n20837), .ZN(n20839) );
  OAI211_X1 U23784 ( .C1(n20943), .C2(n20841), .A(n20840), .B(n20839), .ZN(
        P1_U3136) );
  NOR2_X1 U23785 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20879), .ZN(
        n20867) );
  INV_X1 U23786 ( .A(n20876), .ZN(n20843) );
  NAND2_X1 U23787 ( .A1(n20843), .A2(n11995), .ZN(n20846) );
  OAI22_X1 U23788 ( .A1(n20846), .A2(n20883), .B1(n20845), .B2(n20844), .ZN(
        n20868) );
  AOI22_X1 U23789 ( .A1(n20881), .A2(n20867), .B1(n20880), .B2(n20868), .ZN(
        n20852) );
  OAI21_X1 U23790 ( .B1(n20928), .B2(n20870), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20847) );
  AOI21_X1 U23791 ( .B1(n20847), .B2(n20846), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20850) );
  AOI22_X1 U23792 ( .A1(n20871), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9807), .B2(n20870), .ZN(n20851) );
  OAI211_X1 U23793 ( .C1(n20894), .C2(n20942), .A(n20852), .B(n20851), .ZN(
        P1_U3145) );
  AOI22_X1 U23794 ( .A1(n20896), .A2(n20867), .B1(n20895), .B2(n20868), .ZN(
        n20854) );
  AOI22_X1 U23795 ( .A1(n20871), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n20870), .B2(n9811), .ZN(n20853) );
  OAI211_X1 U23796 ( .C1(n20900), .C2(n20942), .A(n20854), .B(n20853), .ZN(
        P1_U3146) );
  AOI22_X1 U23797 ( .A1(n20902), .A2(n20867), .B1(n20901), .B2(n20868), .ZN(
        n20856) );
  AOI22_X1 U23798 ( .A1(n20871), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n20870), .B2(n9813), .ZN(n20855) );
  OAI211_X1 U23799 ( .C1(n20906), .C2(n20942), .A(n20856), .B(n20855), .ZN(
        P1_U3147) );
  AOI22_X1 U23800 ( .A1(n20908), .A2(n20867), .B1(n20907), .B2(n20868), .ZN(
        n20859) );
  AOI22_X1 U23801 ( .A1(n20871), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n20870), .B2(n20857), .ZN(n20858) );
  OAI211_X1 U23802 ( .C1(n20860), .C2(n20942), .A(n20859), .B(n20858), .ZN(
        P1_U3148) );
  AOI22_X1 U23803 ( .A1(n20914), .A2(n20867), .B1(n20913), .B2(n20868), .ZN(
        n20862) );
  AOI22_X1 U23804 ( .A1(n20871), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n20870), .B2(n20915), .ZN(n20861) );
  OAI211_X1 U23805 ( .C1(n20918), .C2(n20942), .A(n20862), .B(n20861), .ZN(
        P1_U3149) );
  AOI22_X1 U23806 ( .A1(n20920), .A2(n20867), .B1(n20919), .B2(n20868), .ZN(
        n20864) );
  AOI22_X1 U23807 ( .A1(n20871), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n20870), .B2(n20921), .ZN(n20863) );
  OAI211_X1 U23808 ( .C1(n20924), .C2(n20942), .A(n20864), .B(n20863), .ZN(
        P1_U3150) );
  AOI22_X1 U23809 ( .A1(n20926), .A2(n20867), .B1(n20925), .B2(n20868), .ZN(
        n20866) );
  AOI22_X1 U23810 ( .A1(n20871), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n20870), .B2(n9809), .ZN(n20865) );
  OAI211_X1 U23811 ( .C1(n20932), .C2(n20942), .A(n20866), .B(n20865), .ZN(
        P1_U3151) );
  AOI22_X1 U23812 ( .A1(n20936), .A2(n20868), .B1(n20933), .B2(n20867), .ZN(
        n20873) );
  AOI22_X1 U23813 ( .A1(n20871), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n20870), .B2(n20869), .ZN(n20872) );
  OAI211_X1 U23814 ( .C1(n20874), .C2(n20942), .A(n20873), .B(n20872), .ZN(
        P1_U3152) );
  INV_X1 U23815 ( .A(n20877), .ZN(n20934) );
  OR2_X1 U23816 ( .A1(n20876), .A2(n20875), .ZN(n20878) );
  AND2_X1 U23817 ( .A1(n20878), .A2(n20877), .ZN(n20885) );
  OAI22_X1 U23818 ( .A1(n20885), .A2(n20883), .B1(n20879), .B2(n21042), .ZN(
        n20935) );
  AOI22_X1 U23819 ( .A1(n20881), .A2(n20934), .B1(n20880), .B2(n20935), .ZN(
        n20893) );
  OAI21_X1 U23820 ( .B1(n20884), .B2(n20883), .A(n20882), .ZN(n20886) );
  NAND2_X1 U23821 ( .A1(n20886), .A2(n20885), .ZN(n20887) );
  OAI211_X1 U23822 ( .C1(n20890), .C2(n20889), .A(n20888), .B(n20887), .ZN(
        n20939) );
  AOI22_X1 U23823 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20939), .B1(
        n20928), .B2(n9807), .ZN(n20892) );
  OAI211_X1 U23824 ( .C1(n20894), .C2(n20931), .A(n20893), .B(n20892), .ZN(
        P1_U3153) );
  AOI22_X1 U23825 ( .A1(n20896), .A2(n20934), .B1(n20895), .B2(n20935), .ZN(
        n20899) );
  AOI22_X1 U23826 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20939), .B1(
        n20928), .B2(n9811), .ZN(n20898) );
  OAI211_X1 U23827 ( .C1(n20900), .C2(n20931), .A(n20899), .B(n20898), .ZN(
        P1_U3154) );
  AOI22_X1 U23828 ( .A1(n20902), .A2(n20934), .B1(n20901), .B2(n20935), .ZN(
        n20905) );
  AOI22_X1 U23829 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20939), .B1(
        n20928), .B2(n9813), .ZN(n20904) );
  OAI211_X1 U23830 ( .C1(n20906), .C2(n20931), .A(n20905), .B(n20904), .ZN(
        P1_U3155) );
  AOI22_X1 U23831 ( .A1(n20908), .A2(n20934), .B1(n20907), .B2(n20935), .ZN(
        n20911) );
  AOI22_X1 U23832 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20939), .B1(
        n20938), .B2(n20909), .ZN(n20910) );
  OAI211_X1 U23833 ( .C1(n20912), .C2(n20942), .A(n20911), .B(n20910), .ZN(
        P1_U3156) );
  AOI22_X1 U23834 ( .A1(n20914), .A2(n20934), .B1(n20913), .B2(n20935), .ZN(
        n20917) );
  AOI22_X1 U23835 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20939), .B1(
        n20928), .B2(n20915), .ZN(n20916) );
  OAI211_X1 U23836 ( .C1(n20918), .C2(n20931), .A(n20917), .B(n20916), .ZN(
        P1_U3157) );
  AOI22_X1 U23837 ( .A1(n20920), .A2(n20934), .B1(n20919), .B2(n20935), .ZN(
        n20923) );
  AOI22_X1 U23838 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20939), .B1(
        n20928), .B2(n20921), .ZN(n20922) );
  OAI211_X1 U23839 ( .C1(n20924), .C2(n20931), .A(n20923), .B(n20922), .ZN(
        P1_U3158) );
  AOI22_X1 U23840 ( .A1(n20926), .A2(n20934), .B1(n20925), .B2(n20935), .ZN(
        n20930) );
  AOI22_X1 U23841 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20939), .B1(
        n20928), .B2(n9809), .ZN(n20929) );
  OAI211_X1 U23842 ( .C1(n20932), .C2(n20931), .A(n20930), .B(n20929), .ZN(
        P1_U3159) );
  AOI22_X1 U23843 ( .A1(n20936), .A2(n20935), .B1(n20934), .B2(n20933), .ZN(
        n20941) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20939), .B1(
        n20938), .B2(n20937), .ZN(n20940) );
  OAI211_X1 U23845 ( .C1(n20943), .C2(n20942), .A(n20941), .B(n20940), .ZN(
        P1_U3160) );
  OAI221_X1 U23846 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20946), .C1(n21042), 
        .C2(n20945), .A(n20944), .ZN(P1_U3163) );
  AND2_X1 U23847 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21015), .ZN(
        P1_U3164) );
  AND2_X1 U23848 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21015), .ZN(
        P1_U3165) );
  AND2_X1 U23849 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21015), .ZN(
        P1_U3166) );
  AND2_X1 U23850 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21015), .ZN(
        P1_U3167) );
  AND2_X1 U23851 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21015), .ZN(
        P1_U3168) );
  AND2_X1 U23852 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21015), .ZN(
        P1_U3169) );
  AND2_X1 U23853 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21015), .ZN(
        P1_U3170) );
  AND2_X1 U23854 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21015), .ZN(
        P1_U3171) );
  AND2_X1 U23855 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21015), .ZN(
        P1_U3172) );
  AND2_X1 U23856 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21015), .ZN(
        P1_U3173) );
  AND2_X1 U23857 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21015), .ZN(
        P1_U3174) );
  AND2_X1 U23858 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21015), .ZN(
        P1_U3175) );
  AND2_X1 U23859 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21015), .ZN(
        P1_U3176) );
  AND2_X1 U23860 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21015), .ZN(
        P1_U3177) );
  AND2_X1 U23861 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21015), .ZN(
        P1_U3178) );
  AND2_X1 U23862 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21015), .ZN(
        P1_U3179) );
  AND2_X1 U23863 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21015), .ZN(
        P1_U3180) );
  AND2_X1 U23864 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21015), .ZN(
        P1_U3181) );
  AND2_X1 U23865 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21015), .ZN(
        P1_U3182) );
  AND2_X1 U23866 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21015), .ZN(
        P1_U3183) );
  AND2_X1 U23867 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21015), .ZN(
        P1_U3184) );
  AND2_X1 U23868 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21015), .ZN(
        P1_U3185) );
  AND2_X1 U23869 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21015), .ZN(P1_U3186) );
  AND2_X1 U23870 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21015), .ZN(P1_U3187) );
  AND2_X1 U23871 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21015), .ZN(P1_U3188) );
  AND2_X1 U23872 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21015), .ZN(P1_U3189) );
  AND2_X1 U23873 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21015), .ZN(P1_U3190) );
  AND2_X1 U23874 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21015), .ZN(P1_U3191) );
  AND2_X1 U23875 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21015), .ZN(P1_U3192) );
  AND2_X1 U23876 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21015), .ZN(P1_U3193) );
  NOR2_X1 U23877 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20947) );
  OAI22_X1 U23878 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21230), .B1(n20947), 
        .B2(n21190), .ZN(n20948) );
  OAI21_X1 U23879 ( .B1(n21188), .B2(n20948), .A(n21053), .ZN(n20949) );
  OAI221_X1 U23880 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(P1_STATE_REG_0__SCAN_IN), .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20953), .A(n20949), .ZN(P1_U3194) );
  AOI211_X1 U23881 ( .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(n11877), .A(
        n13206), .B(n21190), .ZN(n20954) );
  AOI22_X1 U23882 ( .A1(n21050), .A2(n20954), .B1(n20951), .B2(n20950), .ZN(
        n20958) );
  INV_X1 U23883 ( .A(n20952), .ZN(n20957) );
  OAI21_X1 U23884 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(NA), .A(n20953), .ZN(
        n20955) );
  AOI211_X1 U23885 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20955), .A(n21013), 
        .B(n20954), .ZN(n20956) );
  OAI22_X1 U23886 ( .A1(NA), .A2(n20958), .B1(n20957), .B2(n20956), .ZN(
        P1_U3196) );
  NAND2_X1 U23887 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21013), .ZN(n21003) );
  INV_X1 U23888 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20959) );
  NAND2_X1 U23889 ( .A1(n21013), .A2(n11877), .ZN(n21005) );
  OAI222_X1 U23890 ( .A1(n21003), .A2(n13461), .B1(n20959), .B2(n21013), .C1(
        n20960), .C2(n21005), .ZN(P1_U3197) );
  INV_X1 U23891 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20961) );
  INV_X1 U23892 ( .A(n21003), .ZN(n20988) );
  INV_X1 U23893 ( .A(n20988), .ZN(n21008) );
  OAI222_X1 U23894 ( .A1(n21005), .A2(n20963), .B1(n20961), .B2(n21013), .C1(
        n20960), .C2(n21008), .ZN(P1_U3198) );
  INV_X1 U23895 ( .A(n21005), .ZN(n20985) );
  INV_X1 U23896 ( .A(n20985), .ZN(n21006) );
  OAI222_X1 U23897 ( .A1(n21003), .A2(n20963), .B1(n20962), .B2(n21013), .C1(
        n13706), .C2(n21006), .ZN(P1_U3199) );
  INV_X1 U23898 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20964) );
  OAI222_X1 U23899 ( .A1(n21006), .A2(n20966), .B1(n20964), .B2(n21013), .C1(
        n13706), .C2(n21008), .ZN(P1_U3200) );
  INV_X1 U23900 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20965) );
  OAI222_X1 U23901 ( .A1(n21008), .A2(n20966), .B1(n20965), .B2(n21013), .C1(
        n20968), .C2(n21006), .ZN(P1_U3201) );
  AOI22_X1 U23902 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n21053), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20985), .ZN(n20967) );
  OAI21_X1 U23903 ( .B1(n20968), .B2(n21003), .A(n20967), .ZN(P1_U3202) );
  AOI22_X1 U23904 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21053), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20988), .ZN(n20969) );
  OAI21_X1 U23905 ( .B1(n15127), .B2(n21005), .A(n20969), .ZN(P1_U3203) );
  INV_X1 U23906 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20970) );
  OAI222_X1 U23907 ( .A1(n21006), .A2(n20972), .B1(n20970), .B2(n21013), .C1(
        n15127), .C2(n21003), .ZN(P1_U3204) );
  AOI22_X1 U23908 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n21053), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20985), .ZN(n20971) );
  OAI21_X1 U23909 ( .B1(n20972), .B2(n21003), .A(n20971), .ZN(P1_U3205) );
  AOI22_X1 U23910 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n21053), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20988), .ZN(n20973) );
  OAI21_X1 U23911 ( .B1(n20975), .B2(n21005), .A(n20973), .ZN(P1_U3206) );
  INV_X1 U23912 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20974) );
  OAI222_X1 U23913 ( .A1(n21008), .A2(n20975), .B1(n20974), .B2(n21013), .C1(
        n20977), .C2(n21005), .ZN(P1_U3207) );
  INV_X1 U23914 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20976) );
  OAI222_X1 U23915 ( .A1(n21008), .A2(n20977), .B1(n20976), .B2(n21013), .C1(
        n10074), .C2(n21005), .ZN(P1_U3208) );
  INV_X1 U23916 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20978) );
  OAI222_X1 U23917 ( .A1(n21008), .A2(n10074), .B1(n20978), .B2(n21013), .C1(
        n20979), .C2(n21006), .ZN(P1_U3209) );
  INV_X1 U23918 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20980) );
  OAI222_X1 U23919 ( .A1(n21006), .A2(n10076), .B1(n20980), .B2(n21013), .C1(
        n20979), .C2(n21003), .ZN(P1_U3210) );
  AOI22_X1 U23920 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n21053), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20985), .ZN(n20981) );
  OAI21_X1 U23921 ( .B1(n10076), .B2(n21003), .A(n20981), .ZN(P1_U3211) );
  AOI22_X1 U23922 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21053), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20988), .ZN(n20982) );
  OAI21_X1 U23923 ( .B1(n20983), .B2(n21005), .A(n20982), .ZN(P1_U3212) );
  INV_X1 U23924 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20984) );
  OAI222_X1 U23925 ( .A1(n21006), .A2(n20987), .B1(n20984), .B2(n21013), .C1(
        n20983), .C2(n21003), .ZN(P1_U3213) );
  AOI22_X1 U23926 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21053), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20985), .ZN(n20986) );
  OAI21_X1 U23927 ( .B1(n20987), .B2(n21003), .A(n20986), .ZN(P1_U3214) );
  AOI22_X1 U23928 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21053), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20988), .ZN(n20989) );
  OAI21_X1 U23929 ( .B1(n20990), .B2(n21005), .A(n20989), .ZN(P1_U3215) );
  INV_X1 U23930 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20991) );
  OAI222_X1 U23931 ( .A1(n21006), .A2(n20992), .B1(n20991), .B2(n21013), .C1(
        n20990), .C2(n21003), .ZN(P1_U3216) );
  INV_X1 U23932 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21174) );
  INV_X1 U23933 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20993) );
  OAI222_X1 U23934 ( .A1(n21006), .A2(n21174), .B1(n20993), .B2(n21013), .C1(
        n20992), .C2(n21003), .ZN(P1_U3217) );
  INV_X1 U23935 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20994) );
  OAI222_X1 U23936 ( .A1(n21008), .A2(n21174), .B1(n20994), .B2(n21013), .C1(
        n20995), .C2(n21005), .ZN(P1_U3218) );
  INV_X1 U23937 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20996) );
  OAI222_X1 U23938 ( .A1(n21006), .A2(n21169), .B1(n20996), .B2(n21013), .C1(
        n20995), .C2(n21003), .ZN(P1_U3219) );
  INV_X1 U23939 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20997) );
  OAI222_X1 U23940 ( .A1(n21008), .A2(n21169), .B1(n20997), .B2(n21013), .C1(
        n21187), .C2(n21005), .ZN(P1_U3220) );
  INV_X1 U23941 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20998) );
  OAI222_X1 U23942 ( .A1(n21008), .A2(n21187), .B1(n20998), .B2(n21013), .C1(
        n21000), .C2(n21005), .ZN(P1_U3221) );
  INV_X1 U23943 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20999) );
  OAI222_X1 U23944 ( .A1(n21008), .A2(n21000), .B1(n20999), .B2(n21013), .C1(
        n21163), .C2(n21005), .ZN(P1_U3222) );
  INV_X1 U23945 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21001) );
  OAI222_X1 U23946 ( .A1(n21008), .A2(n21163), .B1(n21001), .B2(n21013), .C1(
        n21079), .C2(n21005), .ZN(P1_U3223) );
  INV_X1 U23947 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21002) );
  OAI222_X1 U23948 ( .A1(n21006), .A2(n21094), .B1(n21002), .B2(n21013), .C1(
        n21079), .C2(n21003), .ZN(P1_U3224) );
  INV_X1 U23949 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21154) );
  INV_X1 U23950 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n21004) );
  OAI222_X1 U23951 ( .A1(n21005), .A2(n21154), .B1(n21004), .B2(n21013), .C1(
        n21094), .C2(n21003), .ZN(P1_U3225) );
  INV_X1 U23952 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21007) );
  OAI222_X1 U23953 ( .A1(n21008), .A2(n21154), .B1(n21007), .B2(n21013), .C1(
        n21165), .C2(n21006), .ZN(P1_U3226) );
  INV_X1 U23954 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21009) );
  AOI22_X1 U23955 ( .A1(n21013), .A2(n21211), .B1(n21009), .B2(n21053), .ZN(
        P1_U3458) );
  INV_X1 U23956 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21156) );
  INV_X1 U23957 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21010) );
  AOI22_X1 U23958 ( .A1(n21013), .A2(n21156), .B1(n21010), .B2(n21053), .ZN(
        P1_U3459) );
  INV_X1 U23959 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21011) );
  AOI22_X1 U23960 ( .A1(n21013), .A2(n21058), .B1(n21011), .B2(n21053), .ZN(
        P1_U3460) );
  INV_X1 U23961 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21057) );
  INV_X1 U23962 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21012) );
  AOI22_X1 U23963 ( .A1(n21013), .A2(n21057), .B1(n21012), .B2(n21053), .ZN(
        P1_U3461) );
  INV_X1 U23964 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21016) );
  INV_X1 U23965 ( .A(n21017), .ZN(n21014) );
  AOI21_X1 U23966 ( .B1(n21016), .B2(n21015), .A(n21014), .ZN(P1_U3464) );
  OAI21_X1 U23967 ( .B1(n21019), .B2(n21018), .A(n21017), .ZN(P1_U3465) );
  INV_X1 U23968 ( .A(n21032), .ZN(n21035) );
  OAI21_X1 U23969 ( .B1(n21022), .B2(n21021), .A(n21020), .ZN(n21031) );
  NOR2_X1 U23970 ( .A1(n21024), .A2(n21023), .ZN(n21029) );
  INV_X1 U23971 ( .A(n13342), .ZN(n21026) );
  OAI22_X1 U23972 ( .A1(n15320), .A2(n21027), .B1(n21026), .B2(n21025), .ZN(
        n21028) );
  AOI211_X1 U23973 ( .C1(n21031), .C2(n21030), .A(n21029), .B(n21028), .ZN(
        n21033) );
  AOI22_X1 U23974 ( .A1(n21035), .A2(n21034), .B1(n21033), .B2(n21032), .ZN(
        P1_U3475) );
  AOI21_X1 U23975 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21036) );
  AOI22_X1 U23976 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21036), .B2(n13461), .ZN(n21038) );
  AOI22_X1 U23977 ( .A1(n21040), .A2(n21038), .B1(n21156), .B2(n21037), .ZN(
        P1_U3481) );
  OAI21_X1 U23978 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21040), .ZN(n21039) );
  OAI21_X1 U23979 ( .B1(n21040), .B2(n21057), .A(n21039), .ZN(P1_U3482) );
  AOI22_X1 U23980 ( .A1(n21013), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21093), 
        .B2(n21053), .ZN(P1_U3483) );
  AOI211_X1 U23981 ( .C1(n21043), .C2(n21172), .A(n21042), .B(n21041), .ZN(
        n21046) );
  OAI21_X1 U23982 ( .B1(n21046), .B2(n21045), .A(n21044), .ZN(n21052) );
  OAI211_X1 U23983 ( .C1(n21050), .C2(n21049), .A(n21048), .B(n21047), .ZN(
        n21051) );
  MUX2_X1 U23984 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(n21052), .S(n21051), 
        .Z(P1_U3485) );
  INV_X1 U23985 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21054) );
  AOI22_X1 U23986 ( .A1(n21013), .A2(n21081), .B1(n21054), .B2(n21053), .ZN(
        P1_U3486) );
  AOI22_X1 U23987 ( .A1(n21222), .A2(keyinput_g1), .B1(keyinput_g16), .B2(
        n21224), .ZN(n21055) );
  OAI221_X1 U23988 ( .B1(n21222), .B2(keyinput_g1), .C1(n21224), .C2(
        keyinput_g16), .A(n21055), .ZN(n21065) );
  AOI22_X1 U23989 ( .A1(n21058), .A2(keyinput_g49), .B1(keyinput_g48), .B2(
        n21057), .ZN(n21056) );
  OAI221_X1 U23990 ( .B1(n21058), .B2(keyinput_g49), .C1(n21057), .C2(
        keyinput_g48), .A(n21056), .ZN(n21064) );
  AOI22_X1 U23991 ( .A1(n21231), .A2(keyinput_g13), .B1(n21154), .B2(
        keyinput_g53), .ZN(n21059) );
  OAI221_X1 U23992 ( .B1(n21231), .B2(keyinput_g13), .C1(n21154), .C2(
        keyinput_g53), .A(n21059), .ZN(n21063) );
  AOI22_X1 U23993 ( .A1(n21061), .A2(keyinput_g9), .B1(keyinput_g50), .B2(
        n21156), .ZN(n21060) );
  OAI221_X1 U23994 ( .B1(n21061), .B2(keyinput_g9), .C1(n21156), .C2(
        keyinput_g50), .A(n21060), .ZN(n21062) );
  NOR4_X1 U23995 ( .A1(n21065), .A2(n21064), .A3(n21063), .A4(n21062), .ZN(
        n21102) );
  AOI22_X1 U23996 ( .A1(n21215), .A2(keyinput_g26), .B1(n21221), .B2(
        keyinput_g25), .ZN(n21066) );
  OAI221_X1 U23997 ( .B1(n21215), .B2(keyinput_g26), .C1(n21221), .C2(
        keyinput_g25), .A(n21066), .ZN(n21075) );
  AOI22_X1 U23998 ( .A1(n21069), .A2(keyinput_g2), .B1(keyinput_g4), .B2(
        n21068), .ZN(n21067) );
  OAI221_X1 U23999 ( .B1(n21069), .B2(keyinput_g2), .C1(n21068), .C2(
        keyinput_g4), .A(n21067), .ZN(n21074) );
  AOI22_X1 U24000 ( .A1(n21187), .A2(keyinput_g58), .B1(keyinput_g45), .B2(
        n21162), .ZN(n21070) );
  OAI221_X1 U24001 ( .B1(n21187), .B2(keyinput_g58), .C1(n21162), .C2(
        keyinput_g45), .A(n21070), .ZN(n21073) );
  AOI22_X1 U24002 ( .A1(n21209), .A2(keyinput_g14), .B1(n21172), .B2(
        keyinput_g44), .ZN(n21071) );
  OAI221_X1 U24003 ( .B1(n21209), .B2(keyinput_g14), .C1(n21172), .C2(
        keyinput_g44), .A(n21071), .ZN(n21072) );
  NOR4_X1 U24004 ( .A1(n21075), .A2(n21074), .A3(n21073), .A4(n21072), .ZN(
        n21101) );
  AOI22_X1 U24005 ( .A1(n21077), .A2(keyinput_g20), .B1(n21174), .B2(
        keyinput_g61), .ZN(n21076) );
  OAI221_X1 U24006 ( .B1(n21077), .B2(keyinput_g20), .C1(n21174), .C2(
        keyinput_g61), .A(n21076), .ZN(n21087) );
  INV_X1 U24007 ( .A(READY1), .ZN(n21205) );
  AOI22_X1 U24008 ( .A1(n21079), .A2(keyinput_g55), .B1(n21205), .B2(
        keyinput_g36), .ZN(n21078) );
  OAI221_X1 U24009 ( .B1(n21079), .B2(keyinput_g55), .C1(n21205), .C2(
        keyinput_g36), .A(n21078), .ZN(n21086) );
  AOI22_X1 U24010 ( .A1(n21081), .A2(keyinput_g0), .B1(n21188), .B2(
        keyinput_g43), .ZN(n21080) );
  OAI221_X1 U24011 ( .B1(n21081), .B2(keyinput_g0), .C1(n21188), .C2(
        keyinput_g43), .A(n21080), .ZN(n21085) );
  AOI22_X1 U24012 ( .A1(n21211), .A2(keyinput_g51), .B1(n21083), .B2(
        keyinput_g6), .ZN(n21082) );
  OAI221_X1 U24013 ( .B1(n21211), .B2(keyinput_g51), .C1(n21083), .C2(
        keyinput_g6), .A(n21082), .ZN(n21084) );
  NOR4_X1 U24014 ( .A1(n21087), .A2(n21086), .A3(n21085), .A4(n21084), .ZN(
        n21100) );
  AOI22_X1 U24015 ( .A1(n21089), .A2(keyinput_g35), .B1(n21175), .B2(
        keyinput_g22), .ZN(n21088) );
  OAI221_X1 U24016 ( .B1(n21089), .B2(keyinput_g35), .C1(n21175), .C2(
        keyinput_g22), .A(n21088), .ZN(n21098) );
  AOI22_X1 U24017 ( .A1(n21163), .A2(keyinput_g56), .B1(n21165), .B2(
        keyinput_g52), .ZN(n21090) );
  OAI221_X1 U24018 ( .B1(n21163), .B2(keyinput_g56), .C1(n21165), .C2(
        keyinput_g52), .A(n21090), .ZN(n21097) );
  AOI22_X1 U24019 ( .A1(n21191), .A2(keyinput_g5), .B1(keyinput_g11), .B2(
        n21171), .ZN(n21091) );
  OAI221_X1 U24020 ( .B1(n21191), .B2(keyinput_g5), .C1(n21171), .C2(
        keyinput_g11), .A(n21091), .ZN(n21096) );
  AOI22_X1 U24021 ( .A1(n21094), .A2(keyinput_g54), .B1(keyinput_g47), .B2(
        n21093), .ZN(n21092) );
  OAI221_X1 U24022 ( .B1(n21094), .B2(keyinput_g54), .C1(n21093), .C2(
        keyinput_g47), .A(n21092), .ZN(n21095) );
  NOR4_X1 U24023 ( .A1(n21098), .A2(n21097), .A3(n21096), .A4(n21095), .ZN(
        n21099) );
  AND4_X1 U24024 ( .A1(n21102), .A2(n21101), .A3(n21100), .A4(n21099), .ZN(
        n21254) );
  OAI22_X1 U24025 ( .A1(DATAI_5_), .A2(keyinput_g27), .B1(keyinput_g30), .B2(
        DATAI_2_), .ZN(n21103) );
  AOI221_X1 U24026 ( .B1(DATAI_5_), .B2(keyinput_g27), .C1(DATAI_2_), .C2(
        keyinput_g30), .A(n21103), .ZN(n21110) );
  OAI22_X1 U24027 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_g63), .B1(
        DATAI_29_), .B2(keyinput_g3), .ZN(n21104) );
  AOI221_X1 U24028 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .C1(
        keyinput_g3), .C2(DATAI_29_), .A(n21104), .ZN(n21109) );
  OAI22_X1 U24029 ( .A1(DATAI_20_), .A2(keyinput_g12), .B1(
        P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .ZN(n21105) );
  AOI221_X1 U24030 ( .B1(DATAI_20_), .B2(keyinput_g12), .C1(keyinput_g42), 
        .C2(P1_D_C_N_REG_SCAN_IN), .A(n21105), .ZN(n21108) );
  OAI22_X1 U24031 ( .A1(DATAI_0_), .A2(keyinput_g32), .B1(NA), .B2(
        keyinput_g34), .ZN(n21106) );
  AOI221_X1 U24032 ( .B1(DATAI_0_), .B2(keyinput_g32), .C1(keyinput_g34), .C2(
        NA), .A(n21106), .ZN(n21107) );
  NAND4_X1 U24033 ( .A1(n21110), .A2(n21109), .A3(n21108), .A4(n21107), .ZN(
        n21139) );
  OAI22_X1 U24034 ( .A1(DATAI_3_), .A2(keyinput_g29), .B1(keyinput_g37), .B2(
        READY2), .ZN(n21111) );
  AOI221_X1 U24035 ( .B1(DATAI_3_), .B2(keyinput_g29), .C1(READY2), .C2(
        keyinput_g37), .A(n21111), .ZN(n21117) );
  OAI22_X1 U24036 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_g62), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .ZN(n21112) );
  AOI221_X1 U24037 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .C1(
        keyinput_g41), .C2(P1_M_IO_N_REG_SCAN_IN), .A(n21112), .ZN(n21116) );
  OAI22_X1 U24038 ( .A1(DATAI_8_), .A2(keyinput_g24), .B1(keyinput_g28), .B2(
        DATAI_4_), .ZN(n21113) );
  AOI221_X1 U24039 ( .B1(DATAI_8_), .B2(keyinput_g24), .C1(DATAI_4_), .C2(
        keyinput_g28), .A(n21113), .ZN(n21115) );
  XNOR2_X1 U24040 ( .A(P1_CODEFETCH_REG_SCAN_IN), .B(keyinput_g40), .ZN(n21114) );
  NAND4_X1 U24041 ( .A1(n21117), .A2(n21116), .A3(n21115), .A4(n21114), .ZN(
        n21138) );
  OAI22_X1 U24042 ( .A1(DATAI_25_), .A2(keyinput_g7), .B1(DATAI_9_), .B2(
        keyinput_g23), .ZN(n21118) );
  AOI221_X1 U24043 ( .B1(DATAI_25_), .B2(keyinput_g7), .C1(keyinput_g23), .C2(
        DATAI_9_), .A(n21118), .ZN(n21127) );
  OAI22_X1 U24044 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(
        P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .ZN(n21119) );
  AOI221_X1 U24045 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(keyinput_g46), 
        .C2(P1_FLUSH_REG_SCAN_IN), .A(n21119), .ZN(n21126) );
  INV_X1 U24046 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21121) );
  OAI22_X1 U24047 ( .A1(n21214), .A2(keyinput_g8), .B1(n21121), .B2(
        keyinput_g38), .ZN(n21120) );
  AOI221_X1 U24048 ( .B1(n21214), .B2(keyinput_g8), .C1(keyinput_g38), .C2(
        n21121), .A(n21120), .ZN(n21125) );
  OAI22_X1 U24049 ( .A1(n21227), .A2(keyinput_g31), .B1(n21123), .B2(
        keyinput_g39), .ZN(n21122) );
  AOI221_X1 U24050 ( .B1(n21227), .B2(keyinput_g31), .C1(keyinput_g39), .C2(
        n21123), .A(n21122), .ZN(n21124) );
  NAND4_X1 U24051 ( .A1(n21127), .A2(n21126), .A3(n21125), .A4(n21124), .ZN(
        n21137) );
  OAI22_X1 U24052 ( .A1(DATAI_11_), .A2(keyinput_g21), .B1(keyinput_g33), .B2(
        HOLD), .ZN(n21128) );
  AOI221_X1 U24053 ( .B1(DATAI_11_), .B2(keyinput_g21), .C1(HOLD), .C2(
        keyinput_g33), .A(n21128), .ZN(n21135) );
  OAI22_X1 U24054 ( .A1(DATAI_14_), .A2(keyinput_g18), .B1(DATAI_13_), .B2(
        keyinput_g19), .ZN(n21129) );
  AOI221_X1 U24055 ( .B1(DATAI_14_), .B2(keyinput_g18), .C1(keyinput_g19), 
        .C2(DATAI_13_), .A(n21129), .ZN(n21134) );
  OAI22_X1 U24056 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_g59), .B1(
        DATAI_22_), .B2(keyinput_g10), .ZN(n21130) );
  AOI221_X1 U24057 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .C1(
        keyinput_g10), .C2(DATAI_22_), .A(n21130), .ZN(n21133) );
  OAI22_X1 U24058 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_g57), .B1(
        DATAI_17_), .B2(keyinput_g15), .ZN(n21131) );
  AOI221_X1 U24059 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .C1(
        keyinput_g15), .C2(DATAI_17_), .A(n21131), .ZN(n21132) );
  NAND4_X1 U24060 ( .A1(n21135), .A2(n21134), .A3(n21133), .A4(n21132), .ZN(
        n21136) );
  NOR4_X1 U24061 ( .A1(n21139), .A2(n21138), .A3(n21137), .A4(n21136), .ZN(
        n21253) );
  OAI22_X1 U24062 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_f57), .B1(
        keyinput_f40), .B2(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21140) );
  AOI221_X1 U24063 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_f40), .A(n21140), .ZN(n21247)
         );
  OAI22_X1 U24064 ( .A1(DATAI_2_), .A2(keyinput_f30), .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_f42), .ZN(n21141) );
  AOI221_X1 U24065 ( .B1(DATAI_2_), .B2(keyinput_f30), .C1(keyinput_f42), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n21141), .ZN(n21246) );
  AOI22_X1 U24066 ( .A1(DATAI_3_), .A2(keyinput_f29), .B1(DATAI_30_), .B2(
        keyinput_f2), .ZN(n21142) );
  OAI221_X1 U24067 ( .B1(DATAI_3_), .B2(keyinput_f29), .C1(DATAI_30_), .C2(
        keyinput_f2), .A(n21142), .ZN(n21149) );
  AOI22_X1 U24068 ( .A1(keyinput_f49), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        DATAI_17_), .B2(keyinput_f15), .ZN(n21143) );
  OAI221_X1 U24069 ( .B1(keyinput_f49), .B2(P1_BYTEENABLE_REG_1__SCAN_IN), 
        .C1(DATAI_17_), .C2(keyinput_f15), .A(n21143), .ZN(n21148) );
  AOI22_X1 U24070 ( .A1(keyinput_f47), .A2(P1_W_R_N_REG_SCAN_IN), .B1(
        P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .ZN(n21144) );
  OAI221_X1 U24071 ( .B1(keyinput_f47), .B2(P1_W_R_N_REG_SCAN_IN), .C1(
        P1_FLUSH_REG_SCAN_IN), .C2(keyinput_f46), .A(n21144), .ZN(n21147) );
  AOI22_X1 U24072 ( .A1(DATAI_15_), .A2(keyinput_f17), .B1(DATAI_12_), .B2(
        keyinput_f20), .ZN(n21145) );
  OAI221_X1 U24073 ( .B1(DATAI_15_), .B2(keyinput_f17), .C1(DATAI_12_), .C2(
        keyinput_f20), .A(n21145), .ZN(n21146) );
  NOR4_X1 U24074 ( .A1(n21149), .A2(n21148), .A3(n21147), .A4(n21146), .ZN(
        n21152) );
  OAI22_X1 U24075 ( .A1(DATAI_28_), .A2(keyinput_f4), .B1(DATAI_22_), .B2(
        keyinput_f10), .ZN(n21150) );
  AOI221_X1 U24076 ( .B1(DATAI_28_), .B2(keyinput_f4), .C1(keyinput_f10), .C2(
        DATAI_22_), .A(n21150), .ZN(n21151) );
  OAI211_X1 U24077 ( .C1(n21154), .C2(keyinput_f53), .A(n21152), .B(n21151), 
        .ZN(n21153) );
  AOI21_X1 U24078 ( .B1(n21154), .B2(keyinput_f53), .A(n21153), .ZN(n21245) );
  AOI22_X1 U24079 ( .A1(n21157), .A2(keyinput_f27), .B1(keyinput_f50), .B2(
        n21156), .ZN(n21155) );
  OAI221_X1 U24080 ( .B1(n21157), .B2(keyinput_f27), .C1(n21156), .C2(
        keyinput_f50), .A(n21155), .ZN(n21243) );
  INV_X1 U24081 ( .A(keyinput_f48), .ZN(n21159) );
  AOI22_X1 U24082 ( .A1(n21160), .A2(keyinput_f3), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(n21159), .ZN(n21158) );
  OAI221_X1 U24083 ( .B1(n21160), .B2(keyinput_f3), .C1(n21159), .C2(
        P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21158), .ZN(n21242) );
  OAI22_X1 U24084 ( .A1(n21163), .A2(keyinput_f56), .B1(n21162), .B2(
        keyinput_f45), .ZN(n21161) );
  AOI221_X1 U24085 ( .B1(n21163), .B2(keyinput_f56), .C1(keyinput_f45), .C2(
        n21162), .A(n21161), .ZN(n21183) );
  AOI22_X1 U24086 ( .A1(n21166), .A2(keyinput_f24), .B1(n21165), .B2(
        keyinput_f52), .ZN(n21164) );
  OAI221_X1 U24087 ( .B1(n21166), .B2(keyinput_f24), .C1(n21165), .C2(
        keyinput_f52), .A(n21164), .ZN(n21179) );
  AOI22_X1 U24088 ( .A1(n21169), .A2(keyinput_f59), .B1(keyinput_f28), .B2(
        n21168), .ZN(n21167) );
  OAI221_X1 U24089 ( .B1(n21169), .B2(keyinput_f59), .C1(n21168), .C2(
        keyinput_f28), .A(n21167), .ZN(n21178) );
  AOI22_X1 U24090 ( .A1(n21172), .A2(keyinput_f44), .B1(keyinput_f11), .B2(
        n21171), .ZN(n21170) );
  OAI221_X1 U24091 ( .B1(n21172), .B2(keyinput_f44), .C1(n21171), .C2(
        keyinput_f11), .A(n21170), .ZN(n21177) );
  AOI22_X1 U24092 ( .A1(n21175), .A2(keyinput_f22), .B1(n21174), .B2(
        keyinput_f61), .ZN(n21173) );
  OAI221_X1 U24093 ( .B1(n21175), .B2(keyinput_f22), .C1(n21174), .C2(
        keyinput_f61), .A(n21173), .ZN(n21176) );
  NOR4_X1 U24094 ( .A1(n21179), .A2(n21178), .A3(n21177), .A4(n21176), .ZN(
        n21182) );
  XNOR2_X1 U24095 ( .A(P1_READREQUEST_REG_SCAN_IN), .B(keyinput_f38), .ZN(
        n21181) );
  XNOR2_X1 U24096 ( .A(keyinput_f35), .B(BS16), .ZN(n21180) );
  NAND4_X1 U24097 ( .A1(n21183), .A2(n21182), .A3(n21181), .A4(n21180), .ZN(
        n21241) );
  AOI22_X1 U24098 ( .A1(DATAI_14_), .A2(keyinput_f18), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_f55), .ZN(n21184) );
  OAI221_X1 U24099 ( .B1(DATAI_14_), .B2(keyinput_f18), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput_f55), .A(n21184), .ZN(n21195)
         );
  AOI22_X1 U24100 ( .A1(DATAI_25_), .A2(keyinput_f7), .B1(DATAI_11_), .B2(
        keyinput_f21), .ZN(n21185) );
  OAI221_X1 U24101 ( .B1(DATAI_25_), .B2(keyinput_f7), .C1(DATAI_11_), .C2(
        keyinput_f21), .A(n21185), .ZN(n21194) );
  AOI22_X1 U24102 ( .A1(n21188), .A2(keyinput_f43), .B1(n21187), .B2(
        keyinput_f58), .ZN(n21186) );
  OAI221_X1 U24103 ( .B1(n21188), .B2(keyinput_f43), .C1(n21187), .C2(
        keyinput_f58), .A(n21186), .ZN(n21193) );
  AOI22_X1 U24104 ( .A1(n21191), .A2(keyinput_f5), .B1(keyinput_f33), .B2(
        n21190), .ZN(n21189) );
  OAI221_X1 U24105 ( .B1(n21191), .B2(keyinput_f5), .C1(n21190), .C2(
        keyinput_f33), .A(n21189), .ZN(n21192) );
  NOR4_X1 U24106 ( .A1(n21195), .A2(n21194), .A3(n21193), .A4(n21192), .ZN(
        n21239) );
  AOI22_X1 U24107 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_f54), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_f63), .ZN(n21196) );
  OAI221_X1 U24108 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_f54), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_f63), .A(n21196), .ZN(n21203)
         );
  AOI22_X1 U24109 ( .A1(DATAI_26_), .A2(keyinput_f6), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_f62), .ZN(n21197) );
  OAI221_X1 U24110 ( .B1(DATAI_26_), .B2(keyinput_f6), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_f62), .A(n21197), .ZN(n21202)
         );
  AOI22_X1 U24111 ( .A1(keyinput_f41), .A2(P1_M_IO_N_REG_SCAN_IN), .B1(
        DATAI_23_), .B2(keyinput_f9), .ZN(n21198) );
  OAI221_X1 U24112 ( .B1(keyinput_f41), .B2(P1_M_IO_N_REG_SCAN_IN), .C1(
        DATAI_23_), .C2(keyinput_f9), .A(n21198), .ZN(n21201) );
  AOI22_X1 U24113 ( .A1(keyinput_f39), .A2(P1_ADS_N_REG_SCAN_IN), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f0), .ZN(n21199) );
  OAI221_X1 U24114 ( .B1(keyinput_f39), .B2(P1_ADS_N_REG_SCAN_IN), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_f0), .A(n21199), .ZN(n21200)
         );
  NOR4_X1 U24115 ( .A1(n21203), .A2(n21202), .A3(n21201), .A4(n21200), .ZN(
        n21238) );
  AOI22_X1 U24116 ( .A1(n21206), .A2(keyinput_f19), .B1(n21205), .B2(
        keyinput_f36), .ZN(n21204) );
  OAI221_X1 U24117 ( .B1(n21206), .B2(keyinput_f19), .C1(n21205), .C2(
        keyinput_f36), .A(n21204), .ZN(n21219) );
  AOI22_X1 U24118 ( .A1(n21209), .A2(keyinput_f14), .B1(keyinput_f32), .B2(
        n21208), .ZN(n21207) );
  OAI221_X1 U24119 ( .B1(n21209), .B2(keyinput_f14), .C1(n21208), .C2(
        keyinput_f32), .A(n21207), .ZN(n21218) );
  INV_X1 U24120 ( .A(READY2), .ZN(n21212) );
  AOI22_X1 U24121 ( .A1(n21212), .A2(keyinput_f37), .B1(keyinput_f51), .B2(
        n21211), .ZN(n21210) );
  OAI221_X1 U24122 ( .B1(n21212), .B2(keyinput_f37), .C1(n21211), .C2(
        keyinput_f51), .A(n21210), .ZN(n21217) );
  AOI22_X1 U24123 ( .A1(n21215), .A2(keyinput_f26), .B1(n21214), .B2(
        keyinput_f8), .ZN(n21213) );
  OAI221_X1 U24124 ( .B1(n21215), .B2(keyinput_f26), .C1(n21214), .C2(
        keyinput_f8), .A(n21213), .ZN(n21216) );
  NOR4_X1 U24125 ( .A1(n21219), .A2(n21218), .A3(n21217), .A4(n21216), .ZN(
        n21237) );
  AOI22_X1 U24126 ( .A1(n21222), .A2(keyinput_f1), .B1(keyinput_f25), .B2(
        n21221), .ZN(n21220) );
  OAI221_X1 U24127 ( .B1(n21222), .B2(keyinput_f1), .C1(n21221), .C2(
        keyinput_f25), .A(n21220), .ZN(n21235) );
  AOI22_X1 U24128 ( .A1(n21225), .A2(keyinput_f12), .B1(keyinput_f16), .B2(
        n21224), .ZN(n21223) );
  OAI221_X1 U24129 ( .B1(n21225), .B2(keyinput_f12), .C1(n21224), .C2(
        keyinput_f16), .A(n21223), .ZN(n21234) );
  AOI22_X1 U24130 ( .A1(n21228), .A2(keyinput_f23), .B1(keyinput_f31), .B2(
        n21227), .ZN(n21226) );
  OAI221_X1 U24131 ( .B1(n21228), .B2(keyinput_f23), .C1(n21227), .C2(
        keyinput_f31), .A(n21226), .ZN(n21233) );
  AOI22_X1 U24132 ( .A1(n21231), .A2(keyinput_f13), .B1(keyinput_f34), .B2(
        n21230), .ZN(n21229) );
  OAI221_X1 U24133 ( .B1(n21231), .B2(keyinput_f13), .C1(n21230), .C2(
        keyinput_f34), .A(n21229), .ZN(n21232) );
  NOR4_X1 U24134 ( .A1(n21235), .A2(n21234), .A3(n21233), .A4(n21232), .ZN(
        n21236) );
  NAND4_X1 U24135 ( .A1(n21239), .A2(n21238), .A3(n21237), .A4(n21236), .ZN(
        n21240) );
  NOR4_X1 U24136 ( .A1(n21243), .A2(n21242), .A3(n21241), .A4(n21240), .ZN(
        n21244) );
  NAND4_X1 U24137 ( .A1(n21247), .A2(n21246), .A3(n21245), .A4(n21244), .ZN(
        n21249) );
  AOI21_X1 U24138 ( .B1(keyinput_f60), .B2(n21249), .A(keyinput_g60), .ZN(
        n21251) );
  INV_X1 U24139 ( .A(keyinput_f60), .ZN(n21248) );
  AOI21_X1 U24140 ( .B1(n21249), .B2(n21248), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n21250) );
  AOI22_X1 U24141 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n21251), .B1(
        keyinput_g60), .B2(n21250), .ZN(n21252) );
  AOI21_X1 U24142 ( .B1(n21254), .B2(n21253), .A(n21252), .ZN(n21257) );
  AOI22_X1 U24143 ( .A1(n21255), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16855), .ZN(n21256) );
  XNOR2_X1 U24144 ( .A(n21257), .B(n21256), .ZN(U355) );
  AND2_X2 U13692 ( .A1(n14595), .A2(n10680), .ZN(n10743) );
  BUF_X2 U11093 ( .A(n17539), .Z(n9648) );
  CLKBUF_X1 U11097 ( .A(n11911), .Z(n12002) );
  CLKBUF_X2 U11113 ( .A(n10444), .Z(n14596) );
  CLKBUF_X1 U11119 ( .A(n14436), .Z(n9640) );
  CLKBUF_X1 U11131 ( .A(n10525), .Z(n10526) );
  CLKBUF_X1 U11135 ( .A(n11333), .Z(n11336) );
  CLKBUF_X1 U11153 ( .A(n11882), .Z(n15302) );
  CLKBUF_X1 U11172 ( .A(n10502), .Z(n10503) );
  CLKBUF_X1 U11180 ( .A(n15572), .Z(n15584) );
  CLKBUF_X1 U11192 ( .A(n11271), .Z(n9663) );
  AND2_X1 U11193 ( .A1(n9824), .A2(n15868), .ZN(n16491) );
  CLKBUF_X1 U11233 ( .A(n16845), .Z(n16850) );
  OR3_X1 U11433 ( .A1(n17713), .A2(n18987), .A3(n18510), .ZN(n21258) );
endmodule

