

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9731, n9732, n9733, n9734, n9735, n9736, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9770, n9771, n9772, n9773, n9774, n9776, n9777, n9778, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065;

  OAI21_X1 U11175 ( .B1(n20423), .B2(n20443), .A(n20660), .ZN(n20445) );
  INV_X1 U11176 ( .A(n20948), .ZN(n20955) );
  INV_X1 U11177 ( .A(n18076), .ZN(n18005) );
  INV_X1 U11178 ( .A(n20927), .ZN(n20954) );
  NOR2_X1 U11179 ( .A1(n20608), .A2(n20655), .ZN(n20699) );
  NAND2_X1 U11180 ( .A1(n13605), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13658) );
  AND4_X1 U11181 ( .A1(n11216), .A2(n11221), .A3(n11217), .A4(n11218), .ZN(
        n10547) );
  OR2_X1 U11182 ( .A1(n13453), .A2(n15172), .ZN(n13454) );
  AND2_X1 U11183 ( .A1(n10426), .A2(n10423), .ZN(n10954) );
  NAND2_X1 U11184 ( .A1(n11776), .A2(n20166), .ZN(n11879) );
  NOR2_X2 U11185 ( .A1(n19375), .A2(n19359), .ZN(n12885) );
  CLKBUF_X1 U11186 ( .A(n16267), .Z(n9761) );
  CLKBUF_X2 U11188 ( .A(n11455), .Z(n12982) );
  NOR2_X1 U11189 ( .A1(n20181), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11456) );
  CLKBUF_X2 U11190 ( .A(n12127), .Z(n13723) );
  INV_X1 U11191 ( .A(n13639), .ZN(n13541) );
  NAND2_X2 U11192 ( .A1(n16374), .A2(n11015), .ZN(n16229) );
  NAND2_X1 U11193 ( .A1(n11179), .A2(n11015), .ZN(n16217) );
  INV_X1 U11194 ( .A(n9732), .ZN(n18335) );
  BUF_X2 U11195 ( .A(n12817), .Z(n18342) );
  NAND2_X1 U11196 ( .A1(n11180), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16221) );
  INV_X4 U11197 ( .A(n13711), .ZN(n13697) );
  AND2_X1 U11200 ( .A1(n12031), .A2(n12041), .ZN(n12127) );
  AND2_X1 U11201 ( .A1(n12042), .A2(n15532), .ZN(n13564) );
  AND2_X1 U11202 ( .A1(n12042), .A2(n15532), .ZN(n9777) );
  CLKBUF_X1 U11203 ( .A(n13610), .Z(n9745) );
  CLKBUF_X1 U11204 ( .A(n19521), .Z(n9731) );
  NOR2_X1 U11205 ( .A1(n19800), .A2(n19489), .ZN(n19521) );
  INV_X1 U11206 ( .A(n12104), .ZN(n13717) );
  AND2_X1 U11207 ( .A1(n12042), .A2(n15532), .ZN(n9776) );
  CLKBUF_X2 U11208 ( .A(n9774), .Z(n13522) );
  INV_X1 U11209 ( .A(n16229), .ZN(n11327) );
  BUF_X1 U11210 ( .A(n12566), .Z(n12664) );
  AND2_X1 U11211 ( .A1(n12458), .A2(n9951), .ZN(n10523) );
  NAND2_X1 U11212 ( .A1(n17289), .A2(n11361), .ZN(n16219) );
  NOR2_X1 U11213 ( .A1(n18524), .A2(n12829), .ZN(n12830) );
  INV_X1 U11215 ( .A(n20166), .ZN(n9742) );
  INV_X1 U11216 ( .A(n11798), .ZN(n11025) );
  NAND2_X1 U11217 ( .A1(n9797), .A2(n9858), .ZN(n10199) );
  INV_X1 U11218 ( .A(n11894), .ZN(n11864) );
  NOR2_X1 U11219 ( .A1(n17484), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12810) );
  CLKBUF_X2 U11220 ( .A(n12743), .Z(n18340) );
  OR2_X1 U11221 ( .A1(n14419), .A2(n14417), .ZN(n20938) );
  INV_X1 U11222 ( .A(n14878), .ZN(n12594) );
  AND2_X1 U11223 ( .A1(n10505), .A2(n10504), .ZN(n15367) );
  BUF_X1 U11224 ( .A(n15537), .Z(n9782) );
  OR2_X1 U11225 ( .A1(n14009), .A2(n14008), .ZN(n10239) );
  AND2_X1 U11226 ( .A1(n10323), .A2(n10321), .ZN(n16661) );
  BUF_X1 U11227 ( .A(n16865), .Z(n16866) );
  NAND2_X1 U11228 ( .A1(n11112), .A2(n11113), .ZN(n11123) );
  INV_X2 U11229 ( .A(n18865), .ZN(n18851) );
  INV_X1 U11230 ( .A(n20938), .ZN(n20959) );
  AND2_X2 U11231 ( .A1(n14740), .A2(n12632), .ZN(n14692) );
  BUF_X1 U11232 ( .A(n12556), .Z(n14391) );
  INV_X1 U11233 ( .A(n21287), .ZN(n21289) );
  AND2_X1 U11234 ( .A1(n16855), .A2(n9820), .ZN(n16684) );
  AND2_X1 U11235 ( .A1(n16855), .A2(n9825), .ZN(n16734) );
  NAND2_X2 U11236 ( .A1(n11701), .A2(n17082), .ZN(n17225) );
  NAND2_X1 U11237 ( .A1(n10440), .A2(n13990), .ZN(n17283) );
  OAI21_X1 U11238 ( .B1(n20138), .B2(n20152), .A(n20660), .ZN(n20186) );
  INV_X1 U11239 ( .A(n20580), .ZN(n20553) );
  INV_X1 U11240 ( .A(n18017), .ZN(n18043) );
  OR3_X1 U11241 ( .A1(n10907), .A2(n10908), .A3(n10424), .ZN(n18391) );
  INV_X1 U11242 ( .A(n10946), .ZN(n19375) );
  NAND2_X1 U11243 ( .A1(n19775), .A2(n19214), .ZN(n19270) );
  INV_X1 U11244 ( .A(n20914), .ZN(n20907) );
  NAND2_X1 U11245 ( .A1(n20526), .A2(n20294), .ZN(n20644) );
  INV_X2 U11246 ( .A(n20863), .ZN(n20862) );
  NOR2_X1 U11247 ( .A1(n12806), .A2(n12805), .ZN(n18510) );
  NOR2_X1 U11248 ( .A1(n12763), .A2(n12762), .ZN(n18524) );
  OR2_X2 U11249 ( .A1(n19787), .A2(n10865), .ZN(n9732) );
  INV_X1 U11250 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21645) );
  OR2_X2 U11251 ( .A1(n12825), .A2(n12824), .ZN(n9733) );
  AND2_X1 U11252 ( .A1(n10134), .A2(n17635), .ZN(n9734) );
  AND2_X2 U11253 ( .A1(n10399), .A2(n10379), .ZN(n9735) );
  INV_X4 U11254 ( .A(n13722), .ZN(n13666) );
  INV_X1 U11255 ( .A(n20166), .ZN(n11889) );
  CLKBUF_X3 U11256 ( .A(n11025), .Z(n20166) );
  INV_X1 U11257 ( .A(n15257), .ZN(n10742) );
  MUX2_X1 U11259 ( .A(n14389), .B(n12566), .S(n14580), .Z(n14395) );
  INV_X2 U11260 ( .A(n16356), .ZN(n9771) );
  NOR2_X2 U11261 ( .A1(n10484), .A2(n10481), .ZN(n12701) );
  AND2_X4 U11262 ( .A1(n12530), .A2(n12529), .ZN(n15557) );
  NAND2_X2 U11263 ( .A1(n11099), .A2(n11098), .ZN(n11127) );
  NAND4_X4 U11264 ( .A1(n12175), .A2(n12174), .A3(n12173), .A4(n12172), .ZN(
        n12184) );
  NOR2_X2 U11265 ( .A1(n12952), .A2(n12951), .ZN(n17143) );
  INV_X1 U11266 ( .A(n9761), .ZN(n9736) );
  NAND2_X1 U11267 ( .A1(n11171), .A2(n17335), .ZN(n16352) );
  AND2_X2 U11268 ( .A1(n11133), .A2(n10776), .ZN(n17281) );
  NOR2_X2 U11269 ( .A1(n12853), .A2(n12943), .ZN(n13096) );
  OR2_X2 U11270 ( .A1(n16408), .A2(n16407), .ZN(n10705) );
  AND2_X4 U11271 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15521) );
  AOI21_X1 U11272 ( .B1(n14467), .B2(n16899), .A(n9882), .ZN(n10830) );
  AND2_X2 U11273 ( .A1(n12839), .A2(n10211), .ZN(n12840) );
  NOR2_X1 U11278 ( .A1(n17484), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9743) );
  NOR2_X1 U11279 ( .A1(n17484), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9744) );
  BUF_X4 U11280 ( .A(n12810), .Z(n18315) );
  NOR2_X2 U11281 ( .A1(n15203), .A2(n12457), .ZN(n12458) );
  AOI21_X2 U11282 ( .B1(n10326), .B2(n9796), .A(n19836), .ZN(n18392) );
  BUF_X8 U11283 ( .A(n13610), .Z(n9746) );
  AND2_X2 U11284 ( .A1(n12042), .A2(n12036), .ZN(n13610) );
  OAI21_X1 U11285 ( .B1(n13156), .B2(n10529), .A(n10527), .ZN(n12393) );
  INV_X1 U11286 ( .A(n12807), .ZN(n9747) );
  NOR2_X2 U11287 ( .A1(n10869), .A2(n10860), .ZN(n10901) );
  NAND2_X2 U11288 ( .A1(n19953), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10869) );
  AND2_X2 U11289 ( .A1(n12197), .A2(n12196), .ZN(n12237) );
  NAND2_X2 U11290 ( .A1(n10199), .A2(n10198), .ZN(n11686) );
  AOI21_X1 U11291 ( .B1(n12995), .B2(n17221), .A(n12996), .ZN(n12997) );
  AND2_X1 U11292 ( .A1(n10078), .A2(n10076), .ZN(n17163) );
  NAND2_X1 U11293 ( .A1(n10316), .A2(n9955), .ZN(n17092) );
  XNOR2_X1 U11294 ( .A(n10179), .B(n12728), .ZN(n12995) );
  AND2_X1 U11295 ( .A1(n10120), .A2(n16743), .ZN(n16745) );
  XNOR2_X1 U11296 ( .A(n9976), .B(n9850), .ZN(n17016) );
  AND2_X1 U11297 ( .A1(n10269), .A2(n10272), .ZN(n16765) );
  NAND2_X2 U11298 ( .A1(n9975), .A2(n11342), .ZN(n10272) );
  OR2_X1 U11299 ( .A1(n17025), .A2(n9977), .ZN(n9976) );
  OR2_X1 U11300 ( .A1(n15084), .A2(n15082), .ZN(n15086) );
  NAND2_X1 U11301 ( .A1(n9983), .A2(n9982), .ZN(n10271) );
  NAND3_X2 U11302 ( .A1(n9788), .A2(n15191), .A3(n9911), .ZN(n10143) );
  NOR2_X1 U11303 ( .A1(n15659), .A2(n15638), .ZN(n15637) );
  NOR3_X1 U11304 ( .A1(n15659), .A2(n10764), .A3(n15638), .ZN(n15623) );
  CLKBUF_X1 U11305 ( .A(n15657), .Z(n15658) );
  CLKBUF_X1 U11306 ( .A(n14762), .Z(n14763) );
  INV_X1 U11307 ( .A(n11290), .ZN(n10549) );
  NAND2_X1 U11308 ( .A1(n15798), .A2(n9861), .ZN(n12010) );
  NAND2_X1 U11309 ( .A1(n10245), .A2(n10243), .ZN(n16434) );
  NOR2_X1 U11310 ( .A1(n15573), .A2(n15574), .ZN(n21381) );
  NOR2_X1 U11311 ( .A1(n13145), .A2(n15575), .ZN(n21539) );
  AND4_X1 U11312 ( .A1(n11223), .A2(n10835), .A3(n11222), .A4(n11215), .ZN(
        n9836) );
  NAND2_X1 U11313 ( .A1(n13555), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13603) );
  NAND2_X1 U11314 ( .A1(n12610), .A2(n12609), .ZN(n14820) );
  AND2_X1 U11315 ( .A1(n11154), .A2(n11152), .ZN(n11265) );
  AND2_X1 U11316 ( .A1(n10108), .A2(n11146), .ZN(n20390) );
  AND2_X1 U11317 ( .A1(n11154), .A2(n11147), .ZN(n11266) );
  NAND2_X1 U11318 ( .A1(n12594), .A2(n10599), .ZN(n14841) );
  INV_X1 U11319 ( .A(n19013), .ZN(n18999) );
  AND2_X1 U11320 ( .A1(n10485), .A2(n14486), .ZN(n12691) );
  CLKBUF_X2 U11321 ( .A(n14171), .Z(n17320) );
  XNOR2_X1 U11322 ( .A(n12297), .B(n12296), .ZN(n13147) );
  AOI22_X1 U11323 ( .A1(n19816), .A2(n19811), .B1(n19810), .B2(n19817), .ZN(
        n19822) );
  INV_X1 U11324 ( .A(n17281), .ZN(n14052) );
  NAND2_X1 U11325 ( .A1(n12393), .A2(n12272), .ZN(n12297) );
  NAND2_X1 U11326 ( .A1(n11817), .A2(n11777), .ZN(n11812) );
  OR2_X1 U11327 ( .A1(n12838), .A2(n12837), .ZN(n12839) );
  INV_X4 U11329 ( .A(n9756), .ZN(n9758) );
  NOR2_X1 U11330 ( .A1(n10842), .A2(n17764), .ZN(n10840) );
  AND2_X1 U11331 ( .A1(n11069), .A2(n11695), .ZN(n11108) );
  INV_X2 U11332 ( .A(n11640), .ZN(n11647) );
  NAND2_X1 U11333 ( .A1(n18399), .A2(n18391), .ZN(n10948) );
  INV_X1 U11335 ( .A(n12186), .ZN(n14961) );
  INV_X1 U11336 ( .A(n12891), .ZN(n18536) );
  AND3_X1 U11338 ( .A1(n11185), .A2(n11184), .A3(n11183), .ZN(n11436) );
  NAND4_X1 U11339 ( .A1(n11199), .A2(n11198), .A3(n11197), .A4(n11196), .ZN(
        n11445) );
  AND3_X1 U11340 ( .A1(n10837), .A2(n9839), .A3(n10806), .ZN(n12178) );
  NOR2_X1 U11341 ( .A1(n12052), .A2(n12051), .ZN(n12068) );
  INV_X1 U11342 ( .A(n11434), .ZN(n11163) );
  INV_X2 U11343 ( .A(n20161), .ZN(n9748) );
  INV_X1 U11344 ( .A(n20181), .ZN(n9749) );
  INV_X1 U11345 ( .A(n16225), .ZN(n11328) );
  NAND2_X2 U11346 ( .A1(n16374), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16225) );
  INV_X1 U11347 ( .A(n16215), .ZN(n11494) );
  INV_X1 U11348 ( .A(n16221), .ZN(n11329) );
  BUF_X2 U11349 ( .A(n15537), .Z(n9781) );
  CLKBUF_X2 U11350 ( .A(n12133), .Z(n13693) );
  CLKBUF_X2 U11351 ( .A(n12743), .Z(n18284) );
  BUF_X2 U11352 ( .A(n12241), .Z(n13647) );
  CLKBUF_X2 U11353 ( .A(n13662), .Z(n13718) );
  INV_X4 U11354 ( .A(n13687), .ZN(n13646) );
  CLKBUF_X1 U11355 ( .A(n13322), .Z(n9773) );
  BUF_X2 U11356 ( .A(n10901), .Z(n18321) );
  INV_X2 U11358 ( .A(n16219), .ZN(n11524) );
  CLKBUF_X3 U11359 ( .A(n16266), .Z(n16377) );
  CLKBUF_X2 U11360 ( .A(n10901), .Z(n18212) );
  INV_X2 U11361 ( .A(n16340), .ZN(n11164) );
  INV_X2 U11362 ( .A(n13231), .ZN(n12160) );
  AND2_X2 U11363 ( .A1(n12031), .A2(n12030), .ZN(n12241) );
  CLKBUF_X2 U11364 ( .A(n12104), .Z(n13614) );
  NOR2_X1 U11365 ( .A1(n10868), .A2(n10860), .ZN(n12817) );
  NAND2_X2 U11366 ( .A1(n12041), .A2(n10744), .ZN(n13687) );
  NAND2_X1 U11367 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10865) );
  NOR2_X4 U11368 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11169) );
  INV_X4 U11369 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11015) );
  AND2_X1 U11370 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15532) );
  AOI21_X1 U11371 ( .B1(n10107), .B2(n10128), .A(n10106), .ZN(n10105) );
  AOI21_X1 U11372 ( .B1(n10127), .B2(n10128), .A(n9808), .ZN(n10421) );
  NOR2_X1 U11373 ( .A1(n10165), .A2(n9993), .ZN(n10149) );
  XNOR2_X1 U11374 ( .A(n10465), .B(n11896), .ZN(n14467) );
  AND2_X1 U11375 ( .A1(n10518), .A2(n10151), .ZN(n17120) );
  AND2_X1 U11376 ( .A1(n17096), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9993) );
  AOI21_X1 U11377 ( .B1(n17054), .B2(n16939), .A(n16739), .ZN(n16740) );
  OAI21_X1 U11378 ( .B1(n16765), .B2(n9920), .A(n10200), .ZN(n17096) );
  XNOR2_X1 U11379 ( .A(n16735), .B(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17054) );
  NAND2_X1 U11380 ( .A1(n16734), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16715) );
  INV_X1 U11381 ( .A(n10638), .ZN(n16646) );
  NAND2_X1 U11382 ( .A1(n10518), .A2(n17091), .ZN(n10128) );
  AND2_X1 U11383 ( .A1(n10314), .A2(n10700), .ZN(n17087) );
  NAND2_X1 U11384 ( .A1(n10272), .A2(n10271), .ZN(n16804) );
  NAND2_X1 U11385 ( .A1(n10272), .A2(n10104), .ZN(n10518) );
  NAND2_X1 U11386 ( .A1(n10118), .A2(n10117), .ZN(n10120) );
  AND2_X1 U11387 ( .A1(n10670), .A2(n10667), .ZN(n10666) );
  INV_X1 U11388 ( .A(n14910), .ZN(n15093) );
  OAI21_X1 U11389 ( .B1(n16783), .B2(n10350), .A(n10347), .ZN(n16792) );
  AOI21_X1 U11390 ( .B1(n16783), .B2(n10355), .A(n16816), .ZN(n16808) );
  NAND2_X1 U11391 ( .A1(n10654), .A2(n10016), .ZN(n10554) );
  NAND2_X1 U11392 ( .A1(n16825), .A2(n11991), .ZN(n16783) );
  NAND2_X1 U11393 ( .A1(n10175), .A2(n10174), .ZN(n14910) );
  NAND2_X1 U11394 ( .A1(n10654), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15126) );
  AND2_X1 U11395 ( .A1(n10271), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10104) );
  AND2_X1 U11396 ( .A1(n14563), .A2(n10668), .ZN(n10667) );
  AND2_X1 U11397 ( .A1(n16709), .A2(n16710), .ZN(n17024) );
  NOR2_X1 U11398 ( .A1(n16709), .A2(n16710), .ZN(n17025) );
  AOI211_X1 U11399 ( .C1(n16978), .C2(n17260), .A(n16977), .B(n16976), .ZN(
        n16982) );
  NAND2_X1 U11400 ( .A1(n15095), .A2(n15257), .ZN(n10654) );
  NAND2_X1 U11401 ( .A1(n10148), .A2(n9910), .ZN(n10234) );
  OR2_X1 U11402 ( .A1(n10516), .A2(n9990), .ZN(n9983) );
  NAND2_X1 U11403 ( .A1(n15142), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15095) );
  AOI21_X1 U11404 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16503), .A(n16389), .ZN(
        n16390) );
  NAND2_X1 U11405 ( .A1(n9988), .A2(n9989), .ZN(n9985) );
  OR2_X1 U11406 ( .A1(n15623), .A2(n15622), .ZN(n16665) );
  AND2_X1 U11407 ( .A1(n10203), .A2(n10779), .ZN(n10126) );
  AND2_X1 U11408 ( .A1(n11341), .A2(n9987), .ZN(n11342) );
  MUX2_X1 U11409 ( .A(n14395), .B(n14394), .S(n14393), .Z(n14509) );
  AND2_X1 U11410 ( .A1(n15191), .A2(n15190), .ZN(n15265) );
  INV_X1 U11411 ( .A(n20492), .ZN(n20509) );
  NAND2_X1 U11412 ( .A1(n10225), .A2(n10224), .ZN(n10228) );
  AND2_X1 U11413 ( .A1(n11338), .A2(n16870), .ZN(n11339) );
  NOR2_X1 U11414 ( .A1(n20422), .A2(n10205), .ZN(n20423) );
  NAND2_X1 U11415 ( .A1(n16413), .A2(n16412), .ZN(n16411) );
  AOI22_X1 U11416 ( .A1(n20428), .A2(n20427), .B1(n20426), .B2(n20425), .ZN(
        n20444) );
  AND2_X1 U11417 ( .A1(n20420), .A2(n20802), .ZN(n20428) );
  OAI211_X1 U11418 ( .C1(n21500), .C2(n21474), .A(n21547), .B(n21473), .ZN(
        n21502) );
  AND2_X1 U11419 ( .A1(n10635), .A2(n11314), .ZN(n10124) );
  XNOR2_X1 U11420 ( .A(n11340), .B(n11894), .ZN(n16867) );
  NAND2_X1 U11421 ( .A1(n10676), .A2(n17229), .ZN(n10675) );
  NAND2_X1 U11422 ( .A1(n16919), .A2(n17228), .ZN(n10150) );
  NAND2_X1 U11423 ( .A1(n10678), .A2(n10679), .ZN(n16901) );
  OAI211_X1 U11424 ( .C1(n21288), .C2(n21474), .A(n21547), .B(n21261), .ZN(
        n21291) );
  AOI22_X1 U11425 ( .A1(n21472), .A2(n21469), .B1(n21467), .B2(n21466), .ZN(
        n21506) );
  OAI211_X1 U11426 ( .C1(n20305), .C2(n20320), .A(n20660), .B(n20304), .ZN(
        n20323) );
  OR2_X1 U11427 ( .A1(n14946), .A2(n14945), .ZN(n14948) );
  NOR2_X2 U11428 ( .A1(n12850), .A2(n10138), .ZN(n17633) );
  OAI211_X1 U11429 ( .C1(n20366), .C2(n20365), .A(n20660), .B(n20364), .ZN(
        n20385) );
  OAI211_X1 U11430 ( .C1(n21569), .C2(n21548), .A(n21547), .B(n21546), .ZN(
        n21573) );
  OAI21_X1 U11431 ( .B1(n10260), .B2(n12430), .A(n17540), .ZN(n10257) );
  XNOR2_X1 U11432 ( .A(n11337), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16870) );
  NAND2_X1 U11433 ( .A1(n16422), .A2(n16237), .ZN(n16418) );
  NAND2_X1 U11434 ( .A1(n16937), .A2(n11894), .ZN(n11734) );
  OAI21_X1 U11435 ( .B1(n21222), .B2(n21207), .A(n21547), .ZN(n21225) );
  OR2_X1 U11436 ( .A1(n10523), .A2(n15257), .ZN(n10399) );
  NAND2_X1 U11437 ( .A1(n20526), .A2(n20801), .ZN(n20580) );
  NAND2_X1 U11438 ( .A1(n12401), .A2(n21023), .ZN(n10369) );
  AND2_X1 U11439 ( .A1(n14335), .A2(n12400), .ZN(n15294) );
  INV_X1 U11440 ( .A(n21132), .ZN(n21135) );
  NAND2_X1 U11441 ( .A1(n10158), .A2(n10156), .ZN(n15202) );
  NOR2_X2 U11442 ( .A1(n20608), .A2(n20450), .ZN(n20470) );
  NOR2_X2 U11443 ( .A1(n20449), .A2(n20450), .ZN(n20508) );
  NOR2_X2 U11444 ( .A1(n20655), .A2(n20396), .ZN(n20417) );
  NOR2_X2 U11445 ( .A1(n20450), .A2(n20396), .ZN(n20246) );
  INV_X1 U11446 ( .A(n20449), .ZN(n20526) );
  INV_X1 U11447 ( .A(n21631), .ZN(n21638) );
  INV_X1 U11448 ( .A(n21381), .ZN(n21437) );
  OR2_X1 U11449 ( .A1(n20199), .A2(n20198), .ZN(n20608) );
  OR2_X1 U11450 ( .A1(n20199), .A2(n20133), .ZN(n20449) );
  NOR2_X2 U11451 ( .A1(n21175), .A2(n21140), .ZN(n21196) );
  NOR2_X2 U11452 ( .A1(n21175), .A2(n21436), .ZN(n21224) );
  NAND2_X1 U11453 ( .A1(n20199), .A2(n20198), .ZN(n20396) );
  NAND2_X1 U11454 ( .A1(n13196), .A2(n13195), .ZN(n14862) );
  NAND2_X1 U11455 ( .A1(n16434), .A2(n16428), .ZN(n16236) );
  NAND2_X1 U11456 ( .A1(n21381), .A2(n21326), .ZN(n21380) );
  AND2_X1 U11457 ( .A1(n9970), .A2(n11313), .ZN(n11317) );
  AND2_X1 U11458 ( .A1(n12454), .A2(n15214), .ZN(n15193) );
  AND2_X1 U11459 ( .A1(n10157), .A2(n10032), .ZN(n10156) );
  NAND2_X1 U11460 ( .A1(n15573), .A2(n13145), .ZN(n21175) );
  CLKBUF_X1 U11461 ( .A(n18718), .Z(n18766) );
  AND2_X1 U11462 ( .A1(n13146), .A2(n13162), .ZN(n14283) );
  NAND2_X1 U11463 ( .A1(n21539), .A2(n21302), .ZN(n21631) );
  NAND2_X1 U11464 ( .A1(n10507), .A2(n10506), .ZN(n10505) );
  NAND2_X1 U11465 ( .A1(n10414), .A2(n12372), .ZN(n15293) );
  NOR2_X1 U11466 ( .A1(n18654), .A2(n17757), .ZN(n17756) );
  NAND2_X1 U11467 ( .A1(n21539), .A2(n21538), .ZN(n21642) );
  NAND3_X1 U11468 ( .A1(n14211), .A2(n10706), .A3(n14212), .ZN(n10245) );
  AND3_X1 U11469 ( .A1(n11272), .A2(n11273), .A3(n9880), .ZN(n10833) );
  OR2_X1 U11470 ( .A1(n18909), .A2(n19120), .ZN(n18819) );
  NOR2_X1 U11471 ( .A1(n13145), .A2(n21229), .ZN(n21303) );
  NOR2_X1 U11472 ( .A1(n11158), .A2(n11157), .ZN(n11159) );
  AND2_X1 U11473 ( .A1(n12368), .A2(n15226), .ZN(n12454) );
  OAI21_X2 U11474 ( .B1(n14180), .B2(n14179), .A(n14198), .ZN(n20817) );
  AND2_X1 U11475 ( .A1(n10812), .A2(n9941), .ZN(n15192) );
  AND2_X1 U11476 ( .A1(n10360), .A2(n10359), .ZN(n18909) );
  NAND2_X1 U11477 ( .A1(n10812), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15226) );
  XNOR2_X1 U11478 ( .A(n10812), .B(n21858), .ZN(n15183) );
  XNOR2_X1 U11479 ( .A(n12369), .B(n12409), .ZN(n13181) );
  AOI22_X1 U11480 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20390), .B1(
        n20487), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11217) );
  INV_X1 U11481 ( .A(n14820), .ZN(n10604) );
  NAND2_X1 U11482 ( .A1(n18877), .A2(n10213), .ZN(n19149) );
  INV_X1 U11483 ( .A(n20363), .ZN(n20359) );
  NAND2_X1 U11484 ( .A1(n10176), .A2(n10747), .ZN(n12375) );
  INV_X1 U11485 ( .A(n20195), .ZN(n20190) );
  NOR2_X1 U11486 ( .A1(n18684), .A2(n17780), .ZN(n17779) );
  AND2_X1 U11487 ( .A1(n12692), .A2(n21047), .ZN(n21030) );
  NAND2_X1 U11488 ( .A1(n12373), .A2(n10033), .ZN(n12374) );
  NAND3_X1 U11489 ( .A1(n10747), .A2(n10017), .A3(n21229), .ZN(n10264) );
  INV_X1 U11490 ( .A(n14841), .ZN(n12610) );
  NAND2_X1 U11491 ( .A1(n10018), .A2(n12298), .ZN(n10033) );
  AND2_X1 U11492 ( .A1(n10747), .A2(n21229), .ZN(n10375) );
  AND2_X1 U11493 ( .A1(n11138), .A2(n14052), .ZN(n11152) );
  AND2_X1 U11494 ( .A1(n10018), .A2(n9904), .ZN(n10017) );
  AND2_X1 U11495 ( .A1(n14176), .A2(n14197), .ZN(n14180) );
  NAND2_X2 U11496 ( .A1(n17734), .A2(n9937), .ZN(n19009) );
  AND2_X1 U11497 ( .A1(n15994), .A2(n14052), .ZN(n11155) );
  NAND2_X1 U11498 ( .A1(n10015), .A2(n10014), .ZN(n10018) );
  NOR2_X2 U11499 ( .A1(n18510), .A2(n19012), .ZN(n18921) );
  CLKBUF_X1 U11500 ( .A(n15564), .Z(n9770) );
  NAND2_X1 U11501 ( .A1(n12691), .A2(n12681), .ZN(n21008) );
  AND2_X1 U11502 ( .A1(n12691), .A2(n15542), .ZN(n15396) );
  OR2_X1 U11503 ( .A1(n12691), .A2(n21051), .ZN(n21047) );
  NAND2_X1 U11504 ( .A1(n13511), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13553) );
  NAND2_X1 U11505 ( .A1(n14175), .A2(n14174), .ZN(n14197) );
  XNOR2_X1 U11506 ( .A(n17283), .B(n14177), .ZN(n14008) );
  AND2_X1 U11507 ( .A1(n11131), .A2(n11133), .ZN(n11146) );
  AND2_X1 U11508 ( .A1(n18481), .A2(n9950), .ZN(n18432) );
  NAND2_X1 U11509 ( .A1(n10023), .A2(n10376), .ZN(n10021) );
  OAI21_X1 U11510 ( .B1(n14171), .B2(n14206), .A(n14170), .ZN(n14175) );
  NOR2_X2 U11511 ( .A1(n19822), .A2(n19836), .ZN(n12934) );
  OR2_X1 U11512 ( .A1(n12297), .A2(n12296), .ZN(n12298) );
  OR2_X2 U11513 ( .A1(n14086), .A2(n17510), .ZN(n20873) );
  XNOR2_X1 U11514 ( .A(n12385), .B(n13154), .ZN(n21139) );
  NAND2_X1 U11515 ( .A1(n11124), .A2(n10265), .ZN(n10402) );
  NOR2_X1 U11516 ( .A1(n10201), .A2(n10344), .ZN(n11134) );
  OR2_X1 U11517 ( .A1(n10557), .A2(n10556), .ZN(n10373) );
  NAND2_X1 U11518 ( .A1(n10526), .A2(n12267), .ZN(n12385) );
  NAND2_X1 U11519 ( .A1(n12293), .A2(n12212), .ZN(n10653) );
  NAND2_X1 U11520 ( .A1(n10025), .A2(n12217), .ZN(n12218) );
  AND2_X1 U11521 ( .A1(n12237), .A2(n12235), .ZN(n12290) );
  XNOR2_X1 U11522 ( .A(n11121), .B(n14313), .ZN(n11122) );
  NOR4_X1 U11523 ( .A1(n17481), .A2(n17536), .A3(n17480), .A4(n17479), .ZN(
        n19802) );
  NAND3_X1 U11524 ( .A1(n9978), .A2(n10098), .A3(n10471), .ZN(n11113) );
  NAND3_X1 U11525 ( .A1(n10054), .A2(n11120), .A3(n11119), .ZN(n14313) );
  NOR2_X1 U11526 ( .A1(n14362), .A2(n14342), .ZN(n10753) );
  NAND2_X1 U11527 ( .A1(n11105), .A2(n11106), .ZN(n11128) );
  AND2_X1 U11528 ( .A1(n11092), .A2(n9973), .ZN(n10344) );
  NOR2_X4 U11529 ( .A1(n19326), .A2(n19812), .ZN(n19214) );
  NAND2_X1 U11530 ( .A1(n12207), .A2(n10519), .ZN(n12235) );
  INV_X1 U11531 ( .A(n14818), .ZN(n12609) );
  INV_X1 U11532 ( .A(n11118), .ZN(n9756) );
  INV_X1 U11533 ( .A(n14957), .ZN(n12578) );
  INV_X2 U11534 ( .A(n18567), .ZN(n9750) );
  AND2_X1 U11535 ( .A1(n12577), .A2(n12576), .ZN(n14957) );
  AND2_X1 U11536 ( .A1(n11385), .A2(n11384), .ZN(n17345) );
  AND2_X1 U11537 ( .A1(n10521), .A2(n10520), .ZN(n10519) );
  OR2_X1 U11538 ( .A1(n13053), .A2(n13052), .ZN(n13055) );
  CLKBUF_X1 U11539 ( .A(n11675), .Z(n17349) );
  OR2_X1 U11540 ( .A1(n13048), .A2(n15698), .ZN(n13053) );
  AND2_X1 U11541 ( .A1(n10155), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10555) );
  NAND2_X1 U11542 ( .A1(n12596), .A2(n21045), .ZN(n12553) );
  AND2_X2 U11543 ( .A1(n9783), .A2(n13864), .ZN(n12638) );
  NAND2_X1 U11544 ( .A1(n10514), .A2(n10512), .ZN(n17285) );
  AOI21_X1 U11545 ( .B1(n9840), .B2(n10044), .A(n20851), .ZN(n10043) );
  INV_X1 U11546 ( .A(n11108), .ZN(n11898) );
  AND2_X1 U11547 ( .A1(n11083), .A2(n11082), .ZN(n11676) );
  NOR2_X2 U11548 ( .A1(n20003), .A2(n14382), .ZN(n19812) );
  OR2_X1 U11549 ( .A1(n10398), .A2(n12202), .ZN(n10395) );
  AND3_X1 U11550 ( .A1(n12499), .A2(n12498), .A3(n12500), .ZN(n12505) );
  AND3_X1 U11551 ( .A1(n12126), .A2(n12125), .A3(n12198), .ZN(n12672) );
  INV_X1 U11552 ( .A(n15522), .ZN(n15538) );
  NAND2_X1 U11553 ( .A1(n12561), .A2(n12586), .ZN(n12562) );
  CLKBUF_X1 U11554 ( .A(n12664), .Z(n9784) );
  CLKBUF_X3 U11555 ( .A(n12664), .Z(n9783) );
  AOI21_X1 U11556 ( .B1(n10069), .B2(n10068), .A(n10071), .ZN(n10066) );
  AND3_X1 U11557 ( .A1(n10381), .A2(n12185), .A3(n12187), .ZN(n14487) );
  BUF_X1 U11558 ( .A(n12187), .Z(n15522) );
  INV_X4 U11559 ( .A(n12566), .ZN(n12561) );
  INV_X2 U11560 ( .A(n14391), .ZN(n13864) );
  AND2_X1 U11561 ( .A1(n12094), .A2(n21106), .ZN(n12202) );
  OR2_X1 U11562 ( .A1(n12518), .A2(n13785), .ZN(n12524) );
  AND2_X1 U11563 ( .A1(n13808), .A2(n10513), .ZN(n10512) );
  NAND2_X1 U11564 ( .A1(n12538), .A2(n12095), .ZN(n15582) );
  INV_X1 U11565 ( .A(n12893), .ZN(n18513) );
  AND2_X1 U11566 ( .A1(n14455), .A2(n14961), .ZN(n10381) );
  AND2_X1 U11567 ( .A1(n10748), .A2(n12178), .ZN(n12187) );
  AND2_X1 U11568 ( .A1(n11684), .A2(n11047), .ZN(n10513) );
  OAI21_X1 U11569 ( .B1(n10073), .B2(n10072), .A(n10074), .ZN(n10067) );
  NAND2_X1 U11570 ( .A1(n11358), .A2(n10832), .ZN(n13808) );
  NAND2_X1 U11571 ( .A1(n11077), .A2(n11074), .ZN(n10191) );
  INV_X1 U11573 ( .A(n11076), .ZN(n14194) );
  AND2_X1 U11574 ( .A1(n13031), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13038) );
  AND2_X1 U11575 ( .A1(n9749), .A2(n9748), .ZN(n10048) );
  OR2_X1 U11576 ( .A1(n12233), .A2(n21645), .ZN(n12305) );
  AND3_X2 U11577 ( .A1(n11336), .A2(n11335), .A3(n11334), .ZN(n11894) );
  NAND2_X1 U11578 ( .A1(n10026), .A2(n12186), .ZN(n10388) );
  NAND3_X4 U11579 ( .A1(n12152), .A2(n12151), .A3(n12150), .ZN(n9762) );
  INV_X1 U11580 ( .A(n11074), .ZN(n11024) );
  OR2_X1 U11581 ( .A1(n10941), .A2(n10940), .ZN(n14380) );
  NAND4_X2 U11582 ( .A1(n12068), .A2(n12067), .A3(n12066), .A4(n12065), .ZN(
        n12186) );
  NAND2_X1 U11583 ( .A1(n11025), .A2(n13989), .ZN(n11076) );
  CLKBUF_X1 U11584 ( .A(n10946), .Z(n18501) );
  NOR2_X2 U11585 ( .A1(n10930), .A2(n10929), .ZN(n19987) );
  OR2_X2 U11586 ( .A1(n12093), .A2(n12092), .ZN(n21106) );
  OR2_X1 U11587 ( .A1(n17872), .A2(n10561), .ZN(n18725) );
  NAND2_X2 U11588 ( .A1(n11023), .A2(n11022), .ZN(n20156) );
  AND4_X1 U11589 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12138) );
  AND4_X1 U11590 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(
        n12080) );
  AND4_X1 U11591 ( .A1(n12164), .A2(n12163), .A3(n12162), .A4(n12161), .ZN(
        n12174) );
  NAND2_X1 U11592 ( .A1(n9794), .A2(n9857), .ZN(n10198) );
  NAND2_X1 U11593 ( .A1(n10220), .A2(n10219), .ZN(n11798) );
  NAND2_X2 U11594 ( .A1(n10673), .A2(n10671), .ZN(n20181) );
  AND4_X1 U11595 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(
        n12066) );
  AND3_X1 U11596 ( .A1(n12064), .A2(n12063), .A3(n12062), .ZN(n12065) );
  NOR2_X1 U11597 ( .A1(n9997), .A2(n9995), .ZN(n9994) );
  AND4_X1 U11598 ( .A1(n12056), .A2(n12055), .A3(n12054), .A4(n12053), .ZN(
        n12067) );
  AND4_X1 U11599 ( .A1(n12168), .A2(n12167), .A3(n12166), .A4(n12165), .ZN(
        n12173) );
  NAND2_X1 U11600 ( .A1(n10791), .A2(n10790), .ZN(n10789) );
  NAND2_X1 U11601 ( .A1(n10672), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10671) );
  NAND2_X1 U11602 ( .A1(n10788), .A2(n10787), .ZN(n10786) );
  INV_X1 U11603 ( .A(n11200), .ZN(n16228) );
  INV_X1 U11604 ( .A(U214), .ZN(n17688) );
  AND2_X1 U11605 ( .A1(n11003), .A2(n11004), .ZN(n10787) );
  AND3_X1 U11606 ( .A1(n11006), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11005), .ZN(n10788) );
  AND3_X1 U11607 ( .A1(n11010), .A2(n11015), .A3(n11007), .ZN(n10790) );
  AND2_X1 U11608 ( .A1(n11009), .A2(n11008), .ZN(n10791) );
  AND3_X1 U11609 ( .A1(n10216), .A2(n10217), .A3(n10215), .ZN(n10214) );
  AND3_X1 U11610 ( .A1(n10223), .A2(n10222), .A3(n11015), .ZN(n10221) );
  INV_X4 U11612 ( .A(n9747), .ZN(n18333) );
  INV_X4 U11613 ( .A(n18239), .ZN(n18341) );
  BUF_X2 U11614 ( .A(n12816), .Z(n18314) );
  CLKBUF_X3 U11615 ( .A(n13322), .Z(n13525) );
  BUF_X2 U11616 ( .A(n12816), .Z(n18344) );
  CLKBUF_X3 U11617 ( .A(n12817), .Z(n18320) );
  NAND2_X2 U11618 ( .A1(n20862), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20778) );
  NAND2_X2 U11619 ( .A1(n16378), .A2(n11015), .ZN(n11252) );
  NAND2_X1 U11620 ( .A1(n10422), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17484) );
  INV_X1 U11621 ( .A(n13687), .ZN(n9751) );
  NOR2_X1 U11622 ( .A1(n10866), .A2(n10865), .ZN(n12807) );
  INV_X1 U11623 ( .A(n16356), .ZN(n9752) );
  INV_X2 U11624 ( .A(n12097), .ZN(n9753) );
  INV_X1 U11625 ( .A(n13711), .ZN(n9754) );
  AND2_X2 U11626 ( .A1(n10405), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12036) );
  NAND2_X1 U11627 ( .A1(n19961), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10866) );
  OR2_X1 U11628 ( .A1(n10859), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10868) );
  NOR3_X2 U11629 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18054) );
  INV_X2 U11630 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12471) );
  INV_X2 U11631 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19953) );
  INV_X1 U11632 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18088) );
  INV_X1 U11633 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17498) );
  INV_X1 U11634 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10405) );
  AND2_X2 U11635 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11171) );
  OR2_X1 U11636 ( .A1(n17136), .A2(n17234), .ZN(n10057) );
  OAI21_X1 U11637 ( .B1(n10060), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n9806), .ZN(n17136) );
  NAND4_X2 U11638 ( .A1(n10378), .A2(n12184), .A3(n12183), .A4(n9905), .ZN(
        n12543) );
  NAND2_X1 U11639 ( .A1(n19987), .A2(n12934), .ZN(n19013) );
  NAND2_X1 U11640 ( .A1(n12934), .A2(n18596), .ZN(n19012) );
  INV_X2 U11641 ( .A(n9734), .ZN(n9755) );
  NAND4_X1 U11642 ( .A1(n10214), .A2(n10999), .A3(n10998), .A4(n10218), .ZN(
        n10219) );
  AND2_X4 U11643 ( .A1(n12471), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12031) );
  INV_X1 U11644 ( .A(n9756), .ZN(n9757) );
  NAND2_X1 U11645 ( .A1(n11115), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10098) );
  INV_X2 U11646 ( .A(n13989), .ZN(n11073) );
  NOR2_X2 U11647 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18000), .ZN(n17986) );
  INV_X1 U11648 ( .A(n16352), .ZN(n16267) );
  NAND3_X4 U11649 ( .A1(n21769), .A2(n17335), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16356) );
  AOI211_X1 U11650 ( .C1(n16967), .C2(n17221), .A(n16966), .B(n16965), .ZN(
        n16968) );
  NAND2_X1 U11651 ( .A1(n16865), .A2(n11339), .ZN(n10109) );
  INV_X1 U11652 ( .A(n11200), .ZN(n9764) );
  OAI211_X1 U11653 ( .C1(n9913), .C2(n16422), .A(n10248), .B(n10247), .ZN(
        n16413) );
  NAND2_X2 U11654 ( .A1(n13493), .A2(n10170), .ZN(n14604) );
  NAND2_X1 U11655 ( .A1(n10639), .A2(n11290), .ZN(n11262) );
  NOR2_X2 U11656 ( .A1(n11151), .A2(n11150), .ZN(n11160) );
  OAI22_X2 U11657 ( .A1(n20451), .A2(n16064), .B1(n20227), .B2(n11149), .ZN(
        n11150) );
  NOR2_X4 U11658 ( .A1(n14284), .A2(n14451), .ZN(n14450) );
  NAND4_X2 U11659 ( .A1(n11161), .A2(n11160), .A3(n11159), .A4(n11162), .ZN(
        n11212) );
  INV_X4 U11660 ( .A(n20965), .ZN(n20952) );
  INV_X4 U11661 ( .A(n16356), .ZN(n16244) );
  INV_X4 U11662 ( .A(n11429), .ZN(n11078) );
  NAND2_X4 U11663 ( .A1(n12031), .A2(n15521), .ZN(n13231) );
  NOR2_X2 U11664 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17832), .ZN(n17820) );
  AND2_X1 U11665 ( .A1(n11171), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9765) );
  INV_X1 U11666 ( .A(n16378), .ZN(n9766) );
  INV_X4 U11667 ( .A(n16289), .ZN(n9767) );
  INV_X2 U11668 ( .A(n16289), .ZN(n9768) );
  NOR2_X2 U11670 ( .A1(n12149), .A2(n12148), .ZN(n12150) );
  NOR2_X2 U11671 ( .A1(n14956), .A2(n10595), .ZN(n14879) );
  NAND2_X2 U11672 ( .A1(n14450), .A2(n20935), .ZN(n14956) );
  NOR2_X2 U11673 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17814), .ZN(n17800) );
  INV_X1 U11674 ( .A(n16356), .ZN(n11172) );
  NOR2_X2 U11675 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17791), .ZN(n17781) );
  INV_X1 U11676 ( .A(n13723), .ZN(n9772) );
  AOI21_X1 U11677 ( .B1(n10242), .B2(n9813), .A(n16365), .ZN(n10451) );
  OR2_X2 U11678 ( .A1(n16401), .A2(n10242), .ZN(n10453) );
  AND2_X1 U11679 ( .A1(n12036), .A2(n15521), .ZN(n13322) );
  NOR2_X2 U11680 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18022), .ZN(n18006) );
  NAND2_X1 U11681 ( .A1(n12553), .A2(n12552), .ZN(n12557) );
  INV_X1 U11682 ( .A(n13636), .ZN(n9774) );
  NAND2_X1 U11683 ( .A1(n12031), .A2(n12042), .ZN(n13636) );
  INV_X1 U11684 ( .A(n12097), .ZN(n9778) );
  INV_X4 U11686 ( .A(n12097), .ZN(n13725) );
  NOR2_X4 U11687 ( .A1(n15823), .A2(n16465), .ZN(n15798) );
  NOR2_X1 U11688 ( .A1(n12566), .A2(n12556), .ZN(n12560) );
  AND2_X1 U11689 ( .A1(n12233), .A2(n12184), .ZN(n10392) );
  OR2_X1 U11690 ( .A1(n12184), .A2(n21645), .ZN(n12304) );
  AOI22_X1 U11691 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19824), .B1(
        n10959), .B2(n10623), .ZN(n10961) );
  NOR2_X1 U11692 ( .A1(n10959), .A2(n10623), .ZN(n10962) );
  NAND2_X1 U11693 ( .A1(n10142), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10141) );
  NAND2_X1 U11694 ( .A1(n9788), .A2(n15191), .ZN(n10524) );
  AND2_X1 U11695 ( .A1(n10384), .A2(n12403), .ZN(n10382) );
  NAND2_X1 U11696 ( .A1(n12491), .A2(n12233), .ZN(n12518) );
  NAND2_X1 U11697 ( .A1(n10237), .A2(n10238), .ZN(n10236) );
  NAND3_X1 U11698 ( .A1(n16894), .A2(n11988), .A3(n10551), .ZN(n10148) );
  INV_X1 U11699 ( .A(n10322), .ZN(n10305) );
  NOR2_X1 U11700 ( .A1(n16649), .A2(n16685), .ZN(n11880) );
  NAND2_X1 U11701 ( .A1(n9793), .A2(n16868), .ZN(n9987) );
  AND4_X1 U11702 ( .A1(n11333), .A2(n11332), .A3(n11331), .A4(n11330), .ZN(
        n11334) );
  AND2_X1 U11703 ( .A1(n11073), .A2(n11798), .ZN(n10075) );
  NOR2_X1 U11704 ( .A1(n12834), .A2(n18513), .ZN(n10134) );
  NOR2_X1 U11705 ( .A1(n19366), .A2(n12854), .ZN(n12884) );
  NAND2_X1 U11706 ( .A1(n12185), .A2(n12184), .ZN(n10398) );
  NAND2_X1 U11707 ( .A1(n15367), .A2(n9866), .ZN(n15353) );
  OR2_X1 U11708 ( .A1(n11802), .A2(n17103), .ZN(n11995) );
  NAND2_X1 U11709 ( .A1(n10311), .A2(n11994), .ZN(n10310) );
  INV_X1 U11710 ( .A(n11993), .ZN(n10311) );
  INV_X1 U11711 ( .A(n10351), .ZN(n10350) );
  AOI21_X1 U11712 ( .B1(n10349), .B2(n10351), .A(n10348), .ZN(n10347) );
  INV_X1 U11713 ( .A(n16794), .ZN(n10348) );
  NOR2_X1 U11714 ( .A1(n20161), .A2(n11058), .ZN(n10068) );
  AND2_X1 U11715 ( .A1(n9749), .A2(n20156), .ZN(n10071) );
  INV_X1 U11716 ( .A(n10191), .ZN(n10069) );
  NAND2_X1 U11717 ( .A1(n10075), .A2(n9748), .ZN(n10072) );
  NAND2_X1 U11718 ( .A1(n20156), .A2(n20851), .ZN(n10074) );
  NAND2_X1 U11719 ( .A1(n20851), .A2(n9749), .ZN(n10073) );
  NAND2_X1 U11720 ( .A1(n10070), .A2(n20156), .ZN(n10065) );
  INV_X1 U11721 ( .A(n11075), .ZN(n10070) );
  NAND2_X1 U11722 ( .A1(n10480), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10420) );
  NAND2_X1 U11723 ( .A1(n12540), .A2(n15582), .ZN(n12205) );
  OR2_X1 U11724 ( .A1(n12286), .A2(n12285), .ZN(n12380) );
  NAND2_X1 U11725 ( .A1(n10388), .A2(n12177), .ZN(n12198) );
  INV_X1 U11726 ( .A(n11243), .ZN(n11454) );
  AND2_X2 U11727 ( .A1(n10979), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11170) );
  INV_X1 U11728 ( .A(n11203), .ZN(n10647) );
  INV_X1 U11729 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16110) );
  NAND2_X1 U11730 ( .A1(n20161), .A2(n20181), .ZN(n11060) );
  NAND2_X1 U11731 ( .A1(n11154), .A2(n11155), .ZN(n11214) );
  NAND2_X1 U11732 ( .A1(n21647), .A2(n21880), .ZN(n14398) );
  NAND2_X1 U11733 ( .A1(n10742), .A2(n9823), .ZN(n10741) );
  NAND2_X1 U11734 ( .A1(n15114), .A2(n10742), .ZN(n10391) );
  AND2_X1 U11735 ( .A1(n12450), .A2(n17539), .ZN(n12451) );
  INV_X1 U11736 ( .A(n17577), .ZN(n10598) );
  OR2_X1 U11737 ( .A1(n12265), .A2(n12264), .ZN(n12386) );
  OR2_X1 U11738 ( .A1(n12195), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12196) );
  NAND2_X1 U11739 ( .A1(n10021), .A2(n9874), .ZN(n10020) );
  NAND2_X1 U11740 ( .A1(n12213), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10025) );
  NAND2_X1 U11741 ( .A1(n12725), .A2(n11871), .ZN(n11873) );
  INV_X1 U11742 ( .A(n11759), .ZN(n10182) );
  INV_X1 U11743 ( .A(n16435), .ZN(n10707) );
  NOR2_X1 U11744 ( .A1(n14300), .A2(n10720), .ZN(n15785) );
  NAND2_X1 U11745 ( .A1(n10722), .A2(n10721), .ZN(n10720) );
  INV_X1 U11746 ( .A(n15810), .ZN(n10721) );
  NAND2_X1 U11747 ( .A1(n14007), .A2(n13989), .ZN(n14349) );
  NOR2_X1 U11748 ( .A1(n20854), .A2(n10286), .ZN(n14007) );
  AND2_X1 U11749 ( .A1(n11058), .A2(n11078), .ZN(n11684) );
  INV_X1 U11750 ( .A(n13014), .ZN(n12016) );
  NAND2_X1 U11751 ( .A1(n10763), .A2(n13000), .ZN(n10762) );
  INV_X1 U11752 ( .A(n15638), .ZN(n10763) );
  NOR2_X1 U11753 ( .A1(n15654), .A2(n15655), .ZN(n15639) );
  NAND2_X1 U11754 ( .A1(n10460), .A2(n10458), .ZN(n16695) );
  NAND2_X1 U11755 ( .A1(n10459), .A2(n9846), .ZN(n10458) );
  OR2_X1 U11756 ( .A1(n9789), .A2(n10229), .ZN(n10224) );
  NAND2_X1 U11757 ( .A1(n10694), .A2(n10226), .ZN(n10225) );
  INV_X1 U11758 ( .A(n10310), .ZN(n10229) );
  NAND2_X1 U11759 ( .A1(n10122), .A2(n11316), .ZN(n16865) );
  NAND2_X1 U11760 ( .A1(n10635), .A2(n11987), .ZN(n10315) );
  INV_X1 U11761 ( .A(n10713), .ZN(n10712) );
  OAI21_X1 U11762 ( .B1(n10715), .B2(n9829), .A(n14263), .ZN(n10713) );
  AND2_X1 U11763 ( .A1(n10193), .A2(n10192), .ZN(n11296) );
  AND2_X1 U11764 ( .A1(n11468), .A2(n11462), .ZN(n10726) );
  NAND2_X1 U11765 ( .A1(n11261), .A2(n10794), .ZN(n10639) );
  AOI21_X1 U11766 ( .B1(n11981), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11097), 
        .ZN(n11098) );
  OR2_X1 U11767 ( .A1(n14349), .A2(n16110), .ZN(n14173) );
  AND2_X1 U11768 ( .A1(n10546), .A2(n19816), .ZN(n17481) );
  INV_X1 U11769 ( .A(n14382), .ZN(n10546) );
  NOR2_X1 U11770 ( .A1(n18938), .A2(n12836), .ZN(n12838) );
  NAND2_X1 U11771 ( .A1(n10531), .A2(n10965), .ZN(n12874) );
  OR2_X1 U11772 ( .A1(n12873), .A2(n10963), .ZN(n10531) );
  INV_X1 U11773 ( .A(n10944), .ZN(n10426) );
  NOR2_X1 U11774 ( .A1(n10948), .A2(n9963), .ZN(n10423) );
  OR2_X1 U11775 ( .A1(n14380), .A2(n10953), .ZN(n9963) );
  NOR2_X1 U11776 ( .A1(n10329), .A2(n12865), .ZN(n12882) );
  NAND2_X1 U11777 ( .A1(n19349), .A2(n10946), .ZN(n10944) );
  NAND2_X1 U11778 ( .A1(n14500), .A2(n14513), .ZN(n14502) );
  INV_X1 U11779 ( .A(n14502), .ZN(n10255) );
  OAI21_X1 U11780 ( .B1(n12534), .B2(n10013), .A(n10486), .ZN(n10485) );
  AOI21_X1 U11781 ( .B1(n10490), .B2(n10489), .A(n10487), .ZN(n10486) );
  INV_X1 U11782 ( .A(n20866), .ZN(n14486) );
  NAND2_X1 U11783 ( .A1(n9890), .A2(n11080), .ZN(n11087) );
  AOI21_X1 U11784 ( .B1(n10292), .B2(n10291), .A(n10290), .ZN(n10289) );
  INV_X1 U11785 ( .A(n16643), .ZN(n10290) );
  INV_X1 U11786 ( .A(n10295), .ZN(n10291) );
  OR2_X1 U11787 ( .A1(n13063), .A2(n10293), .ZN(n10288) );
  NOR2_X1 U11788 ( .A1(n10242), .A2(n16402), .ZN(n10241) );
  NOR2_X1 U11789 ( .A1(n11064), .A2(n20851), .ZN(n10094) );
  NAND2_X1 U11790 ( .A1(n10147), .A2(n9865), .ZN(n16778) );
  NAND2_X1 U11791 ( .A1(n10189), .A2(n9873), .ZN(n10188) );
  AND2_X1 U11792 ( .A1(n15624), .A2(n10734), .ZN(n14431) );
  AND2_X1 U11793 ( .A1(n10736), .A2(n10735), .ZN(n10734) );
  INV_X1 U11794 ( .A(n14429), .ZN(n10735) );
  INV_X1 U11795 ( .A(n10120), .ZN(n16744) );
  NAND2_X1 U11796 ( .A1(n15821), .A2(n11838), .ZN(n16794) );
  NAND2_X1 U11797 ( .A1(n10695), .A2(n10153), .ZN(n16825) );
  NAND2_X1 U11798 ( .A1(n10079), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10078) );
  AOI21_X1 U11799 ( .B1(n15933), .B2(n10717), .A(n9938), .ZN(n10715) );
  NAND2_X1 U11800 ( .A1(n10081), .A2(n11262), .ZN(n11264) );
  INV_X1 U11801 ( .A(n11263), .ZN(n10081) );
  NAND2_X1 U11802 ( .A1(n10080), .A2(n17229), .ZN(n10781) );
  AND2_X2 U11803 ( .A1(n10075), .A2(n10048), .ZN(n11695) );
  OAI21_X1 U11804 ( .B1(n15994), .B2(n14206), .A(n14006), .ZN(n14009) );
  NAND2_X1 U11805 ( .A1(n9840), .A2(n10093), .ZN(n11079) );
  INV_X1 U11806 ( .A(n11064), .ZN(n10093) );
  INV_X1 U11807 ( .A(n10832), .ZN(n13974) );
  AND2_X1 U11808 ( .A1(n20199), .A2(n20133), .ZN(n20357) );
  NOR2_X1 U11809 ( .A1(n12933), .A2(n19006), .ZN(n10850) );
  OR2_X1 U11810 ( .A1(n10564), .A2(n18759), .ZN(n10563) );
  NOR2_X1 U11811 ( .A1(n17935), .A2(n18811), .ZN(n18808) );
  CLKBUF_X1 U11812 ( .A(n12880), .Z(n19177) );
  OR2_X1 U11813 ( .A1(n18938), .A2(n10444), .ZN(n10210) );
  NAND2_X1 U11814 ( .A1(n12837), .A2(n10445), .ZN(n10444) );
  NAND2_X1 U11815 ( .A1(n18938), .A2(n10442), .ZN(n10441) );
  INV_X1 U11816 ( .A(n12837), .ZN(n10442) );
  NOR2_X1 U11817 ( .A1(n17636), .A2(n12932), .ZN(n13089) );
  NAND2_X1 U11818 ( .A1(n17633), .A2(n18920), .ZN(n17636) );
  NOR2_X1 U11819 ( .A1(n19149), .A2(n19024), .ZN(n18656) );
  NAND2_X1 U11820 ( .A1(n18910), .A2(n12917), .ZN(n18877) );
  INV_X1 U11821 ( .A(n12915), .ZN(n12913) );
  NOR2_X1 U11822 ( .A1(n12840), .A2(n19233), .ZN(n12880) );
  INV_X1 U11823 ( .A(n18510), .ZN(n17635) );
  NAND2_X1 U11824 ( .A1(n18911), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18910) );
  OR3_X1 U11825 ( .A1(n11087), .A2(n17348), .A3(n17617), .ZN(n13803) );
  AND2_X1 U11826 ( .A1(n16010), .A2(n13803), .ZN(n20847) );
  NAND2_X1 U11827 ( .A1(n12004), .A2(n12003), .ZN(n13811) );
  NOR2_X1 U11828 ( .A1(n12724), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12726) );
  NAND2_X1 U11829 ( .A1(n9986), .A2(n9984), .ZN(n10269) );
  NAND2_X1 U11830 ( .A1(n9985), .A2(n10270), .ZN(n9984) );
  NAND2_X1 U11831 ( .A1(n16921), .A2(n13884), .ZN(n16933) );
  INV_X1 U11832 ( .A(n10167), .ZN(n10166) );
  OAI21_X1 U11833 ( .B1(n17101), .B2(n17241), .A(n17100), .ZN(n10167) );
  INV_X1 U11834 ( .A(n17241), .ZN(n17260) );
  OAI21_X1 U11835 ( .B1(n18909), .B2(n19190), .A(n9958), .ZN(n9957) );
  NAND2_X1 U11836 ( .A1(n19317), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U11837 ( .A1(n10064), .A2(n10063), .ZN(n10041) );
  INV_X1 U11838 ( .A(n11683), .ZN(n10063) );
  AOI22_X1 U11839 ( .A1(n12510), .A2(n12514), .B1(n12518), .B2(n12516), .ZN(
        n10499) );
  AND2_X1 U11840 ( .A1(n11200), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10178) );
  NOR2_X1 U11841 ( .A1(n11068), .A2(n11067), .ZN(n11069) );
  INV_X1 U11842 ( .A(n10537), .ZN(n10959) );
  OAI21_X1 U11843 ( .B1(n10958), .B2(n10957), .A(n10538), .ZN(n10537) );
  NAND2_X1 U11844 ( .A1(n19803), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10538) );
  AND2_X1 U11845 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10336) );
  AOI21_X1 U11846 ( .B1(n12486), .B2(n12485), .A(n12472), .ZN(n12478) );
  AND2_X1 U11848 ( .A1(n12184), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12491) );
  NAND2_X1 U11849 ( .A1(n10261), .A2(n12204), .ZN(n10520) );
  INV_X1 U11850 ( .A(n12672), .ZN(n10261) );
  OR2_X1 U11851 ( .A1(n12251), .A2(n12250), .ZN(n12437) );
  INV_X1 U11852 ( .A(n13148), .ZN(n10014) );
  INV_X1 U11853 ( .A(n13147), .ZN(n10015) );
  INV_X1 U11854 ( .A(n10558), .ZN(n10023) );
  NOR2_X1 U11855 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21057), .ZN(
        n12477) );
  INV_X1 U11856 ( .A(n10499), .ZN(n10498) );
  OAI21_X1 U11857 ( .B1(n10497), .B2(n9830), .A(n10501), .ZN(n10492) );
  INV_X1 U11858 ( .A(n12525), .ZN(n10501) );
  AOI21_X1 U11859 ( .B1(n10499), .B2(n10500), .A(n9876), .ZN(n10497) );
  OAI21_X1 U11860 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n17596), .A(n12523), 
        .ZN(n12525) );
  AND2_X1 U11861 ( .A1(n16377), .A2(n11015), .ZN(n11200) );
  NAND2_X1 U11862 ( .A1(n10103), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10635) );
  INV_X1 U11863 ( .A(n11315), .ZN(n10103) );
  AND2_X1 U11864 ( .A1(n9927), .A2(n11237), .ZN(n10548) );
  NAND2_X1 U11865 ( .A1(n9980), .A2(n9979), .ZN(n10472) );
  INV_X1 U11866 ( .A(n11111), .ZN(n9980) );
  NAND2_X1 U11867 ( .A1(n11118), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n9979) );
  OAI211_X1 U11868 ( .C1(n11968), .C2(n20734), .A(n11110), .B(n11109), .ZN(
        n11111) );
  INV_X1 U11869 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U11870 ( .A1(n10515), .A2(n11026), .ZN(n10514) );
  NAND2_X1 U11871 ( .A1(n10136), .A2(n10135), .ZN(n12834) );
  INV_X1 U11872 ( .A(n18516), .ZN(n10135) );
  INV_X1 U11873 ( .A(n12833), .ZN(n10136) );
  AND2_X1 U11874 ( .A1(n12478), .A2(n12477), .ZN(n12520) );
  NAND2_X1 U11875 ( .A1(n10030), .A2(n9763), .ZN(n10029) );
  AND2_X1 U11876 ( .A1(n14582), .A2(n10771), .ZN(n10770) );
  INV_X1 U11877 ( .A(n10772), .ZN(n10771) );
  AND2_X1 U11878 ( .A1(n9817), .A2(n14733), .ZN(n10767) );
  OR2_X1 U11879 ( .A1(n15582), .A2(n21645), .ZN(n13737) );
  INV_X1 U11880 ( .A(n13149), .ZN(n13627) );
  INV_X1 U11881 ( .A(n14398), .ZN(n13740) );
  NAND2_X1 U11882 ( .A1(n9841), .A2(n10475), .ZN(n10474) );
  NAND2_X1 U11883 ( .A1(n9841), .A2(n21645), .ZN(n10476) );
  NAND2_X1 U11884 ( .A1(n12295), .A2(n9762), .ZN(n10475) );
  AND3_X1 U11885 ( .A1(n12663), .A2(n12183), .A3(n12536), .ZN(n12542) );
  INV_X1 U11886 ( .A(n14661), .ZN(n10608) );
  INV_X1 U11887 ( .A(n10416), .ZN(n10379) );
  AND2_X1 U11888 ( .A1(n14693), .A2(n10610), .ZN(n10609) );
  INV_X1 U11889 ( .A(n14677), .ZN(n10610) );
  NOR2_X1 U11890 ( .A1(n14794), .A2(n10606), .ZN(n10605) );
  INV_X1 U11891 ( .A(n14785), .ZN(n10606) );
  AND2_X1 U11892 ( .A1(n12593), .A2(n10601), .ZN(n10600) );
  INV_X1 U11893 ( .A(n14870), .ZN(n10601) );
  INV_X1 U11894 ( .A(n12638), .ZN(n12656) );
  OAI211_X1 U11895 ( .C1(n12419), .C2(n10368), .A(n10367), .B(n10366), .ZN(
        n10365) );
  NAND2_X1 U11896 ( .A1(n12420), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10367) );
  NAND2_X1 U11897 ( .A1(n20994), .A2(n12421), .ZN(n10366) );
  INV_X1 U11898 ( .A(n12267), .ZN(n10529) );
  AND2_X1 U11899 ( .A1(n13154), .A2(n10528), .ZN(n10527) );
  NAND2_X1 U11900 ( .A1(n12267), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10528) );
  NOR2_X1 U11901 ( .A1(n15582), .A2(n12185), .ZN(n10489) );
  OAI21_X1 U11902 ( .B1(n12208), .B2(n10036), .A(n10035), .ZN(n10034) );
  NAND2_X1 U11903 ( .A1(n10039), .A2(n12191), .ZN(n10038) );
  NAND2_X1 U11904 ( .A1(n12213), .A2(n9859), .ZN(n10037) );
  NAND2_X1 U11905 ( .A1(n21106), .A2(n12233), .ZN(n12096) );
  INV_X1 U11906 ( .A(n10388), .ZN(n12538) );
  AND3_X2 U11907 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10560) );
  INV_X1 U11908 ( .A(n10027), .ZN(n21510) );
  NAND2_X1 U11909 ( .A1(n10022), .A2(n12319), .ZN(n21229) );
  OAI211_X1 U11910 ( .C1(n10617), .C2(n10653), .A(n21645), .B(n10615), .ZN(
        n10022) );
  INV_X1 U11911 ( .A(n21508), .ZN(n21578) );
  NAND2_X1 U11912 ( .A1(n10299), .A2(n10298), .ZN(n11729) );
  NAND2_X1 U11913 ( .A1(n11358), .A2(n11400), .ZN(n10298) );
  NAND2_X1 U11914 ( .A1(n11387), .A2(n11469), .ZN(n10299) );
  NAND2_X1 U11915 ( .A1(n11877), .A2(n11879), .ZN(n11874) );
  NOR2_X1 U11916 ( .A1(n11859), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10652) );
  NAND2_X1 U11917 ( .A1(n15699), .A2(n10275), .ZN(n10278) );
  OR2_X1 U11918 ( .A1(n11812), .A2(n10642), .ZN(n11830) );
  NAND2_X1 U11919 ( .A1(n10643), .A2(n10803), .ZN(n10642) );
  INV_X1 U11920 ( .A(n10644), .ZN(n10643) );
  INV_X1 U11921 ( .A(n11796), .ZN(n10641) );
  NOR2_X1 U11922 ( .A1(n9785), .A2(n9888), .ZN(n10308) );
  INV_X1 U11923 ( .A(n10308), .ZN(n10306) );
  OAI21_X1 U11924 ( .B1(n11722), .B2(n11889), .A(n11721), .ZN(n11741) );
  NAND2_X1 U11925 ( .A1(n16279), .A2(n10702), .ZN(n10701) );
  NAND2_X1 U11926 ( .A1(n16429), .A2(n10820), .ZN(n16237) );
  AND2_X1 U11927 ( .A1(n13808), .A2(n20850), .ZN(n13962) );
  NAND2_X1 U11928 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10660) );
  NOR2_X1 U11929 ( .A1(n16887), .A2(n10665), .ZN(n10664) );
  NAND2_X1 U11930 ( .A1(n10320), .A2(n10473), .ZN(n10322) );
  AND2_X1 U11931 ( .A1(n9856), .A2(n11886), .ZN(n10473) );
  NAND2_X1 U11932 ( .A1(n16695), .A2(n11868), .ZN(n10323) );
  NAND2_X1 U11933 ( .A1(n10759), .A2(n11950), .ZN(n10758) );
  INV_X1 U11934 ( .A(n15727), .ZN(n10759) );
  NAND2_X1 U11935 ( .A1(n10146), .A2(n10190), .ZN(n9972) );
  AND2_X1 U11936 ( .A1(n9897), .A2(n20054), .ZN(n10190) );
  AND2_X1 U11937 ( .A1(n10097), .A2(n11989), .ZN(n10461) );
  INV_X1 U11938 ( .A(n12013), .ZN(n11950) );
  INV_X1 U11939 ( .A(n9945), .ZN(n9990) );
  NAND2_X1 U11940 ( .A1(n11794), .A2(n11864), .ZN(n11848) );
  INV_X1 U11941 ( .A(n15764), .ZN(n11794) );
  AND2_X1 U11942 ( .A1(n15799), .A2(n11941), .ZN(n10750) );
  INV_X1 U11943 ( .A(n15784), .ZN(n11941) );
  NAND2_X1 U11944 ( .A1(n10725), .A2(n14368), .ZN(n10724) );
  INV_X1 U11945 ( .A(n14358), .ZN(n10725) );
  AND2_X1 U11946 ( .A1(n11929), .A2(n15843), .ZN(n10760) );
  NAND2_X1 U11947 ( .A1(n10728), .A2(n14278), .ZN(n10727) );
  INV_X1 U11948 ( .A(n10729), .ZN(n10728) );
  NAND2_X1 U11949 ( .A1(n10731), .A2(n10730), .ZN(n10729) );
  INV_X1 U11950 ( .A(n14257), .ZN(n10730) );
  INV_X1 U11951 ( .A(n14271), .ZN(n10731) );
  OR2_X1 U11952 ( .A1(n16894), .A2(n10694), .ZN(n10154) );
  NAND2_X1 U11953 ( .A1(n16894), .A2(n11988), .ZN(n10695) );
  AND3_X1 U11954 ( .A1(n11312), .A2(n11311), .A3(n11310), .ZN(n11762) );
  NAND2_X1 U11955 ( .A1(n20054), .A2(n10114), .ZN(n10113) );
  NAND2_X1 U11956 ( .A1(n11864), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10114) );
  INV_X1 U11957 ( .A(n10163), .ZN(n10203) );
  INV_X1 U11958 ( .A(n11264), .ZN(n10778) );
  INV_X1 U11959 ( .A(n14315), .ZN(n10754) );
  INV_X1 U11960 ( .A(n11755), .ZN(n10682) );
  NOR2_X1 U11961 ( .A1(n11202), .A2(n10649), .ZN(n10648) );
  NAND2_X1 U11962 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10646) );
  INV_X1 U11963 ( .A(n14173), .ZN(n14174) );
  AND2_X1 U11964 ( .A1(n20416), .A2(n20253), .ZN(n20296) );
  AND2_X1 U11965 ( .A1(n17281), .A2(n11136), .ZN(n11147) );
  AND3_X1 U11966 ( .A1(n13967), .A2(n14189), .A3(n13994), .ZN(n17336) );
  NOR2_X1 U11967 ( .A1(n10865), .A2(n18072), .ZN(n12809) );
  NOR2_X1 U11968 ( .A1(n10866), .A2(n10868), .ZN(n12731) );
  INV_X1 U11969 ( .A(n12836), .ZN(n10445) );
  OAI21_X1 U11970 ( .B1(n10134), .B2(n17635), .A(n9755), .ZN(n12837) );
  NAND2_X1 U11971 ( .A1(n10209), .A2(n9755), .ZN(n13088) );
  AND2_X1 U11972 ( .A1(n18718), .A2(n10633), .ZN(n18700) );
  AND2_X1 U11973 ( .A1(n18919), .A2(n9795), .ZN(n12848) );
  OAI21_X1 U11974 ( .B1(n18927), .B2(n18926), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12915) );
  NAND2_X1 U11975 ( .A1(n19284), .A2(n12905), .ZN(n12906) );
  AND2_X1 U11976 ( .A1(n9733), .A2(n9969), .ZN(n12900) );
  NOR2_X1 U11977 ( .A1(n19370), .A2(n18399), .ZN(n12856) );
  NAND2_X1 U11978 ( .A1(n18545), .A2(n17477), .ZN(n10956) );
  NAND2_X1 U11979 ( .A1(n12889), .A2(n19779), .ZN(n10439) );
  NOR2_X1 U11980 ( .A1(n10428), .A2(n19987), .ZN(n10427) );
  INV_X1 U11981 ( .A(n17477), .ZN(n10428) );
  NOR2_X1 U11982 ( .A1(n10334), .A2(n10333), .ZN(n10332) );
  OR3_X1 U11983 ( .A1(n21735), .A2(n14400), .A3(n14399), .ZN(n20904) );
  NOR2_X1 U11984 ( .A1(n10173), .A2(n10172), .ZN(n10170) );
  OR2_X1 U11985 ( .A1(n14086), .A2(n14085), .ZN(n14397) );
  NAND2_X1 U11986 ( .A1(n13427), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13453) );
  INV_X1 U11987 ( .A(n14952), .ZN(n10169) );
  NAND2_X1 U11988 ( .A1(n10008), .A2(n12379), .ZN(n14333) );
  NAND2_X1 U11989 ( .A1(n12374), .A2(n9799), .ZN(n10008) );
  NOR2_X1 U11990 ( .A1(n13143), .A2(n10823), .ZN(n13144) );
  AND2_X2 U11991 ( .A1(n9762), .A2(n12177), .ZN(n12566) );
  NAND2_X1 U11992 ( .A1(n10554), .A2(n10389), .ZN(n14500) );
  AND2_X1 U11993 ( .A1(n10391), .A2(n10390), .ZN(n10389) );
  NOR2_X1 U11994 ( .A1(n10739), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10390) );
  NAND2_X1 U11995 ( .A1(n15097), .A2(n9918), .ZN(n14501) );
  NAND2_X1 U11996 ( .A1(n10002), .A2(n15305), .ZN(n10006) );
  NAND2_X1 U11997 ( .A1(n9878), .A2(n10654), .ZN(n10005) );
  NAND2_X1 U11998 ( .A1(n10001), .A2(n10000), .ZN(n10003) );
  AOI21_X1 U11999 ( .B1(n15096), .B2(n15105), .A(n9807), .ZN(n10000) );
  NAND2_X1 U12000 ( .A1(n10554), .A2(n15105), .ZN(n15097) );
  NAND2_X1 U12001 ( .A1(n10007), .A2(n10161), .ZN(n15142) );
  INV_X1 U12002 ( .A(n10162), .ZN(n10161) );
  INV_X1 U12003 ( .A(n12460), .ZN(n10418) );
  INV_X1 U12004 ( .A(n15504), .ZN(n10507) );
  NAND2_X1 U12005 ( .A1(n15394), .A2(n12697), .ZN(n10506) );
  NAND2_X1 U12006 ( .A1(n10812), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10403) );
  NAND2_X1 U12007 ( .A1(n12578), .A2(n10598), .ZN(n10597) );
  NAND2_X1 U12008 ( .A1(n13189), .A2(n10263), .ZN(n12429) );
  NAND2_X1 U12009 ( .A1(n10363), .A2(n10362), .ZN(n17548) );
  INV_X1 U12010 ( .A(n14956), .ZN(n10596) );
  NAND2_X1 U12011 ( .A1(n13156), .A2(n21645), .ZN(n10526) );
  INV_X1 U12012 ( .A(n21462), .ZN(n21326) );
  NOR2_X2 U12013 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21517) );
  INV_X1 U12014 ( .A(n21431), .ZN(n21588) );
  OAI21_X1 U12015 ( .B1(n15558), .B2(n21742), .A(n17530), .ZN(n21114) );
  NAND2_X1 U12016 ( .A1(n12528), .A2(n12527), .ZN(n12529) );
  INV_X1 U12017 ( .A(n12526), .ZN(n12527) );
  NAND4_X1 U12018 ( .A1(n11002), .A2(n11000), .A3(n11001), .A4(n10221), .ZN(
        n10220) );
  NOR2_X1 U12019 ( .A1(n11812), .A2(n11813), .ZN(n11804) );
  AND4_X1 U12020 ( .A1(n11467), .A2(n11466), .A3(n11465), .A4(n11464), .ZN(
        n15958) );
  AND2_X1 U12021 ( .A1(n20059), .A2(n15999), .ZN(n15975) );
  NAND2_X1 U12022 ( .A1(n11129), .A2(n11130), .ZN(n11133) );
  NAND2_X1 U12023 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10051) );
  NAND2_X1 U12024 ( .A1(n10705), .A2(n9798), .ZN(n10240) );
  AND3_X1 U12025 ( .A1(n16164), .A2(n16163), .A3(n16162), .ZN(n16435) );
  AND2_X1 U12026 ( .A1(n11642), .A2(n11641), .ZN(n15810) );
  NOR2_X1 U12027 ( .A1(n10724), .A2(n10723), .ZN(n10722) );
  INV_X1 U12028 ( .A(n16626), .ZN(n10723) );
  CLKBUF_X1 U12029 ( .A(n15785), .Z(n15786) );
  NOR2_X2 U12030 ( .A1(n13803), .A2(n13001), .ZN(n13942) );
  NAND2_X1 U12031 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10053) );
  NAND2_X1 U12032 ( .A1(n9991), .A2(n9945), .ZN(n9989) );
  INV_X1 U12033 ( .A(n13022), .ZN(n12017) );
  OAI21_X1 U12034 ( .B1(n11895), .B2(n11894), .A(n12987), .ZN(n12717) );
  OR2_X1 U12035 ( .A1(n10762), .A2(n14435), .ZN(n10761) );
  NAND2_X1 U12036 ( .A1(n16855), .A2(n9946), .ZN(n16647) );
  INV_X1 U12037 ( .A(n15678), .ZN(n10732) );
  NAND2_X1 U12038 ( .A1(n10461), .A2(n16895), .ZN(n10464) );
  AND4_X1 U12039 ( .A1(n16732), .A2(n11850), .A3(n16727), .A4(n16742), .ZN(
        n11851) );
  NOR2_X1 U12040 ( .A1(n16753), .A2(n10304), .ZN(n11850) );
  NAND2_X1 U12041 ( .A1(n10693), .A2(n16727), .ZN(n10690) );
  NOR2_X1 U12042 ( .A1(n16729), .A2(n16728), .ZN(n10691) );
  NOR2_X1 U12043 ( .A1(n10692), .A2(n10686), .ZN(n10685) );
  NAND2_X1 U12044 ( .A1(n16733), .A2(n16727), .ZN(n10692) );
  NAND2_X1 U12045 ( .A1(n10687), .A2(n10686), .ZN(n10684) );
  AOI21_X1 U12046 ( .B1(n10230), .B2(n10228), .A(n9891), .ZN(n10117) );
  NAND2_X1 U12047 ( .A1(n10234), .A2(n10228), .ZN(n10118) );
  INV_X1 U12048 ( .A(n16856), .ZN(n10060) );
  INV_X1 U12049 ( .A(n15875), .ZN(n10751) );
  NOR2_X1 U12050 ( .A1(n14267), .A2(n10729), .ZN(n14279) );
  OR2_X1 U12051 ( .A1(n14267), .A2(n14271), .ZN(n14273) );
  AND3_X1 U12052 ( .A1(n11502), .A2(n11501), .A3(n11500), .ZN(n14268) );
  NAND2_X1 U12053 ( .A1(n15932), .A2(n10717), .ZN(n10716) );
  CLKBUF_X1 U12054 ( .A(n14261), .Z(n14262) );
  NAND2_X1 U12055 ( .A1(n10718), .A2(n11637), .ZN(n10717) );
  INV_X1 U12056 ( .A(n11762), .ZN(n10718) );
  NAND2_X1 U12057 ( .A1(n9842), .A2(n10150), .ZN(n10040) );
  AND3_X1 U12058 ( .A1(n11478), .A2(n11477), .A3(n11476), .ZN(n15933) );
  NAND2_X1 U12059 ( .A1(n11127), .A2(n11128), .ZN(n10776) );
  OAI21_X1 U12060 ( .B1(n13989), .B2(n10286), .A(n20814), .ZN(n14204) );
  NAND2_X1 U12061 ( .A1(n10286), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14206) );
  NAND2_X1 U12062 ( .A1(n11694), .A2(n11693), .ZN(n17280) );
  AND2_X2 U12063 ( .A1(n10239), .A2(n14178), .ZN(n14179) );
  NOR2_X1 U12064 ( .A1(n20517), .A2(n20516), .ZN(n20522) );
  OR2_X1 U12065 ( .A1(n20817), .A2(n20824), .ZN(n20327) );
  NAND2_X1 U12066 ( .A1(n10674), .A2(n11015), .ZN(n10673) );
  BUF_X1 U12067 ( .A(n11265), .Z(n20616) );
  INV_X1 U12068 ( .A(n20660), .ZN(n20555) );
  NAND2_X1 U12069 ( .A1(n10594), .A2(n18017), .ZN(n10593) );
  INV_X1 U12070 ( .A(n17756), .ZN(n10594) );
  INV_X1 U12071 ( .A(n10572), .ZN(n10570) );
  NOR2_X1 U12072 ( .A1(n10573), .A2(n18043), .ZN(n10572) );
  NOR2_X1 U12073 ( .A1(n18722), .A2(n18017), .ZN(n10573) );
  NAND2_X1 U12074 ( .A1(n10814), .A2(n18761), .ZN(n10568) );
  NAND2_X1 U12075 ( .A1(n18390), .A2(n17465), .ZN(n18353) );
  INV_X1 U12076 ( .A(n18106), .ZN(n18332) );
  INV_X1 U12077 ( .A(n19366), .ZN(n18399) );
  NOR2_X1 U12078 ( .A1(n18540), .A2(n10324), .ZN(n18500) );
  INV_X1 U12079 ( .A(n18509), .ZN(n10325) );
  NAND2_X1 U12080 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12776) );
  OR2_X1 U12081 ( .A1(n17481), .A2(n14383), .ZN(n10545) );
  NOR3_X1 U12082 ( .A1(n14381), .A2(n14380), .A3(n18501), .ZN(n14383) );
  NOR2_X1 U12083 ( .A1(n19366), .A2(n18391), .ZN(n19793) );
  INV_X1 U12084 ( .A(n10846), .ZN(n10856) );
  NAND2_X1 U12085 ( .A1(n10839), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10564) );
  INV_X1 U12086 ( .A(n10579), .ZN(n10578) );
  NOR2_X1 U12087 ( .A1(n18957), .A2(n10577), .ZN(n10576) );
  NOR2_X1 U12088 ( .A1(n18956), .A2(n10582), .ZN(n10581) );
  INV_X1 U12089 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10582) );
  OR2_X1 U12090 ( .A1(n12837), .A2(n10445), .ZN(n10443) );
  INV_X1 U12091 ( .A(n13088), .ZN(n13095) );
  INV_X1 U12092 ( .A(n10209), .ZN(n13086) );
  NOR2_X1 U12093 ( .A1(n12852), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17634) );
  NOR2_X1 U12094 ( .A1(n12850), .A2(n10137), .ZN(n12852) );
  CLKBUF_X1 U12095 ( .A(n18700), .Z(n18707) );
  NOR2_X1 U12096 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12845), .ZN(
        n18753) );
  OAI21_X1 U12097 ( .B1(n12841), .B2(n10456), .A(n9755), .ZN(n12843) );
  INV_X1 U12098 ( .A(n12848), .ZN(n18806) );
  NOR2_X1 U12099 ( .A1(n19143), .A2(n18839), .ZN(n19141) );
  NAND2_X1 U12100 ( .A1(n18919), .A2(n12841), .ZN(n18825) );
  INV_X1 U12101 ( .A(n18939), .ZN(n10625) );
  NAND2_X1 U12102 ( .A1(n10208), .A2(n18974), .ZN(n18970) );
  OAI21_X1 U12103 ( .B1(n18975), .B2(n18976), .A(n19289), .ZN(n10208) );
  XNOR2_X1 U12104 ( .A(n12900), .B(n10407), .ZN(n12901) );
  INV_X1 U12105 ( .A(n18532), .ZN(n10407) );
  AOI21_X1 U12106 ( .B1(n12876), .B2(n12875), .A(n12874), .ZN(n19816) );
  NOR2_X2 U12107 ( .A1(n10875), .A2(n10874), .ZN(n19349) );
  AOI21_X1 U12108 ( .B1(n19807), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n10432) );
  OR2_X1 U12109 ( .A1(n19804), .A2(n19803), .ZN(n10431) );
  NAND2_X1 U12110 ( .A1(n14397), .A2(n14396), .ZN(n21735) );
  INV_X1 U12111 ( .A(n10397), .ZN(n10396) );
  AND2_X1 U12112 ( .A1(n20904), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20956) );
  OR2_X1 U12113 ( .A1(n14419), .A2(n14418), .ZN(n20948) );
  XNOR2_X1 U12114 ( .A(n14404), .B(n14420), .ZN(n14505) );
  NAND2_X1 U12115 ( .A1(n14575), .A2(n21027), .ZN(n10483) );
  INV_X1 U12116 ( .A(n15324), .ZN(n15316) );
  NAND2_X1 U12117 ( .A1(n9885), .A2(n10503), .ZN(n10502) );
  NAND2_X1 U12118 ( .A1(n17559), .A2(n15334), .ZN(n10503) );
  AND2_X1 U12119 ( .A1(n12691), .A2(n12661), .ZN(n21027) );
  OR2_X1 U12120 ( .A1(n12548), .A2(n12547), .ZN(n21012) );
  INV_X1 U12121 ( .A(n21517), .ZN(n21579) );
  INV_X1 U12122 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21389) );
  INV_X1 U12123 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21666) );
  AOI21_X1 U12124 ( .B1(n10669), .B2(n20040), .A(n14561), .ZN(n10668) );
  AND2_X1 U12125 ( .A1(n13122), .A2(n13121), .ZN(n13123) );
  NAND2_X1 U12126 ( .A1(n10297), .A2(n15740), .ZN(n13122) );
  NAND2_X1 U12127 ( .A1(n10288), .A2(n10287), .ZN(n10297) );
  NAND2_X1 U12128 ( .A1(n14438), .A2(n15740), .ZN(n14444) );
  AND2_X1 U12129 ( .A1(n13078), .A2(n13074), .ZN(n16003) );
  INV_X1 U12130 ( .A(n20041), .ZN(n20066) );
  AND2_X1 U12131 ( .A1(n13942), .A2(n20481), .ZN(n20041) );
  XNOR2_X1 U12132 ( .A(n14433), .B(n12704), .ZN(n16388) );
  XNOR2_X1 U12133 ( .A(n10455), .B(n10454), .ZN(n16518) );
  NAND2_X1 U12134 ( .A1(n10452), .A2(n10451), .ZN(n10455) );
  NAND2_X1 U12135 ( .A1(n14189), .A2(n14188), .ZN(n14190) );
  INV_X1 U12136 ( .A(n14187), .ZN(n10047) );
  NAND2_X1 U12137 ( .A1(n16855), .A2(n12007), .ZN(n16735) );
  NAND2_X1 U12138 ( .A1(n16778), .A2(n10698), .ZN(n10700) );
  NAND2_X1 U12139 ( .A1(n16768), .A2(n16769), .ZN(n10314) );
  NAND2_X1 U12140 ( .A1(n16778), .A2(n11995), .ZN(n16768) );
  NAND2_X1 U12141 ( .A1(n10227), .A2(n10231), .ZN(n16777) );
  NAND2_X1 U12142 ( .A1(n10234), .A2(n10310), .ZN(n10227) );
  AOI21_X1 U12143 ( .B1(n20042), .B2(n16935), .A(n16791), .ZN(n10517) );
  INV_X1 U12144 ( .A(n17306), .ZN(n16935) );
  INV_X1 U12145 ( .A(n16933), .ZN(n16924) );
  NAND2_X1 U12146 ( .A1(n13811), .A2(n12022), .ZN(n16921) );
  NOR2_X2 U12147 ( .A1(n13811), .A2(n20854), .ZN(n16899) );
  NAND3_X1 U12148 ( .A1(n20800), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20660), 
        .ZN(n17306) );
  INV_X1 U12149 ( .A(n16899), .ZN(n16942) );
  NAND2_X1 U12150 ( .A1(n12723), .A2(n10799), .ZN(n10179) );
  XNOR2_X1 U12151 ( .A(n12703), .B(n12702), .ZN(n12999) );
  NAND2_X1 U12152 ( .A1(n12984), .A2(n11674), .ZN(n16515) );
  XNOR2_X1 U12153 ( .A(n16641), .B(n16640), .ZN(n16956) );
  OR2_X1 U12154 ( .A1(n14432), .A2(n14431), .ZN(n16950) );
  NAND2_X1 U12155 ( .A1(n9889), .A2(n10082), .ZN(n16993) );
  AOI22_X1 U12156 ( .A1(n16674), .A2(n10087), .B1(n10084), .B2(n10083), .ZN(
        n10082) );
  NAND2_X1 U12157 ( .A1(n16676), .A2(n10089), .ZN(n10088) );
  OAI21_X1 U12158 ( .B1(n16684), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n9805), .ZN(n16994) );
  NAND2_X1 U12159 ( .A1(n16673), .A2(n16672), .ZN(n10090) );
  NAND2_X1 U12160 ( .A1(n10110), .A2(n12005), .ZN(n12008) );
  NAND2_X1 U12161 ( .A1(n10121), .A2(n10696), .ZN(n16755) );
  AND2_X1 U12162 ( .A1(n17081), .A2(n9929), .ZN(n10200) );
  INV_X1 U12163 ( .A(n16804), .ZN(n10316) );
  NAND2_X1 U12164 ( .A1(n10346), .A2(n10351), .ZN(n16793) );
  NAND2_X1 U12165 ( .A1(n16856), .A2(n17167), .ZN(n10076) );
  AND2_X1 U12166 ( .A1(n11897), .A2(n20836), .ZN(n17221) );
  OR2_X1 U12167 ( .A1(n11983), .A2(n11982), .ZN(n17241) );
  INV_X1 U12168 ( .A(n17221), .ZN(n17266) );
  INV_X1 U12169 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17269) );
  OR2_X1 U12170 ( .A1(n17283), .A2(n13993), .ZN(n20133) );
  INV_X1 U12171 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20821) );
  XOR2_X1 U12172 ( .A(n19987), .B(n19349), .Z(n20003) );
  INV_X1 U12173 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19992) );
  NOR2_X1 U12174 ( .A1(n17748), .A2(n18043), .ZN(n12967) );
  INV_X1 U12175 ( .A(n10589), .ZN(n17748) );
  INV_X1 U12176 ( .A(n10972), .ZN(n10973) );
  NOR3_X1 U12177 ( .A1(n10586), .A2(n17751), .A3(n10585), .ZN(n10584) );
  AND2_X1 U12178 ( .A1(n18074), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n10585) );
  NOR2_X1 U12179 ( .A1(n17755), .A2(n19917), .ZN(n10586) );
  NAND2_X1 U12180 ( .A1(n10593), .A2(n10590), .ZN(n10589) );
  INV_X1 U12181 ( .A(n17749), .ZN(n10590) );
  NAND2_X1 U12182 ( .A1(n10592), .A2(n17749), .ZN(n10591) );
  INV_X1 U12183 ( .A(n10593), .ZN(n10592) );
  NAND2_X1 U12184 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18091), .ZN(n18076) );
  INV_X1 U12185 ( .A(n18073), .ZN(n18091) );
  NAND2_X1 U12186 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18279), .ZN(n18252) );
  INV_X1 U12187 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18381) );
  NAND2_X1 U12188 ( .A1(n18481), .A2(n10339), .ZN(n18433) );
  NAND2_X1 U12189 ( .A1(n18481), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n18476) );
  NOR2_X1 U12190 ( .A1(n19375), .A2(n17537), .ZN(n18531) );
  INV_X1 U12191 ( .A(n18392), .ZN(n17537) );
  NAND2_X1 U12192 ( .A1(n18392), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n18540) );
  OR2_X1 U12193 ( .A1(n12940), .A2(n12939), .ZN(n12945) );
  NOR2_X1 U12194 ( .A1(n18861), .A2(n18852), .ZN(n18847) );
  INV_X1 U12195 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18852) );
  NOR3_X1 U12196 ( .A1(n9790), .A2(n18847), .A3(n9960), .ZN(n9959) );
  AND2_X1 U12197 ( .A1(n18852), .A2(n18861), .ZN(n9960) );
  INV_X1 U12198 ( .A(n18859), .ZN(n9961) );
  NOR2_X2 U12199 ( .A1(n19946), .A2(n18901), .ZN(n18865) );
  NAND2_X1 U12200 ( .A1(n18999), .A2(n18877), .ZN(n10360) );
  NAND2_X1 U12201 ( .A1(n18922), .A2(n19177), .ZN(n10359) );
  INV_X1 U12202 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19946) );
  OR2_X1 U12203 ( .A1(n12921), .A2(n12936), .ZN(n12928) );
  NAND2_X1 U12204 ( .A1(n17643), .A2(n17642), .ZN(n17644) );
  AOI21_X1 U12205 ( .B1(n17641), .B2(n19811), .A(n17640), .ZN(n17642) );
  NAND2_X1 U12206 ( .A1(n9965), .A2(n19328), .ZN(n19108) );
  OR2_X1 U12207 ( .A1(n19086), .A2(n19085), .ZN(n19109) );
  NAND2_X1 U12208 ( .A1(n19088), .A2(n19327), .ZN(n19135) );
  NAND2_X1 U12209 ( .A1(n19285), .A2(n19286), .ZN(n19284) );
  INV_X1 U12210 ( .A(n19327), .ZN(n19314) );
  INV_X1 U12211 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19805) );
  INV_X1 U12212 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19806) );
  INV_X1 U12213 ( .A(n12241), .ZN(n13690) );
  INV_X1 U12214 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13348) );
  NOR2_X1 U12215 ( .A1(n12218), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10557) );
  NAND2_X1 U12216 ( .A1(n12663), .A2(n12181), .ZN(n12540) );
  NOR2_X1 U12217 ( .A1(n12510), .A2(n12511), .ZN(n10500) );
  NAND2_X1 U12218 ( .A1(n20331), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10469) );
  NAND2_X1 U12219 ( .A1(n10186), .A2(n10185), .ZN(n11151) );
  NAND2_X1 U12220 ( .A1(n11266), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10186) );
  NAND2_X1 U12221 ( .A1(n20390), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10185) );
  NAND2_X1 U12222 ( .A1(n20487), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10309) );
  AOI22_X1 U12223 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20359), .B1(
        n20424), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11223) );
  NAND2_X1 U12224 ( .A1(n11265), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11219) );
  INV_X1 U12225 ( .A(n16206), .ZN(n11324) );
  NAND2_X1 U12226 ( .A1(n11091), .A2(n11090), .ZN(n9973) );
  AOI21_X1 U12227 ( .B1(n11118), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11072), .ZN(n11093) );
  OAI211_X1 U12228 ( .C1(n11968), .C2(n20732), .A(n11071), .B(n11070), .ZN(
        n11072) );
  NAND2_X1 U12229 ( .A1(n11076), .A2(n20161), .ZN(n11075) );
  NAND2_X1 U12230 ( .A1(n12470), .A2(n12469), .ZN(n12486) );
  OAI21_X1 U12231 ( .B1(n12458), .B2(n10420), .A(n9886), .ZN(n10416) );
  NAND2_X1 U12232 ( .A1(n10812), .A2(n12460), .ZN(n10419) );
  NAND2_X1 U12233 ( .A1(n10742), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10738) );
  AND2_X1 U12234 ( .A1(n12409), .A2(n12422), .ZN(n10384) );
  INV_X1 U12235 ( .A(n12420), .ZN(n10368) );
  NAND2_X1 U12236 ( .A1(n12664), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n12550) );
  NOR2_X1 U12237 ( .A1(n12203), .A2(n10522), .ZN(n10521) );
  NAND2_X1 U12238 ( .A1(n12208), .A2(n12191), .ZN(n10035) );
  AND2_X1 U12239 ( .A1(n12191), .A2(n12209), .ZN(n10036) );
  INV_X1 U12240 ( .A(n12305), .ZN(n12294) );
  INV_X1 U12241 ( .A(n10653), .ZN(n10377) );
  NOR2_X1 U12242 ( .A1(n12234), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10371) );
  NAND2_X1 U12243 ( .A1(n13749), .A2(n12096), .ZN(n12126) );
  NAND2_X1 U12244 ( .A1(n10012), .A2(n10011), .ZN(n12125) );
  NAND2_X1 U12245 ( .A1(n12111), .A2(n12178), .ZN(n10011) );
  NAND2_X1 U12246 ( .A1(n12176), .A2(n10013), .ZN(n10012) );
  NOR2_X1 U12247 ( .A1(n13687), .A2(n9996), .ZN(n9995) );
  INV_X1 U12248 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12275) );
  AOI21_X1 U12249 ( .B1(n9753), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A(n10028), .ZN(n12045) );
  AND3_X1 U12250 ( .A1(n10744), .A2(n15521), .A3(
        P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10028) );
  OR2_X1 U12251 ( .A1(n12318), .A2(n12317), .ZN(n12410) );
  NAND2_X1 U12252 ( .A1(n11779), .A2(n10645), .ZN(n10644) );
  AND2_X1 U12253 ( .A1(n16267), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11305) );
  NOR2_X1 U12254 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16184) );
  NAND2_X1 U12255 ( .A1(n10181), .A2(n11974), .ZN(n10180) );
  INV_X1 U12256 ( .A(n16721), .ZN(n10463) );
  NAND3_X1 U12257 ( .A1(n9972), .A2(n11834), .A3(n16721), .ZN(n10459) );
  NOR2_X1 U12258 ( .A1(n9789), .A2(n10233), .ZN(n10226) );
  AOI22_X1 U12259 ( .A1(n20616), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__5__SCAN_IN), .B2(n11266), .ZN(n11267) );
  NOR2_X1 U12260 ( .A1(n9829), .A2(n10710), .ZN(n10709) );
  INV_X1 U12261 ( .A(n10717), .ZN(n10710) );
  INV_X1 U12262 ( .A(n20054), .ZN(n10238) );
  AOI21_X1 U12263 ( .B1(n20054), .B2(n11864), .A(n11987), .ZN(n10237) );
  NAND2_X1 U12264 ( .A1(n9992), .A2(n11317), .ZN(n11340) );
  NAND2_X1 U12265 ( .A1(n20551), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10193) );
  NAND2_X1 U12266 ( .A1(n11266), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10192) );
  AND2_X1 U12267 ( .A1(n11298), .A2(n11297), .ZN(n9971) );
  AND3_X1 U12268 ( .A1(n11287), .A2(n11286), .A3(n11285), .ZN(n11730) );
  NAND2_X1 U12269 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10300) );
  NAND2_X1 U12270 ( .A1(n11328), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10301) );
  AND2_X1 U12271 ( .A1(n11250), .A2(n11251), .ZN(n10303) );
  AOI22_X1 U12272 ( .A1(n11200), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11329), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10302) );
  NOR2_X1 U12273 ( .A1(n11745), .A2(n11732), .ZN(n11731) );
  NAND2_X1 U12274 ( .A1(n11201), .A2(n10177), .ZN(n10649) );
  NOR2_X1 U12275 ( .A1(n9867), .A2(n10178), .ZN(n10177) );
  INV_X1 U12276 ( .A(n14349), .ZN(n16319) );
  AND2_X1 U12277 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16185) );
  NAND2_X1 U12278 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18088), .ZN(
        n10860) );
  AND2_X1 U12279 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12835), .ZN(
        n12836) );
  AND2_X1 U12280 ( .A1(n10540), .A2(n10539), .ZN(n10958) );
  NAND2_X1 U12281 ( .A1(n19799), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10539) );
  NAND2_X1 U12282 ( .A1(n10542), .A2(n10541), .ZN(n10540) );
  INV_X1 U12283 ( .A(n12859), .ZN(n10541) );
  OAI22_X1 U12284 ( .A1(n19953), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19803), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10957) );
  NAND2_X1 U12285 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19797), .ZN(
        n12859) );
  AOI21_X1 U12286 ( .B1(n10961), .B2(n9860), .A(n10530), .ZN(n10965) );
  AND2_X1 U12287 ( .A1(n19806), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10530) );
  INV_X1 U12288 ( .A(n10947), .ZN(n10328) );
  AOI21_X1 U12289 ( .B1(n18315), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n10336), .ZN(n10335) );
  INV_X1 U12290 ( .A(n10900), .ZN(n10333) );
  INV_X1 U12291 ( .A(n10898), .ZN(n10338) );
  NAND2_X1 U12292 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10337) );
  NAND2_X1 U12293 ( .A1(n14595), .A2(n10773), .ZN(n10772) );
  NAND2_X1 U12294 ( .A1(n12182), .A2(n21106), .ZN(n13749) );
  INV_X1 U12295 ( .A(n13737), .ZN(n13706) );
  AND2_X1 U12296 ( .A1(n10775), .A2(n14660), .ZN(n10774) );
  NOR2_X1 U12297 ( .A1(n14673), .A2(n14691), .ZN(n10775) );
  NAND2_X1 U12298 ( .A1(n13259), .A2(n13258), .ZN(n14863) );
  OR2_X1 U12299 ( .A1(n12333), .A2(n12332), .ZN(n12412) );
  NOR2_X1 U12300 ( .A1(n12232), .A2(n12231), .ZN(n12376) );
  NAND2_X1 U12301 ( .A1(n10812), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12368) );
  NAND2_X1 U12302 ( .A1(n15193), .A2(n15202), .ZN(n10525) );
  NAND2_X1 U12303 ( .A1(n12454), .A2(n10145), .ZN(n15203) );
  INV_X1 U12304 ( .A(n15192), .ZN(n10145) );
  NOR2_X1 U12305 ( .A1(n10385), .A2(n10383), .ZN(n12423) );
  NAND2_X1 U12306 ( .A1(n10176), .A2(n9845), .ZN(n10383) );
  NAND2_X1 U12307 ( .A1(n10747), .A2(n12403), .ZN(n10385) );
  OR2_X1 U12308 ( .A1(n12348), .A2(n12347), .ZN(n12434) );
  NAND2_X1 U12309 ( .A1(n15294), .A2(n12402), .ZN(n10370) );
  INV_X1 U12310 ( .A(n13749), .ZN(n13142) );
  INV_X1 U12311 ( .A(n15557), .ZN(n10490) );
  NAND2_X1 U12312 ( .A1(n14479), .A2(n10488), .ZN(n10487) );
  OR2_X1 U12313 ( .A1(n12535), .A2(n12178), .ZN(n10488) );
  OAI211_X1 U12314 ( .C1(n12437), .C2(n12305), .A(n12289), .B(n12288), .ZN(
        n12296) );
  NAND2_X1 U12315 ( .A1(n12293), .A2(n10612), .ZN(n10619) );
  AND2_X1 U12316 ( .A1(n21201), .A2(n12212), .ZN(n10612) );
  NAND2_X1 U12317 ( .A1(n21201), .A2(n10620), .ZN(n10618) );
  INV_X1 U12318 ( .A(n12218), .ZN(n10620) );
  CLKBUF_X1 U12319 ( .A(n12029), .Z(n12209) );
  NAND2_X1 U12320 ( .A1(n12566), .A2(n12176), .ZN(n14488) );
  NOR2_X1 U12321 ( .A1(n12123), .A2(n12122), .ZN(n12124) );
  INV_X1 U12322 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12050) );
  AND2_X1 U12323 ( .A1(n12300), .A2(n21582), .ZN(n21328) );
  NOR2_X1 U12324 ( .A1(n12159), .A2(n12158), .ZN(n12175) );
  INV_X1 U12325 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12157) );
  OR2_X1 U12326 ( .A1(n13687), .A2(n12143), .ZN(n12146) );
  NOR2_X1 U12327 ( .A1(n12104), .A2(n12275), .ZN(n12148) );
  NAND2_X1 U12328 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12130) );
  INV_X1 U12329 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12141) );
  INV_X1 U12330 ( .A(n21229), .ZN(n15575) );
  NAND2_X1 U12331 ( .A1(n12476), .A2(n12475), .ZN(n12526) );
  OR2_X1 U12332 ( .A1(n12474), .A2(n12473), .ZN(n12476) );
  NOR2_X1 U12333 ( .A1(n10498), .A2(n9830), .ZN(n10496) );
  NAND2_X2 U12334 ( .A1(n12305), .A2(n12304), .ZN(n12528) );
  AND2_X1 U12335 ( .A1(n14484), .A2(n14483), .ZN(n17500) );
  AND2_X1 U12336 ( .A1(n10994), .A2(n10995), .ZN(n10195) );
  AND4_X1 U12337 ( .A1(n10991), .A2(n10990), .A3(n10989), .A4(n10988), .ZN(
        n10992) );
  NOR2_X1 U12338 ( .A1(n11883), .A2(n11882), .ZN(n11892) );
  NOR2_X1 U12339 ( .A1(n11860), .A2(n11859), .ZN(n11861) );
  NAND2_X1 U12340 ( .A1(n16282), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10216) );
  AOI21_X1 U12341 ( .B1(n16340), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n11015), .ZN(n10218) );
  NAND2_X1 U12342 ( .A1(n10656), .A2(n15742), .ZN(n15730) );
  OAI21_X1 U12343 ( .B1(n15758), .B2(n10655), .A(n20059), .ZN(n10656) );
  AND2_X1 U12344 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12019) );
  INV_X1 U12345 ( .A(n11830), .ZN(n11783) );
  AND2_X1 U12346 ( .A1(n9791), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10657) );
  INV_X1 U12347 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16086) );
  NAND2_X1 U12348 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10661) );
  NOR2_X1 U12349 ( .A1(n15851), .A2(n10659), .ZN(n10658) );
  NAND2_X1 U12350 ( .A1(n16651), .A2(n9948), .ZN(n10795) );
  INV_X1 U12351 ( .A(n15621), .ZN(n10764) );
  NOR2_X1 U12352 ( .A1(n13003), .A2(n10737), .ZN(n10736) );
  INV_X1 U12353 ( .A(n15625), .ZN(n10737) );
  OR2_X1 U12354 ( .A1(n13083), .A2(n11894), .ZN(n10181) );
  OAI21_X1 U12355 ( .B1(n11873), .B2(n11894), .A(n16672), .ZN(n10792) );
  NAND2_X1 U12356 ( .A1(n15646), .A2(n11872), .ZN(n11886) );
  NAND2_X1 U12357 ( .A1(n11865), .A2(n11864), .ZN(n11870) );
  INV_X1 U12358 ( .A(n15682), .ZN(n11865) );
  AND2_X1 U12359 ( .A1(n15710), .A2(n15692), .ZN(n10733) );
  AND2_X1 U12360 ( .A1(n16794), .A2(n16785), .ZN(n11994) );
  NOR2_X1 U12361 ( .A1(n17103), .A2(n17091), .ZN(n10785) );
  INV_X1 U12362 ( .A(n16753), .ZN(n10119) );
  INV_X1 U12363 ( .A(n15768), .ZN(n10749) );
  OR2_X1 U12364 ( .A1(n15775), .A2(n11894), .ZN(n11837) );
  NAND2_X1 U12365 ( .A1(n15857), .A2(n9802), .ZN(n15823) );
  AND2_X1 U12366 ( .A1(n9792), .A2(n10099), .ZN(n9802) );
  INV_X1 U12367 ( .A(n15826), .ZN(n10099) );
  NOR2_X1 U12368 ( .A1(n16784), .A2(n10353), .ZN(n10352) );
  INV_X1 U12369 ( .A(n10355), .ZN(n10353) );
  INV_X1 U12370 ( .A(n10352), .ZN(n10349) );
  AND2_X1 U12371 ( .A1(n15903), .A2(n11918), .ZN(n10752) );
  AND2_X1 U12372 ( .A1(n16871), .A2(n16884), .ZN(n16824) );
  NAND2_X1 U12373 ( .A1(n16895), .A2(n10153), .ZN(n10152) );
  INV_X1 U12374 ( .A(n10472), .ZN(n9978) );
  INV_X1 U12375 ( .A(n11123), .ZN(n10265) );
  MUX2_X1 U12376 ( .A(n11729), .B(n11728), .S(n9742), .Z(n11747) );
  NAND2_X1 U12377 ( .A1(n10267), .A2(n10268), .ZN(n10782) );
  NAND2_X1 U12378 ( .A1(n10550), .A2(n11237), .ZN(n10267) );
  AND2_X1 U12379 ( .A1(n11077), .A2(n11078), .ZN(n10044) );
  NAND2_X1 U12380 ( .A1(n10191), .A2(n20181), .ZN(n11406) );
  AND2_X1 U12381 ( .A1(n13808), .A2(n11047), .ZN(n10511) );
  AND2_X1 U12382 ( .A1(n16319), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14177) );
  OR2_X1 U12383 ( .A1(n14349), .A2(n16086), .ZN(n14208) );
  AND2_X1 U12384 ( .A1(n16185), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17289) );
  AOI22_X1 U12385 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11033) );
  NAND2_X1 U12386 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10425) );
  OR2_X2 U12387 ( .A1(n18072), .A2(n10867), .ZN(n18239) );
  NAND2_X1 U12388 ( .A1(n10623), .A2(n10859), .ZN(n10867) );
  INV_X1 U12389 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10623) );
  AOI21_X1 U12390 ( .B1(n18284), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(n9968), .ZN(n12770) );
  AND2_X1 U12391 ( .A1(n12807), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9968) );
  NOR2_X1 U12392 ( .A1(n10860), .A2(n10867), .ZN(n12818) );
  NOR2_X1 U12393 ( .A1(n10869), .A2(n18072), .ZN(n12815) );
  NOR2_X1 U12394 ( .A1(n18773), .A2(n17863), .ZN(n17849) );
  NAND2_X1 U12395 ( .A1(n10581), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10579) );
  NAND2_X1 U12396 ( .A1(n17634), .A2(n9953), .ZN(n10209) );
  NOR2_X1 U12397 ( .A1(n10448), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10447) );
  INV_X1 U12398 ( .A(n10824), .ZN(n10448) );
  NAND2_X1 U12399 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10632) );
  AND2_X1 U12400 ( .A1(n12847), .A2(n19054), .ZN(n10633) );
  NAND2_X1 U12401 ( .A1(n10133), .A2(n10630), .ZN(n10132) );
  INV_X1 U12402 ( .A(n18751), .ZN(n10133) );
  OAI22_X1 U12403 ( .A1(n10961), .A2(n19805), .B1(n10962), .B2(n10960), .ZN(
        n12873) );
  OR2_X1 U12404 ( .A1(n10892), .A2(n10893), .ZN(n10953) );
  INV_X1 U12405 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19799) );
  NAND2_X1 U12406 ( .A1(n19804), .A2(n19803), .ZN(n10435) );
  AND2_X1 U12407 ( .A1(n12531), .A2(n12184), .ZN(n13866) );
  INV_X1 U12408 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14695) );
  INV_X1 U12409 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14460) );
  OR2_X1 U12410 ( .A1(n15110), .A2(n14398), .ZN(n13631) );
  AND2_X1 U12411 ( .A1(n12592), .A2(n12591), .ZN(n14940) );
  AND2_X1 U12412 ( .A1(n13452), .A2(n13451), .ZN(n14716) );
  INV_X1 U12413 ( .A(n15615), .ZN(n15614) );
  NAND2_X1 U12414 ( .A1(n13680), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14402) );
  INV_X1 U12415 ( .A(n13681), .ZN(n13680) );
  INV_X1 U12416 ( .A(n13256), .ZN(n13742) );
  NAND2_X1 U12417 ( .A1(n10770), .A2(n10769), .ZN(n10768) );
  INV_X1 U12418 ( .A(n14568), .ZN(n10769) );
  INV_X1 U12419 ( .A(n13603), .ZN(n13604) );
  INV_X1 U12420 ( .A(n13553), .ZN(n13554) );
  AND2_X1 U12421 ( .A1(n13580), .A2(n13579), .ZN(n14646) );
  OR2_X1 U12422 ( .A1(n15131), .A2(n14398), .ZN(n13580) );
  NOR2_X2 U12423 ( .A1(n13510), .A2(n14695), .ZN(n13511) );
  NAND2_X1 U12424 ( .A1(n13493), .A2(n13492), .ZN(n14689) );
  AND2_X1 U12425 ( .A1(n13426), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13427) );
  INV_X1 U12426 ( .A(n13425), .ZN(n13426) );
  AND2_X1 U12427 ( .A1(n13432), .A2(n13431), .ZN(n14733) );
  NAND2_X1 U12428 ( .A1(n13382), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13425) );
  AND2_X1 U12429 ( .A1(n13381), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13382) );
  INV_X1 U12430 ( .A(n13380), .ZN(n13381) );
  NAND2_X1 U12431 ( .A1(n13317), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13380) );
  INV_X1 U12432 ( .A(n13316), .ZN(n13317) );
  AND2_X1 U12433 ( .A1(n13262), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13356) );
  AND2_X1 U12434 ( .A1(n13261), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13262) );
  INV_X1 U12435 ( .A(n13260), .ZN(n13261) );
  AND2_X1 U12436 ( .A1(n13252), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13211) );
  NAND2_X1 U12437 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n13211), .ZN(
        n13260) );
  INV_X1 U12438 ( .A(n13190), .ZN(n13191) );
  INV_X1 U12439 ( .A(n15060), .ZN(n13182) );
  NAND2_X1 U12440 ( .A1(n13163), .A2(n13335), .ZN(n13172) );
  NOR2_X2 U12441 ( .A1(n14620), .A2(n12653), .ZN(n14578) );
  NAND2_X1 U12442 ( .A1(n15136), .A2(n15081), .ZN(n15084) );
  NOR2_X1 U12443 ( .A1(n9823), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10140) );
  AND2_X1 U12444 ( .A1(n9916), .A2(n14654), .ZN(n10607) );
  AND2_X1 U12445 ( .A1(n12641), .A2(n12640), .ZN(n14661) );
  AND2_X1 U12446 ( .A1(n14692), .A2(n9916), .ZN(n14663) );
  NAND2_X1 U12447 ( .A1(n10143), .A2(n9735), .ZN(n15136) );
  NAND2_X1 U12448 ( .A1(n14692), .A2(n10609), .ZN(n14675) );
  NAND2_X1 U12449 ( .A1(n14692), .A2(n14693), .ZN(n14674) );
  NAND2_X1 U12450 ( .A1(n10523), .A2(n10524), .ZN(n15152) );
  AND2_X1 U12451 ( .A1(n12628), .A2(n12627), .ZN(n14717) );
  NAND2_X1 U12452 ( .A1(n10524), .A2(n12458), .ZN(n15182) );
  AND2_X1 U12453 ( .A1(n12620), .A2(n12619), .ZN(n14757) );
  AND2_X1 U12454 ( .A1(n10603), .A2(n10605), .ZN(n10602) );
  INV_X1 U12455 ( .A(n14767), .ZN(n10603) );
  NAND2_X1 U12456 ( .A1(n10604), .A2(n10605), .ZN(n14787) );
  NOR2_X1 U12457 ( .A1(n14820), .A2(n14794), .ZN(n14795) );
  AND2_X1 U12458 ( .A1(n9809), .A2(n14839), .ZN(n10599) );
  NAND3_X1 U12459 ( .A1(n12578), .A2(n10598), .A3(n14949), .ZN(n10595) );
  AND2_X1 U12460 ( .A1(n17583), .A2(n17556), .ZN(n17563) );
  INV_X1 U12461 ( .A(n14287), .ZN(n12565) );
  OAI21_X1 U12462 ( .B1(n12586), .B2(n12555), .A(n12554), .ZN(n14014) );
  NAND2_X1 U12463 ( .A1(n12438), .A2(n10394), .ZN(n12389) );
  INV_X1 U12464 ( .A(n12386), .ZN(n10394) );
  NAND2_X1 U12465 ( .A1(n12271), .A2(n12270), .ZN(n13154) );
  INV_X1 U12466 ( .A(n12235), .ZN(n12236) );
  INV_X1 U12467 ( .A(n12290), .ZN(n12291) );
  INV_X1 U12468 ( .A(n10747), .ZN(n12373) );
  NOR2_X1 U12469 ( .A1(n12218), .A2(n10559), .ZN(n10262) );
  INV_X1 U12470 ( .A(n12212), .ZN(n10559) );
  NAND2_X1 U12471 ( .A1(n10611), .A2(n12218), .ZN(n10616) );
  NAND2_X1 U12472 ( .A1(n10619), .A2(n10618), .ZN(n10617) );
  NAND2_X1 U12473 ( .A1(n12375), .A2(n15575), .ZN(n10415) );
  INV_X1 U12474 ( .A(n12096), .ZN(n12095) );
  INV_X1 U12475 ( .A(n21384), .ZN(n21540) );
  NAND2_X1 U12476 ( .A1(n15521), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10745) );
  INV_X1 U12477 ( .A(n10744), .ZN(n10746) );
  INV_X1 U12478 ( .A(n10560), .ZN(n15541) );
  OR2_X1 U12479 ( .A1(n9770), .A2(n21139), .ZN(n21360) );
  INV_X1 U12480 ( .A(n21302), .ZN(n21436) );
  OR2_X1 U12481 ( .A1(n9770), .A2(n15604), .ZN(n21462) );
  INV_X1 U12482 ( .A(n21360), .ZN(n21507) );
  NOR2_X1 U12483 ( .A1(n21206), .A2(n21388), .ZN(n21547) );
  AND2_X1 U12484 ( .A1(n9770), .A2(n15604), .ZN(n21302) );
  AND2_X1 U12485 ( .A1(n9770), .A2(n21139), .ZN(n21538) );
  NAND2_X1 U12486 ( .A1(n21000), .A2(n15615), .ZN(n21102) );
  NAND2_X1 U12487 ( .A1(n21000), .A2(n15614), .ZN(n21104) );
  NAND2_X1 U12488 ( .A1(n21644), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17524) );
  OAI21_X1 U12489 ( .B1(n11243), .B2(n11358), .A(n11389), .ZN(n11722) );
  AOI21_X1 U12490 ( .B1(n11378), .B2(n11377), .A(n11376), .ZN(n11402) );
  AND2_X1 U12491 ( .A1(n10651), .A2(n11891), .ZN(n10650) );
  INV_X1 U12492 ( .A(n11882), .ZN(n10651) );
  AND2_X1 U12493 ( .A1(n10289), .A2(n15999), .ZN(n10287) );
  NOR2_X1 U12494 ( .A1(n16655), .A2(n10296), .ZN(n10295) );
  INV_X1 U12495 ( .A(n16667), .ZN(n10296) );
  NOR2_X1 U12496 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n10183) );
  NAND2_X1 U12497 ( .A1(n11874), .A2(n11875), .ZN(n11883) );
  INV_X1 U12498 ( .A(n11873), .ZN(n15646) );
  NAND2_X1 U12499 ( .A1(n11852), .A2(n9912), .ZN(n15662) );
  INV_X1 U12500 ( .A(n10277), .ZN(n10276) );
  OAI21_X1 U12501 ( .B1(n10279), .B2(n16708), .A(n16703), .ZN(n10277) );
  NOR2_X1 U12502 ( .A1(n11830), .A2(n9921), .ZN(n11786) );
  INV_X1 U12503 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U12504 ( .A1(n11783), .A2(n9815), .ZN(n11790) );
  AND2_X1 U12505 ( .A1(n11646), .A2(n11645), .ZN(n15770) );
  NAND2_X1 U12506 ( .A1(n13038), .A2(n9816), .ZN(n13043) );
  NOR2_X1 U12507 ( .A1(n10274), .A2(n10273), .ZN(n15788) );
  INV_X1 U12508 ( .A(n16773), .ZN(n10273) );
  OR2_X1 U12509 ( .A1(n15817), .A2(n16798), .ZN(n20043) );
  NAND2_X1 U12510 ( .A1(n15833), .A2(n16810), .ZN(n15817) );
  NAND2_X1 U12511 ( .A1(n12018), .A2(n9791), .ZN(n13032) );
  NOR2_X1 U12512 ( .A1(n15860), .A2(n16833), .ZN(n15845) );
  OR2_X1 U12513 ( .A1(n15871), .A2(n16845), .ZN(n15860) );
  OR2_X1 U12514 ( .A1(n11763), .A2(n10307), .ZN(n11815) );
  NAND2_X1 U12515 ( .A1(n10308), .A2(n11773), .ZN(n10307) );
  NAND2_X1 U12516 ( .A1(n11827), .A2(n11879), .ZN(n11817) );
  OR2_X1 U12517 ( .A1(n11763), .A2(n10306), .ZN(n11821) );
  NAND2_X1 U12518 ( .A1(n15887), .A2(n16861), .ZN(n15871) );
  AND2_X1 U12519 ( .A1(n15898), .A2(n16878), .ZN(n15887) );
  AND2_X1 U12520 ( .A1(n11770), .A2(n11769), .ZN(n15924) );
  NAND2_X1 U12521 ( .A1(n16932), .A2(n10281), .ZN(n15950) );
  NAND2_X1 U12522 ( .A1(n10285), .A2(n10284), .ZN(n14541) );
  NAND2_X1 U12523 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10284) );
  NAND2_X1 U12524 ( .A1(n15991), .A2(n10286), .ZN(n10285) );
  NOR2_X1 U12525 ( .A1(n14541), .A2(n16002), .ZN(n15973) );
  NAND2_X1 U12526 ( .A1(n16020), .A2(n16019), .ZN(n16026) );
  INV_X1 U12527 ( .A(n10249), .ZN(n10248) );
  OAI21_X1 U12528 ( .B1(n16237), .B2(n9913), .A(n10701), .ZN(n10249) );
  NAND2_X1 U12529 ( .A1(n10244), .A2(n10706), .ZN(n10243) );
  AND2_X1 U12530 ( .A1(n9843), .A2(n10707), .ZN(n10706) );
  AND3_X1 U12531 ( .A1(n11602), .A2(n11601), .A3(n11600), .ZN(n14358) );
  NAND2_X1 U12532 ( .A1(n14305), .A2(n14209), .ZN(n14308) );
  INV_X1 U12533 ( .A(n14208), .ZN(n14209) );
  AND2_X1 U12534 ( .A1(n13965), .A2(n13964), .ZN(n14189) );
  OR2_X1 U12535 ( .A1(n17345), .A2(n17346), .ZN(n13965) );
  NOR2_X1 U12536 ( .A1(n20093), .A2(n14193), .ZN(n14552) );
  AND2_X2 U12537 ( .A1(n13778), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n17305)
         );
  XNOR2_X1 U12538 ( .A(n12712), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13006) );
  NAND2_X1 U12539 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10052) );
  NOR2_X1 U12540 ( .A1(n13055), .A2(n15664), .ZN(n13058) );
  NOR2_X1 U12541 ( .A1(n16769), .A2(n10699), .ZN(n10698) );
  INV_X1 U12542 ( .A(n11995), .ZN(n10699) );
  AND2_X1 U12543 ( .A1(n11995), .A2(n11803), .ZN(n16776) );
  NAND2_X1 U12544 ( .A1(n10694), .A2(n10232), .ZN(n10231) );
  AND2_X1 U12545 ( .A1(n12018), .A2(n10658), .ZN(n13029) );
  NAND2_X1 U12546 ( .A1(n12018), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13027) );
  AND2_X1 U12547 ( .A1(n9854), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10663) );
  INV_X1 U12548 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16887) );
  NAND2_X1 U12549 ( .A1(n12016), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13018) );
  AND4_X1 U12550 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10662) );
  AND2_X1 U12551 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13007) );
  AND2_X1 U12552 ( .A1(n16639), .A2(n12720), .ZN(n12721) );
  NAND2_X1 U12553 ( .A1(n16855), .A2(n10096), .ZN(n10638) );
  AND2_X1 U12554 ( .A1(n9822), .A2(n10637), .ZN(n10096) );
  NOR2_X1 U12555 ( .A1(n16645), .A2(n11974), .ZN(n10637) );
  AND2_X1 U12556 ( .A1(n16662), .A2(n16974), .ZN(n16649) );
  INV_X1 U12557 ( .A(n10181), .ZN(n16651) );
  AND2_X1 U12558 ( .A1(n16648), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10319) );
  OR2_X1 U12559 ( .A1(n15628), .A2(n11894), .ZN(n16662) );
  NOR2_X1 U12560 ( .A1(n10322), .A2(n16685), .ZN(n10321) );
  NAND2_X1 U12561 ( .A1(n11886), .A2(n10792), .ZN(n16676) );
  INV_X1 U12562 ( .A(n16685), .ZN(n10089) );
  NAND2_X1 U12563 ( .A1(n10086), .A2(n10085), .ZN(n10084) );
  NAND2_X1 U12564 ( .A1(n16685), .A2(n16675), .ZN(n10085) );
  INV_X1 U12565 ( .A(n16676), .ZN(n10086) );
  NAND2_X1 U12566 ( .A1(n16676), .A2(n16675), .ZN(n10083) );
  NOR2_X1 U12567 ( .A1(n16676), .A2(n16686), .ZN(n10087) );
  AND2_X1 U12568 ( .A1(n11661), .A2(n11660), .ZN(n15655) );
  CLKBUF_X1 U12569 ( .A(n15639), .Z(n15640) );
  AND2_X1 U12570 ( .A1(n11659), .A2(n11658), .ZN(n15678) );
  AND2_X1 U12571 ( .A1(n16697), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9977) );
  NAND2_X1 U12572 ( .A1(n10756), .A2(n15708), .ZN(n10755) );
  INV_X1 U12573 ( .A(n10758), .ZN(n10756) );
  AND2_X1 U12574 ( .A1(n11653), .A2(n11652), .ZN(n15723) );
  AND2_X1 U12575 ( .A1(n11651), .A2(n11650), .ZN(n12948) );
  INV_X1 U12576 ( .A(n12010), .ZN(n10757) );
  NOR2_X1 U12577 ( .A1(n9954), .A2(n17115), .ZN(n10784) );
  INV_X1 U12578 ( .A(n9985), .ZN(n9982) );
  CLKBUF_X1 U12579 ( .A(n15754), .Z(n15755) );
  NAND2_X1 U12580 ( .A1(n11848), .A2(n12006), .ZN(n16741) );
  NAND2_X1 U12581 ( .A1(n10116), .A2(n10228), .ZN(n10121) );
  OR2_X1 U12582 ( .A1(n10234), .A2(n10230), .ZN(n10116) );
  NAND2_X1 U12583 ( .A1(n10697), .A2(n11997), .ZN(n10696) );
  INV_X1 U12584 ( .A(n10698), .ZN(n10697) );
  AND2_X1 U12585 ( .A1(n17124), .A2(n12958), .ZN(n17112) );
  CLKBUF_X1 U12586 ( .A(n15823), .Z(n15824) );
  NAND2_X1 U12587 ( .A1(n16783), .A2(n10352), .ZN(n10346) );
  NAND2_X1 U12588 ( .A1(n9923), .A2(n16806), .ZN(n10351) );
  INV_X1 U12589 ( .A(n16805), .ZN(n10354) );
  AND2_X1 U12590 ( .A1(n17164), .A2(n12957), .ZN(n17124) );
  NOR2_X1 U12591 ( .A1(n10357), .A2(n10356), .ZN(n10355) );
  INV_X1 U12592 ( .A(n16782), .ZN(n10357) );
  CLKBUF_X1 U12593 ( .A(n14300), .Z(n14301) );
  NAND2_X1 U12594 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10055) );
  CLKBUF_X1 U12595 ( .A(n14276), .Z(n14277) );
  NAND2_X1 U12596 ( .A1(n10207), .A2(n12957), .ZN(n16823) );
  INV_X1 U12597 ( .A(n16856), .ZN(n10207) );
  AND3_X1 U12598 ( .A1(n11544), .A2(n11543), .A3(n11542), .ZN(n14257) );
  AND2_X1 U12599 ( .A1(n17216), .A2(n11708), .ZN(n17176) );
  AND3_X1 U12600 ( .A1(n11523), .A2(n11522), .A3(n11521), .ZN(n14271) );
  INV_X1 U12601 ( .A(n14268), .ZN(n11503) );
  NAND2_X1 U12602 ( .A1(n10754), .A2(n10753), .ZN(n14340) );
  OAI21_X1 U12603 ( .B1(n20054), .B2(n11987), .A(n10113), .ZN(n10112) );
  NAND2_X1 U12604 ( .A1(n20054), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10115) );
  INV_X1 U12605 ( .A(n11317), .ZN(n10194) );
  NAND2_X1 U12606 ( .A1(n10126), .A2(n10125), .ZN(n11316) );
  NAND2_X1 U12607 ( .A1(n10202), .A2(n10780), .ZN(n10125) );
  INV_X1 U12608 ( .A(n10150), .ZN(n10202) );
  NAND2_X1 U12609 ( .A1(n10682), .A2(n10680), .ZN(n10679) );
  INV_X1 U12610 ( .A(n11756), .ZN(n10680) );
  AND3_X1 U12611 ( .A1(n11472), .A2(n11471), .A3(n11470), .ZN(n15943) );
  NAND2_X1 U12612 ( .A1(n9757), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10054) );
  NAND2_X1 U12613 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10050) );
  CLKBUF_X1 U12614 ( .A(n14315), .Z(n14316) );
  NAND2_X1 U12615 ( .A1(n11734), .A2(n15962), .ZN(n16915) );
  CLKBUF_X1 U12616 ( .A(n11980), .Z(n17327) );
  NAND2_X1 U12617 ( .A1(n9766), .A2(n17321), .ZN(n17322) );
  INV_X1 U12618 ( .A(n14175), .ZN(n14172) );
  AND2_X1 U12619 ( .A1(n20817), .A2(n20134), .ZN(n20192) );
  NAND2_X1 U12620 ( .A1(n11021), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11022) );
  NAND2_X1 U12621 ( .A1(n11016), .A2(n11015), .ZN(n11023) );
  AND2_X1 U12622 ( .A1(n20817), .A2(n20824), .ZN(n20801) );
  NOR3_X1 U12623 ( .A1(n20551), .A2(n17300), .A3(n20575), .ZN(n20554) );
  INV_X1 U12624 ( .A(n20176), .ZN(n20179) );
  INV_X1 U12625 ( .A(n20655), .ZN(n20356) );
  INV_X1 U12626 ( .A(n17336), .ZN(n17361) );
  NAND2_X1 U12627 ( .A1(n9981), .A2(n20854), .ZN(n17368) );
  INV_X1 U12628 ( .A(n11087), .ZN(n9981) );
  NAND2_X1 U12629 ( .A1(n12874), .A2(n12860), .ZN(n19814) );
  INV_X1 U12630 ( .A(n10956), .ZN(n12881) );
  NOR2_X1 U12631 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17857), .ZN(n17841) );
  INV_X1 U12632 ( .A(n18771), .ZN(n17863) );
  NOR2_X1 U12633 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17924), .ZN(n17906) );
  NOR2_X1 U12634 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17972), .ZN(n17961) );
  NAND2_X1 U12635 ( .A1(n20004), .A2(n18546), .ZN(n10969) );
  NAND2_X1 U12636 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n10535), .ZN(n10534) );
  NOR2_X1 U12637 ( .A1(n17792), .A2(n10536), .ZN(n10535) );
  NAND2_X1 U12638 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .ZN(n10536) );
  AND2_X1 U12639 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18210), .ZN(n18181) );
  INV_X1 U12640 ( .A(n17466), .ZN(n10543) );
  AND3_X1 U12641 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n18367), .ZN(n17465) );
  NOR2_X1 U12642 ( .A1(n18619), .A2(n10331), .ZN(n10330) );
  NOR2_X1 U12643 ( .A1(n9947), .A2(n10340), .ZN(n10339) );
  INV_X1 U12644 ( .A(n10341), .ZN(n10340) );
  NOR2_X1 U12645 ( .A1(n18565), .A2(n10342), .ZN(n10341) );
  INV_X1 U12646 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n10342) );
  NOR2_X1 U12647 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10457) );
  INV_X1 U12648 ( .A(n12733), .ZN(n18312) );
  INV_X1 U12649 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18694) );
  NOR2_X1 U12650 ( .A1(n17872), .A2(n10563), .ZN(n18734) );
  NAND2_X1 U12651 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18773) );
  NAND2_X1 U12652 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18812) );
  INV_X1 U12653 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18861) );
  INV_X1 U12654 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21906) );
  NAND2_X1 U12655 ( .A1(n10634), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10450) );
  NAND2_X1 U12656 ( .A1(n10628), .A2(n10630), .ZN(n10634) );
  NAND2_X1 U12657 ( .A1(n10631), .A2(n18718), .ZN(n10628) );
  OR2_X1 U12658 ( .A1(n10633), .A2(n18751), .ZN(n10631) );
  NAND2_X1 U12659 ( .A1(n10627), .A2(n10130), .ZN(n18701) );
  INV_X1 U12660 ( .A(n10131), .ZN(n10130) );
  OR2_X1 U12661 ( .A1(n18718), .A2(n10629), .ZN(n10627) );
  OAI21_X1 U12662 ( .B1(n10633), .B2(n10132), .A(n18920), .ZN(n10131) );
  NOR2_X1 U12663 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18920), .ZN(
        n18790) );
  OAI21_X1 U12664 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n9755), .A(
        n12843), .ZN(n12844) );
  AND2_X1 U12665 ( .A1(n9967), .A2(n9966), .ZN(n19088) );
  NAND2_X1 U12666 ( .A1(n19072), .A2(n19073), .ZN(n9966) );
  NAND2_X1 U12667 ( .A1(n19149), .A2(n19811), .ZN(n9967) );
  NOR3_X1 U12668 ( .A1(n19158), .A2(n22014), .A3(n19163), .ZN(n19134) );
  AND2_X1 U12669 ( .A1(n18827), .A2(n18855), .ZN(n18836) );
  NOR2_X1 U12670 ( .A1(n19181), .A2(n19174), .ZN(n19183) );
  NOR2_X1 U12671 ( .A1(n19227), .A2(n18895), .ZN(n19207) );
  NAND2_X1 U12672 ( .A1(n10439), .A2(n10436), .ZN(n19792) );
  AND2_X1 U12673 ( .A1(n12841), .A2(n18920), .ZN(n10129) );
  NAND2_X1 U12674 ( .A1(n18942), .A2(n12912), .ZN(n18927) );
  NAND2_X1 U12675 ( .A1(n18963), .A2(n12908), .ZN(n18950) );
  XNOR2_X1 U12676 ( .A(n12906), .B(n10406), .ZN(n18965) );
  NAND2_X1 U12677 ( .A1(n18965), .A2(n18964), .ZN(n18963) );
  NOR2_X1 U12678 ( .A1(n18987), .A2(n12828), .ZN(n18975) );
  NAND2_X1 U12679 ( .A1(n18975), .A2(n18976), .ZN(n18974) );
  NOR2_X1 U12680 ( .A1(n12826), .A2(n19000), .ZN(n18989) );
  NOR2_X1 U12681 ( .A1(n10956), .A2(n10361), .ZN(n12889) );
  AND2_X1 U12682 ( .A1(n10942), .A2(n19987), .ZN(n10361) );
  NOR2_X1 U12683 ( .A1(n10437), .A2(n19778), .ZN(n19796) );
  NAND2_X1 U12684 ( .A1(n10439), .A2(n10438), .ZN(n10437) );
  INV_X1 U12685 ( .A(n19793), .ZN(n10438) );
  INV_X1 U12686 ( .A(n10865), .ZN(n10422) );
  NOR3_X1 U12687 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19988), .ZN(n19685) );
  INV_X1 U12688 ( .A(n10953), .ZN(n19359) );
  INV_X1 U12689 ( .A(n14380), .ZN(n19363) );
  NOR2_X2 U12690 ( .A1(n10920), .A2(n10919), .ZN(n19366) );
  NAND2_X1 U12691 ( .A1(n19992), .A2(n19347), .ZN(n19421) );
  NOR2_X1 U12692 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20001), .ZN(n18732) );
  INV_X1 U12693 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20900) );
  INV_X1 U12694 ( .A(n20956), .ZN(n20901) );
  INV_X1 U12695 ( .A(n14596), .ZN(n14606) );
  INV_X1 U12696 ( .A(n14959), .ZN(n20974) );
  AND2_X2 U12697 ( .A1(n14016), .A2(n14486), .ZN(n20978) );
  NAND2_X1 U12698 ( .A1(n20978), .A2(n14017), .ZN(n14959) );
  NAND2_X1 U12699 ( .A1(n15066), .A2(n14962), .ZN(n15027) );
  NAND2_X1 U12700 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  NAND2_X1 U12701 ( .A1(n15066), .A2(n14166), .ZN(n15064) );
  INV_X1 U12702 ( .A(n15026), .ZN(n15067) );
  OR3_X1 U12703 ( .A1(n14397), .A2(n14087), .A3(n17521), .ZN(n20982) );
  NAND2_X2 U12704 ( .A1(n20982), .A2(n14160), .ZN(n20985) );
  INV_X1 U12705 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15172) );
  INV_X1 U12706 ( .A(n20873), .ZN(n21001) );
  NAND2_X1 U12707 ( .A1(n14501), .A2(n10254), .ZN(n10251) );
  NAND2_X1 U12708 ( .A1(n10255), .A2(n14503), .ZN(n10250) );
  INV_X1 U12709 ( .A(n15069), .ZN(n10482) );
  OAI21_X1 U12710 ( .B1(n10743), .B2(n10004), .A(n10003), .ZN(n10380) );
  NAND2_X1 U12711 ( .A1(n10554), .A2(n9801), .ZN(n10743) );
  NAND2_X1 U12712 ( .A1(n10005), .A2(n10006), .ZN(n10004) );
  OR3_X1 U12713 ( .A1(n15363), .A2(n15338), .A3(n15335), .ZN(n15324) );
  XNOR2_X1 U12714 ( .A(n10477), .B(n15099), .ZN(n15332) );
  NAND2_X1 U12715 ( .A1(n10479), .A2(n10478), .ZN(n10477) );
  NAND2_X1 U12716 ( .A1(n15097), .A2(n10812), .ZN(n10479) );
  NAND2_X1 U12717 ( .A1(n15098), .A2(n15257), .ZN(n10478) );
  NAND2_X1 U12718 ( .A1(n17561), .A2(n12698), .ZN(n10504) );
  NAND2_X1 U12719 ( .A1(n10417), .A2(n10742), .ZN(n15143) );
  NAND2_X1 U12720 ( .A1(n10523), .A2(n9868), .ZN(n10417) );
  INV_X1 U12721 ( .A(n10505), .ZN(n15388) );
  OR2_X1 U12722 ( .A1(n15374), .A2(n15463), .ZN(n12685) );
  NAND2_X1 U12723 ( .A1(n10158), .A2(n10031), .ZN(n15227) );
  INV_X1 U12724 ( .A(n10032), .ZN(n10404) );
  OR2_X1 U12725 ( .A1(n13791), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17570) );
  NAND2_X1 U12726 ( .A1(n10259), .A2(n12431), .ZN(n17542) );
  NAND2_X1 U12727 ( .A1(n17548), .A2(n12430), .ZN(n10259) );
  INV_X1 U12728 ( .A(n21012), .ZN(n21042) );
  INV_X1 U12729 ( .A(n17570), .ZN(n21051) );
  NAND2_X1 U12730 ( .A1(n10614), .A2(n10613), .ZN(n21327) );
  NAND2_X1 U12731 ( .A1(n10653), .A2(n10621), .ZN(n10613) );
  INV_X1 U12732 ( .A(n10617), .ZN(n10614) );
  INV_X1 U12733 ( .A(n10616), .ZN(n10621) );
  INV_X1 U12734 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21057) );
  OAI21_X1 U12735 ( .B1(n15559), .B2(n17604), .A(n21206), .ZN(n21056) );
  INV_X1 U12736 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17596) );
  OAI21_X1 U12737 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21474), .A(n17591), 
        .ZN(n17597) );
  NOR2_X1 U12738 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n17592) );
  OR2_X1 U12739 ( .A1(n21175), .A2(n21360), .ZN(n21160) );
  OAI21_X1 U12740 ( .B1(n21147), .B2(n21146), .A(n21145), .ZN(n21168) );
  OAI211_X1 U12741 ( .C1(n21349), .C2(n21474), .A(n21391), .B(n21334), .ZN(
        n21352) );
  INV_X1 U12742 ( .A(n21395), .ZN(n21420) );
  OAI22_X1 U12743 ( .A1(n21428), .A2(n21579), .B1(n21432), .B2(n21647), .ZN(
        n21457) );
  OAI211_X1 U12744 ( .C1(n21517), .C2(n21516), .A(n21588), .B(n21515), .ZN(
        n21535) );
  INV_X1 U12745 ( .A(n21543), .ZN(n21572) );
  AND2_X1 U12746 ( .A1(n21114), .A2(n15607), .ZN(n21584) );
  AND2_X1 U12747 ( .A1(n21060), .A2(n21105), .ZN(n21595) );
  AND2_X1 U12748 ( .A1(n21114), .A2(n21063), .ZN(n21596) );
  AND2_X1 U12749 ( .A1(n21114), .A2(n21073), .ZN(n21602) );
  INV_X1 U12750 ( .A(n21402), .ZN(n21607) );
  AND2_X1 U12751 ( .A1(n21114), .A2(n21078), .ZN(n21608) );
  AND2_X1 U12752 ( .A1(n12233), .A2(n21105), .ZN(n21613) );
  AND2_X1 U12753 ( .A1(n21114), .A2(n21085), .ZN(n21614) );
  AND2_X1 U12754 ( .A1(n21114), .A2(n21093), .ZN(n21620) );
  INV_X1 U12755 ( .A(n21642), .ZN(n21628) );
  AND2_X1 U12756 ( .A1(n12182), .A2(n21105), .ZN(n21625) );
  AND2_X1 U12757 ( .A1(n21114), .A2(n21098), .ZN(n21626) );
  OAI21_X1 U12758 ( .B1(n21590), .B2(n21589), .A(n21588), .ZN(n21639) );
  INV_X1 U12759 ( .A(n21417), .ZN(n21633) );
  AND2_X1 U12760 ( .A1(n21114), .A2(n21109), .ZN(n21636) );
  NAND3_X1 U12761 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21645), .A3(n15557), 
        .ZN(n17530) );
  OR2_X1 U12762 ( .A1(n17524), .A2(n21645), .ZN(n20866) );
  INV_X2 U12763 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21647) );
  INV_X1 U12764 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21644) );
  NAND2_X1 U12765 ( .A1(n21661), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21746) );
  NAND2_X1 U12766 ( .A1(n10294), .A2(n9814), .ZN(n14437) );
  NAND2_X1 U12767 ( .A1(n13063), .A2(n10295), .ZN(n10294) );
  INV_X1 U12768 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15739) );
  NAND2_X1 U12769 ( .A1(n20847), .A2(n13076), .ZN(n16009) );
  AND2_X1 U12770 ( .A1(n11806), .A2(n11809), .ZN(n15821) );
  NAND2_X1 U12771 ( .A1(n14324), .A2(n11462), .ZN(n15959) );
  INV_X1 U12772 ( .A(n15975), .ZN(n16015) );
  INV_X1 U12773 ( .A(n15740), .ZN(n20038) );
  AND2_X1 U12774 ( .A1(n16009), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20031) );
  NAND2_X1 U12775 ( .A1(n10283), .A2(n10282), .ZN(n16002) );
  NAND2_X1 U12776 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U12777 ( .A1(n10286), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10283) );
  NOR2_X1 U12778 ( .A1(n20077), .A2(n20078), .ZN(n20075) );
  INV_X1 U12779 ( .A(n20076), .ZN(n16497) );
  AND2_X1 U12780 ( .A1(n13995), .A2(n17372), .ZN(n20082) );
  INV_X2 U12781 ( .A(n20082), .ZN(n16503) );
  NAND2_X1 U12782 ( .A1(n20082), .A2(n20181), .ZN(n20076) );
  NAND2_X1 U12783 ( .A1(n10246), .A2(n16391), .ZN(n16519) );
  NAND2_X1 U12784 ( .A1(n16396), .A2(n10240), .ZN(n16403) );
  AND2_X1 U12785 ( .A1(n14552), .A2(n17305), .ZN(n16615) );
  NOR2_X2 U12786 ( .A1(n20093), .A2(n14192), .ZN(n16618) );
  NAND2_X1 U12787 ( .A1(n10719), .A2(n10722), .ZN(n15809) );
  INV_X1 U12788 ( .A(n14300), .ZN(n10719) );
  AND2_X1 U12789 ( .A1(n16625), .A2(n20085), .ZN(n16637) );
  OR2_X1 U12790 ( .A1(n16618), .A2(n14552), .ZN(n16634) );
  INV_X1 U12791 ( .A(n20133), .ZN(n20198) );
  INV_X1 U12792 ( .A(n16625), .ZN(n22058) );
  INV_X1 U12793 ( .A(n16634), .ZN(n22062) );
  INV_X1 U12794 ( .A(n13977), .ZN(n14053) );
  NAND2_X1 U12795 ( .A1(n13878), .A2(n20853), .ZN(n20132) );
  OAI21_X1 U12796 ( .B1(n13876), .B2(n13875), .A(n13958), .ZN(n13878) );
  INV_X1 U12797 ( .A(n20101), .ZN(n20130) );
  INV_X1 U12798 ( .A(n13942), .ZN(n13857) );
  NAND2_X1 U12799 ( .A1(n13958), .A2(n13857), .ZN(n13907) );
  INV_X1 U12800 ( .A(n16921), .ZN(n16930) );
  NAND2_X1 U12801 ( .A1(n10187), .A2(n16639), .ZN(n10465) );
  NAND2_X1 U12802 ( .A1(n10188), .A2(n16638), .ZN(n10187) );
  XNOR2_X1 U12803 ( .A(n10638), .B(n12987), .ZN(n14473) );
  INV_X1 U12804 ( .A(n16684), .ZN(n16694) );
  INV_X1 U12805 ( .A(n16715), .ZN(n16714) );
  NAND2_X1 U12806 ( .A1(n10462), .A2(n11851), .ZN(n16724) );
  NAND2_X1 U12807 ( .A1(n10464), .A2(n9863), .ZN(n10462) );
  OAI21_X1 U12808 ( .B1(n10693), .B2(n10691), .A(n10690), .ZN(n10689) );
  INV_X1 U12809 ( .A(n10313), .ZN(n10312) );
  OAI21_X1 U12810 ( .B1(n17089), .B2(n17241), .A(n17088), .ZN(n10313) );
  NAND2_X1 U12811 ( .A1(n10060), .A2(n10059), .ZN(n17138) );
  NAND2_X1 U12812 ( .A1(n16823), .A2(n10077), .ZN(n17162) );
  NAND2_X1 U12813 ( .A1(n10078), .A2(n17155), .ZN(n10077) );
  NAND2_X1 U12814 ( .A1(n16858), .A2(n16857), .ZN(n10049) );
  INV_X1 U12815 ( .A(n10711), .ZN(n14264) );
  AOI21_X1 U12816 ( .B1(n10716), .B2(n10715), .A(n9829), .ZN(n10711) );
  OR2_X1 U12817 ( .A1(n15932), .A2(n15933), .ZN(n10714) );
  INV_X1 U12818 ( .A(n10781), .ZN(n16908) );
  AND2_X1 U12819 ( .A1(n11697), .A2(n17225), .ZN(n17254) );
  CLKBUF_X1 U12820 ( .A(n16938), .Z(n17261) );
  OR2_X1 U12821 ( .A1(n11983), .A2(n11696), .ZN(n17082) );
  INV_X1 U12822 ( .A(n10776), .ZN(n11135) );
  NAND2_X1 U12823 ( .A1(n17281), .A2(n13988), .ZN(n10440) );
  INV_X2 U12824 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21769) );
  INV_X1 U12825 ( .A(n20824), .ZN(n20134) );
  NAND2_X1 U12826 ( .A1(n10095), .A2(n13975), .ZN(n17355) );
  OAI21_X1 U12827 ( .B1(n20225), .B2(n20808), .A(n20222), .ZN(n20245) );
  INV_X1 U12828 ( .A(n20271), .ZN(n20290) );
  OAI22_X1 U12829 ( .A1(n20298), .A2(n17300), .B1(n20297), .B2(n20303), .ZN(
        n20321) );
  OAI211_X1 U12830 ( .C1(n20350), .C2(n20329), .A(n20328), .B(n20660), .ZN(
        n20353) );
  AND2_X1 U12831 ( .A1(n20357), .A2(n20294), .ZN(n20351) );
  AND2_X1 U12832 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20330), .ZN(
        n20350) );
  OAI21_X1 U12833 ( .B1(n20388), .B2(n20489), .A(n20360), .ZN(n20383) );
  AOI211_X2 U12834 ( .C1(n17300), .C2(n20393), .A(n20552), .B(n20391), .ZN(
        n20411) );
  OAI211_X1 U12835 ( .C1(n20457), .C2(n20453), .A(n20660), .B(n20452), .ZN(
        n20475) );
  OAI21_X1 U12836 ( .B1(n20457), .B2(n20456), .A(n20455), .ZN(n20474) );
  AND2_X1 U12837 ( .A1(n20486), .A2(n20660), .ZN(n20492) );
  OAI21_X1 U12838 ( .B1(n20513), .B2(n20489), .A(n20488), .ZN(n20507) );
  INV_X1 U12839 ( .A(n20541), .ZN(n20544) );
  AOI21_X1 U12840 ( .B1(n17300), .B2(n20518), .A(n20522), .ZN(n20543) );
  AOI211_X2 U12841 ( .C1(n17300), .C2(n20556), .A(n20552), .B(n20554), .ZN(
        n20576) );
  NAND2_X1 U12842 ( .A1(n17304), .A2(n17303), .ZN(n20605) );
  OAI21_X1 U12843 ( .B1(n11266), .B2(n17300), .A(n20814), .ZN(n17302) );
  OAI21_X1 U12844 ( .B1(n20550), .B2(n20808), .A(n17308), .ZN(n20602) );
  OAI21_X1 U12845 ( .B1(n11266), .B2(n20615), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17308) );
  NAND2_X1 U12846 ( .A1(n20618), .A2(n20617), .ZN(n20646) );
  INV_X1 U12847 ( .A(n20369), .ZN(n20662) );
  INV_X1 U12848 ( .A(n20702), .ZN(n20709) );
  OAI21_X1 U12849 ( .B1(n20654), .B2(n20808), .A(n20651), .ZN(n20707) );
  INV_X1 U12850 ( .A(n20699), .ZN(n20713) );
  NAND3_X1 U12851 ( .A1(n17365), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17617) );
  INV_X1 U12852 ( .A(n20850), .ZN(n20844) );
  INV_X1 U12853 ( .A(n17617), .ZN(n17372) );
  AND2_X1 U12854 ( .A1(n10286), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17375) );
  INV_X1 U12855 ( .A(n13877), .ZN(n20853) );
  INV_X1 U12856 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20732) );
  INV_X1 U12857 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20734) );
  NAND2_X1 U12858 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20728), .ZN(n20863) );
  NOR2_X1 U12859 ( .A1(n19813), .A2(n18598), .ZN(n20004) );
  INV_X1 U12860 ( .A(n12934), .ZN(n17734) );
  INV_X1 U12861 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17764) );
  NAND2_X1 U12862 ( .A1(n10574), .A2(n10847), .ZN(n10571) );
  NAND2_X1 U12863 ( .A1(n10570), .A2(n10574), .ZN(n10569) );
  INV_X1 U12864 ( .A(n18713), .ZN(n10574) );
  OAI21_X1 U12865 ( .B1(n17822), .B2(n18722), .A(n10572), .ZN(n10575) );
  NOR2_X1 U12866 ( .A1(n17809), .A2(n18722), .ZN(n17808) );
  AND2_X1 U12867 ( .A1(n17822), .A2(n18017), .ZN(n17809) );
  INV_X1 U12868 ( .A(n18055), .ZN(n18081) );
  NOR4_X1 U12869 ( .A1(n19898), .A2(n19896), .A3(n19894), .A4(n17847), .ZN(
        n17836) );
  NAND2_X1 U12870 ( .A1(n10567), .A2(n10566), .ZN(n17831) );
  INV_X1 U12871 ( .A(n10568), .ZN(n10565) );
  NAND2_X1 U12872 ( .A1(n17851), .A2(n10814), .ZN(n17839) );
  NOR2_X1 U12873 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17878), .ZN(n17861) );
  NOR2_X1 U12874 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17898), .ZN(n17886) );
  INV_X1 U12875 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17950) );
  NOR2_X1 U12876 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18046), .ZN(n18032) );
  NAND2_X1 U12877 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n18143), .ZN(n18130) );
  INV_X1 U12878 ( .A(n18130), .ZN(n18140) );
  NOR2_X1 U12879 ( .A1(n18170), .A2(n10532), .ZN(n18143) );
  NAND2_X1 U12880 ( .A1(n10533), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n10532) );
  INV_X1 U12881 ( .A(n10534), .ZN(n10533) );
  NOR2_X1 U12882 ( .A1(n18170), .A2(n10534), .ZN(n18148) );
  NOR3_X1 U12883 ( .A1(n18170), .A2(n21800), .A3(n10536), .ZN(n18151) );
  NOR2_X1 U12884 ( .A1(n18170), .A2(n10536), .ZN(n18157) );
  NAND2_X1 U12885 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18183), .ZN(n18170) );
  AND2_X1 U12886 ( .A1(n19375), .A2(n18181), .ZN(n18183) );
  NOR3_X1 U12887 ( .A1(n9832), .A2(n18195), .A3(n18224), .ZN(n18210) );
  INV_X1 U12888 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n18224) );
  NAND2_X1 U12889 ( .A1(n18265), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n18249) );
  NOR2_X1 U12890 ( .A1(n18252), .A2(n17900), .ZN(n18265) );
  NAND2_X1 U12891 ( .A1(n18364), .A2(n9819), .ZN(n17463) );
  AND2_X1 U12892 ( .A1(n18364), .A2(n9944), .ZN(n18279) );
  NAND2_X1 U12893 ( .A1(n18364), .A2(n17464), .ZN(n18354) );
  INV_X1 U12894 ( .A(n18353), .ZN(n18364) );
  INV_X1 U12895 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18371) );
  AND2_X1 U12896 ( .A1(n10545), .A2(n10544), .ZN(n18390) );
  NOR3_X1 U12897 ( .A1(n19349), .A2(n19987), .A3(n19836), .ZN(n10544) );
  INV_X1 U12898 ( .A(n18409), .ZN(n18405) );
  NAND2_X1 U12899 ( .A1(n18421), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n18417) );
  NOR2_X1 U12900 ( .A1(n18616), .A2(n18427), .ZN(n18421) );
  OR2_X1 U12901 ( .A1(n18614), .A2(n18426), .ZN(n18427) );
  NOR2_X1 U12902 ( .A1(n18601), .A2(n18464), .ZN(n18460) );
  NOR2_X2 U12903 ( .A1(n18399), .A2(n18523), .ZN(n18463) );
  AND2_X1 U12904 ( .A1(n18500), .A2(n18395), .ZN(n18481) );
  NOR2_X1 U12905 ( .A1(n12753), .A2(n12752), .ZN(n18516) );
  INV_X1 U12906 ( .A(n18531), .ZN(n18523) );
  INV_X1 U12907 ( .A(n18538), .ZN(n18528) );
  NOR2_X1 U12908 ( .A1(n18590), .A2(n18530), .ZN(n18529) );
  AND4_X1 U12909 ( .A1(n12784), .A2(n12783), .A3(n12782), .A4(n12781), .ZN(
        n12785) );
  INV_X1 U12910 ( .A(n17536), .ZN(n10326) );
  INV_X1 U12911 ( .A(n10545), .ZN(n17535) );
  AND2_X1 U12912 ( .A1(n19793), .A2(n18392), .ZN(n18537) );
  NOR2_X1 U12913 ( .A1(n19793), .A2(n18523), .ZN(n18538) );
  NOR3_X1 U12914 ( .A1(n18545), .A2(n19986), .A3(n18598), .ZN(n18568) );
  CLKBUF_X1 U12915 ( .A(n18648), .Z(n18637) );
  NOR2_X2 U12916 ( .A1(n18598), .A2(n19828), .ZN(n18649) );
  INV_X1 U12917 ( .A(n18644), .ZN(n18651) );
  INV_X1 U12918 ( .A(n18656), .ZN(n19020) );
  INV_X1 U12919 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n22029) );
  NAND2_X1 U12920 ( .A1(n10562), .A2(n10826), .ZN(n10561) );
  INV_X1 U12921 ( .A(n10563), .ZN(n10562) );
  INV_X1 U12922 ( .A(n18819), .ZN(n18794) );
  INV_X1 U12923 ( .A(n18957), .ZN(n10580) );
  INV_X1 U12924 ( .A(n10211), .ZN(n18933) );
  NAND2_X1 U12925 ( .A1(n10212), .A2(n10441), .ZN(n18934) );
  INV_X1 U12926 ( .A(n19369), .ZN(n19659) );
  NOR2_X1 U12927 ( .A1(n18957), .A2(n18956), .ZN(n18941) );
  INV_X1 U12928 ( .A(n19009), .ZN(n18980) );
  INV_X1 U12929 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19006) );
  INV_X1 U12930 ( .A(n19012), .ZN(n19003) );
  AOI21_X1 U12931 ( .B1(n13134), .B2(n19240), .A(n13109), .ZN(n13110) );
  OAI21_X1 U12932 ( .B1(n13091), .B2(n13089), .A(n13090), .ZN(n13092) );
  NAND2_X1 U12933 ( .A1(n17634), .A2(n18655), .ZN(n17490) );
  NOR2_X1 U12934 ( .A1(n19031), .A2(n10408), .ZN(n19023) );
  OR2_X1 U12935 ( .A1(n19314), .A2(n10409), .ZN(n10408) );
  AND2_X1 U12936 ( .A1(n19326), .A2(n12851), .ZN(n10409) );
  INV_X1 U12937 ( .A(n17633), .ZN(n18671) );
  NAND2_X1 U12938 ( .A1(n10412), .A2(n10410), .ZN(n19031) );
  AOI21_X1 U12939 ( .B1(n19019), .B2(n19073), .A(n10411), .ZN(n10410) );
  OR2_X1 U12940 ( .A1(n18656), .A2(n19307), .ZN(n10412) );
  NAND2_X1 U12941 ( .A1(n19040), .A2(n19021), .ZN(n10411) );
  NAND2_X1 U12942 ( .A1(n18718), .A2(n12847), .ZN(n18708) );
  OR3_X1 U12943 ( .A1(n18752), .A2(n18741), .A3(n19084), .ZN(n18719) );
  INV_X1 U12944 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19127) );
  INV_X1 U12945 ( .A(n12843), .ZN(n18805) );
  INV_X1 U12946 ( .A(n18877), .ZN(n19203) );
  INV_X1 U12947 ( .A(n19117), .ZN(n19292) );
  NAND2_X1 U12948 ( .A1(n18990), .A2(n12904), .ZN(n19285) );
  AOI21_X2 U12949 ( .B1(n12879), .B2(n12878), .A(n19836), .ZN(n19327) );
  AOI211_X1 U12950 ( .C1(n12870), .C2(n19817), .A(n12869), .B(n17479), .ZN(
        n12879) );
  INV_X1 U12951 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19797) );
  INV_X1 U12952 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19803) );
  NOR2_X1 U12953 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19805), .ZN(
        n19604) );
  CLKBUF_X1 U12954 ( .A(n18088), .Z(n19967) );
  AOI211_X1 U12955 ( .C1(n19985), .C2(n19823), .A(n19348), .B(n17482), .ZN(
        n19968) );
  INV_X1 U12956 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19824) );
  NOR2_X1 U12957 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20002) );
  NOR2_X1 U12958 ( .A1(n19826), .A2(n10429), .ZN(n19837) );
  NAND2_X1 U12959 ( .A1(n10430), .A2(n9862), .ZN(n10429) );
  INV_X1 U12960 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19937) );
  OAI211_X1 U12961 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19861), .B(n19922), .ZN(n19986) );
  INV_X1 U12962 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19861) );
  NAND2_X1 U12963 ( .A1(n19861), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19999) );
  AND2_X1 U12964 ( .A1(n13759), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15615)
         );
  INV_X1 U12965 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21968) );
  OR2_X1 U12966 ( .A1(n17307), .A2(n13779), .ZN(n17654) );
  CLKBUF_X1 U12967 ( .A(n17722), .Z(n17721) );
  NAND2_X1 U12968 ( .A1(n21740), .A2(n10396), .ZN(n21741) );
  AND4_X1 U12969 ( .A1(n20920), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20921) );
  AOI21_X1 U12970 ( .B1(n14513), .B2(n14514), .A(n14511), .ZN(n10484) );
  NAND2_X1 U12971 ( .A1(n10483), .A2(n10482), .ZN(n10481) );
  OAI21_X1 U12972 ( .B1(n14560), .B2(n14559), .A(n10666), .ZN(P2_U2824) );
  NAND2_X1 U12973 ( .A1(n14562), .A2(n16003), .ZN(n10670) );
  NOR2_X1 U12974 ( .A1(n13124), .A2(n13123), .ZN(n13126) );
  AOI21_X1 U12975 ( .B1(n14560), .B2(n14444), .A(n14443), .ZN(n14445) );
  OAI21_X1 U12976 ( .B1(n16515), .B2(n20085), .A(n16514), .ZN(n16516) );
  NOR2_X1 U12977 ( .A1(n16510), .A2(n16513), .ZN(n16514) );
  NAND2_X1 U12978 ( .A1(n16953), .A2(n16939), .ZN(n10102) );
  AOI21_X1 U12979 ( .B1(n16952), .B2(n16935), .A(n16644), .ZN(n10101) );
  AND2_X1 U12980 ( .A1(n12008), .A2(n16735), .ZN(n12027) );
  NAND2_X1 U12981 ( .A1(n10266), .A2(n16939), .ZN(n16764) );
  OAI211_X1 U12982 ( .C1(n16771), .C2(n16911), .A(n10553), .B(n10552), .ZN(
        P2_U2997) );
  AOI21_X1 U12983 ( .B1(n17083), .B2(n16935), .A(n16770), .ZN(n10553) );
  OAI21_X1 U12984 ( .B1(n17110), .B2(n16942), .A(n10105), .ZN(P2_U2999) );
  INV_X1 U12985 ( .A(n10517), .ZN(n10106) );
  AND2_X1 U12986 ( .A1(n17092), .A2(n16939), .ZN(n10107) );
  NAND2_X1 U12987 ( .A1(n17120), .A2(n16939), .ZN(n16802) );
  NAND2_X1 U12988 ( .A1(n16847), .A2(n10061), .ZN(P2_U3004) );
  INV_X1 U12989 ( .A(n10062), .ZN(n10061) );
  OAI21_X1 U12990 ( .B1(n17174), .B2(n16942), .A(n16846), .ZN(n10062) );
  AOI21_X1 U12991 ( .B1(n10669), .B2(n12994), .A(n12993), .ZN(n12998) );
  NAND2_X1 U12992 ( .A1(n12992), .A2(n12991), .ZN(n12993) );
  NAND2_X1 U12993 ( .A1(n10318), .A2(n17262), .ZN(n10317) );
  INV_X1 U12994 ( .A(n16969), .ZN(n10318) );
  OAI211_X1 U12995 ( .C1(n16994), .C2(n17234), .A(n10092), .B(n10091), .ZN(
        P2_U3020) );
  INV_X1 U12996 ( .A(n16992), .ZN(n10091) );
  NAND2_X1 U12997 ( .A1(n16993), .A2(n17221), .ZN(n10092) );
  NAND2_X1 U12998 ( .A1(n10149), .A2(n10164), .ZN(P2_U3030) );
  NAND2_X1 U12999 ( .A1(n17102), .A2(n17103), .ZN(n10164) );
  NAND2_X1 U13000 ( .A1(n10168), .A2(n10166), .ZN(n10165) );
  OAI21_X1 U13001 ( .B1(n17110), .B2(n17266), .A(n10421), .ZN(P2_U3031) );
  AND2_X1 U13002 ( .A1(n17092), .A2(n17262), .ZN(n10127) );
  NOR4_X1 U13003 ( .A1(n10975), .A2(n12970), .A3(n10974), .A4(n10973), .ZN(
        n10976) );
  NAND2_X1 U13004 ( .A1(n10587), .A2(n10583), .ZN(P3_U2642) );
  AND2_X1 U13005 ( .A1(n17754), .A2(n10584), .ZN(n10583) );
  INV_X1 U13006 ( .A(n10977), .ZN(n10588) );
  NOR2_X1 U13007 ( .A1(n12945), .A2(n12944), .ZN(n12946) );
  NAND2_X1 U13008 ( .A1(n9962), .A2(n9956), .ZN(P3_U2817) );
  INV_X1 U13009 ( .A(n18853), .ZN(n9962) );
  NOR3_X1 U13010 ( .A1(n9961), .A2(n9959), .A3(n9957), .ZN(n9956) );
  NOR2_X1 U13011 ( .A1(n12928), .A2(n12927), .ZN(n12929) );
  OR3_X1 U13012 ( .A1(n18670), .A2(n19171), .A3(n18661), .ZN(n17649) );
  AOI21_X1 U13013 ( .B1(n9964), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n9847), .ZN(n19104) );
  NAND2_X1 U13014 ( .A1(n19108), .A2(n19101), .ZN(n9964) );
  OR3_X1 U13015 ( .A1(n19841), .A2(n19840), .A3(n19839), .ZN(n19842) );
  OR2_X1 U13016 ( .A1(n17654), .A2(n17688), .ZN(U212) );
  CLKBUF_X3 U13017 ( .A(n12731), .Z(n17439) );
  INV_X1 U13018 ( .A(n12184), .ZN(n14455) );
  NAND2_X4 U13019 ( .A1(n10748), .A2(n12184), .ZN(n12586) );
  CLKBUF_X3 U13020 ( .A(n12808), .Z(n18334) );
  NOR2_X1 U13021 ( .A1(n19787), .A2(n10868), .ZN(n12743) );
  XOR2_X1 U13022 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n10851), .Z(
        n10855) );
  INV_X1 U13023 ( .A(n12818), .ZN(n12733) );
  AND2_X1 U13024 ( .A1(n12594), .A2(n10600), .ZN(n14851) );
  NAND2_X1 U13025 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10662), .ZN(
        n13014) );
  INV_X1 U13026 ( .A(n10766), .ZN(n14734) );
  NAND2_X1 U13027 ( .A1(n12374), .A2(n12375), .ZN(n13145) );
  INV_X1 U13028 ( .A(n18343), .ZN(n18267) );
  OR2_X1 U13029 ( .A1(n11768), .A2(n11767), .ZN(n9785) );
  INV_X1 U13030 ( .A(n11442), .ZN(n11640) );
  NAND2_X1 U13031 ( .A1(n14447), .A2(n14449), .ZN(n14448) );
  NAND2_X1 U13032 ( .A1(n15798), .A2(n10750), .ZN(n15767) );
  NAND2_X1 U13033 ( .A1(n10757), .A2(n11950), .ZN(n12011) );
  AND2_X1 U13034 ( .A1(n13493), .A2(n9849), .ZN(n14631) );
  AND2_X1 U13035 ( .A1(n13493), .A2(n10775), .ZN(n14659) );
  AND2_X1 U13036 ( .A1(n14762), .A2(n10767), .ZN(n9786) );
  NAND2_X1 U13037 ( .A1(n15798), .A2(n15799), .ZN(n15782) );
  NAND2_X1 U13038 ( .A1(n11783), .A2(n9915), .ZN(n9787) );
  AND3_X2 U13039 ( .A1(n10525), .A2(n9853), .A3(n12453), .ZN(n9788) );
  INV_X1 U13040 ( .A(n10694), .ZN(n10153) );
  NAND2_X1 U13041 ( .A1(n16776), .A2(n11997), .ZN(n9789) );
  OR2_X1 U13042 ( .A1(n18846), .A2(n17935), .ZN(n9790) );
  AND2_X1 U13043 ( .A1(n10658), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9791) );
  INV_X1 U13044 ( .A(n10364), .ZN(n17551) );
  NAND2_X1 U13045 ( .A1(n15226), .A2(n10159), .ZN(n15224) );
  AND2_X1 U13046 ( .A1(n10760), .A2(n15858), .ZN(n9792) );
  AND2_X1 U13047 ( .A1(n16870), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9793) );
  NAND2_X1 U13048 ( .A1(n10182), .A2(n11761), .ZN(n11763) );
  AND3_X1 U13049 ( .A1(n10980), .A2(n11015), .A3(n10983), .ZN(n9794) );
  NAND2_X1 U13050 ( .A1(n14211), .A2(n14212), .ZN(n16020) );
  AND2_X1 U13051 ( .A1(n12841), .A2(n10213), .ZN(n9795) );
  INV_X4 U13052 ( .A(n11163), .ZN(n20854) );
  OR3_X1 U13053 ( .A1(n17535), .A2(n18546), .A3(n18596), .ZN(n9796) );
  AND3_X1 U13054 ( .A1(n10987), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10984), .ZN(n9797) );
  AND2_X1 U13055 ( .A1(n10704), .A2(n16321), .ZN(n9798) );
  AND2_X1 U13056 ( .A1(n12375), .A2(n12424), .ZN(n9799) );
  AND2_X1 U13057 ( .A1(n10197), .A2(n10198), .ZN(n9800) );
  AND2_X1 U13058 ( .A1(n10391), .A2(n10740), .ZN(n9801) );
  AND4_X1 U13059 ( .A1(n10879), .A2(n10878), .A3(n10877), .A4(n10876), .ZN(
        n9803) );
  AND4_X1 U13060 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n9804) );
  NAND2_X1 U13061 ( .A1(n12293), .A2(n10262), .ZN(n10558) );
  AND2_X1 U13062 ( .A1(n16669), .A2(n10090), .ZN(n9805) );
  AND2_X1 U13063 ( .A1(n16804), .A2(n10056), .ZN(n9806) );
  NAND2_X1 U13064 ( .A1(n15183), .A2(n12459), .ZN(n10387) );
  OR2_X1 U13065 ( .A1(n10742), .A2(n15314), .ZN(n9807) );
  OR2_X1 U13066 ( .A1(n17109), .A2(n9914), .ZN(n9808) );
  AND2_X1 U13067 ( .A1(n10600), .A2(n14852), .ZN(n9809) );
  INV_X1 U13068 ( .A(n12234), .ZN(n10400) );
  AND2_X1 U13069 ( .A1(n11289), .A2(n11864), .ZN(n9810) );
  AND2_X1 U13070 ( .A1(n10684), .A2(n10689), .ZN(n9811) );
  NAND2_X1 U13071 ( .A1(n10694), .A2(n10551), .ZN(n9812) );
  NOR3_X1 U13072 ( .A1(n13055), .A2(n10660), .A3(n10661), .ZN(n13064) );
  OAI21_X1 U13073 ( .B1(n10279), .B2(n10280), .A(n16747), .ZN(n15741) );
  NAND2_X1 U13074 ( .A1(n12594), .A2(n12593), .ZN(n14869) );
  NAND2_X1 U13075 ( .A1(n10596), .A2(n12578), .ZN(n14955) );
  NOR2_X1 U13076 ( .A1(n16391), .A2(n16338), .ZN(n9813) );
  MUX2_X1 U13077 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13006), .S(
        n10286), .Z(n20059) );
  INV_X1 U13078 ( .A(n20059), .ZN(n10279) );
  OR2_X1 U13079 ( .A1(n20059), .A2(n16655), .ZN(n9814) );
  AND2_X1 U13080 ( .A1(n9915), .A2(n11791), .ZN(n9815) );
  AND2_X1 U13081 ( .A1(n12019), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9816) );
  AND2_X1 U13082 ( .A1(n13387), .A2(n13406), .ZN(n9817) );
  AND2_X1 U13083 ( .A1(n17464), .A2(n10543), .ZN(n9818) );
  AND2_X1 U13084 ( .A1(n9818), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n9819) );
  AND2_X1 U13085 ( .A1(n11347), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9820) );
  AND2_X1 U13086 ( .A1(n9820), .A2(n16943), .ZN(n9821) );
  AND2_X1 U13087 ( .A1(n9821), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9822) );
  NAND2_X1 U13088 ( .A1(n15128), .A2(n15118), .ZN(n9823) );
  AND4_X1 U13089 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n9824) );
  AND2_X1 U13090 ( .A1(n12007), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9825) );
  AND2_X1 U13091 ( .A1(n10330), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9826) );
  AND2_X1 U13092 ( .A1(n10785), .A2(n10784), .ZN(n9827) );
  AND2_X1 U13093 ( .A1(n9827), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9828) );
  OR2_X2 U13094 ( .A1(n20992), .A2(n14290), .ZN(n21006) );
  INV_X1 U13095 ( .A(n12809), .ZN(n18106) );
  AND2_X2 U13096 ( .A1(n16244), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11189) );
  INV_X1 U13097 ( .A(n12815), .ZN(n10931) );
  AND2_X1 U13098 ( .A1(n18718), .A2(n18751), .ZN(n18752) );
  NAND2_X1 U13099 ( .A1(n15257), .A2(n15478), .ZN(n10032) );
  AND4_X1 U13100 ( .A1(n14447), .A2(n14449), .A3(n13182), .A4(n10169), .ZN(
        n14861) );
  NAND2_X1 U13101 ( .A1(n16026), .A2(n16025), .ZN(n16439) );
  INV_X1 U13102 ( .A(n10398), .ZN(n12438) );
  AND2_X1 U13103 ( .A1(n11637), .A2(n11864), .ZN(n9829) );
  NAND2_X1 U13104 ( .A1(n16855), .A2(n9821), .ZN(n16669) );
  AND2_X1 U13105 ( .A1(n12518), .A2(n12520), .ZN(n9830) );
  NAND2_X1 U13106 ( .A1(n9840), .A2(n10094), .ZN(n11426) );
  NOR2_X1 U13107 ( .A1(n14300), .A2(n10724), .ZN(n14366) );
  INV_X1 U13108 ( .A(n10242), .ZN(n16396) );
  NAND2_X1 U13109 ( .A1(n15182), .A2(n15183), .ZN(n15151) );
  AND2_X1 U13110 ( .A1(n12016), .A2(n10664), .ZN(n13017) );
  NOR2_X1 U13111 ( .A1(n12010), .A2(n10758), .ZN(n15707) );
  NOR2_X1 U13112 ( .A1(n17872), .A2(n18796), .ZN(n10844) );
  AND3_X1 U13113 ( .A1(n10378), .A2(n12183), .A3(n10026), .ZN(n12531) );
  OAI211_X1 U13114 ( .C1(n10191), .C2(n20161), .A(n11075), .B(n20181), .ZN(
        n11394) );
  NAND2_X1 U13115 ( .A1(n13493), .A2(n10774), .ZN(n9831) );
  OR2_X1 U13116 ( .A1(n18249), .A2(n18235), .ZN(n9832) );
  AND2_X1 U13117 ( .A1(n18481), .A2(n10341), .ZN(n9833) );
  AND2_X1 U13118 ( .A1(n13493), .A2(n10171), .ZN(n9834) );
  OR2_X1 U13119 ( .A1(n14187), .A2(n11059), .ZN(n9835) );
  AND2_X1 U13120 ( .A1(n18421), .A2(n10330), .ZN(n9837) );
  AND2_X4 U13121 ( .A1(n12030), .A2(n12036), .ZN(n9838) );
  AND4_X1 U13122 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n12105), .ZN(
        n9839) );
  NOR2_X1 U13123 ( .A1(n13011), .A2(n16920), .ZN(n13012) );
  AND2_X1 U13124 ( .A1(n11063), .A2(n11062), .ZN(n9840) );
  NAND2_X1 U13125 ( .A1(n14762), .A2(n13387), .ZN(n14744) );
  AND2_X1 U13126 ( .A1(n12383), .A2(n12384), .ZN(n9841) );
  INV_X1 U13127 ( .A(n12177), .ZN(n10748) );
  INV_X1 U13128 ( .A(n15224), .ZN(n10158) );
  NAND2_X1 U13129 ( .A1(n10415), .A2(n12369), .ZN(n15573) );
  AND2_X1 U13130 ( .A1(n11264), .A2(n10781), .ZN(n9842) );
  AND2_X1 U13131 ( .A1(n16025), .A2(n10808), .ZN(n9843) );
  AND2_X1 U13132 ( .A1(n14191), .A2(n11437), .ZN(n11442) );
  OR2_X1 U13133 ( .A1(n16963), .A2(n20065), .ZN(n9844) );
  AND2_X1 U13134 ( .A1(n11991), .A2(n10358), .ZN(n10551) );
  AND2_X1 U13135 ( .A1(n21229), .A2(n12409), .ZN(n9845) );
  OR2_X1 U13136 ( .A1(n11851), .A2(n10463), .ZN(n9846) );
  NAND2_X1 U13137 ( .A1(n10636), .A2(n11315), .ZN(n16893) );
  AND2_X1 U13138 ( .A1(n19102), .A2(n19239), .ZN(n9847) );
  AND2_X1 U13139 ( .A1(n15722), .A2(n15710), .ZN(n15691) );
  AND2_X1 U13140 ( .A1(n10750), .A2(n10749), .ZN(n9848) );
  AND2_X1 U13141 ( .A1(n10774), .A2(n14646), .ZN(n9849) );
  INV_X1 U13142 ( .A(n12133), .ZN(n13713) );
  INV_X1 U13143 ( .A(n11479), .ZN(n11637) );
  OR2_X1 U13144 ( .A1(n16700), .A2(n16699), .ZN(n9850) );
  NAND2_X1 U13145 ( .A1(n11776), .A2(n11764), .ZN(n11771) );
  INV_X2 U13146 ( .A(n19987), .ZN(n18596) );
  AND4_X1 U13147 ( .A1(n14862), .A2(n14938), .A3(n14864), .A4(n14865), .ZN(
        n9851) );
  AND4_X1 U13148 ( .A1(n11260), .A2(n11259), .A3(n11258), .A4(n11257), .ZN(
        n9852) );
  OR2_X1 U13149 ( .A1(n11812), .A2(n10644), .ZN(n11800) );
  XNOR2_X1 U13150 ( .A(n12984), .B(n12983), .ZN(n14551) );
  INV_X1 U13151 ( .A(n14551), .ZN(n10669) );
  XNOR2_X1 U13152 ( .A(n12710), .B(n12709), .ZN(n16017) );
  NAND2_X1 U13153 ( .A1(n10278), .A2(n16708), .ZN(n15684) );
  AND2_X1 U13154 ( .A1(n15205), .A2(n15213), .ZN(n9853) );
  INV_X1 U13155 ( .A(n14605), .ZN(n10773) );
  NAND2_X1 U13156 ( .A1(n13063), .A2(n16667), .ZN(n13067) );
  AND2_X1 U13157 ( .A1(n12178), .A2(n12177), .ZN(n12183) );
  AND2_X1 U13158 ( .A1(n10664), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9854) );
  INV_X1 U13159 ( .A(n12208), .ZN(n10039) );
  AND2_X1 U13160 ( .A1(n16855), .A2(n9822), .ZN(n9855) );
  AND2_X1 U13161 ( .A1(n10792), .A2(n16698), .ZN(n9856) );
  AND2_X1 U13162 ( .A1(n10982), .A2(n10981), .ZN(n9857) );
  AND2_X1 U13163 ( .A1(n10986), .A2(n10985), .ZN(n9858) );
  AND2_X1 U13164 ( .A1(n12208), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9859) );
  OR2_X1 U13165 ( .A1(n10962), .A2(n19805), .ZN(n9860) );
  NAND2_X1 U13166 ( .A1(n14762), .A2(n9817), .ZN(n10766) );
  AND2_X1 U13167 ( .A1(n9848), .A2(n15752), .ZN(n9861) );
  NOR2_X1 U13168 ( .A1(n19825), .A2(n19980), .ZN(n9862) );
  AND2_X1 U13169 ( .A1(n11834), .A2(n9972), .ZN(n9863) );
  AND2_X1 U13170 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9864) );
  AND2_X1 U13171 ( .A1(n10310), .A2(n16776), .ZN(n9865) );
  OR2_X1 U13172 ( .A1(n21008), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9866) );
  AND2_X1 U13173 ( .A1(n11329), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n9867) );
  NOR2_X1 U13174 ( .A1(n10953), .A2(n12854), .ZN(n19779) );
  AND2_X1 U13175 ( .A1(n10524), .A2(n10418), .ZN(n9868) );
  AND2_X1 U13176 ( .A1(n16647), .A2(n16645), .ZN(n9869) );
  OR2_X1 U13177 ( .A1(n11213), .A2(n11143), .ZN(n9870) );
  NAND2_X1 U13178 ( .A1(n16855), .A2(n11347), .ZN(n16693) );
  AND2_X1 U13179 ( .A1(n13631), .A2(n13630), .ZN(n9871) );
  OR2_X1 U13180 ( .A1(n12524), .A2(n12526), .ZN(n9872) );
  INV_X1 U13181 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20831) );
  AND2_X1 U13182 ( .A1(n10795), .A2(n12720), .ZN(n9873) );
  AND2_X1 U13183 ( .A1(n10373), .A2(n10400), .ZN(n9874) );
  INV_X1 U13184 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18796) );
  NAND2_X1 U13185 ( .A1(n10370), .A2(n10369), .ZN(n10364) );
  NAND2_X1 U13186 ( .A1(n12008), .A2(n10777), .ZN(n9875) );
  AND2_X1 U13187 ( .A1(n12517), .A2(n12516), .ZN(n9876) );
  OR2_X1 U13188 ( .A1(n16660), .A2(n10319), .ZN(n9877) );
  INV_X1 U13189 ( .A(n10386), .ZN(n12663) );
  OAI21_X1 U13190 ( .B1(n10388), .B2(n12233), .A(n12202), .ZN(n10386) );
  INV_X1 U13191 ( .A(n14691), .ZN(n13492) );
  AND2_X1 U13192 ( .A1(n10016), .A2(n15305), .ZN(n9878) );
  NAND2_X1 U13193 ( .A1(n10525), .A2(n9853), .ZN(n9879) );
  INV_X1 U13194 ( .A(n10740), .ZN(n10739) );
  AND2_X1 U13195 ( .A1(n9901), .A2(n10741), .ZN(n10740) );
  INV_X1 U13196 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18930) );
  NAND2_X1 U13197 ( .A1(n19009), .A2(n18732), .ZN(n18692) );
  AND4_X1 U13198 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n9880) );
  AND4_X1 U13199 ( .A1(n11294), .A2(n11293), .A3(n11292), .A4(n11291), .ZN(
        n9881) );
  OR2_X1 U13200 ( .A1(n14472), .A2(n14471), .ZN(n9882) );
  OR2_X1 U13201 ( .A1(n17108), .A2(n17091), .ZN(n9883) );
  INV_X1 U13202 ( .A(n10172), .ZN(n10171) );
  NAND2_X1 U13203 ( .A1(n9849), .A2(n14630), .ZN(n10172) );
  INV_X1 U13204 ( .A(n10233), .ZN(n10232) );
  NAND2_X1 U13205 ( .A1(n10310), .A2(n10551), .ZN(n10233) );
  AND2_X1 U13206 ( .A1(n10032), .A2(n10403), .ZN(n9884) );
  OR2_X1 U13207 ( .A1(n21008), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9885) );
  AND2_X1 U13208 ( .A1(n10738), .A2(n10419), .ZN(n9886) );
  AND2_X1 U13209 ( .A1(n10196), .A2(n10199), .ZN(n9887) );
  NAND2_X1 U13210 ( .A1(n11764), .A2(n11772), .ZN(n9888) );
  NAND2_X1 U13211 ( .A1(n10288), .A2(n10289), .ZN(n14560) );
  NAND2_X1 U13212 ( .A1(n11073), .A2(n11025), .ZN(n11077) );
  INV_X1 U13213 ( .A(n16895), .ZN(n11988) );
  OR2_X1 U13214 ( .A1(n16674), .A2(n10088), .ZN(n9889) );
  INV_X1 U13215 ( .A(n16733), .ZN(n10693) );
  AND2_X1 U13216 ( .A1(n11024), .A2(n20851), .ZN(n9890) );
  NAND2_X1 U13217 ( .A1(n10696), .A2(n10119), .ZN(n9891) );
  INV_X1 U13218 ( .A(n12518), .ZN(n12521) );
  NAND2_X1 U13219 ( .A1(n15722), .A2(n10733), .ZN(n15677) );
  INV_X1 U13220 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16920) );
  NOR2_X1 U13221 ( .A1(n15243), .A2(n10404), .ZN(n9892) );
  AND3_X1 U13222 ( .A1(n10881), .A2(n10880), .A3(n10883), .ZN(n9893) );
  NAND2_X1 U13223 ( .A1(n10144), .A2(n10742), .ZN(n15105) );
  INV_X1 U13224 ( .A(n15105), .ZN(n10002) );
  AND2_X1 U13225 ( .A1(n16783), .A2(n16782), .ZN(n9894) );
  AND3_X1 U13226 ( .A1(n10338), .A2(n10897), .A3(n10337), .ZN(n9895) );
  INV_X1 U13227 ( .A(n18239), .ZN(n12819) );
  AND2_X1 U13228 ( .A1(n10951), .A2(n10328), .ZN(n9896) );
  AND2_X1 U13229 ( .A1(n11989), .A2(n11987), .ZN(n9897) );
  AND2_X1 U13230 ( .A1(n11989), .A2(n10236), .ZN(n9898) );
  AND2_X1 U13231 ( .A1(n12185), .A2(n12465), .ZN(n9899) );
  NAND2_X1 U13232 ( .A1(n10139), .A2(n10141), .ZN(n10016) );
  INV_X1 U13233 ( .A(n10016), .ZN(n15096) );
  AND2_X1 U13234 ( .A1(n11720), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16910) );
  INV_X1 U13235 ( .A(n16910), .ZN(n10780) );
  AND2_X1 U13236 ( .A1(n10682), .A2(n15962), .ZN(n9900) );
  INV_X1 U13237 ( .A(n12431), .ZN(n10260) );
  AND2_X1 U13238 ( .A1(n10742), .A2(n12462), .ZN(n9901) );
  AND2_X1 U13239 ( .A1(n10752), .A2(n10751), .ZN(n9902) );
  AND2_X1 U13240 ( .A1(n11996), .A2(n11992), .ZN(n9903) );
  AND2_X1 U13241 ( .A1(n12298), .A2(n10382), .ZN(n9904) );
  AND2_X1 U13242 ( .A1(n10026), .A2(n21106), .ZN(n9905) );
  AND2_X1 U13243 ( .A1(n11880), .A2(n10180), .ZN(n9906) );
  AND2_X1 U13244 ( .A1(n12198), .A2(n12185), .ZN(n9907) );
  AND2_X1 U13245 ( .A1(n10372), .A2(n10376), .ZN(n9908) );
  AND2_X1 U13246 ( .A1(n10443), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9909) );
  INV_X1 U13247 ( .A(n11341), .ZN(n9991) );
  OR3_X1 U13248 ( .A1(n11340), .A2(n11894), .A3(n17191), .ZN(n11341) );
  INV_X1 U13249 ( .A(n10387), .ZN(n10480) );
  INV_X1 U13250 ( .A(n10688), .ZN(n10687) );
  NAND2_X1 U13251 ( .A1(n10693), .A2(n16729), .ZN(n10688) );
  AND2_X1 U13252 ( .A1(n11994), .A2(n11992), .ZN(n9910) );
  NAND2_X1 U13253 ( .A1(n10420), .A2(n15257), .ZN(n9911) );
  INV_X1 U13254 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10622) );
  NAND2_X1 U13255 ( .A1(n18017), .A2(n10825), .ZN(n17851) );
  INV_X1 U13256 ( .A(n20065), .ZN(n20040) );
  AND2_X1 U13257 ( .A1(n13038), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13037) );
  INV_X1 U13258 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10659) );
  INV_X1 U13259 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U13260 ( .A1(n11731), .A2(n11747), .ZN(n11759) );
  NAND2_X1 U13261 ( .A1(n16026), .A2(n9843), .ZN(n16433) );
  AND2_X1 U13262 ( .A1(n13064), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13114) );
  NOR2_X1 U13263 ( .A1(n14300), .A2(n14358), .ZN(n14357) );
  NAND2_X1 U13264 ( .A1(n15857), .A2(n9792), .ZN(n15822) );
  OR2_X1 U13265 ( .A1(n11983), .A2(n20840), .ZN(n17234) );
  INV_X1 U13266 ( .A(n17234), .ZN(n17262) );
  NAND2_X1 U13267 ( .A1(n15902), .A2(n15903), .ZN(n14352) );
  INV_X1 U13268 ( .A(n11813), .ZN(n10645) );
  AOI22_X1 U13269 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n19799), .B2(n19961), .ZN(
        n12871) );
  INV_X1 U13270 ( .A(n12871), .ZN(n10542) );
  INV_X1 U13271 ( .A(n10556), .ZN(n10376) );
  NOR2_X1 U13272 ( .A1(n12376), .A2(n12305), .ZN(n10556) );
  AND2_X1 U13273 ( .A1(n10652), .A2(n11853), .ZN(n9912) );
  NOR2_X1 U13274 ( .A1(n12020), .A2(n15739), .ZN(n12711) );
  AND2_X1 U13275 ( .A1(n15902), .A2(n9902), .ZN(n15857) );
  OR2_X1 U13276 ( .A1(n16279), .A2(n10702), .ZN(n9913) );
  AND2_X1 U13277 ( .A1(n15798), .A2(n9848), .ZN(n15751) );
  NAND2_X1 U13278 ( .A1(n14879), .A2(n14880), .ZN(n14878) );
  NAND2_X1 U13279 ( .A1(n15842), .A2(n15843), .ZN(n15829) );
  NAND2_X1 U13280 ( .A1(n10754), .A2(n11906), .ZN(n14341) );
  NAND2_X1 U13281 ( .A1(n10714), .A2(n10717), .ZN(n14275) );
  NOR2_X1 U13282 ( .A1(n12010), .A2(n10755), .ZN(n15694) );
  NOR2_X1 U13283 ( .A1(n14340), .A2(n15919), .ZN(n15902) );
  AND2_X1 U13284 ( .A1(n15857), .A2(n15858), .ZN(n15842) );
  AND2_X1 U13285 ( .A1(n12711), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13045) );
  AND2_X1 U13286 ( .A1(n12016), .A2(n9854), .ZN(n13020) );
  AND2_X1 U13287 ( .A1(n12594), .A2(n9809), .ZN(n14838) );
  NAND2_X1 U13288 ( .A1(n12303), .A2(n12302), .ZN(n21201) );
  INV_X1 U13289 ( .A(n21201), .ZN(n10611) );
  NAND2_X1 U13290 ( .A1(n15902), .A2(n10752), .ZN(n14351) );
  AND2_X1 U13291 ( .A1(n20042), .A2(n17260), .ZN(n9914) );
  INV_X1 U13292 ( .A(n10279), .ZN(n10275) );
  AND2_X1 U13293 ( .A1(n12018), .A2(n10657), .ZN(n13031) );
  INV_X1 U13294 ( .A(n10510), .ZN(n11677) );
  AND2_X1 U13295 ( .A1(n11782), .A2(n10641), .ZN(n9915) );
  NAND2_X1 U13296 ( .A1(n14281), .A2(n13162), .ZN(n14447) );
  AND2_X1 U13297 ( .A1(n10609), .A2(n10608), .ZN(n9916) );
  OR3_X1 U13298 ( .A1(n13055), .A2(n10661), .A3(n13061), .ZN(n9917) );
  AND2_X1 U13299 ( .A1(n12463), .A2(n15305), .ZN(n9918) );
  INV_X1 U13300 ( .A(n16019), .ZN(n10244) );
  OR2_X1 U13301 ( .A1(n17280), .A2(n10064), .ZN(n9919) );
  NOR2_X1 U13302 ( .A1(n17262), .A2(n17080), .ZN(n9920) );
  INV_X1 U13303 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13042) );
  NAND2_X1 U13304 ( .A1(n9815), .A2(n10640), .ZN(n9921) );
  INV_X1 U13305 ( .A(n10280), .ZN(n15758) );
  NOR2_X1 U13306 ( .A1(n15777), .A2(n16759), .ZN(n10280) );
  INV_X1 U13307 ( .A(n10274), .ZN(n15804) );
  OR2_X1 U13308 ( .A1(n20043), .A2(n20037), .ZN(n10274) );
  OR2_X1 U13309 ( .A1(n16321), .A2(n16407), .ZN(n9922) );
  INV_X1 U13310 ( .A(n16816), .ZN(n10358) );
  OR2_X1 U13311 ( .A1(n16816), .A2(n10354), .ZN(n9923) );
  INV_X1 U13312 ( .A(n16815), .ZN(n10356) );
  OR2_X1 U13313 ( .A1(n19206), .A2(n19100), .ZN(n9924) );
  AND2_X1 U13314 ( .A1(n16298), .A2(n16319), .ZN(n9925) );
  NOR2_X1 U13315 ( .A1(n14956), .A2(n10597), .ZN(n9926) );
  NAND2_X1 U13316 ( .A1(n10514), .A2(n10511), .ZN(n10510) );
  AND2_X1 U13317 ( .A1(n11211), .A2(n11469), .ZN(n9927) );
  AND2_X1 U13318 ( .A1(n11211), .A2(n11237), .ZN(n9928) );
  OR2_X1 U13319 ( .A1(n17082), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9929) );
  AND2_X1 U13320 ( .A1(n9912), .A2(n10183), .ZN(n9930) );
  AND2_X1 U13321 ( .A1(n10733), .A2(n10732), .ZN(n9931) );
  AND2_X1 U13322 ( .A1(n10767), .A2(n14716), .ZN(n9932) );
  AND2_X1 U13323 ( .A1(n9816), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9933) );
  AND2_X1 U13324 ( .A1(n10565), .A2(n17851), .ZN(n9934) );
  INV_X1 U13325 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16800) );
  AND2_X1 U13326 ( .A1(n16848), .A2(n16824), .ZN(n9935) );
  INV_X1 U13327 ( .A(n10293), .ZN(n10292) );
  NAND2_X1 U13328 ( .A1(n9814), .A2(n10275), .ZN(n10293) );
  NAND2_X1 U13329 ( .A1(n13142), .A2(n14487), .ZN(n12544) );
  AND2_X1 U13330 ( .A1(n18364), .A2(n9818), .ZN(n9936) );
  NAND2_X1 U13331 ( .A1(n9852), .A2(n9804), .ZN(n11469) );
  INV_X1 U13332 ( .A(n11469), .ZN(n10794) );
  NAND2_X1 U13333 ( .A1(n12565), .A2(n12564), .ZN(n14284) );
  INV_X1 U13334 ( .A(n19120), .ZN(n10213) );
  NOR2_X1 U13335 ( .A1(n18725), .A2(n18694), .ZN(n18691) );
  OR2_X1 U13336 ( .A1(n19984), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n9937) );
  INV_X1 U13337 ( .A(n16183), .ZN(n16372) );
  AND2_X1 U13338 ( .A1(n11481), .A2(n11480), .ZN(n9938) );
  INV_X1 U13339 ( .A(n9755), .ZN(n18920) );
  OR2_X1 U13340 ( .A1(n13055), .A2(n10661), .ZN(n9939) );
  INV_X1 U13341 ( .A(n10630), .ZN(n10629) );
  NOR2_X1 U13342 ( .A1(n18741), .A2(n10632), .ZN(n10630) );
  INV_X1 U13343 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n19233) );
  INV_X1 U13344 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n9996) );
  AND2_X1 U13345 ( .A1(n11894), .A2(n11987), .ZN(n9940) );
  OR2_X1 U13346 ( .A1(n15236), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9941) );
  AND2_X1 U13347 ( .A1(n10398), .A2(n21739), .ZN(n9942) );
  AND2_X1 U13348 ( .A1(n10650), .A2(n11875), .ZN(n9943) );
  AND2_X1 U13349 ( .A1(n9819), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U13350 ( .A1(n10580), .A2(n10581), .ZN(n17942) );
  INV_X1 U13351 ( .A(n20062), .ZN(n15999) );
  AND3_X1 U13352 ( .A1(n12958), .A2(n12957), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n9945) );
  AND2_X1 U13353 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18028) );
  INV_X1 U13354 ( .A(n20800), .ZN(n20808) );
  NOR2_X2 U13355 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20800) );
  INV_X1 U13356 ( .A(n16747), .ZN(n10655) );
  NAND2_X1 U13357 ( .A1(n15973), .A2(n15976), .ZN(n15966) );
  INV_X1 U13358 ( .A(n15966), .ZN(n10281) );
  AND2_X2 U13359 ( .A1(n10978), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17324) );
  AND2_X1 U13360 ( .A1(n9822), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9946) );
  NAND2_X1 U13361 ( .A1(n18440), .A2(n10818), .ZN(n9947) );
  OR2_X1 U13362 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9948) );
  INV_X1 U13363 ( .A(n10783), .ZN(n10270) );
  NAND2_X1 U13364 ( .A1(n10785), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10783) );
  INV_X1 U13365 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n9998) );
  INV_X1 U13366 ( .A(n10206), .ZN(n10059) );
  NAND2_X1 U13367 ( .A1(n12957), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10206) );
  OR2_X1 U13368 ( .A1(n17872), .A2(n10564), .ZN(n9949) );
  AND2_X1 U13369 ( .A1(n10339), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n9950) );
  AND2_X1 U13370 ( .A1(n22032), .A2(n21858), .ZN(n9951) );
  OR2_X1 U13371 ( .A1(n9990), .A2(n10783), .ZN(n9952) );
  INV_X1 U13372 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18594) );
  INV_X1 U13373 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10331) );
  INV_X1 U13374 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18060) );
  NOR2_X1 U13375 ( .A1(n17950), .A2(n17943), .ZN(n18834) );
  AND2_X1 U13376 ( .A1(n18655), .A2(n17631), .ZN(n9953) );
  INV_X1 U13377 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10406) );
  NAND2_X1 U13378 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n9954) );
  AND2_X1 U13379 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n9955) );
  INV_X1 U13380 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20814) );
  AOI21_X1 U13381 ( .B1(n17483), .B2(n17477), .A(n10800), .ZN(n17536) );
  OR2_X1 U13382 ( .A1(n19801), .A2(n19802), .ZN(n10434) );
  NOR4_X2 U13383 ( .A1(n19317), .A2(n20004), .A3(n18067), .A4(n19833), .ZN(
        n18073) );
  AOI22_X2 U13384 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20175), .ZN(n20665) );
  NOR2_X2 U13385 ( .A1(n17305), .A2(n17306), .ZN(n20175) );
  NAND2_X2 U13386 ( .A1(n17733), .A2(n20003), .ZN(n18545) );
  NOR2_X4 U13387 ( .A1(n19270), .A2(n18596), .ZN(n19811) );
  NAND3_X1 U13388 ( .A1(n19098), .A2(n19099), .A3(n9924), .ZN(n9965) );
  INV_X1 U13389 ( .A(n9969), .ZN(n12891) );
  XNOR2_X1 U13390 ( .A(n9969), .B(n10622), .ZN(n19001) );
  XNOR2_X1 U13391 ( .A(n18532), .B(n9969), .ZN(n12827) );
  OR2_X2 U13392 ( .A1(n12774), .A2(n12773), .ZN(n9969) );
  NAND4_X1 U13393 ( .A1(n9881), .A2(n11296), .A3(n11295), .A4(n9971), .ZN(
        n9970) );
  INV_X1 U13394 ( .A(n9973), .ZN(n11094) );
  OAI211_X1 U13395 ( .C1(n17095), .C2(n17094), .A(n17093), .B(n9974), .ZN(
        P2_U3029) );
  NAND3_X1 U13396 ( .A1(n17102), .A2(n17094), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9974) );
  OAI21_X2 U13397 ( .B1(n17092), .B2(n17234), .A(n9883), .ZN(n17102) );
  INV_X1 U13398 ( .A(n16865), .ZN(n9975) );
  AND2_X2 U13399 ( .A1(n16695), .A2(n16722), .ZN(n16709) );
  INV_X2 U13400 ( .A(n11686), .ZN(n20851) );
  OR2_X1 U13401 ( .A1(n10516), .A2(n9952), .ZN(n9986) );
  NAND3_X1 U13402 ( .A1(n9793), .A2(n16868), .A3(n9945), .ZN(n9988) );
  INV_X1 U13403 ( .A(n10184), .ZN(n9992) );
  NAND2_X2 U13404 ( .A1(n10549), .A2(n11289), .ZN(n10184) );
  NAND2_X1 U13405 ( .A1(n12049), .A2(n9994), .ZN(n12052) );
  OAI22_X1 U13406 ( .A1(n13636), .A2(n9999), .B1(n13711), .B2(n9998), .ZN(
        n9997) );
  INV_X1 U13407 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n9999) );
  NAND2_X2 U13408 ( .A1(n10744), .A2(n15521), .ZN(n13711) );
  XNOR2_X2 U13409 ( .A(n12237), .B(n12236), .ZN(n13156) );
  OR2_X1 U13410 ( .A1(n10002), .A2(n10654), .ZN(n10001) );
  NAND3_X1 U13411 ( .A1(n9788), .A2(n15191), .A3(n10480), .ZN(n10007) );
  NAND2_X2 U13412 ( .A1(n15253), .A2(n12451), .ZN(n15191) );
  NAND2_X1 U13413 ( .A1(n14333), .A2(n14332), .ZN(n14335) );
  OAI21_X1 U13414 ( .B1(n12543), .B2(n9899), .A(n12544), .ZN(n10010) );
  NAND2_X1 U13415 ( .A1(n12537), .A2(n10009), .ZN(n12189) );
  INV_X1 U13416 ( .A(n10010), .ZN(n10009) );
  NAND2_X2 U13417 ( .A1(n12672), .A2(n12188), .ZN(n12537) );
  INV_X1 U13418 ( .A(n12178), .ZN(n10013) );
  INV_X2 U13419 ( .A(n10033), .ZN(n10176) );
  NAND2_X1 U13420 ( .A1(n10374), .A2(n10377), .ZN(n10024) );
  NAND3_X2 U13421 ( .A1(n10019), .A2(n10020), .A3(n10160), .ZN(n10747) );
  NAND3_X1 U13422 ( .A1(n9908), .A2(n12234), .A3(n10024), .ZN(n10019) );
  INV_X2 U13423 ( .A(n12182), .ZN(n10026) );
  OR2_X2 U13424 ( .A1(n12047), .A2(n12048), .ZN(n12182) );
  NAND2_X1 U13425 ( .A1(n12292), .A2(n12291), .ZN(n10027) );
  NAND3_X1 U13426 ( .A1(n12293), .A2(n10027), .A3(n21645), .ZN(n10413) );
  NAND2_X1 U13427 ( .A1(n10027), .A2(n12293), .ZN(n21384) );
  NOR2_X4 U13428 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10744) );
  NAND4_X1 U13429 ( .A1(n12180), .A2(n10816), .A3(n12205), .A4(n10029), .ZN(
        n12680) );
  NAND4_X1 U13430 ( .A1(n9907), .A2(n12126), .A3(n12125), .A4(n15538), .ZN(
        n10030) );
  AND2_X1 U13431 ( .A1(n15237), .A2(n10032), .ZN(n10031) );
  OAI211_X2 U13432 ( .C1(n12213), .C2(n10038), .A(n10037), .B(n10034), .ZN(
        n21172) );
  NAND2_X1 U13433 ( .A1(n10040), .A2(n11314), .ZN(n10401) );
  NAND2_X1 U13434 ( .A1(n10124), .A2(n10040), .ZN(n10123) );
  OAI21_X1 U13435 ( .B1(n16910), .B2(n10040), .A(n16909), .ZN(n17235) );
  NAND2_X1 U13436 ( .A1(n10042), .A2(n10041), .ZN(n10046) );
  NAND3_X1 U13437 ( .A1(n10067), .A2(n10066), .A3(n10065), .ZN(n10042) );
  NAND2_X1 U13438 ( .A1(n10043), .A2(n11079), .ZN(n11690) );
  NAND2_X1 U13439 ( .A1(n10045), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11086) );
  NAND2_X1 U13440 ( .A1(n10046), .A2(n11690), .ZN(n10045) );
  NAND2_X4 U13441 ( .A1(n10109), .A2(n11342), .ZN(n16855) );
  NAND2_X1 U13442 ( .A1(n10047), .A2(n11695), .ZN(n14188) );
  MUX2_X1 U13443 ( .A(n11683), .B(n13974), .S(n11695), .Z(n11685) );
  NAND2_X2 U13444 ( .A1(n16855), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16856) );
  AND2_X1 U13445 ( .A1(n10049), .A2(n16856), .ZN(n17175) );
  NAND3_X1 U13446 ( .A1(n10050), .A2(n11900), .A3(n11899), .ZN(n14317) );
  NAND3_X1 U13447 ( .A1(n10051), .A2(n11955), .A3(n11954), .ZN(n15708) );
  NAND3_X1 U13448 ( .A1(n10052), .A2(n11973), .A3(n11972), .ZN(n13000) );
  NAND3_X1 U13449 ( .A1(n10053), .A2(n11979), .A3(n11978), .ZN(n12704) );
  NAND3_X1 U13450 ( .A1(n10055), .A2(n11925), .A3(n11924), .ZN(n15843) );
  NAND3_X1 U13451 ( .A1(n11024), .A2(n11058), .A3(n11358), .ZN(n10515) );
  NAND2_X2 U13452 ( .A1(n9887), .A2(n9800), .ZN(n11358) );
  NAND2_X1 U13453 ( .A1(n10206), .A2(n10058), .ZN(n10056) );
  NAND2_X1 U13454 ( .A1(n17135), .A2(n10057), .ZN(P2_U3033) );
  INV_X1 U13455 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10058) );
  INV_X1 U13456 ( .A(n11695), .ZN(n10064) );
  INV_X1 U13457 ( .A(n16856), .ZN(n10079) );
  INV_X1 U13458 ( .A(n11720), .ZN(n10080) );
  XNOR2_X2 U13459 ( .A(n11290), .B(n11289), .ZN(n11720) );
  NAND2_X2 U13460 ( .A1(n16938), .A2(n11247), .ZN(n11263) );
  INV_X1 U13461 ( .A(n11079), .ZN(n10095) );
  NAND2_X1 U13462 ( .A1(n10695), .A2(n10097), .ZN(n16873) );
  OAI21_X1 U13463 ( .B1(n11758), .B2(n10238), .A(n10237), .ZN(n10097) );
  NAND2_X1 U13464 ( .A1(n10098), .A2(n10471), .ZN(n10470) );
  NAND2_X1 U13465 ( .A1(n15694), .A2(n15695), .ZN(n15674) );
  NAND3_X1 U13466 ( .A1(n10102), .A2(n10101), .A3(n10100), .ZN(P2_U2985) );
  OR2_X1 U13467 ( .A1(n16956), .A2(n16942), .ZN(n10100) );
  NOR2_X2 U13468 ( .A1(n16646), .A2(n9869), .ZN(n16953) );
  NAND3_X1 U13469 ( .A1(n11720), .A2(n10194), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11315) );
  AND2_X2 U13470 ( .A1(n10108), .A2(n11147), .ZN(n20331) );
  AND2_X2 U13471 ( .A1(n10108), .A2(n11155), .ZN(n20299) );
  NAND2_X1 U13472 ( .A1(n11152), .A2(n10108), .ZN(n20363) );
  AND2_X2 U13473 ( .A1(n14199), .A2(n15986), .ZN(n10108) );
  NAND3_X1 U13474 ( .A1(n10272), .A2(n10271), .A3(n9828), .ZN(n10110) );
  NAND3_X1 U13475 ( .A1(n10272), .A2(n10271), .A3(n9827), .ZN(n16756) );
  NAND2_X1 U13476 ( .A1(n11758), .A2(n11894), .ZN(n10146) );
  OAI211_X1 U13477 ( .C1(n11758), .C2(n10115), .A(n10112), .B(n10111), .ZN(
        n16894) );
  NAND2_X1 U13478 ( .A1(n11758), .A2(n9940), .ZN(n10111) );
  XNOR2_X2 U13479 ( .A(n10184), .B(n11317), .ZN(n11758) );
  NAND2_X1 U13480 ( .A1(n10123), .A2(n10315), .ZN(n10122) );
  NAND3_X1 U13481 ( .A1(n18919), .A2(n9795), .A3(n18714), .ZN(n12846) );
  NAND2_X2 U13482 ( .A1(n10129), .A2(n10624), .ZN(n18919) );
  INV_X1 U13483 ( .A(n10449), .ZN(n10137) );
  NAND2_X1 U13484 ( .A1(n10449), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10138) );
  NAND3_X1 U13485 ( .A1(n10143), .A2(n9735), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10139) );
  NAND3_X1 U13486 ( .A1(n10143), .A2(n9735), .A3(n12461), .ZN(n15114) );
  NAND3_X1 U13487 ( .A1(n10143), .A2(n9735), .A3(n10140), .ZN(n10144) );
  INV_X1 U13488 ( .A(n15338), .ZN(n10142) );
  NAND3_X1 U13489 ( .A1(n10148), .A2(n9812), .A3(n9910), .ZN(n10147) );
  NAND2_X1 U13490 ( .A1(n10150), .A2(n11264), .ZN(n16907) );
  NAND2_X1 U13491 ( .A1(n16804), .A2(n17115), .ZN(n10151) );
  NAND3_X1 U13492 ( .A1(n10154), .A2(n16824), .A3(n10152), .ZN(n16851) );
  NAND3_X1 U13493 ( .A1(n10154), .A2(n9935), .A3(n10152), .ZN(n16854) );
  NAND3_X1 U13494 ( .A1(n12544), .A2(n12543), .A3(n21060), .ZN(n10155) );
  NAND2_X1 U13495 ( .A1(n15257), .A2(n12367), .ZN(n10157) );
  NAND2_X1 U13496 ( .A1(n15257), .A2(n15463), .ZN(n10159) );
  INV_X4 U13497 ( .A(n10812), .ZN(n15257) );
  NAND3_X1 U13498 ( .A1(n10558), .A2(n10377), .A3(n10371), .ZN(n10160) );
  OAI21_X1 U13499 ( .B1(n12458), .B2(n10387), .A(n15257), .ZN(n10162) );
  INV_X1 U13500 ( .A(n11758), .ZN(n11314) );
  OAI21_X1 U13501 ( .B1(n10781), .B2(n16910), .A(n11758), .ZN(n10163) );
  NAND3_X1 U13502 ( .A1(n16778), .A2(n17097), .A3(n17221), .ZN(n10168) );
  NAND3_X1 U13503 ( .A1(n14447), .A2(n14449), .A3(n13182), .ZN(n14953) );
  INV_X1 U13504 ( .A(n9871), .ZN(n10173) );
  INV_X1 U13505 ( .A(n14581), .ZN(n10174) );
  OR2_X1 U13506 ( .A1(n14596), .A2(n14595), .ZN(n10175) );
  NOR2_X2 U13507 ( .A1(n11763), .A2(n9785), .ZN(n11776) );
  NAND2_X1 U13508 ( .A1(n11852), .A2(n9930), .ZN(n11877) );
  NOR2_X2 U13509 ( .A1(n14199), .A2(n14171), .ZN(n11154) );
  INV_X1 U13510 ( .A(n10188), .ZN(n16641) );
  NAND3_X1 U13511 ( .A1(n10323), .A2(n9906), .A3(n10305), .ZN(n10189) );
  NAND2_X1 U13512 ( .A1(n10189), .A2(n10795), .ZN(n12718) );
  NAND2_X1 U13513 ( .A1(n10992), .A2(n11015), .ZN(n10197) );
  NAND2_X2 U13514 ( .A1(n10197), .A2(n10196), .ZN(n11434) );
  NAND3_X1 U13515 ( .A1(n10195), .A2(n10997), .A3(n10996), .ZN(n10196) );
  INV_X2 U13516 ( .A(n11434), .ZN(n20146) );
  NAND2_X1 U13517 ( .A1(n11084), .A2(n20146), .ZN(n11068) );
  NOR2_X2 U13518 ( .A1(n11686), .A2(n10286), .ZN(n11084) );
  NAND3_X1 U13519 ( .A1(n10549), .A2(n11317), .A3(n9810), .ZN(n11337) );
  AND2_X4 U13520 ( .A1(n11171), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16378) );
  INV_X1 U13521 ( .A(n10508), .ZN(n10201) );
  NAND2_X1 U13522 ( .A1(n10204), .A2(n9870), .ZN(n11144) );
  NAND2_X1 U13523 ( .A1(n20424), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10204) );
  OAI21_X1 U13524 ( .B1(n20424), .B2(n20800), .A(n20814), .ZN(n10205) );
  AND2_X2 U13525 ( .A1(n11024), .A2(n11080), .ZN(n11417) );
  AND4_X2 U13526 ( .A1(n9748), .A2(n11078), .A3(n20181), .A4(n20156), .ZN(
        n11080) );
  NAND2_X2 U13527 ( .A1(n11038), .A2(n11037), .ZN(n20161) );
  NAND3_X1 U13528 ( .A1(n17137), .A2(n16939), .A3(n17138), .ZN(n16822) );
  NOR2_X1 U13529 ( .A1(n19001), .A2(n19008), .ZN(n19000) );
  NOR2_X2 U13530 ( .A1(n18970), .A2(n18969), .ZN(n18968) );
  NAND3_X1 U13531 ( .A1(n10210), .A2(n9909), .A3(n10441), .ZN(n10211) );
  AND2_X1 U13532 ( .A1(n10210), .A2(n10443), .ZN(n10212) );
  AOI21_X2 U13533 ( .B1(n18806), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12844), .ZN(n18799) );
  NAND2_X1 U13534 ( .A1(n16266), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10215) );
  NAND2_X1 U13535 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10217) );
  NAND2_X1 U13536 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10222) );
  NAND2_X1 U13537 ( .A1(n16282), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10223) );
  INV_X1 U13538 ( .A(n10231), .ZN(n10230) );
  NAND2_X1 U13539 ( .A1(n11758), .A2(n10237), .ZN(n10235) );
  NAND2_X1 U13540 ( .A1(n10235), .A2(n9898), .ZN(n10694) );
  NAND2_X1 U13541 ( .A1(n10239), .A2(n14010), .ZN(n20824) );
  AND2_X2 U13542 ( .A1(n10241), .A2(n10240), .ZN(n16401) );
  OAI21_X2 U13543 ( .B1(n16408), .B2(n9922), .A(n10703), .ZN(n10242) );
  AND2_X2 U13544 ( .A1(n14210), .A2(n14308), .ZN(n14212) );
  NAND2_X2 U13545 ( .A1(n14198), .A2(n14197), .ZN(n14211) );
  NAND3_X1 U13546 ( .A1(n16519), .A2(n16497), .A3(n16520), .ZN(n16393) );
  NAND2_X1 U13547 ( .A1(n10453), .A2(n9813), .ZN(n16520) );
  NAND2_X1 U13548 ( .A1(n10453), .A2(n16397), .ZN(n10246) );
  NAND3_X1 U13549 ( .A1(n16422), .A2(n16279), .A3(n16237), .ZN(n10247) );
  NAND2_X2 U13550 ( .A1(n16424), .A2(n16423), .ZN(n16422) );
  XNOR2_X2 U13551 ( .A(n16236), .B(n10820), .ZN(n16424) );
  NAND2_X1 U13552 ( .A1(n11134), .A2(n10776), .ZN(n11126) );
  NAND3_X1 U13553 ( .A1(n10252), .A2(n10251), .A3(n10250), .ZN(n14519) );
  NAND3_X1 U13554 ( .A1(n10253), .A2(n14502), .A3(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10252) );
  NAND2_X1 U13555 ( .A1(n14501), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10253) );
  AND2_X1 U13556 ( .A1(n14503), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10254) );
  NAND2_X1 U13557 ( .A1(n10258), .A2(n10256), .ZN(n15253) );
  INV_X1 U13558 ( .A(n10257), .ZN(n10256) );
  NAND3_X1 U13559 ( .A1(n10363), .A2(n10362), .A3(n12431), .ZN(n10258) );
  NAND2_X2 U13560 ( .A1(n21172), .A2(n12290), .ZN(n12293) );
  AND2_X4 U13561 ( .A1(n10264), .A2(n12366), .ZN(n10812) );
  XNOR2_X1 U13562 ( .A(n10264), .B(n12432), .ZN(n13249) );
  AND2_X1 U13563 ( .A1(n10264), .A2(n12424), .ZN(n10263) );
  NAND2_X1 U13564 ( .A1(n10266), .A2(n17262), .ZN(n17078) );
  NOR2_X1 U13565 ( .A1(n16757), .A2(n16758), .ZN(n10266) );
  XNOR2_X2 U13566 ( .A(n11263), .B(n11262), .ZN(n16919) );
  NAND2_X1 U13567 ( .A1(n11212), .A2(n11211), .ZN(n10268) );
  NAND3_X1 U13568 ( .A1(n10550), .A2(n11212), .A3(n9928), .ZN(n11261) );
  NAND3_X1 U13569 ( .A1(n11261), .A2(n16936), .A3(n10782), .ZN(n16938) );
  NAND2_X1 U13570 ( .A1(n10278), .A2(n10276), .ZN(n15665) );
  INV_X2 U13571 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n10286) );
  NAND3_X1 U13572 ( .A1(n11995), .A2(n9903), .A3(n11994), .ZN(n10304) );
  MUX2_X1 U13573 ( .A(n11805), .B(n9742), .S(n11804), .Z(n11806) );
  INV_X1 U13574 ( .A(n11180), .ZN(n16183) );
  AND2_X4 U13575 ( .A1(n11170), .A2(n17335), .ZN(n11180) );
  OAI21_X1 U13576 ( .B1(n11513), .B2(n20363), .A(n10309), .ZN(n11158) );
  AND2_X2 U13577 ( .A1(n11153), .A2(n11152), .ZN(n20487) );
  AND2_X2 U13578 ( .A1(n11125), .A2(n17320), .ZN(n11153) );
  OAI21_X1 U13579 ( .B1(n17087), .B2(n17266), .A(n10312), .ZN(n17090) );
  NAND2_X1 U13580 ( .A1(n16968), .A2(n10317), .ZN(P2_U3018) );
  NAND2_X1 U13581 ( .A1(n11868), .A2(n11869), .ZN(n10320) );
  NOR2_X1 U13582 ( .A1(n16661), .A2(n9877), .ZN(n16650) );
  NOR2_X1 U13583 ( .A1(n12780), .A2(n12779), .ZN(n12786) );
  OR2_X2 U13584 ( .A1(n16416), .A2(n16281), .ZN(n10813) );
  NAND2_X1 U13585 ( .A1(n18799), .A2(n19127), .ZN(n18798) );
  INV_X1 U13586 ( .A(n10801), .ZN(n10704) );
  NOR2_X1 U13587 ( .A1(n18989), .A2(n18988), .ZN(n18987) );
  NAND2_X1 U13588 ( .A1(n20454), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11220) );
  NAND3_X1 U13589 ( .A1(n9824), .A2(P3_EAX_REG_0__SCAN_IN), .A3(n10325), .ZN(
        n10324) );
  NAND2_X1 U13590 ( .A1(n19355), .A2(n10945), .ZN(n12855) );
  NAND2_X1 U13591 ( .A1(n12855), .A2(n10948), .ZN(n10327) );
  NAND3_X1 U13592 ( .A1(n9896), .A2(n10950), .A3(n10327), .ZN(n12865) );
  AND2_X1 U13593 ( .A1(n10952), .A2(n10953), .ZN(n10329) );
  NAND2_X1 U13594 ( .A1(n18421), .A2(n9826), .ZN(n18409) );
  NAND3_X1 U13595 ( .A1(n9895), .A2(n10899), .A3(n10332), .ZN(n12854) );
  NAND3_X1 U13596 ( .A1(n10895), .A2(n10335), .A3(n10896), .ZN(n10334) );
  AND2_X2 U13597 ( .A1(n10345), .A2(n10343), .ZN(n11124) );
  NAND2_X1 U13598 ( .A1(n10508), .A2(n10344), .ZN(n10343) );
  NAND3_X1 U13599 ( .A1(n10508), .A2(n11128), .A3(n11127), .ZN(n10345) );
  NAND2_X1 U13600 ( .A1(n11094), .A2(n11093), .ZN(n10508) );
  NAND2_X2 U13601 ( .A1(n10677), .A2(n10675), .ZN(n16895) );
  INV_X2 U13602 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19961) );
  NAND3_X1 U13603 ( .A1(n9803), .A2(n10882), .A3(n9893), .ZN(n10946) );
  NOR2_X2 U13604 ( .A1(n19012), .A2(n17635), .ZN(n18922) );
  NAND2_X2 U13605 ( .A1(n12889), .A2(n12888), .ZN(n19326) );
  NAND4_X1 U13606 ( .A1(n12417), .A2(n10370), .A3(n10369), .A4(n12418), .ZN(
        n10362) );
  INV_X1 U13607 ( .A(n10365), .ZN(n10363) );
  AND2_X1 U13608 ( .A1(n10558), .A2(n21645), .ZN(n10374) );
  NAND2_X1 U13609 ( .A1(n10558), .A2(n10557), .ZN(n10372) );
  NAND2_X2 U13610 ( .A1(n10176), .A2(n10375), .ZN(n12369) );
  INV_X1 U13611 ( .A(n12490), .ZN(n10378) );
  XNOR2_X1 U13612 ( .A(n10380), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15313) );
  NAND2_X1 U13613 ( .A1(n12185), .A2(n9763), .ZN(n12199) );
  NAND3_X1 U13614 ( .A1(n10176), .A2(n9845), .A3(n10747), .ZN(n12404) );
  AND2_X2 U13615 ( .A1(n12029), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12030) );
  NAND2_X1 U13616 ( .A1(n10388), .A2(n21106), .ZN(n14165) );
  NAND2_X1 U13617 ( .A1(n10392), .A2(n12185), .ZN(n10393) );
  NAND3_X1 U13618 ( .A1(n14488), .A2(n10393), .A3(n12667), .ZN(n12203) );
  NOR2_X1 U13619 ( .A1(n12443), .A2(n10398), .ZN(n12444) );
  NAND3_X1 U13620 ( .A1(n12673), .A2(n12201), .A3(n10395), .ZN(n10522) );
  OAI21_X1 U13621 ( .B1(n10398), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U13622 ( .A1(n10401), .A2(n11316), .ZN(n10636) );
  NAND2_X2 U13623 ( .A1(n10402), .A2(n11114), .ZN(n14312) );
  OAI21_X1 U13624 ( .B1(n15362), .B2(n20873), .A(n15134), .ZN(P1_U2975) );
  OAI21_X1 U13625 ( .B1(n15323), .B2(n20873), .A(n15094), .ZN(P1_U2971) );
  NAND2_X1 U13626 ( .A1(n10413), .A2(n12295), .ZN(n13148) );
  OAI21_X1 U13627 ( .B1(n21384), .B2(n10476), .A(n10474), .ZN(n14293) );
  NAND3_X1 U13628 ( .A1(n10415), .A2(n12424), .A3(n12369), .ZN(n10414) );
  NAND3_X1 U13629 ( .A1(n10910), .A2(n10909), .A3(n10425), .ZN(n10424) );
  NAND2_X1 U13630 ( .A1(n18545), .A2(n10427), .ZN(n12883) );
  NAND3_X1 U13631 ( .A1(n10433), .A2(n10432), .A3(n10431), .ZN(n10430) );
  NAND3_X1 U13632 ( .A1(n10435), .A2(n19800), .A3(n10434), .ZN(n10433) );
  INV_X1 U13633 ( .A(n19778), .ZN(n10436) );
  INV_X2 U13634 ( .A(n19792), .ZN(n19775) );
  AOI22_X1 U13635 ( .A1(n19796), .A2(n19967), .B1(n19794), .B2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19963) );
  NAND2_X2 U13636 ( .A1(n18798), .A2(n9755), .ZN(n18718) );
  AND3_X2 U13637 ( .A1(n10626), .A2(n18952), .A3(n10625), .ZN(n18938) );
  NAND3_X1 U13638 ( .A1(n10450), .A2(n10446), .A3(n10447), .ZN(n10449) );
  OR2_X2 U13639 ( .A1(n18700), .A2(n18920), .ZN(n10446) );
  NAND3_X1 U13640 ( .A1(n10450), .A2(n10824), .A3(n10446), .ZN(n18685) );
  NAND2_X1 U13641 ( .A1(n16401), .A2(n9813), .ZN(n10452) );
  INV_X1 U13642 ( .A(n16387), .ZN(n10454) );
  NAND3_X1 U13643 ( .A1(n12842), .A2(n19174), .A3(n19163), .ZN(n10456) );
  NAND2_X2 U13644 ( .A1(n12840), .A2(n19233), .ZN(n12841) );
  AND2_X4 U13645 ( .A1(n10457), .A2(n9864), .ZN(n18313) );
  NAND3_X1 U13646 ( .A1(n9846), .A2(n10461), .A3(n16895), .ZN(n10460) );
  NAND2_X1 U13647 ( .A1(n20487), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10466) );
  NAND2_X1 U13648 ( .A1(n20454), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10467) );
  AND2_X2 U13649 ( .A1(n11153), .A2(n11147), .ZN(n20454) );
  NAND2_X1 U13650 ( .A1(n20424), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10468) );
  AND2_X2 U13651 ( .A1(n11153), .A2(n11155), .ZN(n20424) );
  NAND2_X1 U13652 ( .A1(n10470), .A2(n10472), .ZN(n11112) );
  INV_X1 U13653 ( .A(n11107), .ZN(n10471) );
  NAND2_X4 U13654 ( .A1(n10560), .A2(n17498), .ZN(n13722) );
  NAND2_X1 U13655 ( .A1(n12396), .A2(n14293), .ZN(n12398) );
  NOR2_X2 U13656 ( .A1(n12700), .A2(n14513), .ZN(n14511) );
  NAND2_X1 U13657 ( .A1(n10493), .A2(n10491), .ZN(n10495) );
  INV_X1 U13658 ( .A(n10492), .ZN(n10491) );
  NAND2_X1 U13659 ( .A1(n10494), .A2(n10496), .ZN(n10493) );
  INV_X1 U13660 ( .A(n12515), .ZN(n10494) );
  NAND2_X1 U13661 ( .A1(n10495), .A2(n9872), .ZN(n12530) );
  NOR2_X2 U13662 ( .A1(n15353), .A2(n10502), .ZN(n15337) );
  AND2_X2 U13663 ( .A1(n10509), .A2(n11288), .ZN(n11289) );
  NAND2_X1 U13664 ( .A1(n10833), .A2(n10834), .ZN(n10509) );
  NAND4_X1 U13665 ( .A1(n17368), .A2(n17285), .A3(n9835), .A4(n11426), .ZN(
        n11065) );
  INV_X1 U13666 ( .A(n11339), .ZN(n10516) );
  NAND3_X2 U13667 ( .A1(n11212), .A2(n10548), .A3(n10550), .ZN(n11290) );
  NAND2_X2 U13668 ( .A1(n10547), .A2(n9836), .ZN(n10550) );
  OR2_X1 U13669 ( .A1(n17087), .A2(n16942), .ZN(n10552) );
  NAND2_X2 U13670 ( .A1(n12189), .A2(n10555), .ZN(n12208) );
  NAND2_X1 U13671 ( .A1(n15550), .A2(n10558), .ZN(n15520) );
  NAND2_X1 U13672 ( .A1(n10653), .A2(n12218), .ZN(n15550) );
  NAND2_X2 U13673 ( .A1(n10560), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12104) );
  NAND2_X1 U13674 ( .A1(n10568), .A2(n18017), .ZN(n10567) );
  OAI21_X1 U13676 ( .B1(n17822), .B2(n10571), .A(n10569), .ZN(n17801) );
  INV_X1 U13677 ( .A(n10575), .ZN(n17802) );
  NAND2_X1 U13678 ( .A1(n10578), .A2(n10576), .ZN(n17935) );
  INV_X1 U13679 ( .A(n18834), .ZN(n10577) );
  NOR2_X1 U13680 ( .A1(n10579), .A2(n18957), .ZN(n10852) );
  NAND3_X1 U13681 ( .A1(n10591), .A2(n10589), .A3(n10588), .ZN(n10587) );
  NAND2_X1 U13682 ( .A1(n10604), .A2(n10602), .ZN(n14769) );
  AND2_X2 U13683 ( .A1(n14692), .A2(n10607), .ZN(n14640) );
  NAND3_X1 U13684 ( .A1(n10616), .A2(n10619), .A3(n10618), .ZN(n10615) );
  OAI21_X1 U13685 ( .B1(n15332), .B2(n20873), .A(n15104), .ZN(P1_U2972) );
  OAI211_X1 U13686 ( .C1(n17651), .C2(n18655), .A(n17649), .B(n17650), .ZN(
        P3_U2834) );
  INV_X1 U13687 ( .A(n12880), .ZN(n10624) );
  NOR2_X1 U13688 ( .A1(n12880), .A2(n18826), .ZN(n18918) );
  INV_X1 U13689 ( .A(n12841), .ZN(n18826) );
  NAND2_X1 U13690 ( .A1(n10626), .A2(n18952), .ZN(n18940) );
  OAI21_X1 U13691 ( .B1(n18953), .B2(n18954), .A(n21839), .ZN(n10626) );
  NAND2_X1 U13692 ( .A1(n11783), .A2(n11782), .ZN(n11795) );
  NAND4_X1 U13693 ( .A1(n10648), .A2(n11210), .A3(n10647), .A4(n10646), .ZN(
        n11243) );
  NAND2_X1 U13694 ( .A1(n11874), .A2(n9943), .ZN(n12724) );
  NAND2_X1 U13695 ( .A1(n11852), .A2(n11853), .ZN(n11860) );
  NAND3_X1 U13696 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13011) );
  NAND2_X1 U13697 ( .A1(n13038), .A2(n9933), .ZN(n12020) );
  NAND2_X1 U13698 ( .A1(n12016), .A2(n10663), .ZN(n13022) );
  INV_X1 U13699 ( .A(n11417), .ZN(n11082) );
  NAND4_X1 U13700 ( .A1(n11046), .A2(n11045), .A3(n11043), .A4(n11044), .ZN(
        n10672) );
  NAND4_X1 U13701 ( .A1(n11041), .A2(n11040), .A3(n11039), .A4(n11042), .ZN(
        n10674) );
  INV_X1 U13702 ( .A(n16903), .ZN(n10676) );
  NAND2_X1 U13703 ( .A1(n11757), .A2(n16901), .ZN(n10677) );
  NAND2_X1 U13704 ( .A1(n11734), .A2(n9900), .ZN(n10678) );
  NAND2_X2 U13705 ( .A1(n10681), .A2(n15935), .ZN(n16903) );
  NAND2_X1 U13706 ( .A1(n11720), .A2(n11894), .ZN(n10681) );
  NAND2_X1 U13707 ( .A1(n16744), .A2(n16742), .ZN(n16730) );
  OAI211_X1 U13708 ( .C1(n16744), .C2(n10688), .A(n9811), .B(n10683), .ZN(
        n17056) );
  NAND2_X1 U13709 ( .A1(n16744), .A2(n10685), .ZN(n10683) );
  INV_X1 U13710 ( .A(n16742), .ZN(n10686) );
  OAI21_X1 U13711 ( .B1(n17056), .B2(n17266), .A(n17055), .ZN(P2_U3025) );
  NAND2_X1 U13712 ( .A1(n16418), .A2(n16417), .ZN(n16416) );
  INV_X1 U13713 ( .A(n16417), .ZN(n10702) );
  NAND2_X1 U13714 ( .A1(n10801), .A2(n16322), .ZN(n10703) );
  XNOR2_X2 U13715 ( .A(n16299), .B(n9925), .ZN(n16408) );
  INV_X1 U13716 ( .A(n10705), .ZN(n16406) );
  NAND2_X1 U13717 ( .A1(n15932), .A2(n10709), .ZN(n10708) );
  NAND2_X1 U13718 ( .A1(n10708), .A2(n10712), .ZN(n14261) );
  NAND2_X1 U13719 ( .A1(n14324), .A2(n10726), .ZN(n15942) );
  NAND2_X2 U13720 ( .A1(n14322), .A2(n14321), .ZN(n14324) );
  INV_X1 U13721 ( .A(n14276), .ZN(n11583) );
  OR2_X2 U13722 ( .A1(n14267), .A2(n10727), .ZN(n14276) );
  NAND2_X1 U13723 ( .A1(n15722), .A2(n9931), .ZN(n15654) );
  NAND2_X1 U13724 ( .A1(n15624), .A2(n10736), .ZN(n14430) );
  NAND2_X1 U13725 ( .A1(n15624), .A2(n15625), .ZN(n13002) );
  AND2_X1 U13726 ( .A1(n11798), .A2(n20181), .ZN(n14191) );
  NAND2_X1 U13727 ( .A1(n10744), .A2(n12042), .ZN(n12097) );
  AND2_X2 U13728 ( .A1(n10744), .A2(n12030), .ZN(n12132) );
  OAI21_X1 U13729 ( .B1(n15521), .B2(n10746), .A(n10745), .ZN(n15533) );
  NAND2_X1 U13730 ( .A1(n10807), .A2(n12124), .ZN(n12177) );
  NOR3_X4 U13731 ( .A1(n15659), .A2(n10761), .A3(n10764), .ZN(n14433) );
  OR3_X1 U13732 ( .A1(n15659), .A2(n10762), .A3(n10764), .ZN(n14434) );
  OAI21_X1 U13733 ( .B1(n12182), .B2(n12178), .A(n21106), .ZN(n12665) );
  NAND2_X1 U13734 ( .A1(n10765), .A2(n13144), .ZN(n13146) );
  NAND3_X1 U13735 ( .A1(n12374), .A2(n12375), .A3(n13335), .ZN(n10765) );
  NAND2_X1 U13736 ( .A1(n14762), .A2(n9932), .ZN(n14706) );
  NAND2_X1 U13737 ( .A1(n14607), .A2(n10770), .ZN(n14566) );
  NOR2_X1 U13738 ( .A1(n14604), .A2(n14605), .ZN(n14596) );
  NOR2_X1 U13739 ( .A1(n14604), .A2(n10772), .ZN(n14581) );
  NOR2_X2 U13740 ( .A1(n14604), .A2(n10768), .ZN(n14567) );
  AND2_X1 U13741 ( .A1(n16735), .A2(n17262), .ZN(n10777) );
  NAND2_X1 U13742 ( .A1(n10780), .A2(n10778), .ZN(n10779) );
  AND2_X1 U13743 ( .A1(n10782), .A2(n11261), .ZN(n16937) );
  NAND2_X2 U13744 ( .A1(n11169), .A2(n17335), .ZN(n16289) );
  INV_X4 U13745 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17335) );
  NAND2_X2 U13746 ( .A1(n10789), .A2(n10786), .ZN(n13989) );
  NAND2_X1 U13747 ( .A1(n10793), .A2(n16698), .ZN(n16674) );
  OAI21_X1 U13748 ( .B1(n16695), .B2(n11869), .A(n11868), .ZN(n10793) );
  OAI21_X2 U13749 ( .B1(n14211), .B2(n14212), .A(n16020), .ZN(n20199) );
  INV_X1 U13750 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12029) );
  INV_X1 U13751 ( .A(n16236), .ZN(n16429) );
  NAND2_X2 U13752 ( .A1(n12416), .A2(n12415), .ZN(n20994) );
  INV_X1 U13753 ( .A(n13024), .ZN(n12018) );
  INV_X1 U13754 ( .A(n11719), .ZN(n11986) );
  NOR2_X1 U13755 ( .A1(n17368), .A2(n17617), .ZN(n13005) );
  OR2_X1 U13756 ( .A1(n12423), .A2(n12422), .ZN(n13189) );
  OR2_X1 U13757 ( .A1(n16388), .A2(n20066), .ZN(n13125) );
  INV_X1 U13758 ( .A(n13564), .ZN(n12222) );
  NAND2_X1 U13759 ( .A1(n11474), .A2(n11473), .ZN(n15932) );
  CLKBUF_X1 U13760 ( .A(n15942), .Z(n15961) );
  INV_X1 U13761 ( .A(n15942), .ZN(n11474) );
  OAI21_X1 U13762 ( .B1(n16017), .B2(n17306), .A(n12715), .ZN(n12716) );
  NAND2_X1 U13763 ( .A1(n15785), .A2(n10805), .ZN(n15769) );
  OR2_X1 U13764 ( .A1(n15034), .A2(n13749), .ZN(n13760) );
  OR2_X1 U13765 ( .A1(n14431), .A2(n11673), .ZN(n11674) );
  NAND2_X1 U13766 ( .A1(n14431), .A2(n11673), .ZN(n12984) );
  AOI22_X1 U13767 ( .A1(n16267), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11027) );
  XNOR2_X1 U13768 ( .A(n13148), .B(n13147), .ZN(n15564) );
  AND2_X1 U13769 ( .A1(n20978), .A2(n21106), .ZN(n20975) );
  NOR2_X1 U13770 ( .A1(n14056), .A2(n9942), .ZN(n14164) );
  INV_X2 U13771 ( .A(n14164), .ZN(n20988) );
  NAND2_X1 U13772 ( .A1(n15576), .A2(n13784), .ZN(n15252) );
  INV_X2 U13773 ( .A(n15252), .ZN(n21000) );
  AND2_X1 U13774 ( .A1(n16872), .A2(n16885), .ZN(n11989) );
  OR2_X1 U13775 ( .A1(n13760), .A2(n15614), .ZN(n15037) );
  NAND2_X1 U13776 ( .A1(n13748), .A2(n14486), .ZN(n15034) );
  INV_X2 U13777 ( .A(n15034), .ZN(n15066) );
  OR3_X1 U13778 ( .A1(n14511), .A2(n14510), .A3(n14503), .ZN(n10796) );
  OR2_X1 U13779 ( .A1(n14437), .A2(n13072), .ZN(n10797) );
  OR2_X1 U13780 ( .A1(n16964), .A2(n20066), .ZN(n10798) );
  AND2_X1 U13781 ( .A1(n12722), .A2(n12721), .ZN(n10799) );
  OR2_X1 U13782 ( .A1(n17478), .A2(n19990), .ZN(n10800) );
  AND2_X1 U13783 ( .A1(n16299), .A2(n9925), .ZN(n10801) );
  AND3_X1 U13784 ( .A1(n12078), .A2(n12077), .A3(n12076), .ZN(n10802) );
  OR2_X1 U13785 ( .A1(n20166), .A2(n11780), .ZN(n10803) );
  OR2_X1 U13786 ( .A1(n20166), .A2(n16421), .ZN(n10804) );
  INV_X1 U13787 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12061) );
  INV_X1 U13788 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11773) );
  NAND2_X1 U13789 ( .A1(n11644), .A2(n11643), .ZN(n10805) );
  AND2_X1 U13790 ( .A1(n12099), .A2(n12098), .ZN(n10806) );
  AND4_X1 U13791 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(
        n10807) );
  NOR2_X1 U13792 ( .A1(n16440), .A2(n16140), .ZN(n10808) );
  INV_X2 U13793 ( .A(n19999), .ZN(n19928) );
  OR2_X1 U13794 ( .A1(n14392), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10809) );
  OR3_X1 U13795 ( .A1(n14514), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14513), .ZN(n10810) );
  INV_X1 U13796 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14503) );
  OR2_X1 U13797 ( .A1(n16515), .A2(n20065), .ZN(n10811) );
  INV_X1 U13798 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13034) );
  INV_X1 U13799 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16842) );
  INV_X1 U13800 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11774) );
  NAND2_X1 U13801 ( .A1(n12365), .A2(n12364), .ZN(n12422) );
  OR2_X1 U13802 ( .A1(n10855), .A2(n17849), .ZN(n10814) );
  XNOR2_X1 U13803 ( .A(n12968), .B(n12967), .ZN(n10815) );
  NAND2_X1 U13804 ( .A1(n12179), .A2(n12562), .ZN(n10816) );
  AND2_X1 U13805 ( .A1(n18390), .A2(n18501), .ZN(n18387) );
  INV_X2 U13806 ( .A(n18387), .ZN(n18379) );
  OR2_X1 U13807 ( .A1(n11983), .A2(n11680), .ZN(n17256) );
  INV_X1 U13808 ( .A(n17256), .ZN(n12994) );
  NAND2_X1 U13809 ( .A1(n10279), .A2(n15999), .ZN(n15740) );
  OR2_X1 U13810 ( .A1(n11245), .A2(n14524), .ZN(n10817) );
  INV_X1 U13811 ( .A(n13362), .ZN(n13335) );
  INV_X1 U13812 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11348) );
  INV_X2 U13813 ( .A(n21746), .ZN(n21734) );
  AND2_X1 U13814 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .ZN(n10818) );
  OR3_X1 U13815 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n18740), .ZN(n10819) );
  XOR2_X1 U13816 ( .A(n16253), .B(n16256), .Z(n10820) );
  NAND3_X1 U13817 ( .A1(n11582), .A2(n11581), .A3(n11580), .ZN(n10821) );
  AND2_X1 U13818 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10822) );
  AND2_X1 U13819 ( .A1(n13173), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10823) );
  NOR2_X1 U13820 ( .A1(n21106), .A2(n21647), .ZN(n13183) );
  INV_X1 U13821 ( .A(n13183), .ZN(n13149) );
  AND2_X1 U13822 ( .A1(n14552), .A2(n17307), .ZN(n16616) );
  OR2_X1 U13823 ( .A1(n9755), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10824) );
  OR2_X1 U13824 ( .A1(n17895), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10825) );
  INV_X1 U13825 ( .A(n14215), .ZN(n20989) );
  AND2_X1 U13826 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10826) );
  NOR2_X1 U13827 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17600), .ZN(n20979) );
  INV_X1 U13828 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12549) );
  AND3_X1 U13829 ( .A1(n13137), .A2(n13136), .A3(n10831), .ZN(n10827) );
  OR2_X1 U13830 ( .A1(n12981), .A2(n12980), .ZN(P3_U2640) );
  AND2_X1 U13831 ( .A1(n12853), .A2(n12943), .ZN(n10829) );
  AND2_X1 U13832 ( .A1(n20800), .A2(n17366), .ZN(n20033) );
  OR2_X1 U13833 ( .A1(n13135), .A2(n19013), .ZN(n10831) );
  NAND2_X1 U13834 ( .A1(n11434), .A2(n11686), .ZN(n10832) );
  INV_X1 U13835 ( .A(n11358), .ZN(n11387) );
  INV_X1 U13836 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17365) );
  AND4_X1 U13837 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(
        n10834) );
  AND2_X1 U13838 ( .A1(n11220), .A2(n11219), .ZN(n10835) );
  AND4_X1 U13839 ( .A1(n12137), .A2(n12136), .A3(n12135), .A4(n12134), .ZN(
        n10836) );
  AND2_X1 U13840 ( .A1(n12110), .A2(n12109), .ZN(n10837) );
  INV_X1 U13841 ( .A(n11684), .ZN(n11067) );
  INV_X1 U13842 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13685) );
  INV_X1 U13843 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U13844 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12099) );
  INV_X1 U13845 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U13846 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20299), .B1(
        n20331), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U13847 ( .A1(n11889), .A2(n14181), .ZN(n11721) );
  AND2_X1 U13848 ( .A1(n17366), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11089) );
  XNOR2_X1 U13849 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12485) );
  OR2_X1 U13850 ( .A1(n12363), .A2(n12362), .ZN(n12433) );
  NAND2_X1 U13851 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12062) );
  OAI21_X1 U13852 ( .B1(n11861), .B2(n10804), .A(n11879), .ZN(n11862) );
  MUX2_X1 U13853 ( .A(n11727), .B(P2_EBX_REG_3__SCAN_IN), .S(n11889), .Z(
        n11732) );
  NAND2_X1 U13854 ( .A1(n14194), .A2(n20156), .ZN(n11026) );
  AOI22_X1 U13855 ( .A1(n16282), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11032) );
  INV_X1 U13856 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12254) );
  INV_X1 U13857 ( .A(n12437), .ZN(n12443) );
  INV_X1 U13858 ( .A(n14286), .ZN(n12564) );
  INV_X1 U13859 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13532) );
  NAND2_X1 U13860 ( .A1(n11358), .A2(n11388), .ZN(n11389) );
  INV_X1 U13861 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U13862 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11046) );
  INV_X1 U13863 ( .A(n14353), .ZN(n11918) );
  AND2_X1 U13864 ( .A1(n11409), .A2(n11408), .ZN(n13959) );
  OR4_X1 U13865 ( .A1(n12520), .A2(n12503), .A3(n12509), .A4(n12516), .ZN(
        n12487) );
  NOR2_X1 U13866 ( .A1(n13722), .A2(n12157), .ZN(n12158) );
  AND2_X1 U13867 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13297) );
  INV_X1 U13868 ( .A(n13141), .ZN(n13143) );
  AND2_X1 U13869 ( .A1(n15375), .A2(n15374), .ZN(n15460) );
  OR2_X1 U13870 ( .A1(n12420), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12418) );
  AND2_X1 U13871 ( .A1(n12176), .A2(n9763), .ZN(n12188) );
  OR2_X1 U13872 ( .A1(n12518), .A2(n13532), .ZN(n12270) );
  INV_X1 U13873 ( .A(n11363), .ZN(n11364) );
  INV_X1 U13874 ( .A(n15676), .ZN(n11961) );
  INV_X1 U13875 ( .A(n15830), .ZN(n11929) );
  OR2_X1 U13876 ( .A1(n16276), .A2(n16280), .ZN(n16314) );
  AND2_X1 U13877 ( .A1(n12717), .A2(n16638), .ZN(n12719) );
  AND2_X1 U13878 ( .A1(n11667), .A2(n11666), .ZN(n13003) );
  OR2_X1 U13879 ( .A1(n17204), .A2(n17188), .ZN(n17046) );
  INV_X1 U13880 ( .A(n18738), .ZN(n10854) );
  INV_X1 U13881 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21810) );
  INV_X1 U13882 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n21817) );
  INV_X1 U13883 ( .A(n13107), .ZN(n13090) );
  INV_X1 U13884 ( .A(n19814), .ZN(n17478) );
  INV_X1 U13885 ( .A(n14940), .ZN(n12593) );
  NAND2_X1 U13886 ( .A1(n13356), .A2(n13297), .ZN(n13316) );
  AOI21_X1 U13887 ( .B1(n13188), .B2(n13335), .A(n13187), .ZN(n14952) );
  OR2_X1 U13888 ( .A1(n21008), .A2(n12684), .ZN(n15374) );
  NAND2_X1 U13889 ( .A1(n21060), .A2(n12186), .ZN(n13785) );
  INV_X1 U13890 ( .A(n21142), .ZN(n21173) );
  INV_X1 U13891 ( .A(n15567), .ZN(n21430) );
  INV_X1 U13892 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21468) );
  INV_X1 U13893 ( .A(n11892), .ZN(n11885) );
  NAND2_X1 U13894 ( .A1(n11855), .A2(n11879), .ZN(n11852) );
  INV_X1 U13895 ( .A(n13031), .ZN(n13035) );
  INV_X1 U13896 ( .A(n11977), .ZN(n12707) );
  AND2_X1 U13897 ( .A1(n16297), .A2(n16296), .ZN(n16315) );
  AND2_X1 U13898 ( .A1(n11887), .A2(n16673), .ZN(n16685) );
  NOR2_X1 U13899 ( .A1(n11870), .A2(n11348), .ZN(n16700) );
  NAND2_X1 U13900 ( .A1(n15735), .A2(n11864), .ZN(n11835) );
  AND2_X1 U13901 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12957) );
  AND2_X1 U13902 ( .A1(n14169), .A2(n14200), .ZN(n20548) );
  INV_X1 U13903 ( .A(n20151), .ZN(n20180) );
  INV_X1 U13904 ( .A(n13108), .ZN(n13109) );
  INV_X1 U13905 ( .A(n19183), .ZN(n19158) );
  INV_X1 U13906 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19303) );
  OR2_X1 U13907 ( .A1(n19962), .A2(n19845), .ZN(n19347) );
  INV_X1 U13908 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14708) );
  NOR2_X1 U13909 ( .A1(n14505), .A2(n21644), .ZN(n14405) );
  NAND2_X1 U13910 ( .A1(n20904), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14456) );
  AND2_X1 U13911 ( .A1(n14402), .A2(n13682), .ZN(n14583) );
  AND2_X1 U13912 ( .A1(n12608), .A2(n12607), .ZN(n14818) );
  NAND2_X1 U13913 ( .A1(n10026), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13362) );
  INV_X1 U13914 ( .A(n13472), .ZN(n14707) );
  AND2_X1 U13915 ( .A1(n13335), .A2(n13282), .ZN(n14848) );
  NOR2_X1 U13916 ( .A1(n13251), .A2(n20900), .ZN(n13252) );
  NAND2_X1 U13917 ( .A1(n17592), .A2(n21645), .ZN(n13791) );
  NAND2_X1 U13918 ( .A1(n12184), .A2(n21060), .ZN(n12556) );
  INV_X1 U13919 ( .A(n17500), .ZN(n15552) );
  INV_X1 U13920 ( .A(n13145), .ZN(n15574) );
  INV_X1 U13921 ( .A(n21539), .ZN(n21514) );
  AND2_X1 U13922 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21114), .ZN(n21105) );
  OR2_X1 U13923 ( .A1(n11411), .A2(n11401), .ZN(n11403) );
  NOR2_X1 U13924 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17366) );
  INV_X1 U13925 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15664) );
  INV_X1 U13926 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15698) );
  INV_X1 U13927 ( .A(n11852), .ZN(n11789) );
  INV_X1 U13928 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15851) );
  INV_X1 U13929 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16494) );
  OR2_X1 U13930 ( .A1(n14310), .A2(n10244), .ZN(n14346) );
  AND2_X1 U13931 ( .A1(n11669), .A2(n11668), .ZN(n14429) );
  INV_X1 U13932 ( .A(n17348), .ZN(n13963) );
  AOI21_X1 U13933 ( .B1(n16438), .B2(n16935), .A(n12024), .ZN(n12025) );
  OR2_X1 U13934 ( .A1(n11847), .A2(n12005), .ZN(n16727) );
  OR2_X1 U13935 ( .A1(n11983), .A2(n17346), .ZN(n11701) );
  OR2_X1 U13936 ( .A1(n11845), .A2(n16857), .ZN(n16849) );
  INV_X1 U13937 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17253) );
  INV_X1 U13938 ( .A(n20801), .ZN(n20264) );
  NOR3_X1 U13939 ( .A1(n20390), .A2(n17300), .A3(n20421), .ZN(n20391) );
  INV_X1 U13940 ( .A(n20192), .ZN(n20450) );
  OR2_X1 U13941 ( .A1(n20817), .A2(n20134), .ZN(n20655) );
  OAI211_X1 U13942 ( .C1(n10542), .C2(n12859), .A(n10965), .B(n10964), .ZN(
        n12860) );
  NOR2_X1 U13943 ( .A1(n18394), .A2(n18393), .ZN(n18395) );
  NOR2_X1 U13944 ( .A1(n18735), .A2(n10853), .ZN(n18693) );
  NOR2_X1 U13945 ( .A1(n19006), .A2(n18770), .ZN(n18771) );
  INV_X1 U13946 ( .A(n17982), .ZN(n17993) );
  NAND2_X1 U13947 ( .A1(n12846), .A2(n10819), .ZN(n12847) );
  INV_X1 U13948 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n19163) );
  XNOR2_X1 U13949 ( .A(n12827), .B(n19303), .ZN(n18988) );
  INV_X1 U13950 ( .A(n19326), .ZN(n19794) );
  INV_X2 U13951 ( .A(n9732), .ZN(n18039) );
  INV_X1 U13952 ( .A(n19514), .ZN(n19489) );
  INV_X1 U13953 ( .A(n19839), .ZN(n19680) );
  INV_X1 U13954 ( .A(n20925), .ZN(n20945) );
  AND2_X1 U13955 ( .A1(n14405), .A2(n20904), .ZN(n20914) );
  OR2_X1 U13956 ( .A1(n20914), .A2(n14454), .ZN(n20950) );
  INV_X1 U13957 ( .A(n20978), .ZN(n14943) );
  INV_X1 U13958 ( .A(n15037), .ZN(n15029) );
  NOR2_X1 U13959 ( .A1(n14948), .A2(n14877), .ZN(n14939) );
  AND2_X1 U13960 ( .A1(n15066), .A2(n14165), .ZN(n15026) );
  INV_X1 U13961 ( .A(n21006), .ZN(n15178) );
  NAND2_X1 U13962 ( .A1(n13191), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13251) );
  NAND2_X1 U13963 ( .A1(n13185), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13190) );
  NAND2_X1 U13964 ( .A1(n15557), .A2(n14486), .ZN(n14086) );
  NAND2_X1 U13965 ( .A1(n20873), .A2(n13792), .ZN(n15173) );
  AND2_X1 U13966 ( .A1(n17559), .A2(n12676), .ZN(n21035) );
  OAI22_X1 U13967 ( .A1(n15613), .A2(n15608), .B1(n21329), .B2(n21203), .ZN(
        n21110) );
  OAI211_X1 U13968 ( .C1(n21517), .C2(n21117), .A(n21588), .B(n21116), .ZN(
        n21136) );
  INV_X1 U13969 ( .A(n21160), .ZN(n21167) );
  OAI21_X1 U13970 ( .B1(n21180), .B2(n21179), .A(n21178), .ZN(n21197) );
  OAI21_X1 U13971 ( .B1(n21541), .B2(n21203), .A(n21202), .ZN(n21223) );
  OAI22_X1 U13972 ( .A1(n21264), .A2(n21263), .B1(n21262), .B2(n21541), .ZN(
        n21290) );
  OAI211_X1 U13973 ( .C1(n21301), .C2(n21517), .A(n21588), .B(n21300), .ZN(
        n21322) );
  INV_X1 U13974 ( .A(n21315), .ZN(n21351) );
  OAI211_X1 U13975 ( .C1(n21517), .C2(n21359), .A(n21588), .B(n21358), .ZN(
        n21377) );
  NOR2_X2 U13976 ( .A1(n21437), .A2(n21360), .ZN(n21419) );
  OAI21_X1 U13977 ( .B1(n21435), .B2(n21434), .A(n21433), .ZN(n21458) );
  NOR2_X2 U13978 ( .A1(n21514), .A2(n21462), .ZN(n21534) );
  AND2_X1 U13979 ( .A1(n12184), .A2(n21105), .ZN(n21583) );
  AND2_X1 U13980 ( .A1(n10013), .A2(n21105), .ZN(n21601) );
  INV_X1 U13981 ( .A(n21408), .ZN(n21619) );
  OAI21_X1 U13982 ( .B1(n21587), .B2(n21647), .A(n21581), .ZN(n21635) );
  NAND2_X1 U13983 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21653) );
  INV_X1 U13984 ( .A(n21653), .ZN(n21739) );
  INV_X1 U13985 ( .A(n21709), .ZN(n21705) );
  NAND2_X1 U13986 ( .A1(n11403), .A2(n11402), .ZN(n17348) );
  INV_X1 U13987 ( .A(n16009), .ZN(n20057) );
  NOR2_X1 U13988 ( .A1(n14350), .A2(n16024), .ZN(n16495) );
  NOR2_X1 U13989 ( .A1(n14361), .A2(n16156), .ZN(n16493) );
  AND2_X1 U13990 ( .A1(n16458), .A2(n16450), .ZN(n16451) );
  AND2_X1 U13991 ( .A1(n13843), .A2(n13842), .ZN(n22063) );
  INV_X1 U13992 ( .A(n13907), .ZN(n13955) );
  AND2_X1 U13993 ( .A1(n13005), .A2(n13963), .ZN(n14556) );
  INV_X1 U13994 ( .A(n16911), .ZN(n16939) );
  INV_X1 U13995 ( .A(n16693), .ZN(n16706) );
  AND2_X1 U13996 ( .A1(n14351), .A2(n14354), .ZN(n17183) );
  NAND2_X1 U13997 ( .A1(n11432), .A2(n17372), .ZN(n11983) );
  NAND2_X1 U13998 ( .A1(n20143), .A2(n20142), .ZN(n20185) );
  OAI21_X1 U13999 ( .B1(n20193), .B2(n20808), .A(n20191), .ZN(n20216) );
  OAI21_X1 U14000 ( .B1(n17300), .B2(n20263), .A(n20262), .ZN(n20289) );
  NOR2_X2 U14001 ( .A1(n20396), .A2(n20264), .ZN(n20322) );
  OAI22_X1 U14002 ( .A1(n20334), .A2(n20333), .B1(n17300), .B2(n20332), .ZN(
        n20352) );
  NOR2_X2 U14003 ( .A1(n20396), .A2(n20327), .ZN(n20384) );
  INV_X1 U14004 ( .A(n20425), .ZN(n20421) );
  NAND2_X1 U14005 ( .A1(n12015), .A2(n12014), .ZN(n20660) );
  OAI21_X1 U14006 ( .B1(n20575), .B2(n20814), .A(n20558), .ZN(n20577) );
  NOR2_X2 U14007 ( .A1(n20608), .A2(n20327), .ZN(n20604) );
  INV_X1 U14008 ( .A(n20327), .ZN(n20294) );
  INV_X1 U14009 ( .A(n20257), .ZN(n20652) );
  INV_X1 U14010 ( .A(n20629), .ZN(n20684) );
  NOR2_X2 U14011 ( .A1(n17307), .A2(n17306), .ZN(n20176) );
  AND2_X1 U14012 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17270) );
  NOR2_X1 U14013 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19995) );
  AND2_X1 U14014 ( .A1(n17483), .A2(n12881), .ZN(n19813) );
  NOR2_X1 U14015 ( .A1(n17752), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10975) );
  INV_X1 U14016 ( .A(n18090), .ZN(n18080) );
  NOR2_X1 U14017 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17947), .ZN(n17930) );
  INV_X1 U14018 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20001) );
  NOR2_X2 U14019 ( .A1(n19829), .A2(n10969), .ZN(n18055) );
  NOR2_X1 U14020 ( .A1(n18605), .A2(n18459), .ZN(n18453) );
  INV_X1 U14021 ( .A(n18444), .ZN(n18471) );
  NOR2_X1 U14022 ( .A1(n18577), .A2(n18499), .ZN(n18495) );
  INV_X1 U14023 ( .A(n19349), .ZN(n18546) );
  NAND2_X1 U14024 ( .A1(n19985), .A2(n19814), .ZN(n18598) );
  INV_X1 U14025 ( .A(n18610), .ZN(n18648) );
  NAND2_X1 U14026 ( .A1(n18660), .A2(n18661), .ZN(n18659) );
  NOR2_X1 U14027 ( .A1(n19113), .A2(n18741), .ZN(n19077) );
  INV_X1 U14028 ( .A(n19116), .ZN(n19113) );
  INV_X1 U14029 ( .A(n19421), .ZN(n19632) );
  INV_X1 U14030 ( .A(n17634), .ZN(n18670) );
  INV_X1 U14031 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21959) );
  INV_X1 U14032 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19070) );
  INV_X1 U14033 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n22014) );
  NOR2_X2 U14034 ( .A1(n18510), .A2(n19297), .ZN(n19239) );
  NOR2_X1 U14035 ( .A1(n12858), .A2(n12866), .ZN(n19810) );
  NOR2_X1 U14036 ( .A1(n19317), .A2(n19327), .ZN(n19325) );
  NOR2_X1 U14037 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19937), .ZN(
        n19962) );
  AND2_X1 U14038 ( .A1(n19680), .A2(n19400), .ZN(n19373) );
  INV_X1 U14039 ( .A(n19504), .ZN(n19508) );
  INV_X1 U14040 ( .A(n19725), .ZN(n19681) );
  AND2_X1 U14041 ( .A1(n19680), .A2(n19686), .ZN(n19711) );
  INV_X1 U14042 ( .A(n19623), .ZN(n19757) );
  NOR2_X1 U14043 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19937), .ZN(n19839) );
  NOR2_X1 U14044 ( .A1(n19841), .A2(n20001), .ZN(n19985) );
  INV_X1 U14045 ( .A(n19981), .ZN(n19990) );
  INV_X1 U14046 ( .A(n17305), .ZN(n17307) );
  INV_X1 U14047 ( .A(U212), .ZN(n17687) );
  OR2_X1 U14048 ( .A1(n14086), .A2(n12543), .ZN(n14056) );
  INV_X1 U14049 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21880) );
  AOI21_X1 U14050 ( .B1(n14575), .B2(n20954), .A(n14574), .ZN(n14576) );
  INV_X1 U14051 ( .A(n20950), .ZN(n20962) );
  OR2_X1 U14052 ( .A1(n13760), .A2(n15615), .ZN(n15033) );
  AND2_X1 U14053 ( .A1(n14061), .A2(n14060), .ZN(n21108) );
  AND2_X1 U14054 ( .A1(n14083), .A2(n14082), .ZN(n21072) );
  NAND2_X1 U14055 ( .A1(n20980), .A2(n12184), .ZN(n14153) );
  INV_X2 U14056 ( .A(n20979), .ZN(n14160) );
  OR2_X1 U14057 ( .A1(n14056), .A2(n14055), .ZN(n14242) );
  OAI21_X1 U14058 ( .B1(n14798), .B2(n14783), .A(n14782), .ZN(n15223) );
  INV_X1 U14059 ( .A(n21027), .ZN(n21054) );
  INV_X1 U14060 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21509) );
  OR2_X1 U14061 ( .A1(n21175), .A2(n21462), .ZN(n21132) );
  AOI22_X1 U14062 ( .A1(n21143), .A2(n21146), .B1(n21388), .B2(n21144), .ZN(
        n21171) );
  INV_X1 U14063 ( .A(n21174), .ZN(n21200) );
  NAND2_X1 U14064 ( .A1(n21303), .A2(n21326), .ZN(n21245) );
  NAND2_X1 U14065 ( .A1(n21303), .A2(n21507), .ZN(n21287) );
  NAND2_X1 U14066 ( .A1(n21303), .A2(n21538), .ZN(n21325) );
  AOI22_X1 U14067 ( .A1(n21394), .A2(n21390), .B1(n21388), .B2(n21387), .ZN(
        n21423) );
  NAND2_X1 U14068 ( .A1(n21381), .A2(n21538), .ZN(n21461) );
  INV_X1 U14069 ( .A(n21602), .ZN(n21485) );
  INV_X1 U14070 ( .A(n21636), .ZN(n21505) );
  NAND2_X1 U14071 ( .A1(n21539), .A2(n21507), .ZN(n21543) );
  INV_X1 U14072 ( .A(n21621), .ZN(n21566) );
  INV_X1 U14073 ( .A(n21489), .ZN(n21618) );
  INV_X1 U14074 ( .A(n21496), .ZN(n21632) );
  INV_X1 U14075 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21474) );
  NOR2_X1 U14076 ( .A1(n21734), .A2(n20871), .ZN(n21724) );
  INV_X1 U14077 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21661) );
  INV_X1 U14078 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20481) );
  OR2_X1 U14079 ( .A1(n13958), .A2(n17367), .ZN(n20065) );
  INV_X1 U14080 ( .A(n20031), .ZN(n20073) );
  NAND2_X1 U14081 ( .A1(n20084), .A2(n14194), .ZN(n16625) );
  AND2_X1 U14082 ( .A1(n14190), .A2(n17372), .ZN(n20084) );
  NAND2_X1 U14083 ( .A1(n20084), .A2(n9749), .ZN(n20085) );
  NAND2_X1 U14084 ( .A1(n13879), .A2(n11084), .ZN(n13977) );
  NAND2_X1 U14085 ( .A1(n10286), .A2(n17270), .ZN(n20845) );
  NAND2_X1 U14086 ( .A1(n20132), .A2(n20845), .ZN(n20101) );
  INV_X1 U14087 ( .A(n14556), .ZN(n13958) );
  AOI21_X1 U14088 ( .B1(n12027), .B2(n16939), .A(n12026), .ZN(n12028) );
  NAND2_X1 U14089 ( .A1(n12009), .A2(n20854), .ZN(n16911) );
  AOI21_X1 U14090 ( .B1(n16438), .B2(n17260), .A(n12964), .ZN(n12965) );
  INV_X1 U14091 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20812) );
  INV_X1 U14092 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17362) );
  NAND2_X1 U14093 ( .A1(n20192), .A2(n20357), .ZN(n20220) );
  AND2_X1 U14094 ( .A1(n20256), .A2(n20255), .ZN(n20271) );
  NAND2_X1 U14095 ( .A1(n20357), .A2(n20801), .ZN(n20287) );
  INV_X1 U14096 ( .A(n20351), .ZN(n20347) );
  INV_X1 U14097 ( .A(n20384), .ZN(n20361) );
  NAND2_X1 U14098 ( .A1(n20357), .A2(n20356), .ZN(n20415) );
  INV_X1 U14099 ( .A(n20417), .ZN(n20448) );
  INV_X1 U14100 ( .A(n20470), .ZN(n20478) );
  INV_X1 U14101 ( .A(n20508), .ZN(n20505) );
  NAND2_X1 U14102 ( .A1(n20479), .A2(n20801), .ZN(n20541) );
  INV_X1 U14103 ( .A(n20686), .ZN(n20630) );
  INV_X1 U14104 ( .A(n20698), .ZN(n20638) );
  INV_X1 U14105 ( .A(n20674), .ZN(n20626) );
  INV_X1 U14106 ( .A(n20586), .ZN(n20671) );
  NAND2_X1 U14107 ( .A1(n20526), .A2(n20356), .ZN(n20702) );
  AOI21_X1 U14108 ( .B1(n17370), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n17369), 
        .ZN(n17612) );
  INV_X1 U14109 ( .A(n20792), .ZN(n20715) );
  INV_X1 U14110 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20728) );
  CLKBUF_X1 U14111 ( .A(n20782), .Z(n20777) );
  NAND2_X1 U14112 ( .A1(n19946), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19841) );
  INV_X1 U14113 ( .A(n18067), .ZN(n10977) );
  INV_X1 U14114 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18759) );
  INV_X1 U14115 ( .A(n18074), .ZN(n18059) );
  INV_X1 U14116 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18956) );
  NOR2_X1 U14117 ( .A1(n18103), .A2(n18102), .ZN(n18129) );
  INV_X1 U14118 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18370) );
  INV_X1 U14119 ( .A(n18537), .ZN(n18525) );
  OR2_X1 U14120 ( .A1(n19946), .A2(n19848), .ZN(n18559) );
  OR2_X1 U14121 ( .A1(n19982), .A2(n18568), .ZN(n18567) );
  INV_X1 U14122 ( .A(n18568), .ZN(n18593) );
  AOI211_X1 U14123 ( .C1(n19990), .C2(n18596), .A(n18595), .B(n18598), .ZN(
        n18610) );
  INV_X1 U14124 ( .A(n18649), .ZN(n18646) );
  INV_X1 U14125 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n19136) );
  INV_X1 U14126 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18895) );
  INV_X1 U14127 ( .A(n19002), .ZN(n18994) );
  NAND2_X1 U14128 ( .A1(n19685), .A2(n19632), .ZN(n19369) );
  INV_X1 U14129 ( .A(n13111), .ZN(n13112) );
  INV_X1 U14130 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21877) );
  INV_X1 U14131 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n19227) );
  INV_X1 U14132 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19251) );
  NAND2_X1 U14133 ( .A1(n19810), .A2(n19327), .ZN(n19297) );
  INV_X1 U14134 ( .A(n17470), .ZN(n19984) );
  INV_X1 U14135 ( .A(n19713), .ZN(n19399) );
  INV_X1 U14136 ( .A(n19769), .ZN(n19416) );
  INV_X1 U14137 ( .A(n19438), .ZN(n19445) );
  INV_X1 U14138 ( .A(n19481), .ZN(n19488) );
  INV_X1 U14139 ( .A(n19549), .ZN(n19556) );
  INV_X1 U14140 ( .A(n19599), .ZN(n19597) );
  INV_X1 U14141 ( .A(n19643), .ZN(n19653) );
  INV_X1 U14142 ( .A(n19732), .ZN(n19697) );
  OR2_X1 U14143 ( .A1(n19800), .A2(n19656), .ZN(n19762) );
  INV_X1 U14144 ( .A(n19985), .ZN(n19836) );
  INV_X1 U14145 ( .A(n19934), .ZN(n19931) );
  INV_X1 U14146 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19869) );
  INV_X1 U14147 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19894) );
  INV_X1 U14148 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n21883) );
  NOR2_X1 U14149 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13779), .ZN(n17722)
         );
  INV_X1 U14150 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20775) );
  OAI211_X1 U14151 ( .C1(n12999), .C2(n16911), .A(n12730), .B(n12729), .ZN(
        P2_U2983) );
  NAND4_X1 U14152 ( .A1(n15615), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n13768), .A4(
        n13767), .ZN(U214) );
  NAND2_X1 U14153 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18028), .ZN(
        n18957) );
  NAND3_X1 U14154 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17943) );
  NAND2_X1 U14155 ( .A1(n18847), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18811) );
  INV_X1 U14156 ( .A(n18812), .ZN(n10838) );
  NAND2_X1 U14157 ( .A1(n18808), .A2(n10838), .ZN(n17872) );
  INV_X1 U14158 ( .A(n18773), .ZN(n10839) );
  NAND2_X1 U14159 ( .A1(n18691), .A2(n10822), .ZN(n18682) );
  NOR2_X2 U14160 ( .A1(n18682), .A2(n22029), .ZN(n18663) );
  NAND2_X1 U14161 ( .A1(n18663), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10842) );
  NAND2_X1 U14162 ( .A1(n10840), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12933) );
  XOR2_X1 U14163 ( .A(n10850), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12968) );
  INV_X1 U14164 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21895) );
  INV_X1 U14165 ( .A(n10840), .ZN(n17624) );
  NOR2_X1 U14166 ( .A1(n19006), .A2(n17624), .ZN(n12935) );
  INV_X1 U14167 ( .A(n12935), .ZN(n10841) );
  AOI21_X1 U14168 ( .B1(n21895), .B2(n10841), .A(n10850), .ZN(n17749) );
  OR2_X1 U14169 ( .A1(n19006), .A2(n10842), .ZN(n10843) );
  AOI21_X1 U14170 ( .B1(n17764), .B2(n10843), .A(n12935), .ZN(n18654) );
  INV_X1 U14171 ( .A(n18663), .ZN(n18662) );
  NOR2_X1 U14172 ( .A1(n19006), .A2(n18662), .ZN(n10845) );
  OAI21_X1 U14173 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n10845), .A(
        n10843), .ZN(n18673) );
  INV_X1 U14174 ( .A(n18673), .ZN(n17768) );
  INV_X1 U14175 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18735) );
  INV_X1 U14176 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18747) );
  INV_X1 U14177 ( .A(n10844), .ZN(n18770) );
  NAND2_X1 U14178 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17849), .ZN(
        n10849) );
  NOR2_X1 U14179 ( .A1(n18747), .A2(n10849), .ZN(n10848) );
  INV_X1 U14180 ( .A(n10848), .ZN(n10853) );
  NAND2_X1 U14181 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18693), .ZN(
        n10846) );
  NAND3_X1 U14182 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n10856), .ZN(n18665) );
  AOI21_X1 U14183 ( .B1(n22029), .B2(n18665), .A(n10845), .ZN(n18684) );
  INV_X1 U14184 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18710) );
  AOI22_X1 U14185 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n10856), .B1(
        n10846), .B2(n18710), .ZN(n18713) );
  OAI21_X1 U14186 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18693), .A(
        n10846), .ZN(n10847) );
  INV_X1 U14187 ( .A(n10847), .ZN(n18722) );
  AOI21_X1 U14188 ( .B1(n18747), .B2(n10849), .A(n10848), .ZN(n18750) );
  OAI21_X1 U14189 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17849), .A(
        n10849), .ZN(n18761) );
  INV_X1 U14190 ( .A(n18761), .ZN(n17840) );
  NAND2_X1 U14191 ( .A1(n10850), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10851) );
  INV_X4 U14192 ( .A(n10855), .ZN(n18017) );
  NAND2_X1 U14193 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10852), .ZN(
        n17982) );
  NAND2_X1 U14194 ( .A1(n18834), .A2(n17993), .ZN(n17944) );
  NOR2_X1 U14195 ( .A1(n18811), .A2(n17944), .ZN(n18810) );
  NAND2_X1 U14196 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18810), .ZN(
        n17895) );
  NOR2_X1 U14197 ( .A1(n18750), .A2(n17831), .ZN(n17830) );
  OR2_X1 U14198 ( .A1(n17830), .A2(n18043), .ZN(n17821) );
  AOI21_X1 U14199 ( .B1(n18735), .B2(n10853), .A(n18693), .ZN(n18738) );
  NAND2_X1 U14200 ( .A1(n17821), .A2(n10854), .ZN(n17822) );
  NOR2_X1 U14201 ( .A1(n17801), .A2(n18043), .ZN(n17789) );
  INV_X1 U14202 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18695) );
  NAND2_X1 U14203 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n10856), .ZN(
        n10858) );
  INV_X1 U14204 ( .A(n18665), .ZN(n10857) );
  AOI21_X1 U14205 ( .B1(n18695), .B2(n10858), .A(n10857), .ZN(n18698) );
  NOR2_X1 U14206 ( .A1(n17789), .A2(n18698), .ZN(n17788) );
  NOR2_X1 U14207 ( .A1(n17788), .A2(n18043), .ZN(n17780) );
  NOR2_X1 U14208 ( .A1(n17779), .A2(n18043), .ZN(n17767) );
  NOR2_X1 U14209 ( .A1(n17768), .A2(n17767), .ZN(n17766) );
  NOR2_X1 U14210 ( .A1(n17766), .A2(n18043), .ZN(n17757) );
  NOR4_X4 U14211 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n19946), .ZN(n18067) );
  INV_X1 U14212 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19988) );
  NAND2_X1 U14213 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19981) );
  INV_X1 U14214 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10859) );
  INV_X2 U14215 ( .A(n12733), .ZN(n18345) );
  AOI22_X1 U14216 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U14217 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U14218 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10862) );
  NAND2_X2 U14219 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U14220 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10861) );
  NAND4_X1 U14221 ( .A1(n10864), .A2(n10863), .A3(n10862), .A4(n10861), .ZN(
        n10875) );
  AOI22_X1 U14222 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10873) );
  NOR2_X2 U14223 ( .A1(n19787), .A2(n10869), .ZN(n12808) );
  AOI22_X1 U14224 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10872) );
  NOR2_X2 U14225 ( .A1(n10866), .A2(n10867), .ZN(n18343) );
  INV_X2 U14226 ( .A(n18267), .ZN(n18297) );
  NOR2_X2 U14227 ( .A1(n19787), .A2(n10867), .ZN(n12768) );
  BUF_X4 U14228 ( .A(n12768), .Z(n18322) );
  AOI22_X1 U14229 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10871) );
  NOR2_X2 U14230 ( .A1(n10868), .A2(n18072), .ZN(n12816) );
  AOI22_X1 U14231 ( .A1(n18314), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10870) );
  NAND4_X1 U14232 ( .A1(n10873), .A2(n10872), .A3(n10871), .A4(n10870), .ZN(
        n10874) );
  AOI22_X1 U14233 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18343), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U14234 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10878) );
  INV_X4 U14235 ( .A(n10931), .ZN(n18268) );
  AOI22_X1 U14236 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18212), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U14237 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U14238 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U14239 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U14240 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U14241 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U14242 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10887) );
  INV_X2 U14243 ( .A(n18106), .ZN(n17456) );
  AOI22_X1 U14244 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U14245 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U14246 ( .A1(n18315), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10884) );
  NAND4_X1 U14247 ( .A1(n10887), .A2(n10886), .A3(n10885), .A4(n10884), .ZN(
        n10893) );
  AOI22_X1 U14248 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U14249 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U14250 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U14251 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10888) );
  NAND4_X1 U14252 ( .A1(n10891), .A2(n10890), .A3(n10889), .A4(n10888), .ZN(
        n10892) );
  AOI22_X1 U14253 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U14254 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U14255 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10894) );
  OAI21_X1 U14256 ( .B1(n18239), .B2(n18381), .A(n10894), .ZN(n10898) );
  AOI22_X1 U14257 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U14258 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U14259 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U14260 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U14261 ( .A1(n18314), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U14262 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10902) );
  OAI21_X1 U14263 ( .B1(n10931), .B2(n21810), .A(n10902), .ZN(n10908) );
  AOI22_X1 U14264 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U14265 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U14266 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U14267 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10903) );
  NAND4_X1 U14268 ( .A1(n10906), .A2(n10905), .A3(n10904), .A4(n10903), .ZN(
        n10907) );
  INV_X1 U14269 ( .A(n18391), .ZN(n19370) );
  AOI22_X1 U14270 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U14271 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10913) );
  INV_X2 U14272 ( .A(n18267), .ZN(n17455) );
  AOI22_X1 U14273 ( .A1(n18314), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U14274 ( .A1(n18315), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10911) );
  NAND4_X1 U14275 ( .A1(n10914), .A2(n10913), .A3(n10912), .A4(n10911), .ZN(
        n10920) );
  AOI22_X1 U14276 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U14277 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U14278 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U14279 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10915) );
  NAND4_X1 U14280 ( .A1(n10918), .A2(n10917), .A3(n10916), .A4(n10915), .ZN(
        n10919) );
  NAND2_X1 U14281 ( .A1(n19779), .A2(n12856), .ZN(n14381) );
  NOR2_X1 U14282 ( .A1(n10944), .A2(n14381), .ZN(n10942) );
  AOI22_X1 U14283 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U14284 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U14285 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17456), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U14286 ( .A1(n18315), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10921) );
  NAND4_X1 U14287 ( .A1(n10924), .A2(n10923), .A3(n10922), .A4(n10921), .ZN(
        n10930) );
  AOI22_X1 U14288 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17439), .ZN(n10928) );
  AOI22_X1 U14289 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18039), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U14290 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18312), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U14291 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10925) );
  NAND4_X1 U14292 ( .A1(n10928), .A2(n10927), .A3(n10926), .A4(n10925), .ZN(
        n10929) );
  AOI22_X1 U14293 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17439), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U14294 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U14295 ( .A1(n18314), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U14296 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10932) );
  NAND4_X1 U14297 ( .A1(n10935), .A2(n10934), .A3(n10933), .A4(n10932), .ZN(
        n10941) );
  AOI22_X1 U14298 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U14299 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U14300 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U14301 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10936) );
  NAND4_X1 U14302 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(
        n10940) );
  NOR3_X2 U14303 ( .A1(n12854), .A2(n18391), .A3(n14380), .ZN(n10949) );
  NAND4_X1 U14304 ( .A1(n12885), .A2(n19366), .A3(n10949), .A4(n18546), .ZN(
        n18595) );
  NAND2_X1 U14305 ( .A1(n10954), .A2(n12854), .ZN(n12864) );
  NAND2_X1 U14306 ( .A1(n18595), .A2(n12864), .ZN(n17733) );
  INV_X1 U14307 ( .A(n18595), .ZN(n18597) );
  NAND2_X1 U14308 ( .A1(n18597), .A2(n18596), .ZN(n17477) );
  NOR2_X1 U14309 ( .A1(n19349), .A2(n18596), .ZN(n10943) );
  OAI21_X1 U14310 ( .B1(n19375), .B2(n19793), .A(n10943), .ZN(n12867) );
  OAI21_X1 U14311 ( .B1(n12884), .B2(n10949), .A(n12867), .ZN(n10952) );
  AOI22_X1 U14312 ( .A1(n19359), .A2(n10944), .B1(n19363), .B2(n19793), .ZN(
        n10951) );
  INV_X1 U14313 ( .A(n12854), .ZN(n19355) );
  NAND2_X1 U14314 ( .A1(n19349), .A2(n18596), .ZN(n10945) );
  AOI21_X1 U14315 ( .B1(n18501), .B2(n10948), .A(n19363), .ZN(n10947) );
  NOR2_X1 U14316 ( .A1(n12854), .A2(n10948), .ZN(n12877) );
  OAI21_X1 U14317 ( .B1(n10949), .B2(n12877), .A(n19349), .ZN(n10950) );
  NAND2_X1 U14318 ( .A1(n10954), .A2(n12882), .ZN(n12888) );
  INV_X1 U14319 ( .A(n12888), .ZN(n10955) );
  NAND2_X1 U14320 ( .A1(n12889), .A2(n10955), .ZN(n17483) );
  XNOR2_X1 U14321 ( .A(n10958), .B(n10957), .ZN(n10963) );
  NAND2_X1 U14322 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19824), .ZN(
        n10960) );
  NAND2_X1 U14323 ( .A1(n10542), .A2(n12859), .ZN(n10964) );
  NAND2_X1 U14324 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18596), .ZN(n10966) );
  AOI211_X4 U14325 ( .C1(n19988), .C2(n19981), .A(n10969), .B(n10966), .ZN(
        n18090) );
  NAND2_X1 U14326 ( .A1(n18054), .A2(n18371), .ZN(n18046) );
  INV_X1 U14327 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18356) );
  NAND2_X1 U14328 ( .A1(n18032), .A2(n18356), .ZN(n18022) );
  INV_X1 U14329 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18003) );
  NAND2_X1 U14330 ( .A1(n18006), .A2(n18003), .ZN(n18000) );
  INV_X1 U14331 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18309) );
  NAND2_X1 U14332 ( .A1(n17986), .A2(n18309), .ZN(n17972) );
  INV_X1 U14333 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17955) );
  NAND2_X1 U14334 ( .A1(n17961), .A2(n17955), .ZN(n17947) );
  INV_X1 U14335 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17925) );
  NAND2_X1 U14336 ( .A1(n17930), .A2(n17925), .ZN(n17924) );
  INV_X1 U14337 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17900) );
  NAND2_X1 U14338 ( .A1(n17906), .A2(n17900), .ZN(n17898) );
  INV_X1 U14339 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n18235) );
  NAND2_X1 U14340 ( .A1(n17886), .A2(n18235), .ZN(n17878) );
  INV_X1 U14341 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n18195) );
  NAND2_X1 U14342 ( .A1(n17861), .A2(n18195), .ZN(n17857) );
  INV_X1 U14343 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18182) );
  NAND2_X1 U14344 ( .A1(n17841), .A2(n18182), .ZN(n17832) );
  INV_X1 U14345 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n18097) );
  NAND2_X1 U14346 ( .A1(n17820), .A2(n18097), .ZN(n17814) );
  INV_X1 U14347 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17792) );
  NAND2_X1 U14348 ( .A1(n17800), .A2(n17792), .ZN(n17791) );
  INV_X1 U14349 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17773) );
  NAND2_X1 U14350 ( .A1(n17781), .A2(n17773), .ZN(n17772) );
  NOR2_X2 U14351 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17772), .ZN(n17758) );
  INV_X1 U14352 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n18098) );
  NAND2_X1 U14353 ( .A1(n17758), .A2(n18098), .ZN(n10971) );
  NAND2_X1 U14354 ( .A1(n18090), .A2(n10971), .ZN(n17752) );
  INV_X1 U14355 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19913) );
  NAND2_X2 U14356 ( .A1(n19928), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19922) );
  AOI211_X1 U14357 ( .C1(n19986), .C2(n19987), .A(n19990), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n10970) );
  INV_X1 U14358 ( .A(n10970), .ZN(n19829) );
  INV_X1 U14359 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19911) );
  INV_X1 U14360 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19906) );
  INV_X1 U14361 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19904) );
  INV_X1 U14362 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19902) );
  INV_X1 U14363 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19898) );
  INV_X1 U14364 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19896) );
  INV_X1 U14365 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19889) );
  INV_X1 U14366 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19885) );
  INV_X1 U14367 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19882) );
  INV_X1 U14368 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19872) );
  NAND3_X1 U14369 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n18040) );
  NOR3_X1 U14370 ( .A1(n19872), .A2(n19869), .A3(n18040), .ZN(n17992) );
  NAND4_X1 U14371 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17992), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n17959) );
  NAND2_X1 U14372 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n17941) );
  NOR3_X1 U14373 ( .A1(n19882), .A2(n17959), .A3(n17941), .ZN(n17933) );
  NAND2_X1 U14374 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17933), .ZN(n17918) );
  NOR2_X1 U14375 ( .A1(n19885), .A2(n17918), .ZN(n17910) );
  NAND2_X1 U14376 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17910), .ZN(n17890) );
  NOR2_X1 U14377 ( .A1(n19889), .A2(n17890), .ZN(n17871) );
  NAND3_X1 U14378 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_17__SCAN_IN), 
        .A3(n17871), .ZN(n17847) );
  NAND2_X1 U14379 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n17836), .ZN(n17818) );
  OR2_X1 U14380 ( .A1(n19902), .A2(n17818), .ZN(n17811) );
  NOR2_X1 U14381 ( .A1(n19904), .A2(n17811), .ZN(n17799) );
  INV_X1 U14382 ( .A(n17799), .ZN(n17787) );
  NOR2_X1 U14383 ( .A1(n19906), .A2(n17787), .ZN(n17793) );
  NAND2_X1 U14384 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17793), .ZN(n17778) );
  NOR2_X1 U14385 ( .A1(n19911), .A2(n17778), .ZN(n10967) );
  NAND2_X1 U14386 ( .A1(n18055), .A2(n10967), .ZN(n17765) );
  NOR2_X1 U14387 ( .A1(n19913), .A2(n17765), .ZN(n17761) );
  NAND3_X1 U14388 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n17761), .ZN(n12972) );
  NOR2_X1 U14389 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n12972), .ZN(n12970) );
  NAND3_X2 U14390 ( .A1(n20002), .A2(n19992), .A3(n20001), .ZN(n19328) );
  INV_X4 U14391 ( .A(n19328), .ZN(n19317) );
  NOR2_X1 U14392 ( .A1(n19841), .A2(n19680), .ZN(n19833) );
  NAND2_X1 U14393 ( .A1(n18091), .A2(n18081), .ZN(n18089) );
  NAND2_X1 U14394 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n10968) );
  AND2_X1 U14395 ( .A1(n18091), .A2(n10967), .ZN(n17777) );
  INV_X1 U14396 ( .A(n18089), .ZN(n17889) );
  AOI21_X1 U14397 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n17777), .A(n17889), 
        .ZN(n17771) );
  AOI21_X1 U14398 ( .B1(n18089), .B2(n10968), .A(n17771), .ZN(n17755) );
  INV_X1 U14399 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19921) );
  INV_X1 U14400 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12938) );
  OAI22_X1 U14401 ( .A1(n17755), .A2(n19921), .B1(n12938), .B2(n18076), .ZN(
        n10974) );
  AOI211_X4 U14402 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18596), .A(n10970), .B(
        n10969), .ZN(n18074) );
  NOR2_X1 U14403 ( .A1(n18080), .A2(n10971), .ZN(n12969) );
  OAI21_X1 U14404 ( .B1(n18074), .B2(n12969), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n10972) );
  OAI21_X1 U14405 ( .B1(n10815), .B2(n10977), .A(n10976), .ZN(P3_U2641) );
  INV_X1 U14406 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16066) );
  AOI22_X1 U14407 ( .A1(n16267), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10983) );
  AND2_X4 U14408 ( .A1(n17324), .A2(n11361), .ZN(n16340) );
  AND2_X4 U14409 ( .A1(n17324), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16266) );
  AOI22_X1 U14410 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U14411 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10981) );
  INV_X1 U14412 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10979) );
  AND2_X4 U14413 ( .A1(n11170), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11179) );
  AOI22_X1 U14414 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U14415 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U14416 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U14417 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16244), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U14418 ( .A1(n16267), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U14419 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U14420 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U14421 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10989) );
  INV_X2 U14422 ( .A(n16352), .ZN(n16282) );
  AOI22_X1 U14423 ( .A1(n16267), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U14424 ( .A1(n16267), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U14425 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11172), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10993) );
  AND2_X1 U14426 ( .A1(n10993), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10996) );
  AOI22_X1 U14427 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U14428 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14429 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14430 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16244), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14431 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U14432 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16244), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U14433 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U14434 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U14435 ( .A1(n16282), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U14436 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U14437 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U14438 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11179), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U14439 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U14440 ( .A1(n16282), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11007) );
  AOI22_X1 U14441 ( .A1(n11180), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U14442 ( .A1(n11798), .A2(n13989), .ZN(n11074) );
  AOI22_X1 U14443 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U14444 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14445 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11172), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U14446 ( .A1(n16282), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11011) );
  NAND4_X1 U14447 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(
        n11016) );
  AOI22_X1 U14448 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U14449 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14450 ( .A1(n16282), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14451 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11017) );
  NAND4_X1 U14452 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11021) );
  AOI22_X1 U14453 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U14454 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16244), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14455 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11028) );
  NAND4_X1 U14456 ( .A1(n11030), .A2(n11029), .A3(n11028), .A4(n11027), .ZN(
        n11031) );
  NAND2_X1 U14457 ( .A1(n11031), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11038) );
  AOI22_X1 U14458 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14459 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11172), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11034) );
  NAND4_X1 U14460 ( .A1(n11035), .A2(n11034), .A3(n11033), .A4(n11032), .ZN(
        n11036) );
  NAND2_X1 U14461 ( .A1(n11036), .A2(n11015), .ZN(n11037) );
  AOI22_X1 U14462 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U14463 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n16340), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11041) );
  AOI22_X1 U14464 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9771), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U14465 ( .A1(n16267), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U14466 ( .A1(n16267), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16378), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11045) );
  AOI22_X1 U14467 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11172), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U14468 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11043) );
  INV_X1 U14469 ( .A(n11060), .ZN(n11047) );
  INV_X1 U14470 ( .A(n20156), .ZN(n11058) );
  AOI22_X1 U14471 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11051) );
  AOI22_X1 U14472 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U14473 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9752), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U14474 ( .A1(n16282), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11048) );
  NAND4_X1 U14475 ( .A1(n11051), .A2(n11050), .A3(n11049), .A4(n11048), .ZN(
        n11057) );
  AOI22_X1 U14476 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14477 ( .A1(n11179), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11180), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14478 ( .A1(n9768), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9752), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14479 ( .A1(n16282), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11052) );
  NAND4_X1 U14480 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11056) );
  MUX2_X2 U14481 ( .A(n11057), .B(n11056), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11429) );
  NAND2_X1 U14482 ( .A1(n11684), .A2(n13974), .ZN(n14187) );
  NAND2_X1 U14483 ( .A1(n14191), .A2(n11073), .ZN(n11059) );
  NAND2_X1 U14484 ( .A1(n11076), .A2(n20156), .ZN(n11063) );
  NAND2_X1 U14485 ( .A1(n11073), .A2(n9748), .ZN(n11061) );
  NAND2_X1 U14486 ( .A1(n11061), .A2(n11060), .ZN(n11062) );
  NAND4_X1 U14487 ( .A1(n9748), .A2(n11429), .A3(n11025), .A4(n20181), .ZN(
        n11064) );
  AND2_X2 U14488 ( .A1(n11065), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11118) );
  INV_X1 U14489 ( .A(n11068), .ZN(n11066) );
  NAND2_X1 U14490 ( .A1(n11108), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11071) );
  NAND2_X1 U14491 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11070) );
  INV_X1 U14492 ( .A(n11093), .ZN(n11092) );
  NAND2_X1 U14493 ( .A1(n11076), .A2(n11434), .ZN(n11683) );
  INV_X1 U14494 ( .A(n11077), .ZN(n11081) );
  NAND2_X2 U14495 ( .A1(n11080), .A2(n11081), .ZN(n17352) );
  NAND3_X1 U14496 ( .A1(n17352), .A2(n11078), .A3(n11163), .ZN(n11083) );
  NAND2_X1 U14497 ( .A1(n11676), .A2(n11084), .ZN(n11085) );
  NAND2_X1 U14498 ( .A1(n11086), .A2(n11085), .ZN(n11095) );
  NAND2_X1 U14499 ( .A1(n11095), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11091) );
  NAND2_X1 U14500 ( .A1(n11087), .A2(n11426), .ZN(n11675) );
  INV_X1 U14501 ( .A(n11675), .ZN(n11088) );
  NAND2_X1 U14502 ( .A1(n11088), .A2(n9835), .ZN(n11980) );
  AOI21_X1 U14503 ( .B1(n11980), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11089), 
        .ZN(n11090) );
  BUF_X2 U14504 ( .A(n11095), .Z(n11115) );
  NAND2_X1 U14505 ( .A1(n11115), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11099) );
  INV_X1 U14506 ( .A(n17285), .ZN(n11981) );
  NAND2_X1 U14507 ( .A1(n17366), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11096) );
  NAND2_X1 U14508 ( .A1(n11898), .A2(n11096), .ZN(n11097) );
  INV_X1 U14509 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n16008) );
  INV_X1 U14510 ( .A(n17366), .ZN(n11101) );
  NAND2_X1 U14511 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11100) );
  AND2_X1 U14512 ( .A1(n11101), .A2(n11100), .ZN(n11103) );
  NAND2_X1 U14513 ( .A1(n11108), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11102) );
  OAI211_X1 U14514 ( .C1(n11968), .C2(n16008), .A(n11103), .B(n11102), .ZN(
        n11104) );
  AOI21_X1 U14515 ( .B1(n11118), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11104), .ZN(n11106) );
  INV_X1 U14516 ( .A(n11115), .ZN(n11105) );
  OAI21_X1 U14517 ( .B1(n20821), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n17365), 
        .ZN(n11107) );
  NAND2_X1 U14518 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11110) );
  NAND2_X1 U14519 ( .A1(n11108), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11109) );
  NAND2_X1 U14520 ( .A1(n11115), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11117) );
  NAND2_X1 U14521 ( .A1(n17366), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11116) );
  NAND2_X1 U14522 ( .A1(n11117), .A2(n11116), .ZN(n11121) );
  INV_X4 U14523 ( .A(n11898), .ZN(n12705) );
  AOI22_X1 U14524 ( .A1(n12705), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11120) );
  INV_X1 U14525 ( .A(n11968), .ZN(n11977) );
  NAND2_X1 U14526 ( .A1(n11977), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11119) );
  XNOR2_X2 U14527 ( .A(n14312), .B(n11122), .ZN(n14199) );
  INV_X1 U14528 ( .A(n14199), .ZN(n11125) );
  XNOR2_X2 U14529 ( .A(n11124), .B(n11123), .ZN(n14171) );
  INV_X1 U14530 ( .A(n11126), .ZN(n11131) );
  INV_X1 U14531 ( .A(n11127), .ZN(n11130) );
  INV_X1 U14532 ( .A(n11128), .ZN(n11129) );
  AND2_X2 U14533 ( .A1(n11153), .A2(n11146), .ZN(n20517) );
  INV_X1 U14534 ( .A(n20517), .ZN(n11132) );
  AND2_X2 U14535 ( .A1(n11154), .A2(n11146), .ZN(n11271) );
  INV_X1 U14536 ( .A(n11271), .ZN(n20658) );
  INV_X1 U14537 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16051) );
  OAI22_X1 U14538 ( .A1(n16066), .A2(n11132), .B1(n20658), .B2(n16051), .ZN(
        n11141) );
  INV_X1 U14539 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16065) );
  AND2_X2 U14540 ( .A1(n14199), .A2(n17320), .ZN(n11148) );
  INV_X1 U14541 ( .A(n11134), .ZN(n11136) );
  NAND2_X1 U14542 ( .A1(n11148), .A2(n11147), .ZN(n20195) );
  NAND2_X1 U14543 ( .A1(n11136), .A2(n11135), .ZN(n11137) );
  AND2_X4 U14544 ( .A1(n11126), .A2(n11137), .ZN(n15994) );
  INV_X1 U14545 ( .A(n15994), .ZN(n11138) );
  INV_X1 U14546 ( .A(n11265), .ZN(n11139) );
  INV_X1 U14547 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16061) );
  OAI22_X1 U14548 ( .A1(n16065), .A2(n20195), .B1(n11139), .B2(n16061), .ZN(
        n11140) );
  NOR2_X1 U14549 ( .A1(n11141), .A2(n11140), .ZN(n11162) );
  AND2_X2 U14550 ( .A1(n11148), .A2(n11155), .ZN(n20141) );
  INV_X1 U14551 ( .A(n14171), .ZN(n15986) );
  AOI22_X1 U14552 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20141), .B1(
        n20331), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11142) );
  INV_X1 U14553 ( .A(n11142), .ZN(n11145) );
  INV_X1 U14554 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11143) );
  NAND2_X1 U14555 ( .A1(n11148), .A2(n11146), .ZN(n11213) );
  INV_X1 U14556 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16052) );
  NOR2_X1 U14557 ( .A1(n11145), .A2(n11144), .ZN(n11161) );
  INV_X2 U14558 ( .A(n20454), .ZN(n20451) );
  INV_X1 U14559 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16064) );
  NAND2_X1 U14560 ( .A1(n11148), .A2(n11152), .ZN(n20227) );
  INV_X1 U14561 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11149) );
  INV_X1 U14562 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11513) );
  INV_X1 U14563 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16060) );
  INV_X1 U14564 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U14565 ( .A1(n20299), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11156) );
  OAI211_X1 U14566 ( .C1(n11515), .C2(n11214), .A(n11156), .B(n20146), .ZN(
        n11157) );
  INV_X1 U14567 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11484) );
  INV_X4 U14568 ( .A(n11164), .ZN(n16374) );
  INV_X1 U14569 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16030) );
  OAI22_X1 U14570 ( .A1(n9764), .A2(n11484), .B1(n16225), .B2(n16030), .ZN(
        n11167) );
  INV_X1 U14571 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11165) );
  INV_X1 U14572 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16028) );
  OAI22_X1 U14573 ( .A1(n16229), .A2(n11165), .B1(n16219), .B2(n16028), .ZN(
        n11166) );
  NOR2_X1 U14574 ( .A1(n11167), .A2(n11166), .ZN(n11185) );
  AND2_X1 U14575 ( .A1(n21769), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11168) );
  AND2_X2 U14576 ( .A1(n16184), .A2(n11168), .ZN(n16203) );
  AND2_X2 U14577 ( .A1(n16184), .A2(n11169), .ZN(n16204) );
  AOI22_X1 U14578 ( .A1(n16203), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11176) );
  AND2_X2 U14579 ( .A1(n11170), .A2(n16184), .ZN(n16205) );
  INV_X1 U14580 ( .A(n11171), .ZN(n17286) );
  INV_X1 U14581 ( .A(n17286), .ZN(n14545) );
  AND2_X2 U14582 ( .A1(n16184), .A2(n14545), .ZN(n16202) );
  AOI22_X1 U14583 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11175) );
  NAND2_X1 U14584 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11174) );
  AND2_X2 U14585 ( .A1(n17289), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16206) );
  NAND2_X1 U14586 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11173) );
  NAND4_X1 U14587 ( .A1(n11176), .A2(n11175), .A3(n11174), .A4(n11173), .ZN(
        n11178) );
  INV_X2 U14588 ( .A(n11305), .ZN(n16153) );
  INV_X1 U14589 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11485) );
  INV_X1 U14590 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16029) );
  OAI22_X1 U14591 ( .A1(n16153), .A2(n11485), .B1(n11252), .B2(n16029), .ZN(
        n11177) );
  NOR2_X1 U14592 ( .A1(n11178), .A2(n11177), .ZN(n11184) );
  INV_X1 U14593 ( .A(n11179), .ZN(n16182) );
  INV_X1 U14594 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16027) );
  NAND2_X2 U14595 ( .A1(n16377), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16109) );
  INV_X1 U14596 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16038) );
  OAI22_X1 U14597 ( .A1(n16217), .A2(n16027), .B1(n16109), .B2(n16038), .ZN(
        n11182) );
  INV_X1 U14598 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16044) );
  INV_X1 U14600 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16042) );
  OAI22_X1 U14601 ( .A1(n16221), .A2(n16044), .B1(n16215), .B2(n16042), .ZN(
        n11181) );
  NOR2_X1 U14602 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  INV_X1 U14603 ( .A(n11436), .ZN(n11186) );
  AND2_X1 U14604 ( .A1(n20854), .A2(n11186), .ZN(n11238) );
  AOI22_X1 U14605 ( .A1(n11329), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11199) );
  INV_X1 U14606 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16050) );
  OAI22_X1 U14607 ( .A1(n16217), .A2(n16050), .B1(n16215), .B2(n16064), .ZN(
        n11188) );
  INV_X1 U14608 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n21861) );
  OAI22_X1 U14609 ( .A1(n16109), .A2(n16061), .B1(n11324), .B2(n21861), .ZN(
        n11187) );
  NOR2_X1 U14610 ( .A1(n11188), .A2(n11187), .ZN(n11198) );
  AOI22_X1 U14611 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14612 ( .A1(n16203), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11192) );
  NAND2_X1 U14613 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11191) );
  NAND2_X1 U14614 ( .A1(n11524), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11190) );
  NAND4_X1 U14615 ( .A1(n11193), .A2(n11192), .A3(n11191), .A4(n11190), .ZN(
        n11195) );
  OAI22_X1 U14616 ( .A1(n16153), .A2(n11515), .B1(n11252), .B2(n16052), .ZN(
        n11194) );
  NOR2_X1 U14617 ( .A1(n11195), .A2(n11194), .ZN(n11197) );
  AOI22_X1 U14618 ( .A1(n11328), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11200), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11196) );
  NAND2_X1 U14619 ( .A1(n11238), .A2(n11445), .ZN(n11244) );
  INV_X1 U14620 ( .A(n16217), .ZN(n11249) );
  NAND2_X1 U14621 ( .A1(n11249), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11201) );
  INV_X1 U14622 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16096) );
  INV_X1 U14623 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16108) );
  OAI22_X1 U14624 ( .A1(n16225), .A2(n16096), .B1(n16215), .B2(n16108), .ZN(
        n11203) );
  INV_X1 U14625 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16105) );
  OAI22_X1 U14626 ( .A1(n16109), .A2(n16105), .B1(n11324), .B2(n16110), .ZN(
        n11202) );
  AOI22_X1 U14627 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n16202), .B1(
        n16203), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14628 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n16205), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U14629 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11205) );
  NAND2_X1 U14630 ( .A1(n11524), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11204) );
  NAND4_X1 U14631 ( .A1(n11207), .A2(n11206), .A3(n11205), .A4(n11204), .ZN(
        n11209) );
  INV_X1 U14632 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11536) );
  INV_X1 U14633 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16097) );
  OAI22_X1 U14634 ( .A1(n11536), .A2(n16153), .B1(n11252), .B2(n16097), .ZN(
        n11208) );
  NOR2_X1 U14635 ( .A1(n11209), .A2(n11208), .ZN(n11210) );
  NAND2_X1 U14636 ( .A1(n11244), .A2(n11454), .ZN(n11211) );
  INV_X2 U14637 ( .A(n20227), .ZN(n20221) );
  INV_X2 U14638 ( .A(n11213), .ZN(n20259) );
  AOI22_X1 U14639 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20221), .B1(
        n20259), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11218) );
  INV_X1 U14640 ( .A(n11214), .ZN(n20551) );
  AOI22_X1 U14641 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20551), .B1(
        n20517), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14642 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n11271), .B1(
        n11266), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14643 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20190), .B1(
        n20141), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14644 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n16202), .B1(
        n16203), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14645 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n16205), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11226) );
  NAND2_X1 U14646 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11225) );
  NAND2_X1 U14647 ( .A1(n11524), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11224) );
  NAND4_X1 U14648 ( .A1(n11227), .A2(n11226), .A3(n11225), .A4(n11224), .ZN(
        n11229) );
  INV_X1 U14649 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11556) );
  INV_X1 U14650 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16074) );
  OAI22_X1 U14651 ( .A1(n11556), .A2(n16153), .B1(n11252), .B2(n16074), .ZN(
        n11228) );
  NOR2_X1 U14652 ( .A1(n11229), .A2(n11228), .ZN(n11236) );
  INV_X1 U14653 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11230) );
  INV_X1 U14654 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16085) );
  OAI22_X1 U14655 ( .A1(n16229), .A2(n11230), .B1(n16215), .B2(n16085), .ZN(
        n11232) );
  INV_X1 U14656 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16082) );
  OAI22_X1 U14657 ( .A1(n16109), .A2(n16082), .B1(n11324), .B2(n16086), .ZN(
        n11231) );
  NOR2_X1 U14658 ( .A1(n11232), .A2(n11231), .ZN(n11235) );
  AOI22_X1 U14659 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11249), .B1(
        n11328), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14660 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11200), .B1(
        n11329), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11233) );
  NAND4_X1 U14661 ( .A1(n11236), .A2(n11235), .A3(n11234), .A4(n11233), .ZN(
        n11463) );
  OR2_X1 U14662 ( .A1(n20146), .A2(n11463), .ZN(n11237) );
  INV_X1 U14663 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14524) );
  INV_X1 U14664 ( .A(n11238), .ZN(n13881) );
  NAND2_X1 U14665 ( .A1(n13881), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13880) );
  INV_X1 U14666 ( .A(n11445), .ZN(n11239) );
  XNOR2_X1 U14667 ( .A(n11239), .B(n11436), .ZN(n11240) );
  NOR2_X1 U14668 ( .A1(n13880), .A2(n11240), .ZN(n11242) );
  INV_X1 U14669 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21897) );
  AND2_X1 U14670 ( .A1(n13880), .A2(n11240), .ZN(n11241) );
  OR2_X1 U14671 ( .A1(n11242), .A2(n11241), .ZN(n13999) );
  NOR2_X1 U14672 ( .A1(n21897), .A2(n13999), .ZN(n13998) );
  NOR2_X1 U14673 ( .A1(n11242), .A2(n13998), .ZN(n11245) );
  XNOR2_X1 U14674 ( .A(n14524), .B(n11245), .ZN(n14520) );
  XNOR2_X1 U14675 ( .A(n11244), .B(n11243), .ZN(n14521) );
  OAI21_X1 U14676 ( .B1(n14520), .B2(n14521), .A(n10817), .ZN(n11246) );
  XNOR2_X1 U14677 ( .A(n11246), .B(n17253), .ZN(n16936) );
  NAND2_X1 U14678 ( .A1(n11246), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11247) );
  INV_X1 U14679 ( .A(n16109), .ZN(n11248) );
  AOI22_X1 U14680 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11249), .B1(
        n11248), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11251) );
  AOI22_X1 U14681 ( .A1(n11494), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11524), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11250) );
  INV_X1 U14682 ( .A(n11252), .ZN(n11253) );
  AOI22_X1 U14683 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11305), .B1(
        n11253), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14684 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n16203), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11259) );
  INV_X1 U14685 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16133) );
  NAND2_X1 U14686 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11255) );
  NAND2_X1 U14687 ( .A1(n16202), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11254) );
  OAI211_X1 U14688 ( .C1(n11324), .C2(n16133), .A(n11255), .B(n11254), .ZN(
        n11256) );
  INV_X1 U14689 ( .A(n11256), .ZN(n11258) );
  NAND2_X1 U14690 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11257) );
  INV_X1 U14691 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U14692 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20221), .B1(
        n20141), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14693 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20359), .B1(
        n20259), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14694 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20390), .B1(
        n20551), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U14695 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20299), .B1(
        n20190), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14696 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n11271), .B1(
        n20517), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11272) );
  INV_X1 U14697 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16144) );
  INV_X1 U14698 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11274) );
  OAI22_X1 U14699 ( .A1(n16225), .A2(n16144), .B1(n16229), .B2(n11274), .ZN(
        n11276) );
  INV_X1 U14700 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16159) );
  INV_X1 U14701 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11592) );
  OAI22_X1 U14702 ( .A1(n16221), .A2(n16159), .B1(n16228), .B2(n11592), .ZN(
        n11275) );
  NOR2_X1 U14703 ( .A1(n11276), .A2(n11275), .ZN(n11287) );
  AOI22_X1 U14704 ( .A1(n16203), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14705 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11279) );
  NAND2_X1 U14706 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11278) );
  NAND2_X1 U14707 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11277) );
  NAND4_X1 U14708 ( .A1(n11280), .A2(n11279), .A3(n11278), .A4(n11277), .ZN(
        n11282) );
  INV_X1 U14709 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11594) );
  INV_X1 U14710 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16143) );
  OAI22_X1 U14711 ( .A1(n16153), .A2(n11594), .B1(n11252), .B2(n16143), .ZN(
        n11281) );
  NOR2_X1 U14712 ( .A1(n11282), .A2(n11281), .ZN(n11286) );
  INV_X1 U14713 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16141) );
  INV_X1 U14714 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16152) );
  OAI22_X1 U14715 ( .A1(n16217), .A2(n16141), .B1(n16109), .B2(n16152), .ZN(
        n11284) );
  INV_X1 U14716 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16157) );
  INV_X1 U14717 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16142) );
  OAI22_X1 U14718 ( .A1(n16215), .A2(n16157), .B1(n16219), .B2(n16142), .ZN(
        n11283) );
  NOR2_X1 U14719 ( .A1(n11284), .A2(n11283), .ZN(n11285) );
  NAND2_X1 U14720 ( .A1(n11730), .A2(n20854), .ZN(n11288) );
  INV_X1 U14721 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U14722 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20190), .B1(
        n20141), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14723 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20221), .B1(
        n20259), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11293) );
  AOI22_X1 U14724 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20299), .B1(
        n20331), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14725 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20359), .B1(
        n20390), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14726 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20454), .B1(
        n20424), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11298) );
  AOI22_X1 U14727 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20487), .B1(
        n20517), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U14728 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20616), .B1(
        n11271), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11295) );
  INV_X1 U14729 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16341) );
  INV_X1 U14730 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17312) );
  OAI22_X1 U14731 ( .A1(n16341), .A2(n16109), .B1(n16225), .B2(n17312), .ZN(
        n11300) );
  INV_X1 U14732 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11613) );
  INV_X1 U14733 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16355) );
  OAI22_X1 U14734 ( .A1(n11613), .A2(n16228), .B1(n16229), .B2(n16355), .ZN(
        n11299) );
  NOR2_X1 U14735 ( .A1(n11300), .A2(n11299), .ZN(n11312) );
  AOI22_X1 U14736 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n16202), .B1(
        n16203), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14737 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n16205), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U14738 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11302) );
  NAND2_X1 U14739 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11301) );
  NAND4_X1 U14740 ( .A1(n11304), .A2(n11303), .A3(n11302), .A4(n11301), .ZN(
        n11307) );
  INV_X1 U14741 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16342) );
  INV_X1 U14742 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11612) );
  OAI22_X1 U14743 ( .A1(n16342), .A2(n11252), .B1(n16153), .B2(n11612), .ZN(
        n11306) );
  NOR2_X1 U14744 ( .A1(n11307), .A2(n11306), .ZN(n11311) );
  INV_X1 U14745 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16351) );
  INV_X1 U14746 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16176) );
  OAI22_X1 U14747 ( .A1(n16351), .A2(n16217), .B1(n16221), .B2(n16176), .ZN(
        n11309) );
  INV_X1 U14748 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16339) );
  INV_X1 U14749 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16165) );
  OAI22_X1 U14750 ( .A1(n16339), .A2(n16215), .B1(n16219), .B2(n16165), .ZN(
        n11308) );
  NOR2_X1 U14751 ( .A1(n11309), .A2(n11308), .ZN(n11310) );
  NAND2_X1 U14752 ( .A1(n11762), .A2(n20854), .ZN(n11313) );
  AOI22_X1 U14753 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n16203), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14754 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n16205), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11320) );
  NAND2_X1 U14755 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11319) );
  NAND2_X1 U14756 ( .A1(n11524), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11318) );
  NAND4_X1 U14757 ( .A1(n11321), .A2(n11320), .A3(n11319), .A4(n11318), .ZN(
        n11323) );
  INV_X1 U14758 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11631) );
  INV_X1 U14759 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16227) );
  OAI22_X1 U14760 ( .A1(n11631), .A2(n16153), .B1(n11252), .B2(n16227), .ZN(
        n11322) );
  NOR2_X1 U14761 ( .A1(n11323), .A2(n11322), .ZN(n11336) );
  INV_X1 U14762 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n21759) );
  INV_X1 U14763 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16216) );
  OAI22_X1 U14764 ( .A1(n16109), .A2(n21759), .B1(n16215), .B2(n16216), .ZN(
        n11326) );
  INV_X1 U14765 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16230) );
  OAI22_X1 U14766 ( .A1(n16217), .A2(n16230), .B1(n11324), .B2(n16494), .ZN(
        n11325) );
  NOR2_X1 U14767 ( .A1(n11326), .A2(n11325), .ZN(n11335) );
  NAND2_X1 U14768 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U14769 ( .A1(n11328), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11332) );
  NAND2_X1 U14770 ( .A1(n11200), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11331) );
  NAND2_X1 U14771 ( .A1(n11329), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11330) );
  INV_X1 U14772 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17190) );
  NAND2_X1 U14773 ( .A1(n16867), .A2(n17190), .ZN(n11338) );
  INV_X1 U14774 ( .A(n16867), .ZN(n16868) );
  INV_X1 U14775 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17191) );
  AND4_X1 U14776 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11345) );
  NAND3_X1 U14777 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12959) );
  INV_X1 U14778 ( .A(n12959), .ZN(n11343) );
  AND4_X1 U14779 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(n11343), .ZN(n11344) );
  NAND3_X1 U14780 ( .A1(n11345), .A2(n11344), .A3(n12957), .ZN(n17045) );
  NAND3_X1 U14781 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11346) );
  NOR2_X1 U14782 ( .A1(n17045), .A2(n11346), .ZN(n11347) );
  AND2_X1 U14783 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16943) );
  INV_X1 U14784 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16974) );
  INV_X1 U14785 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16645) );
  MUX2_X1 U14786 ( .A(n20831), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11365) );
  NAND2_X1 U14787 ( .A1(n17269), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11363) );
  NAND2_X1 U14788 ( .A1(n11365), .A2(n11364), .ZN(n11350) );
  NAND2_X1 U14789 ( .A1(n20831), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11349) );
  NAND2_X1 U14790 ( .A1(n11350), .A2(n11349), .ZN(n11360) );
  XNOR2_X1 U14791 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11359) );
  NAND2_X1 U14792 ( .A1(n11360), .A2(n11359), .ZN(n11352) );
  NAND2_X1 U14793 ( .A1(n20821), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11351) );
  NAND2_X1 U14794 ( .A1(n11352), .A2(n11351), .ZN(n11356) );
  XNOR2_X1 U14795 ( .A(n11015), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11353) );
  XNOR2_X1 U14796 ( .A(n11356), .B(n11353), .ZN(n11399) );
  MUX2_X1 U14797 ( .A(n11463), .B(n11399), .S(n11358), .Z(n11726) );
  INV_X1 U14798 ( .A(n11353), .ZN(n11355) );
  NOR2_X1 U14799 ( .A1(n11015), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11354) );
  AOI21_X1 U14800 ( .B1(n11356), .B2(n11355), .A(n11354), .ZN(n11375) );
  INV_X1 U14801 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17534) );
  NOR2_X1 U14802 ( .A1(n17534), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11357) );
  NAND2_X1 U14803 ( .A1(n11375), .A2(n11357), .ZN(n11400) );
  AND2_X1 U14804 ( .A1(n11726), .A2(n11729), .ZN(n11391) );
  XNOR2_X1 U14805 ( .A(n11360), .B(n11359), .ZN(n11388) );
  INV_X1 U14806 ( .A(n11388), .ZN(n11398) );
  NAND2_X1 U14807 ( .A1(n13974), .A2(n11398), .ZN(n11370) );
  INV_X1 U14808 ( .A(n11365), .ZN(n11390) );
  NAND2_X1 U14809 ( .A1(n11361), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11362) );
  NAND2_X1 U14810 ( .A1(n11363), .A2(n11362), .ZN(n11410) );
  OAI21_X1 U14811 ( .B1(n11390), .B2(n11410), .A(n11387), .ZN(n11369) );
  NAND2_X1 U14812 ( .A1(n20854), .A2(n11410), .ZN(n11367) );
  XNOR2_X1 U14813 ( .A(n11365), .B(n11364), .ZN(n11401) );
  INV_X1 U14814 ( .A(n11401), .ZN(n11366) );
  NAND3_X1 U14815 ( .A1(n11367), .A2(n11366), .A3(n11686), .ZN(n11368) );
  AND3_X1 U14816 ( .A1(n11370), .A2(n11369), .A3(n11368), .ZN(n11373) );
  NOR2_X1 U14817 ( .A1(n11084), .A2(n20854), .ZN(n11371) );
  MUX2_X1 U14818 ( .A(n11371), .B(n11387), .S(n11398), .Z(n11372) );
  OAI21_X1 U14819 ( .B1(n11373), .B2(n11372), .A(n11399), .ZN(n11374) );
  OAI21_X1 U14820 ( .B1(n11391), .B2(n11387), .A(n11374), .ZN(n11381) );
  INV_X1 U14821 ( .A(n11375), .ZN(n11378) );
  NAND2_X1 U14822 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17362), .ZN(
        n11377) );
  NOR2_X1 U14823 ( .A1(n17362), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11376) );
  INV_X1 U14824 ( .A(n11400), .ZN(n11379) );
  AOI21_X1 U14825 ( .B1(n11387), .B2(n11379), .A(n10286), .ZN(n11380) );
  NAND3_X1 U14826 ( .A1(n11381), .A2(n11402), .A3(n11380), .ZN(n11385) );
  INV_X1 U14827 ( .A(n11402), .ZN(n11383) );
  NOR2_X1 U14828 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11382) );
  AOI21_X1 U14829 ( .B1(n11383), .B2(n11084), .A(n11382), .ZN(n11384) );
  AOI21_X1 U14830 ( .B1(n17345), .B2(n11686), .A(n9748), .ZN(n11424) );
  INV_X1 U14831 ( .A(n17345), .ZN(n11386) );
  NAND2_X1 U14832 ( .A1(n11386), .A2(n20146), .ZN(n13876) );
  MUX2_X1 U14833 ( .A(n11436), .B(n11410), .S(n11358), .Z(n11735) );
  OAI21_X1 U14834 ( .B1(n11735), .B2(n11390), .A(n11722), .ZN(n11392) );
  NAND2_X1 U14835 ( .A1(n11392), .A2(n11391), .ZN(n11393) );
  AND2_X1 U14836 ( .A1(n11393), .A2(n11402), .ZN(n20841) );
  NAND2_X1 U14837 ( .A1(n20851), .A2(n20854), .ZN(n11404) );
  NOR2_X1 U14838 ( .A1(n17352), .A2(n11404), .ZN(n11433) );
  NAND2_X1 U14839 ( .A1(n20841), .A2(n11433), .ZN(n11422) );
  NAND2_X1 U14840 ( .A1(n20854), .A2(n20161), .ZN(n11395) );
  NAND2_X1 U14841 ( .A1(n11395), .A2(n11686), .ZN(n11396) );
  NAND2_X1 U14842 ( .A1(n11396), .A2(n20156), .ZN(n11397) );
  OAI21_X1 U14843 ( .B1(n11394), .B2(n11397), .A(n11078), .ZN(n11409) );
  NAND3_X1 U14844 ( .A1(n11400), .A2(n11399), .A3(n11398), .ZN(n11411) );
  NOR2_X1 U14845 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20725) );
  INV_X1 U14846 ( .A(n20725), .ZN(n20011) );
  NAND3_X1 U14847 ( .A1(n20728), .A2(n20778), .A3(n20011), .ZN(n13877) );
  NAND2_X1 U14848 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20850) );
  NOR2_X1 U14849 ( .A1(n13877), .A2(n20844), .ZN(n13809) );
  NAND3_X1 U14850 ( .A1(n11417), .A2(n13963), .A3(n13809), .ZN(n11407) );
  INV_X1 U14851 ( .A(n11404), .ZN(n11405) );
  NAND2_X1 U14852 ( .A1(n11406), .A2(n11405), .ZN(n11691) );
  AND2_X1 U14853 ( .A1(n11407), .A2(n11691), .ZN(n11408) );
  NOR2_X1 U14854 ( .A1(n11411), .A2(n11410), .ZN(n11412) );
  NOR2_X1 U14855 ( .A1(n17348), .A2(n11412), .ZN(n11415) );
  INV_X1 U14856 ( .A(n17289), .ZN(n11413) );
  AND2_X1 U14857 ( .A1(n11413), .A2(n17362), .ZN(n13972) );
  NAND2_X1 U14858 ( .A1(n16109), .A2(n13972), .ZN(n11414) );
  INV_X1 U14859 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n17273) );
  NAND2_X1 U14860 ( .A1(n11414), .A2(n17273), .ZN(n17271) );
  MUX2_X1 U14861 ( .A(n11415), .B(n17271), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20835) );
  NOR2_X1 U14862 ( .A1(n17352), .A2(n20854), .ZN(n11416) );
  NAND2_X1 U14863 ( .A1(n20835), .A2(n11416), .ZN(n11421) );
  MUX2_X1 U14864 ( .A(n11417), .B(n11429), .S(n20854), .Z(n11419) );
  NOR2_X1 U14865 ( .A1(n17348), .A2(n20844), .ZN(n11418) );
  NAND2_X1 U14866 ( .A1(n11419), .A2(n11418), .ZN(n11420) );
  NAND4_X1 U14867 ( .A1(n11422), .A2(n13959), .A3(n11421), .A4(n11420), .ZN(
        n11423) );
  AOI21_X1 U14868 ( .B1(n11424), .B2(n13876), .A(n11423), .ZN(n11431) );
  INV_X1 U14869 ( .A(n13809), .ZN(n11425) );
  OR2_X1 U14870 ( .A1(n13876), .A2(n11425), .ZN(n11428) );
  INV_X1 U14871 ( .A(n11426), .ZN(n11427) );
  NAND2_X1 U14872 ( .A1(n11428), .A2(n11427), .ZN(n13961) );
  NAND2_X1 U14873 ( .A1(n13961), .A2(n11429), .ZN(n11430) );
  NAND2_X1 U14874 ( .A1(n11431), .A2(n11430), .ZN(n11432) );
  INV_X1 U14875 ( .A(n11433), .ZN(n20840) );
  AND2_X1 U14876 ( .A1(n11434), .A2(n20814), .ZN(n11437) );
  NAND2_X1 U14877 ( .A1(n11437), .A2(n11025), .ZN(n11479) );
  MUX2_X1 U14878 ( .A(n20181), .B(n17269), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11435) );
  NOR2_X1 U14879 ( .A1(n11434), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11455) );
  NAND2_X1 U14880 ( .A1(n11455), .A2(n14194), .ZN(n11453) );
  OAI211_X2 U14881 ( .C1(n11436), .C2(n11479), .A(n11435), .B(n11453), .ZN(
        n14042) );
  NAND2_X1 U14882 ( .A1(n11442), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11441) );
  INV_X1 U14883 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14020) );
  NAND2_X1 U14884 ( .A1(n9749), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11438) );
  OAI211_X1 U14885 ( .C1(n20854), .C2(n14020), .A(n11438), .B(n20814), .ZN(
        n11439) );
  INV_X1 U14886 ( .A(n11439), .ZN(n11440) );
  NAND2_X1 U14887 ( .A1(n11441), .A2(n11440), .ZN(n14041) );
  NAND2_X1 U14888 ( .A1(n14042), .A2(n14041), .ZN(n14043) );
  AOI22_X1 U14889 ( .A1(n11455), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n11456), .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U14890 ( .A1(n11442), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11443) );
  NAND2_X1 U14891 ( .A1(n11444), .A2(n11443), .ZN(n11449) );
  XNOR2_X1 U14892 ( .A(n14043), .B(n11449), .ZN(n14027) );
  NAND2_X1 U14893 ( .A1(n11445), .A2(n11025), .ZN(n11724) );
  INV_X1 U14894 ( .A(n11724), .ZN(n11447) );
  NOR2_X1 U14895 ( .A1(n14194), .A2(n9749), .ZN(n11446) );
  AOI21_X1 U14896 ( .B1(n11447), .B2(n20854), .A(n11446), .ZN(n11448) );
  MUX2_X2 U14897 ( .A(n20831), .B(n11448), .S(n20814), .Z(n14026) );
  NAND2_X1 U14898 ( .A1(n14027), .A2(n14026), .ZN(n14029) );
  INV_X1 U14899 ( .A(n11449), .ZN(n11450) );
  NAND2_X1 U14900 ( .A1(n14043), .A2(n11450), .ZN(n11451) );
  NAND2_X1 U14901 ( .A1(n14029), .A2(n11451), .ZN(n11461) );
  NAND2_X1 U14902 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11452) );
  OAI211_X1 U14903 ( .C1(n11479), .C2(n11454), .A(n11453), .B(n11452), .ZN(
        n11459) );
  XNOR2_X1 U14904 ( .A(n11461), .B(n11459), .ZN(n14322) );
  AOI22_X1 U14905 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n11456), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n11458) );
  NAND2_X1 U14906 ( .A1(n11647), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11457) );
  AND2_X1 U14907 ( .A1(n11458), .A2(n11457), .ZN(n14321) );
  INV_X1 U14908 ( .A(n11459), .ZN(n11460) );
  NAND2_X1 U14909 ( .A1(n11461), .A2(n11460), .ZN(n11462) );
  AOI22_X1 U14910 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11467) );
  NAND2_X1 U14911 ( .A1(n11647), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U14912 ( .A1(n11637), .A2(n11463), .ZN(n11465) );
  NAND2_X1 U14913 ( .A1(n11670), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11464) );
  INV_X1 U14914 ( .A(n15958), .ZN(n11468) );
  AOI22_X1 U14915 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n11456), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11472) );
  NAND2_X1 U14916 ( .A1(n11647), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U14917 ( .A1(n11637), .A2(n11469), .ZN(n11470) );
  INV_X1 U14918 ( .A(n15943), .ZN(n11473) );
  AOI22_X1 U14919 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n11456), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11478) );
  NAND2_X1 U14920 ( .A1(n11647), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11477) );
  INV_X1 U14921 ( .A(n11730), .ZN(n11475) );
  NAND2_X1 U14922 ( .A1(n11637), .A2(n11475), .ZN(n11476) );
  AOI22_X1 U14923 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n11456), .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14924 ( .A1(n11647), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14925 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n11456), .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n11483) );
  NAND2_X1 U14926 ( .A1(n11647), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11482) );
  NAND2_X1 U14927 ( .A1(n11483), .A2(n11482), .ZN(n14263) );
  INV_X1 U14928 ( .A(n14261), .ZN(n11504) );
  AOI22_X1 U14929 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n11502) );
  OAI22_X1 U14930 ( .A1(n16225), .A2(n16038), .B1(n16109), .B2(n16028), .ZN(
        n11487) );
  OAI22_X1 U14931 ( .A1(n16221), .A2(n11485), .B1(n16229), .B2(n11484), .ZN(
        n11486) );
  NOR2_X1 U14932 ( .A1(n11487), .A2(n11486), .ZN(n11499) );
  AOI22_X1 U14933 ( .A1(n16203), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14934 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11490) );
  NAND2_X1 U14935 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11489) );
  NAND2_X1 U14936 ( .A1(n11524), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11488) );
  NAND4_X1 U14937 ( .A1(n11491), .A2(n11490), .A3(n11489), .A4(n11488), .ZN(
        n11493) );
  OAI22_X1 U14938 ( .A1(n16153), .A2(n16030), .B1(n11252), .B2(n16042), .ZN(
        n11492) );
  NOR2_X1 U14939 ( .A1(n11493), .A2(n11492), .ZN(n11498) );
  AOI22_X1 U14940 ( .A1(n11494), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16206), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11497) );
  OAI22_X1 U14941 ( .A1(n16217), .A2(n16029), .B1(n16228), .B2(n16027), .ZN(
        n11495) );
  INV_X1 U14942 ( .A(n11495), .ZN(n11496) );
  NAND4_X1 U14943 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n16498) );
  NAND2_X1 U14944 ( .A1(n11637), .A2(n16498), .ZN(n11501) );
  NAND2_X1 U14945 ( .A1(n11647), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U14946 ( .A1(n11504), .A2(n11503), .ZN(n14267) );
  AOI22_X1 U14947 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11523) );
  OAI22_X1 U14948 ( .A1(n16217), .A2(n16052), .B1(n16109), .B2(n16051), .ZN(
        n11506) );
  OAI22_X1 U14949 ( .A1(n16215), .A2(n16060), .B1(n16219), .B2(n21861), .ZN(
        n11505) );
  NOR2_X1 U14950 ( .A1(n11506), .A2(n11505), .ZN(n11520) );
  AOI22_X1 U14951 ( .A1(n16203), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14952 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11509) );
  NAND2_X1 U14953 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14954 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11507) );
  NAND4_X1 U14955 ( .A1(n11510), .A2(n11509), .A3(n11508), .A4(n11507), .ZN(
        n11512) );
  INV_X1 U14956 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16053) );
  OAI22_X1 U14957 ( .A1(n16153), .A2(n16053), .B1(n11252), .B2(n16064), .ZN(
        n11511) );
  NOR2_X1 U14958 ( .A1(n11512), .A2(n11511), .ZN(n11519) );
  OAI22_X1 U14959 ( .A1(n16225), .A2(n16061), .B1(n16229), .B2(n11513), .ZN(
        n11514) );
  INV_X1 U14960 ( .A(n11514), .ZN(n11518) );
  OAI22_X1 U14961 ( .A1(n16221), .A2(n11515), .B1(n16228), .B2(n16050), .ZN(
        n11516) );
  INV_X1 U14962 ( .A(n11516), .ZN(n11517) );
  NAND4_X1 U14963 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(
        n16021) );
  NAND2_X1 U14964 ( .A1(n11637), .A2(n16021), .ZN(n11522) );
  NAND2_X1 U14965 ( .A1(n11647), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14966 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14967 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n16203), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14968 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n16205), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11527) );
  NAND2_X1 U14969 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11526) );
  NAND2_X1 U14970 ( .A1(n11524), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11525) );
  NAND4_X1 U14971 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11530) );
  OAI22_X1 U14972 ( .A1(n16108), .A2(n11252), .B1(n16153), .B2(n16096), .ZN(
        n11529) );
  NOR2_X1 U14973 ( .A1(n11530), .A2(n11529), .ZN(n11541) );
  INV_X1 U14974 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16104) );
  OAI22_X1 U14975 ( .A1(n16217), .A2(n16097), .B1(n16215), .B2(n16104), .ZN(
        n11534) );
  INV_X1 U14976 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11532) );
  NAND2_X1 U14977 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11531) );
  OAI21_X1 U14978 ( .B1(n16229), .B2(n11532), .A(n11531), .ZN(n11533) );
  NOR2_X1 U14979 ( .A1(n11534), .A2(n11533), .ZN(n11540) );
  INV_X1 U14980 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16094) );
  OAI22_X1 U14981 ( .A1(n16105), .A2(n16225), .B1(n16109), .B2(n16094), .ZN(
        n11535) );
  INV_X1 U14982 ( .A(n11535), .ZN(n11539) );
  INV_X1 U14983 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16095) );
  OAI22_X1 U14984 ( .A1(n16095), .A2(n16228), .B1(n16221), .B2(n11536), .ZN(
        n11537) );
  INV_X1 U14985 ( .A(n11537), .ZN(n11538) );
  NAND4_X1 U14986 ( .A1(n11541), .A2(n11540), .A3(n11539), .A4(n11538), .ZN(
        n16477) );
  NAND2_X1 U14987 ( .A1(n11637), .A2(n16477), .ZN(n11543) );
  NAND2_X1 U14988 ( .A1(n11647), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11542) );
  INV_X1 U14989 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20748) );
  AOI22_X1 U14990 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11563) );
  INV_X1 U14991 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11545) );
  OAI22_X1 U14992 ( .A1(n11545), .A2(n16109), .B1(n16217), .B2(n16074), .ZN(
        n11547) );
  INV_X1 U14993 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16081) );
  OAI22_X1 U14994 ( .A1(n16081), .A2(n16215), .B1(n16219), .B2(n16086), .ZN(
        n11546) );
  NOR2_X1 U14995 ( .A1(n11547), .A2(n11546), .ZN(n11561) );
  AOI22_X1 U14996 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n16204), .B1(
        n16203), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14997 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n16205), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U14998 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11549) );
  NAND2_X1 U14999 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11548) );
  NAND4_X1 U15000 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11553) );
  INV_X1 U15001 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16073) );
  OAI22_X1 U15002 ( .A1(n16085), .A2(n11252), .B1(n16153), .B2(n16073), .ZN(
        n11552) );
  NOR2_X1 U15003 ( .A1(n11553), .A2(n11552), .ZN(n11560) );
  INV_X1 U15004 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11554) );
  OAI22_X1 U15005 ( .A1(n11554), .A2(n16229), .B1(n16225), .B2(n16082), .ZN(
        n11555) );
  INV_X1 U15006 ( .A(n11555), .ZN(n11559) );
  INV_X1 U15007 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16072) );
  OAI22_X1 U15008 ( .A1(n16072), .A2(n16228), .B1(n16221), .B2(n11556), .ZN(
        n11557) );
  INV_X1 U15009 ( .A(n11557), .ZN(n11558) );
  NAND4_X1 U15010 ( .A1(n11561), .A2(n11560), .A3(n11559), .A4(n11558), .ZN(
        n16489) );
  NAND2_X1 U15011 ( .A1(n11637), .A2(n16489), .ZN(n11562) );
  OAI211_X1 U15012 ( .C1(n11640), .C2(n20748), .A(n11563), .B(n11562), .ZN(
        n14278) );
  AOI22_X1 U15013 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n11582) );
  INV_X1 U15014 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16118) );
  INV_X1 U15015 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16121) );
  OAI22_X1 U15016 ( .A1(n16118), .A2(n16109), .B1(n16217), .B2(n16121), .ZN(
        n11565) );
  INV_X1 U15017 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16128) );
  OAI22_X1 U15018 ( .A1(n16128), .A2(n16215), .B1(n16219), .B2(n16133), .ZN(
        n11564) );
  NOR2_X1 U15019 ( .A1(n11565), .A2(n11564), .ZN(n11579) );
  AOI22_X1 U15020 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n16204), .B1(
        n16203), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U15021 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n16205), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U15022 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11567) );
  INV_X1 U15023 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n21882) );
  NAND2_X1 U15024 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11566) );
  NAND4_X1 U15025 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n11571) );
  INV_X1 U15026 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16132) );
  INV_X1 U15027 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16120) );
  OAI22_X1 U15028 ( .A1(n16132), .A2(n11252), .B1(n16153), .B2(n16120), .ZN(
        n11570) );
  NOR2_X1 U15029 ( .A1(n11571), .A2(n11570), .ZN(n11578) );
  INV_X1 U15030 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11572) );
  INV_X1 U15031 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16129) );
  OAI22_X1 U15032 ( .A1(n11572), .A2(n16229), .B1(n16225), .B2(n16129), .ZN(
        n11573) );
  INV_X1 U15033 ( .A(n11573), .ZN(n11577) );
  INV_X1 U15034 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16119) );
  INV_X1 U15035 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11574) );
  OAI22_X1 U15036 ( .A1(n16119), .A2(n16228), .B1(n16221), .B2(n11574), .ZN(
        n11575) );
  INV_X1 U15037 ( .A(n11575), .ZN(n11576) );
  NAND4_X1 U15038 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n16484) );
  NAND2_X1 U15039 ( .A1(n11637), .A2(n16484), .ZN(n11581) );
  NAND2_X1 U15040 ( .A1(n11647), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U15041 ( .A1(n11583), .A2(n10821), .ZN(n14300) );
  AOI22_X1 U15042 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U15043 ( .A1(n16203), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U15044 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11586) );
  NAND2_X1 U15045 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11585) );
  NAND2_X1 U15046 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11584) );
  NAND4_X1 U15047 ( .A1(n11587), .A2(n11586), .A3(n11585), .A4(n11584), .ZN(
        n11589) );
  OAI22_X1 U15048 ( .A1(n16153), .A2(n16144), .B1(n11252), .B2(n16157), .ZN(
        n11588) );
  NOR2_X1 U15049 ( .A1(n11589), .A2(n11588), .ZN(n11599) );
  INV_X1 U15050 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16151) );
  OAI22_X1 U15051 ( .A1(n16217), .A2(n16143), .B1(n16215), .B2(n16151), .ZN(
        n11591) );
  INV_X1 U15052 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16156) );
  OAI22_X1 U15053 ( .A1(n16225), .A2(n16152), .B1(n16219), .B2(n16156), .ZN(
        n11590) );
  NOR2_X1 U15054 ( .A1(n11591), .A2(n11590), .ZN(n11598) );
  OAI22_X1 U15055 ( .A1(n16109), .A2(n16142), .B1(n16229), .B2(n11592), .ZN(
        n11593) );
  INV_X1 U15056 ( .A(n11593), .ZN(n11597) );
  OAI22_X1 U15057 ( .A1(n16221), .A2(n11594), .B1(n16228), .B2(n16141), .ZN(
        n11595) );
  INV_X1 U15058 ( .A(n11595), .ZN(n11596) );
  NAND4_X1 U15059 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n16479) );
  NAND2_X1 U15060 ( .A1(n11637), .A2(n16479), .ZN(n11601) );
  NAND2_X1 U15061 ( .A1(n11647), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11600) );
  INV_X1 U15062 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n15813) );
  AOI22_X1 U15063 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U15064 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n16203), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U15065 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n16205), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11605) );
  NAND2_X1 U15066 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11604) );
  NAND2_X1 U15067 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11603) );
  NAND4_X1 U15068 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11608) );
  OAI22_X1 U15069 ( .A1(n16339), .A2(n11252), .B1(n16153), .B2(n17312), .ZN(
        n11607) );
  NOR2_X1 U15070 ( .A1(n11608), .A2(n11607), .ZN(n11618) );
  OAI22_X1 U15071 ( .A1(n16217), .A2(n16342), .B1(n16215), .B2(n21796), .ZN(
        n11610) );
  INV_X1 U15072 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16174) );
  OAI22_X1 U15073 ( .A1(n16228), .A2(n16351), .B1(n16219), .B2(n16174), .ZN(
        n11609) );
  NOR2_X1 U15074 ( .A1(n11610), .A2(n11609), .ZN(n11617) );
  OAI22_X1 U15075 ( .A1(n16341), .A2(n16225), .B1(n16109), .B2(n16165), .ZN(
        n11611) );
  INV_X1 U15076 ( .A(n11611), .ZN(n11616) );
  OAI22_X1 U15077 ( .A1(n11613), .A2(n16229), .B1(n16221), .B2(n11612), .ZN(
        n11614) );
  INV_X1 U15078 ( .A(n11614), .ZN(n11615) );
  NAND4_X1 U15079 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n16472) );
  NAND2_X1 U15080 ( .A1(n11637), .A2(n16472), .ZN(n11619) );
  OAI211_X1 U15081 ( .C1(n15813), .C2(n11640), .A(n11620), .B(n11619), .ZN(
        n14368) );
  INV_X1 U15082 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n16789) );
  AOI22_X1 U15083 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11639) );
  INV_X1 U15084 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16224) );
  OAI22_X1 U15085 ( .A1(n16227), .A2(n16217), .B1(n16109), .B2(n16224), .ZN(
        n11622) );
  INV_X1 U15086 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16211) );
  OAI22_X1 U15087 ( .A1(n16211), .A2(n16215), .B1(n16219), .B2(n16494), .ZN(
        n11621) );
  NOR2_X1 U15088 ( .A1(n11622), .A2(n11621), .ZN(n11636) );
  AOI22_X1 U15089 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n16204), .B1(
        n16203), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U15090 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n16205), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U15091 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11624) );
  NAND2_X1 U15092 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11623) );
  NAND4_X1 U15093 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11628) );
  INV_X1 U15094 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16220) );
  OAI22_X1 U15095 ( .A1(n16216), .A2(n11252), .B1(n16153), .B2(n16220), .ZN(
        n11627) );
  NOR2_X1 U15096 ( .A1(n11628), .A2(n11627), .ZN(n11635) );
  INV_X1 U15097 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11629) );
  OAI22_X1 U15098 ( .A1(n11629), .A2(n16229), .B1(n16225), .B2(n21759), .ZN(
        n11630) );
  INV_X1 U15099 ( .A(n11630), .ZN(n11634) );
  OAI22_X1 U15100 ( .A1(n16230), .A2(n16228), .B1(n16221), .B2(n11631), .ZN(
        n11632) );
  INV_X1 U15101 ( .A(n11632), .ZN(n11633) );
  NAND4_X1 U15102 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n16456) );
  NAND2_X1 U15103 ( .A1(n11637), .A2(n16456), .ZN(n11638) );
  OAI211_X1 U15104 ( .C1(n11640), .C2(n16789), .A(n11639), .B(n11638), .ZN(
        n16626) );
  AOI22_X1 U15105 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n11642) );
  NAND2_X1 U15106 ( .A1(n11647), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U15107 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n11644) );
  NAND2_X1 U15108 ( .A1(n11647), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U15109 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n11646) );
  NAND2_X1 U15110 ( .A1(n11647), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11645) );
  NOR2_X2 U15111 ( .A1(n15769), .A2(n15770), .ZN(n15754) );
  AOI22_X1 U15112 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n11649) );
  NAND2_X1 U15113 ( .A1(n11647), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11648) );
  NAND2_X1 U15114 ( .A1(n11649), .A2(n11648), .ZN(n15756) );
  NAND2_X1 U15115 ( .A1(n15754), .A2(n15756), .ZN(n12949) );
  AOI22_X1 U15116 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n11651) );
  NAND2_X1 U15117 ( .A1(n11647), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11650) );
  OR2_X2 U15118 ( .A1(n12949), .A2(n12948), .ZN(n15724) );
  AOI22_X1 U15119 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n11653) );
  NAND2_X1 U15120 ( .A1(n11647), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11652) );
  NOR2_X4 U15121 ( .A1(n15724), .A2(n15723), .ZN(n15722) );
  AOI22_X1 U15122 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11655) );
  NAND2_X1 U15123 ( .A1(n11647), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U15124 ( .A1(n11655), .A2(n11654), .ZN(n15710) );
  AOI22_X1 U15125 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11657) );
  NAND2_X1 U15126 ( .A1(n11647), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11656) );
  NAND2_X1 U15127 ( .A1(n11657), .A2(n11656), .ZN(n15692) );
  AOI22_X1 U15128 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n11659) );
  NAND2_X1 U15129 ( .A1(n11647), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U15130 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n11661) );
  NAND2_X1 U15131 ( .A1(n11647), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U15132 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11663) );
  NAND2_X1 U15133 ( .A1(n11647), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11662) );
  NAND2_X1 U15134 ( .A1(n11663), .A2(n11662), .ZN(n15641) );
  AND2_X2 U15135 ( .A1(n15639), .A2(n15641), .ZN(n15624) );
  AOI22_X1 U15136 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11665) );
  NAND2_X1 U15137 ( .A1(n11647), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U15138 ( .A1(n11665), .A2(n11664), .ZN(n15625) );
  AOI22_X1 U15139 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n11667) );
  NAND2_X1 U15140 ( .A1(n11647), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U15141 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n11669) );
  NAND2_X1 U15142 ( .A1(n11647), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U15143 ( .A1(n12982), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n11670), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n11672) );
  NAND2_X1 U15144 ( .A1(n11647), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11671) );
  NAND2_X1 U15145 ( .A1(n11672), .A2(n11671), .ZN(n11673) );
  NAND2_X1 U15146 ( .A1(n17349), .A2(n20146), .ZN(n11679) );
  INV_X1 U15147 ( .A(n11676), .ZN(n11678) );
  NAND2_X1 U15148 ( .A1(n11678), .A2(n11677), .ZN(n17347) );
  AND2_X1 U15149 ( .A1(n11679), .A2(n17347), .ZN(n11680) );
  NAND2_X1 U15150 ( .A1(n20033), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14469) );
  NAND2_X1 U15151 ( .A1(n11078), .A2(n20854), .ZN(n11681) );
  NOR2_X1 U15152 ( .A1(n11681), .A2(n9742), .ZN(n11682) );
  NAND2_X1 U15153 ( .A1(n11677), .A2(n11682), .ZN(n17346) );
  NAND2_X1 U15154 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14018) );
  NOR2_X1 U15155 ( .A1(n14524), .A2(n14018), .ZN(n11704) );
  INV_X1 U15156 ( .A(n11704), .ZN(n14523) );
  NAND2_X1 U15157 ( .A1(n14524), .A2(n14018), .ZN(n14522) );
  INV_X1 U15158 ( .A(n14522), .ZN(n11702) );
  AOI21_X1 U15159 ( .B1(n11701), .B2(n14523), .A(n11702), .ZN(n11697) );
  INV_X1 U15160 ( .A(n13808), .ZN(n13807) );
  OAI21_X1 U15161 ( .B1(n11685), .B2(n13807), .A(n11684), .ZN(n11689) );
  OAI22_X1 U15162 ( .A1(n13808), .A2(n9748), .B1(n11078), .B2(n11686), .ZN(
        n11687) );
  INV_X1 U15163 ( .A(n11687), .ZN(n11688) );
  AND3_X1 U15164 ( .A1(n11690), .A2(n11689), .A3(n11688), .ZN(n11694) );
  NAND2_X1 U15165 ( .A1(n11394), .A2(n20146), .ZN(n14544) );
  NAND2_X1 U15166 ( .A1(n14544), .A2(n11691), .ZN(n11692) );
  NAND2_X1 U15167 ( .A1(n11692), .A2(n20156), .ZN(n11693) );
  NOR2_X1 U15168 ( .A1(n17280), .A2(n11695), .ZN(n11696) );
  NOR3_X1 U15169 ( .A1(n17253), .A2(n17229), .A3(n17228), .ZN(n17213) );
  AND2_X1 U15170 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17213), .ZN(
        n11705) );
  NAND2_X1 U15171 ( .A1(n17254), .A2(n11705), .ZN(n17204) );
  NAND2_X1 U15172 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17188) );
  INV_X1 U15173 ( .A(n17045), .ZN(n12007) );
  NAND2_X1 U15174 ( .A1(n12007), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11711) );
  NOR2_X1 U15175 ( .A1(n17046), .A2(n11711), .ZN(n17033) );
  INV_X1 U15176 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21939) );
  INV_X1 U15177 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17032) );
  NOR2_X1 U15178 ( .A1(n21939), .A2(n17032), .ZN(n11709) );
  AND2_X1 U15179 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n11709), .ZN(
        n11698) );
  NAND2_X1 U15180 ( .A1(n17033), .A2(n11698), .ZN(n16998) );
  NAND2_X1 U15181 ( .A1(n16943), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11699) );
  OR2_X1 U15182 ( .A1(n16998), .A2(n11699), .ZN(n16959) );
  INV_X1 U15183 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11974) );
  NOR3_X1 U15184 ( .A1(n16959), .A2(n16645), .A3(n11974), .ZN(n12990) );
  INV_X1 U15185 ( .A(n17046), .ZN(n11700) );
  INV_X1 U15186 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16857) );
  NAND2_X1 U15187 ( .A1(n11700), .A2(n16857), .ZN(n17179) );
  INV_X1 U15188 ( .A(n11701), .ZN(n17080) );
  NAND2_X1 U15189 ( .A1(n17080), .A2(n11702), .ZN(n11703) );
  INV_X1 U15190 ( .A(n20033), .ZN(n20051) );
  NAND2_X1 U15191 ( .A1(n11983), .A2(n20051), .ZN(n14525) );
  OAI211_X1 U15192 ( .C1(n11704), .C2(n17082), .A(n11703), .B(n14525), .ZN(
        n17255) );
  INV_X1 U15193 ( .A(n11705), .ZN(n11706) );
  AND2_X1 U15194 ( .A1(n17225), .A2(n11706), .ZN(n11707) );
  NOR2_X1 U15195 ( .A1(n17255), .A2(n11707), .ZN(n17216) );
  NAND2_X1 U15196 ( .A1(n17225), .A2(n17188), .ZN(n11708) );
  NAND2_X1 U15197 ( .A1(n17179), .A2(n17176), .ZN(n12952) );
  INV_X1 U15198 ( .A(n12952), .ZN(n17168) );
  INV_X1 U15199 ( .A(n17225), .ZN(n14049) );
  NAND2_X1 U15200 ( .A1(n17168), .A2(n14049), .ZN(n12985) );
  INV_X1 U15201 ( .A(n12985), .ZN(n11717) );
  NOR3_X1 U15202 ( .A1(n16645), .A2(n11974), .A3(n16974), .ZN(n11716) );
  INV_X1 U15203 ( .A(n11709), .ZN(n17020) );
  NOR2_X1 U15204 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17020), .ZN(
        n11710) );
  AND2_X1 U15205 ( .A1(n17033), .A2(n11710), .ZN(n17009) );
  NAND2_X1 U15206 ( .A1(n17225), .A2(n11711), .ZN(n11712) );
  NAND2_X1 U15207 ( .A1(n17176), .A2(n11712), .ZN(n17049) );
  AND2_X1 U15208 ( .A1(n17225), .A2(n17020), .ZN(n11713) );
  OR2_X1 U15209 ( .A1(n17049), .A2(n11713), .ZN(n17011) );
  OR2_X1 U15210 ( .A1(n17009), .A2(n17011), .ZN(n17000) );
  INV_X1 U15211 ( .A(n17000), .ZN(n11714) );
  NAND2_X1 U15212 ( .A1(n11714), .A2(n16943), .ZN(n11715) );
  NAND2_X1 U15213 ( .A1(n12985), .A2(n11715), .ZN(n16975) );
  OAI211_X1 U15214 ( .C1(n11717), .C2(n11716), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n16975), .ZN(n12986) );
  OAI21_X1 U15215 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12990), .A(
        n12986), .ZN(n11718) );
  OAI211_X1 U15216 ( .C1(n16515), .C2(n17256), .A(n14469), .B(n11718), .ZN(
        n11719) );
  INV_X1 U15217 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14181) );
  NOR2_X1 U15218 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11723) );
  NAND2_X1 U15219 ( .A1(n9742), .A2(n11723), .ZN(n11725) );
  NAND2_X1 U15220 ( .A1(n11725), .A2(n11724), .ZN(n11736) );
  NAND2_X1 U15221 ( .A1(n11741), .A2(n11736), .ZN(n11745) );
  INV_X1 U15222 ( .A(n11726), .ZN(n11727) );
  INV_X1 U15223 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11728) );
  MUX2_X1 U15224 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n11730), .S(n20166), .Z(
        n11760) );
  XNOR2_X1 U15225 ( .A(n11759), .B(n11760), .ZN(n15935) );
  NAND2_X1 U15226 ( .A1(n16903), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11757) );
  INV_X1 U15227 ( .A(n11731), .ZN(n11749) );
  NAND2_X1 U15228 ( .A1(n11745), .A2(n11732), .ZN(n11733) );
  NAND2_X1 U15229 ( .A1(n11749), .A2(n11733), .ZN(n15962) );
  INV_X1 U15230 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13996) );
  MUX2_X1 U15231 ( .A(n13996), .B(n11735), .S(n20166), .Z(n13882) );
  NOR2_X1 U15232 ( .A1(n13882), .A2(n14020), .ZN(n11738) );
  INV_X1 U15233 ( .A(n11736), .ZN(n11742) );
  NAND3_X1 U15234 ( .A1(n11889), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11737) );
  AND2_X1 U15235 ( .A1(n11742), .A2(n11737), .ZN(n15990) );
  NAND2_X1 U15236 ( .A1(n11738), .A2(n15990), .ZN(n14001) );
  NAND2_X1 U15237 ( .A1(n14001), .A2(n21897), .ZN(n11740) );
  INV_X1 U15238 ( .A(n11738), .ZN(n13883) );
  INV_X1 U15239 ( .A(n15990), .ZN(n11739) );
  NAND2_X1 U15240 ( .A1(n13883), .A2(n11739), .ZN(n14000) );
  AND2_X1 U15241 ( .A1(n11740), .A2(n14000), .ZN(n14527) );
  INV_X1 U15242 ( .A(n11741), .ZN(n11743) );
  NAND2_X1 U15243 ( .A1(n11743), .A2(n11742), .ZN(n11744) );
  NAND2_X1 U15244 ( .A1(n11745), .A2(n11744), .ZN(n15979) );
  XNOR2_X1 U15245 ( .A(n15979), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14526) );
  NOR2_X1 U15246 ( .A1(n15979), .A2(n14524), .ZN(n11746) );
  AOI21_X1 U15247 ( .B1(n14527), .B2(n14526), .A(n11746), .ZN(n11751) );
  INV_X1 U15248 ( .A(n11747), .ZN(n11748) );
  NAND2_X1 U15249 ( .A1(n11749), .A2(n11748), .ZN(n11750) );
  NAND2_X1 U15250 ( .A1(n11759), .A2(n11750), .ZN(n16916) );
  AND2_X1 U15251 ( .A1(n16916), .A2(n17228), .ZN(n11752) );
  AOI21_X1 U15252 ( .B1(n11751), .B2(n17253), .A(n11752), .ZN(n11756) );
  INV_X1 U15253 ( .A(n11751), .ZN(n16928) );
  INV_X1 U15254 ( .A(n11752), .ZN(n11753) );
  NAND3_X1 U15255 ( .A1(n16928), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n11753), .ZN(n11754) );
  OAI21_X1 U15256 ( .B1(n16916), .B2(n17228), .A(n11754), .ZN(n11755) );
  INV_X1 U15257 ( .A(n11760), .ZN(n11761) );
  MUX2_X1 U15258 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11762), .S(n20166), .Z(
        n11768) );
  XNOR2_X1 U15259 ( .A(n11763), .B(n11768), .ZN(n20054) );
  MUX2_X1 U15260 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n11894), .S(n20166), .Z(
        n11767) );
  NAND2_X1 U15261 ( .A1(n9742), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11764) );
  INV_X1 U15262 ( .A(n11776), .ZN(n11770) );
  INV_X1 U15263 ( .A(n11764), .ZN(n11765) );
  NAND2_X1 U15264 ( .A1(n11770), .A2(n11765), .ZN(n11766) );
  NAND2_X1 U15265 ( .A1(n11771), .A2(n11766), .ZN(n15905) );
  NOR2_X1 U15266 ( .A1(n15905), .A2(n11894), .ZN(n11818) );
  NAND2_X1 U15267 ( .A1(n11818), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16872) );
  OAI21_X1 U15268 ( .B1(n11763), .B2(n11768), .A(n11767), .ZN(n11769) );
  NAND2_X1 U15269 ( .A1(n15924), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16885) );
  INV_X1 U15270 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11772) );
  INV_X1 U15271 ( .A(n11815), .ZN(n11775) );
  NAND2_X1 U15272 ( .A1(n11775), .A2(n11774), .ZN(n11827) );
  INV_X1 U15273 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n16485) );
  NOR2_X1 U15274 ( .A1(n20166), .A2(n16485), .ZN(n11826) );
  INV_X1 U15275 ( .A(n11826), .ZN(n11777) );
  INV_X1 U15276 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11778) );
  NOR2_X1 U15277 ( .A1(n20166), .A2(n11778), .ZN(n11813) );
  OAI21_X1 U15278 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n11889), .ZN(n11779) );
  INV_X1 U15279 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11780) );
  INV_X1 U15280 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11781) );
  NOR2_X1 U15281 ( .A1(n20166), .A2(n11781), .ZN(n11829) );
  INV_X1 U15282 ( .A(n11829), .ZN(n11782) );
  INV_X1 U15283 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11784) );
  NOR2_X1 U15284 ( .A1(n20166), .A2(n11784), .ZN(n11796) );
  NAND2_X1 U15285 ( .A1(n9742), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11791) );
  INV_X1 U15286 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11785) );
  NAND2_X1 U15287 ( .A1(n11786), .A2(n11785), .ZN(n11855) );
  INV_X1 U15288 ( .A(n11786), .ZN(n11787) );
  NAND3_X1 U15289 ( .A1(n11787), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n11889), 
        .ZN(n11788) );
  AND2_X1 U15290 ( .A1(n11789), .A2(n11788), .ZN(n15735) );
  INV_X1 U15291 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17044) );
  NAND2_X1 U15292 ( .A1(n11835), .A2(n17044), .ZN(n16731) );
  INV_X1 U15293 ( .A(n11791), .ZN(n11792) );
  NAND2_X1 U15294 ( .A1(n9787), .A2(n11792), .ZN(n11793) );
  NAND2_X1 U15295 ( .A1(n11790), .A2(n11793), .ZN(n15764) );
  INV_X1 U15296 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12006) );
  NAND2_X1 U15297 ( .A1(n11795), .A2(n11796), .ZN(n11797) );
  NAND2_X1 U15298 ( .A1(n9787), .A2(n11797), .ZN(n15775) );
  INV_X1 U15299 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12955) );
  NAND2_X1 U15300 ( .A1(n11837), .A2(n12955), .ZN(n16743) );
  AND2_X1 U15301 ( .A1(n16741), .A2(n16743), .ZN(n11998) );
  NAND2_X1 U15302 ( .A1(n9742), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11799) );
  XNOR2_X1 U15303 ( .A(n11790), .B(n11799), .ZN(n15748) );
  NAND2_X1 U15304 ( .A1(n15748), .A2(n11864), .ZN(n11847) );
  INV_X1 U15305 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12005) );
  NAND2_X1 U15306 ( .A1(n11847), .A2(n12005), .ZN(n11999) );
  AND2_X1 U15307 ( .A1(n11998), .A2(n11999), .ZN(n16729) );
  NAND3_X1 U15308 ( .A1(n11800), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n11889), 
        .ZN(n11801) );
  OAI211_X1 U15309 ( .C1(n11800), .C2(P2_EBX_REG_16__SCAN_IN), .A(n11801), .B(
        n11879), .ZN(n15801) );
  OR2_X1 U15310 ( .A1(n15801), .A2(n11894), .ZN(n11802) );
  INV_X1 U15311 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17103) );
  NAND2_X1 U15312 ( .A1(n11802), .A2(n17103), .ZN(n11803) );
  NAND2_X1 U15313 ( .A1(n11889), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11805) );
  INV_X1 U15314 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n16476) );
  NAND2_X1 U15315 ( .A1(n11804), .A2(n16476), .ZN(n11809) );
  NAND2_X1 U15316 ( .A1(n15821), .A2(n11864), .ZN(n11807) );
  INV_X1 U15317 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17115) );
  NAND2_X1 U15318 ( .A1(n11807), .A2(n17115), .ZN(n16796) );
  INV_X1 U15319 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n21962) );
  NOR2_X1 U15320 ( .A1(n20166), .A2(n21962), .ZN(n11808) );
  NAND2_X1 U15321 ( .A1(n11809), .A2(n11808), .ZN(n11810) );
  NAND2_X1 U15322 ( .A1(n11810), .A2(n11800), .ZN(n20035) );
  OR2_X1 U15323 ( .A1(n20035), .A2(n11894), .ZN(n11811) );
  INV_X1 U15324 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17091) );
  NAND2_X1 U15325 ( .A1(n11811), .A2(n17091), .ZN(n16786) );
  XNOR2_X1 U15326 ( .A(n11812), .B(n10645), .ZN(n15837) );
  NAND2_X1 U15327 ( .A1(n15837), .A2(n11864), .ZN(n11841) );
  NAND2_X1 U15328 ( .A1(n11841), .A2(n10058), .ZN(n16805) );
  AND3_X1 U15329 ( .A1(n16796), .A2(n16786), .A3(n16805), .ZN(n11993) );
  NOR2_X1 U15330 ( .A1(n20166), .A2(n11774), .ZN(n11814) );
  AND2_X1 U15331 ( .A1(n11815), .A2(n11814), .ZN(n11816) );
  NOR2_X1 U15332 ( .A1(n11817), .A2(n11816), .ZN(n15868) );
  NAND2_X1 U15333 ( .A1(n15868), .A2(n11864), .ZN(n11843) );
  INV_X1 U15334 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17155) );
  NAND2_X1 U15335 ( .A1(n11843), .A2(n17155), .ZN(n16828) );
  INV_X1 U15336 ( .A(n11818), .ZN(n11819) );
  NAND2_X1 U15337 ( .A1(n11819), .A2(n17191), .ZN(n16871) );
  INV_X1 U15338 ( .A(n15924), .ZN(n11820) );
  NAND2_X1 U15339 ( .A1(n11820), .A2(n17190), .ZN(n16884) );
  NAND2_X1 U15340 ( .A1(n11889), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11822) );
  MUX2_X1 U15341 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n11822), .S(n11821), .Z(
        n11823) );
  NAND2_X1 U15342 ( .A1(n11823), .A2(n11879), .ZN(n15877) );
  OR2_X1 U15343 ( .A1(n15877), .A2(n11894), .ZN(n11824) );
  INV_X1 U15344 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17167) );
  NAND2_X1 U15345 ( .A1(n11824), .A2(n17167), .ZN(n16838) );
  NAND2_X1 U15346 ( .A1(n9742), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11825) );
  XNOR2_X1 U15347 ( .A(n11771), .B(n11825), .ZN(n15892) );
  NAND2_X1 U15348 ( .A1(n15892), .A2(n11864), .ZN(n11845) );
  NAND2_X1 U15349 ( .A1(n11845), .A2(n16857), .ZN(n16848) );
  NAND4_X1 U15350 ( .A1(n16828), .A2(n16824), .A3(n16838), .A4(n16848), .ZN(
        n11990) );
  NAND2_X1 U15351 ( .A1(n11827), .A2(n11826), .ZN(n11828) );
  AND2_X1 U15352 ( .A1(n11812), .A2(n11828), .ZN(n15854) );
  AOI21_X1 U15353 ( .B1(n15854), .B2(n11864), .A(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16816) );
  NOR2_X1 U15354 ( .A1(n11990), .A2(n16816), .ZN(n11832) );
  NAND2_X1 U15355 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  NAND2_X1 U15356 ( .A1(n11795), .A2(n11831), .ZN(n11839) );
  INV_X1 U15357 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17094) );
  OAI21_X1 U15358 ( .B1(n11839), .B2(n11894), .A(n17094), .ZN(n11997) );
  AND4_X1 U15359 ( .A1(n16776), .A2(n11993), .A3(n11832), .A4(n11997), .ZN(
        n11833) );
  AND3_X1 U15360 ( .A1(n16731), .A2(n16729), .A3(n11833), .ZN(n11834) );
  INV_X1 U15361 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11987) );
  INV_X1 U15362 ( .A(n11835), .ZN(n11836) );
  NAND2_X1 U15363 ( .A1(n11836), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16732) );
  NOR2_X1 U15364 ( .A1(n11837), .A2(n12955), .ZN(n16753) );
  AND2_X1 U15365 ( .A1(n11864), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11838) );
  OR3_X1 U15366 ( .A1(n20035), .A2(n11894), .A3(n17091), .ZN(n16785) );
  INV_X1 U15367 ( .A(n11839), .ZN(n15792) );
  AND2_X1 U15368 ( .A1(n11864), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11840) );
  NAND2_X1 U15369 ( .A1(n15792), .A2(n11840), .ZN(n11996) );
  INV_X1 U15370 ( .A(n11841), .ZN(n11842) );
  NAND2_X1 U15371 ( .A1(n11842), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16806) );
  OR2_X1 U15372 ( .A1(n11843), .A2(n17155), .ZN(n16829) );
  NAND2_X1 U15373 ( .A1(n11864), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11844) );
  OR2_X1 U15374 ( .A1(n15877), .A2(n11844), .ZN(n16837) );
  AND2_X1 U15375 ( .A1(n16837), .A2(n16849), .ZN(n16826) );
  AND2_X1 U15376 ( .A1(n16829), .A2(n16826), .ZN(n16782) );
  AND2_X1 U15377 ( .A1(n11864), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11846) );
  NAND2_X1 U15378 ( .A1(n15854), .A2(n11846), .ZN(n16815) );
  AND3_X1 U15379 ( .A1(n16806), .A2(n16782), .A3(n16815), .ZN(n11992) );
  INV_X1 U15380 ( .A(n11848), .ZN(n11849) );
  NAND2_X1 U15381 ( .A1(n11849), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16742) );
  NAND2_X1 U15382 ( .A1(n9742), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11853) );
  INV_X1 U15383 ( .A(n11853), .ZN(n11854) );
  NAND2_X1 U15384 ( .A1(n11855), .A2(n11854), .ZN(n11856) );
  NAND2_X1 U15385 ( .A1(n11860), .A2(n11856), .ZN(n15714) );
  OR2_X1 U15386 ( .A1(n15714), .A2(n11894), .ZN(n11866) );
  NAND2_X1 U15387 ( .A1(n11866), .A2(n17032), .ZN(n16721) );
  INV_X1 U15388 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11857) );
  NOR2_X1 U15389 ( .A1(n20166), .A2(n11857), .ZN(n11859) );
  INV_X1 U15390 ( .A(n11859), .ZN(n11858) );
  XNOR2_X1 U15391 ( .A(n11860), .B(n11858), .ZN(n15704) );
  NAND2_X1 U15392 ( .A1(n15704), .A2(n11864), .ZN(n16696) );
  AND2_X1 U15393 ( .A1(n16696), .A2(n21939), .ZN(n11869) );
  INV_X1 U15394 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16421) );
  INV_X1 U15395 ( .A(n11862), .ZN(n11863) );
  NAND2_X1 U15396 ( .A1(n15662), .A2(n11863), .ZN(n15682) );
  OR2_X1 U15397 ( .A1(n11866), .A2(n17032), .ZN(n16722) );
  AOI21_X1 U15398 ( .B1(n21939), .B2(n16722), .A(n16696), .ZN(n11867) );
  NOR2_X1 U15399 ( .A1(n16700), .A2(n11867), .ZN(n11868) );
  NAND2_X1 U15400 ( .A1(n11870), .A2(n11348), .ZN(n16698) );
  INV_X1 U15401 ( .A(n11874), .ZN(n12725) );
  OAI211_X1 U15402 ( .C1(n15662), .C2(P2_EBX_REG_25__SCAN_IN), .A(
        P2_EBX_REG_26__SCAN_IN), .B(n9742), .ZN(n11871) );
  AND2_X1 U15403 ( .A1(n11864), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11872) );
  INV_X1 U15404 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16672) );
  NAND2_X1 U15405 ( .A1(n9742), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11875) );
  INV_X1 U15406 ( .A(n11875), .ZN(n11876) );
  NAND2_X1 U15407 ( .A1(n11877), .A2(n11876), .ZN(n11878) );
  NAND2_X1 U15408 ( .A1(n11883), .A2(n11878), .ZN(n15628) );
  NAND2_X1 U15409 ( .A1(n11879), .A2(n11864), .ZN(n11887) );
  INV_X1 U15410 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16673) );
  INV_X1 U15411 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11881) );
  NOR2_X1 U15412 ( .A1(n20166), .A2(n11881), .ZN(n11882) );
  NAND2_X1 U15413 ( .A1(n11883), .A2(n11882), .ZN(n11884) );
  NAND2_X1 U15414 ( .A1(n11885), .A2(n11884), .ZN(n13083) );
  INV_X1 U15415 ( .A(n11886), .ZN(n11888) );
  NOR2_X1 U15416 ( .A1(n11887), .A2(n16673), .ZN(n16686) );
  NOR2_X1 U15417 ( .A1(n11888), .A2(n16686), .ZN(n12720) );
  INV_X1 U15418 ( .A(n12720), .ZN(n16660) );
  NAND2_X1 U15419 ( .A1(n9742), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11891) );
  XNOR2_X1 U15420 ( .A(n11892), .B(n11891), .ZN(n11890) );
  OAI21_X1 U15421 ( .B1(n11890), .B2(n11894), .A(n16645), .ZN(n16638) );
  INV_X1 U15422 ( .A(n11890), .ZN(n14441) );
  NAND3_X1 U15423 ( .A1(n14441), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11864), .ZN(n16639) );
  NAND2_X1 U15424 ( .A1(n11889), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11893) );
  XOR2_X1 U15425 ( .A(n11893), .B(n12724), .Z(n11895) );
  INV_X1 U15426 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12987) );
  INV_X1 U15427 ( .A(n11895), .ZN(n13119) );
  NAND3_X1 U15428 ( .A1(n13119), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n11864), .ZN(n12722) );
  NAND2_X1 U15429 ( .A1(n12717), .A2(n12722), .ZN(n11896) );
  INV_X1 U15430 ( .A(n11983), .ZN(n11897) );
  NOR2_X1 U15431 ( .A1(n17352), .A2(n11358), .ZN(n20836) );
  INV_X1 U15432 ( .A(n14312), .ZN(n11902) );
  AOI22_X1 U15433 ( .A1(n12705), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11900) );
  NAND2_X1 U15434 ( .A1(n11977), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11899) );
  AND2_X1 U15435 ( .A1(n14317), .A2(n14313), .ZN(n11901) );
  NAND2_X1 U15436 ( .A1(n11902), .A2(n11901), .ZN(n14315) );
  INV_X1 U15437 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n16904) );
  NAND2_X1 U15438 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11904) );
  NAND2_X1 U15439 ( .A1(n12705), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11903) );
  OAI211_X1 U15440 ( .C1(n12707), .C2(n16904), .A(n11904), .B(n11903), .ZN(
        n11905) );
  AOI21_X1 U15441 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11905), .ZN(n14362) );
  INV_X1 U15442 ( .A(n14362), .ZN(n11906) );
  INV_X1 U15443 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n21812) );
  NAND2_X1 U15444 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11908) );
  NAND2_X1 U15445 ( .A1(n12705), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11907) );
  OAI211_X1 U15446 ( .C1(n11968), .C2(n21812), .A(n11908), .B(n11907), .ZN(
        n11909) );
  AOI21_X1 U15447 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11909), .ZN(n14342) );
  INV_X1 U15448 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20741) );
  NAND2_X1 U15449 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11911) );
  NAND2_X1 U15450 ( .A1(n12705), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11910) );
  OAI211_X1 U15451 ( .C1(n11968), .C2(n20741), .A(n11911), .B(n11910), .ZN(
        n11912) );
  AOI21_X1 U15452 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11912), .ZN(n15919) );
  INV_X1 U15453 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20743) );
  NAND2_X1 U15454 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11914) );
  AOI22_X1 U15455 ( .A1(n12705), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11913) );
  OAI211_X1 U15456 ( .C1(n20743), .C2(n12707), .A(n11914), .B(n11913), .ZN(
        n15903) );
  INV_X1 U15457 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20745) );
  NAND2_X1 U15458 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11916) );
  NAND2_X1 U15459 ( .A1(n12705), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11915) );
  OAI211_X1 U15460 ( .C1(n11968), .C2(n20745), .A(n11916), .B(n11915), .ZN(
        n11917) );
  AOI21_X1 U15461 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11917), .ZN(n14353) );
  INV_X1 U15462 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n16841) );
  NAND2_X1 U15463 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11920) );
  NAND2_X1 U15464 ( .A1(n12705), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11919) );
  OAI211_X1 U15465 ( .C1(n11968), .C2(n16841), .A(n11920), .B(n11919), .ZN(
        n11921) );
  AOI21_X1 U15466 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11921), .ZN(n15875) );
  NAND2_X1 U15467 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11923) );
  AOI22_X1 U15468 ( .A1(n12705), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11922) );
  OAI211_X1 U15469 ( .C1(n20748), .C2(n12707), .A(n11923), .B(n11922), .ZN(
        n15858) );
  INV_X1 U15470 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U15471 ( .A1(n12705), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11925) );
  NAND2_X1 U15472 ( .A1(n11977), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11924) );
  INV_X1 U15473 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16809) );
  NAND2_X1 U15474 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11927) );
  NAND2_X1 U15475 ( .A1(n12705), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11926) );
  OAI211_X1 U15476 ( .C1(n12707), .C2(n16809), .A(n11927), .B(n11926), .ZN(
        n11928) );
  AOI21_X1 U15477 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11928), .ZN(n15830) );
  NAND2_X1 U15478 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11931) );
  NAND2_X1 U15479 ( .A1(n12705), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11930) );
  OAI211_X1 U15480 ( .C1(n12707), .C2(n15813), .A(n11931), .B(n11930), .ZN(
        n11932) );
  AOI21_X1 U15481 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11932), .ZN(n15826) );
  NAND2_X1 U15482 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11934) );
  NAND2_X1 U15483 ( .A1(n12705), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11933) );
  OAI211_X1 U15484 ( .C1(n11968), .C2(n16789), .A(n11934), .B(n11933), .ZN(
        n11935) );
  AOI21_X1 U15485 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11935), .ZN(n16465) );
  INV_X1 U15486 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20755) );
  NAND2_X1 U15487 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11937) );
  AOI22_X1 U15488 ( .A1(n12705), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11936) );
  OAI211_X1 U15489 ( .C1(n20755), .C2(n12707), .A(n11937), .B(n11936), .ZN(
        n15799) );
  INV_X1 U15490 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20757) );
  NAND2_X1 U15491 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U15492 ( .A1(n12705), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11938) );
  OAI211_X1 U15493 ( .C1(n11968), .C2(n20757), .A(n11939), .B(n11938), .ZN(
        n11940) );
  AOI21_X1 U15494 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11940), .ZN(n15784) );
  INV_X1 U15495 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15772) );
  NAND2_X1 U15496 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11943) );
  NAND2_X1 U15497 ( .A1(n12705), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11942) );
  OAI211_X1 U15498 ( .C1(n11968), .C2(n15772), .A(n11943), .B(n11942), .ZN(
        n11944) );
  AOI21_X1 U15499 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11944), .ZN(n15768) );
  INV_X1 U15500 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20760) );
  NAND2_X1 U15501 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11946) );
  AOI22_X1 U15502 ( .A1(n12705), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11945) );
  OAI211_X1 U15503 ( .C1(n20760), .C2(n12707), .A(n11946), .B(n11945), .ZN(
        n15752) );
  INV_X1 U15504 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20762) );
  NAND2_X1 U15505 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U15506 ( .A1(n12705), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11947) );
  OAI211_X1 U15507 ( .C1(n12707), .C2(n20762), .A(n11948), .B(n11947), .ZN(
        n11949) );
  AOI21_X1 U15508 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11949), .ZN(n12013) );
  INV_X1 U15509 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20764) );
  NAND2_X1 U15510 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U15511 ( .A1(n12705), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11951) );
  OAI211_X1 U15512 ( .C1(n11968), .C2(n20764), .A(n11952), .B(n11951), .ZN(
        n11953) );
  AOI21_X1 U15513 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11953), .ZN(n15727) );
  AOI22_X1 U15514 ( .A1(n12705), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11955) );
  NAND2_X1 U15515 ( .A1(n11977), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11954) );
  INV_X1 U15516 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20767) );
  NAND2_X1 U15517 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11957) );
  AOI22_X1 U15518 ( .A1(n12705), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11956) );
  OAI211_X1 U15519 ( .C1(n20767), .C2(n12707), .A(n11957), .B(n11956), .ZN(
        n15695) );
  INV_X1 U15520 ( .A(n15674), .ZN(n11962) );
  INV_X1 U15521 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20769) );
  NAND2_X1 U15522 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11959) );
  NAND2_X1 U15523 ( .A1(n12705), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11958) );
  OAI211_X1 U15524 ( .C1(n12707), .C2(n20769), .A(n11959), .B(n11958), .ZN(
        n11960) );
  AOI21_X1 U15525 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11960), .ZN(n15676) );
  NAND2_X1 U15526 ( .A1(n11962), .A2(n11961), .ZN(n15657) );
  INV_X1 U15527 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n21909) );
  NAND2_X1 U15528 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U15529 ( .A1(n12705), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11963) );
  OAI211_X1 U15530 ( .C1(n12707), .C2(n21909), .A(n11964), .B(n11963), .ZN(
        n11965) );
  AOI21_X1 U15531 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11965), .ZN(n15661) );
  OR2_X2 U15532 ( .A1(n15657), .A2(n15661), .ZN(n15659) );
  INV_X1 U15533 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n16677) );
  NAND2_X1 U15534 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11967) );
  NAND2_X1 U15535 ( .A1(n12705), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11966) );
  OAI211_X1 U15536 ( .C1(n11968), .C2(n16677), .A(n11967), .B(n11966), .ZN(
        n11969) );
  AOI21_X1 U15537 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11969), .ZN(n15638) );
  INV_X1 U15538 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20774) );
  NAND2_X1 U15539 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11971) );
  AOI22_X1 U15540 ( .A1(n12705), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11970) );
  OAI211_X1 U15541 ( .C1(n20774), .C2(n12707), .A(n11971), .B(n11970), .ZN(
        n15621) );
  AOI22_X1 U15542 ( .A1(n12705), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11973) );
  NAND2_X1 U15543 ( .A1(n11977), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11972) );
  INV_X1 U15544 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20776) );
  AOI22_X1 U15545 ( .A1(n12705), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11975) );
  OAI21_X1 U15546 ( .B1(n12707), .B2(n20776), .A(n11975), .ZN(n11976) );
  AOI21_X1 U15547 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11976), .ZN(n14435) );
  AOI22_X1 U15548 ( .A1(n12705), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11979) );
  NAND2_X1 U15549 ( .A1(n11977), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11978) );
  AOI21_X1 U15550 ( .B1(n17327), .B2(n20854), .A(n11981), .ZN(n11982) );
  NOR2_X1 U15551 ( .A1(n16388), .A2(n17241), .ZN(n11984) );
  AOI21_X1 U15552 ( .B1(n14467), .B2(n17221), .A(n11984), .ZN(n11985) );
  OAI211_X1 U15553 ( .C1(n14473), .C2(n17234), .A(n11986), .B(n11985), .ZN(
        P2_U3016) );
  INV_X1 U15554 ( .A(n11990), .ZN(n11991) );
  NAND2_X1 U15555 ( .A1(n11997), .A2(n11996), .ZN(n16769) );
  NAND2_X1 U15556 ( .A1(n16730), .A2(n11998), .ZN(n12001) );
  NAND2_X1 U15557 ( .A1(n16727), .A2(n11999), .ZN(n12000) );
  XNOR2_X1 U15558 ( .A(n12001), .B(n12000), .ZN(n12966) );
  MUX2_X1 U15559 ( .A(n20841), .B(n20835), .S(n20146), .Z(n12004) );
  NAND2_X1 U15560 ( .A1(n20851), .A2(n17372), .ZN(n12002) );
  NOR2_X1 U15561 ( .A1(n17352), .A2(n12002), .ZN(n12003) );
  AND2_X1 U15562 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12958) );
  INV_X1 U15563 ( .A(n13811), .ZN(n12009) );
  INV_X1 U15564 ( .A(n12011), .ZN(n12012) );
  AOI21_X1 U15565 ( .B1(n12013), .B2(n12010), .A(n12012), .ZN(n16438) );
  NAND2_X1 U15566 ( .A1(n17375), .A2(n17362), .ZN(n12015) );
  OAI21_X1 U15567 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n10286), .ZN(n17611) );
  OR2_X1 U15568 ( .A1(n17611), .A2(n17270), .ZN(n12014) );
  NAND2_X1 U15569 ( .A1(n12017), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13024) );
  AND2_X1 U15570 ( .A1(n12020), .A2(n15739), .ZN(n12021) );
  OR2_X1 U15571 ( .A1(n12021), .A2(n12711), .ZN(n15742) );
  NOR2_X1 U15572 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13971) );
  OR2_X1 U15573 ( .A1(n20800), .A2(n13971), .ZN(n17268) );
  NAND2_X1 U15574 ( .A1(n17268), .A2(n10286), .ZN(n12022) );
  NAND2_X1 U15575 ( .A1(n20481), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13068) );
  NAND2_X1 U15576 ( .A1(n14206), .A2(n13068), .ZN(n13884) );
  INV_X1 U15577 ( .A(n20033), .ZN(n16877) );
  NOR2_X1 U15578 ( .A1(n16877), .A2(n20762), .ZN(n12962) );
  AOI21_X1 U15579 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12962), .ZN(n12023) );
  OAI21_X1 U15580 ( .B1(n15742), .B2(n16933), .A(n12023), .ZN(n12024) );
  INV_X1 U15581 ( .A(n12025), .ZN(n12026) );
  OAI21_X1 U15582 ( .B1(n12966), .B2(n16942), .A(n12028), .ZN(P2_U2994) );
  AND2_X2 U15583 ( .A1(n12030), .A2(n15532), .ZN(n12133) );
  AOI22_X1 U15584 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12133), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12035) );
  NOR2_X2 U15585 ( .A1(n12029), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12041) );
  AOI22_X1 U15586 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15587 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12132), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12033) );
  NOR2_X4 U15588 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15589 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9774), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12032) );
  NAND4_X1 U15590 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12032), .ZN(
        n12048) );
  INV_X1 U15591 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12039) );
  AND2_X2 U15592 ( .A1(n12036), .A2(n12041), .ZN(n13662) );
  NAND2_X1 U15593 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12038) );
  NAND2_X1 U15594 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12037) );
  OAI211_X1 U15595 ( .C1(n12104), .C2(n12039), .A(n12038), .B(n12037), .ZN(
        n12040) );
  INV_X1 U15596 ( .A(n12040), .ZN(n12046) );
  AOI22_X1 U15597 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12044) );
  NAND2_X1 U15598 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12043) );
  NAND4_X1 U15599 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12047) );
  NAND2_X1 U15600 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12049) );
  NOR2_X1 U15601 ( .A1(n12104), .A2(n12050), .ZN(n12051) );
  NAND2_X1 U15602 ( .A1(n13322), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12056) );
  NAND2_X1 U15603 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12055) );
  NAND2_X1 U15604 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12054) );
  NAND2_X1 U15605 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12053) );
  NAND2_X1 U15606 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12060) );
  NAND2_X1 U15607 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12059) );
  NAND2_X1 U15608 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12058) );
  NAND2_X1 U15609 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12057) );
  NAND2_X1 U15610 ( .A1(n12133), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12064) );
  NAND2_X1 U15611 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12063) );
  AOI22_X1 U15612 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12132), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15613 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12133), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15614 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9774), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15615 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12069) );
  NAND2_X1 U15616 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12074) );
  NAND2_X1 U15617 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12073) );
  OAI211_X1 U15618 ( .C1(n12104), .C2(n12322), .A(n12074), .B(n12073), .ZN(
        n12075) );
  INV_X1 U15619 ( .A(n12075), .ZN(n12079) );
  AOI22_X1 U15620 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12078) );
  NAND2_X1 U15621 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12077) );
  AOI22_X1 U15622 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12076) );
  AND3_X2 U15623 ( .A1(n12080), .A2(n12079), .A3(n10802), .ZN(n12181) );
  NAND2_X1 U15624 ( .A1(n14961), .A2(n12182), .ZN(n12094) );
  INV_X1 U15625 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13518) );
  NAND2_X1 U15626 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12082) );
  NAND2_X1 U15627 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12081) );
  OAI211_X1 U15628 ( .C1(n13614), .C2(n13518), .A(n12082), .B(n12081), .ZN(
        n12083) );
  INV_X1 U15629 ( .A(n12083), .ZN(n12087) );
  AOI22_X1 U15630 ( .A1(n9753), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15631 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9777), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12085) );
  NAND2_X1 U15632 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12084) );
  NAND4_X1 U15633 ( .A1(n12087), .A2(n12086), .A3(n12085), .A4(n12084), .ZN(
        n12093) );
  AOI22_X1 U15634 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9774), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15635 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15636 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12132), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U15637 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12133), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12088) );
  NAND4_X1 U15638 ( .A1(n12091), .A2(n12090), .A3(n12089), .A4(n12088), .ZN(
        n12092) );
  INV_X2 U15639 ( .A(n12181), .ZN(n12233) );
  AND2_X2 U15640 ( .A1(n12181), .A2(n12186), .ZN(n12176) );
  NAND2_X1 U15641 ( .A1(n12182), .A2(n12186), .ZN(n12111) );
  AOI22_X1 U15642 ( .A1(n9774), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13725), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15643 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12108) );
  INV_X1 U15644 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12102) );
  NAND2_X1 U15645 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12101) );
  NAND2_X1 U15646 ( .A1(n12133), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12100) );
  OAI211_X1 U15647 ( .C1(n13722), .C2(n12102), .A(n12101), .B(n12100), .ZN(
        n12103) );
  INV_X1 U15648 ( .A(n12103), .ZN(n12107) );
  AOI22_X1 U15649 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9777), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12106) );
  NAND2_X1 U15650 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12105) );
  AOI22_X1 U15651 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15652 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13525), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15653 ( .A1(n15537), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15654 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12132), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15655 ( .A1(n13322), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12133), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15656 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12127), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15657 ( .A1(n9774), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9777), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12118) );
  NAND2_X1 U15658 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12117) );
  AOI22_X1 U15659 ( .A1(n9778), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9754), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12116) );
  NAND3_X1 U15660 ( .A1(n12118), .A2(n12117), .A3(n12116), .ZN(n12123) );
  INV_X1 U15661 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12121) );
  NAND2_X1 U15662 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12120) );
  NAND2_X1 U15663 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12119) );
  OAI211_X1 U15664 ( .C1(n12104), .C2(n12121), .A(n12120), .B(n12119), .ZN(
        n12122) );
  NAND2_X1 U15665 ( .A1(n9774), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12131) );
  NAND2_X1 U15666 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12129) );
  NAND2_X1 U15667 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12128) );
  NAND2_X1 U15668 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12137) );
  NAND2_X1 U15669 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12136) );
  NAND2_X1 U15670 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12135) );
  NAND2_X1 U15671 ( .A1(n12133), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12134) );
  AND2_X2 U15672 ( .A1(n12138), .A2(n10836), .ZN(n12152) );
  NAND2_X1 U15673 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12140) );
  NAND2_X1 U15674 ( .A1(n13322), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12139) );
  OAI211_X1 U15675 ( .C1(n13722), .C2(n12141), .A(n12140), .B(n12139), .ZN(
        n12142) );
  INV_X1 U15676 ( .A(n12142), .ZN(n12151) );
  NAND2_X1 U15677 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12147) );
  INV_X1 U15678 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12143) );
  NAND2_X1 U15679 ( .A1(n9778), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12145) );
  NAND2_X1 U15680 ( .A1(n9776), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12144) );
  NAND4_X1 U15681 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12149) );
  NAND3_X4 U15682 ( .A1(n12152), .A2(n12151), .A3(n12150), .ZN(n21060) );
  NAND2_X1 U15683 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12156) );
  NAND2_X1 U15684 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12155) );
  NAND2_X1 U15685 ( .A1(n9778), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12154) );
  NAND2_X1 U15686 ( .A1(n13564), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12153) );
  NAND4_X1 U15687 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12159) );
  NAND2_X1 U15688 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12164) );
  NAND2_X1 U15689 ( .A1(n9774), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12163) );
  NAND2_X1 U15690 ( .A1(n12241), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12162) );
  NAND2_X1 U15691 ( .A1(n12127), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12161) );
  NAND2_X1 U15692 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12168) );
  NAND2_X1 U15693 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12167) );
  NAND2_X1 U15694 ( .A1(n13322), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12166) );
  NAND2_X1 U15695 ( .A1(n12133), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12165) );
  NAND2_X1 U15696 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12170) );
  NAND2_X1 U15697 ( .A1(n9745), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12169) );
  OAI211_X1 U15698 ( .C1(n12104), .C2(n12254), .A(n12170), .B(n12169), .ZN(
        n12171) );
  INV_X1 U15699 ( .A(n12171), .ZN(n12172) );
  NAND2_X1 U15700 ( .A1(n12184), .A2(n10013), .ZN(n12667) );
  INV_X1 U15701 ( .A(n12203), .ZN(n12180) );
  INV_X1 U15702 ( .A(n12183), .ZN(n12179) );
  NAND2_X1 U15703 ( .A1(n12680), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12193) );
  NAND2_X1 U15704 ( .A1(n14961), .A2(n12181), .ZN(n12490) );
  XNOR2_X1 U15705 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12465) );
  NAND2_X1 U15706 ( .A1(n12193), .A2(n12208), .ZN(n12213) );
  NAND2_X1 U15707 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12215) );
  OAI21_X1 U15708 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n12215), .ZN(n21386) );
  NAND2_X1 U15709 ( .A1(n17524), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12210) );
  OAI21_X1 U15710 ( .B1(n13791), .B2(n21386), .A(n12210), .ZN(n12190) );
  INV_X1 U15711 ( .A(n12190), .ZN(n12191) );
  INV_X1 U15712 ( .A(n17524), .ZN(n12192) );
  MUX2_X1 U15713 ( .A(n12192), .B(n13791), .S(n21509), .Z(n12194) );
  NAND3_X1 U15714 ( .A1(n12193), .A2(n12208), .A3(n12194), .ZN(n12197) );
  INV_X1 U15715 ( .A(n12194), .ZN(n12195) );
  INV_X1 U15716 ( .A(n12198), .ZN(n12200) );
  NAND2_X1 U15717 ( .A1(n12200), .A2(n12199), .ZN(n12204) );
  INV_X1 U15718 ( .A(n17592), .ZN(n15601) );
  NOR2_X1 U15719 ( .A1(n15601), .A2(n21645), .ZN(n12201) );
  NAND2_X1 U15720 ( .A1(n15522), .A2(n10026), .ZN(n12673) );
  NAND2_X1 U15721 ( .A1(n12205), .A2(n12184), .ZN(n12206) );
  NAND2_X1 U15722 ( .A1(n12206), .A2(n21060), .ZN(n12207) );
  NAND2_X1 U15723 ( .A1(n12210), .A2(n12209), .ZN(n12211) );
  NAND2_X1 U15724 ( .A1(n10039), .A2(n12211), .ZN(n12212) );
  INV_X1 U15725 ( .A(n13791), .ZN(n12301) );
  INV_X1 U15726 ( .A(n12215), .ZN(n12214) );
  NAND2_X1 U15727 ( .A1(n12214), .A2(n21389), .ZN(n21424) );
  NAND2_X1 U15728 ( .A1(n12215), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12216) );
  NAND2_X1 U15729 ( .A1(n21424), .A2(n12216), .ZN(n15609) );
  AOI22_X1 U15730 ( .A1(n12301), .A2(n15609), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17524), .ZN(n12217) );
  NAND2_X1 U15731 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12220) );
  NAND2_X1 U15732 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12219) );
  OAI211_X1 U15733 ( .C1(n13614), .C2(n13238), .A(n12220), .B(n12219), .ZN(
        n12221) );
  INV_X1 U15734 ( .A(n12221), .ZN(n12226) );
  AOI22_X1 U15735 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15736 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9777), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12224) );
  NAND2_X1 U15737 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12223) );
  NAND4_X1 U15738 ( .A1(n12226), .A2(n12225), .A3(n12224), .A4(n12223), .ZN(
        n12232) );
  INV_X1 U15739 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n22000) );
  AOI22_X1 U15740 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15741 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12229) );
  INV_X1 U15742 ( .A(n9838), .ZN(n13639) );
  AOI22_X1 U15743 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15744 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12227) );
  NAND4_X1 U15745 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(
        n12231) );
  OAI22_X1 U15746 ( .A1(n12518), .A2(n13238), .B1(n12376), .B2(n12304), .ZN(
        n12234) );
  INV_X1 U15747 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13709) );
  NAND2_X1 U15748 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12239) );
  NAND2_X1 U15749 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12238) );
  OAI211_X1 U15750 ( .C1(n13614), .C2(n13709), .A(n12239), .B(n12238), .ZN(
        n12240) );
  INV_X1 U15751 ( .A(n12240), .ZN(n12245) );
  AOI22_X1 U15752 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15753 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12243) );
  NAND2_X1 U15754 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12242) );
  NAND4_X1 U15755 ( .A1(n12245), .A2(n12244), .A3(n12243), .A4(n12242), .ZN(
        n12251) );
  AOI22_X1 U15756 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13525), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15757 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15758 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9753), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15759 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12246) );
  NAND4_X1 U15760 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12250) );
  NAND2_X1 U15761 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12253) );
  NAND2_X1 U15762 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12252) );
  OAI211_X1 U15763 ( .C1(n13722), .C2(n12254), .A(n12253), .B(n12252), .ZN(
        n12255) );
  INV_X1 U15764 ( .A(n12255), .ZN(n12259) );
  AOI22_X1 U15765 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12258) );
  AOI22_X1 U15766 ( .A1(n9753), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12257) );
  NAND2_X1 U15767 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12256) );
  NAND4_X1 U15768 ( .A1(n12259), .A2(n12258), .A3(n12257), .A4(n12256), .ZN(
        n12265) );
  AOI22_X1 U15769 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15770 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15771 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9782), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15772 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9777), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12260) );
  NAND4_X1 U15773 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12264) );
  XNOR2_X1 U15774 ( .A(n12443), .B(n12386), .ZN(n12266) );
  NAND2_X1 U15775 ( .A1(n12266), .A2(n12294), .ZN(n12267) );
  NAND2_X1 U15776 ( .A1(n9763), .A2(n12386), .ZN(n12268) );
  OAI211_X1 U15777 ( .C1(n12443), .C2(n12233), .A(n12268), .B(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n12269) );
  INV_X1 U15778 ( .A(n12269), .ZN(n12271) );
  NAND2_X1 U15779 ( .A1(n12294), .A2(n12437), .ZN(n12272) );
  INV_X1 U15780 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13203) );
  OR2_X1 U15781 ( .A1(n12518), .A2(n13203), .ZN(n12289) );
  INV_X1 U15782 ( .A(n12304), .ZN(n12287) );
  NAND2_X1 U15783 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12274) );
  NAND2_X1 U15784 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12273) );
  OAI211_X1 U15785 ( .C1(n13722), .C2(n12275), .A(n12274), .B(n12273), .ZN(
        n12276) );
  INV_X1 U15786 ( .A(n12276), .ZN(n12280) );
  AOI22_X1 U15787 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15788 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12278) );
  NAND2_X1 U15789 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12277) );
  NAND4_X1 U15790 ( .A1(n12280), .A2(n12279), .A3(n12278), .A4(n12277), .ZN(
        n12286) );
  AOI22_X1 U15791 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15792 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15793 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15794 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12281) );
  NAND4_X1 U15795 ( .A1(n12284), .A2(n12283), .A3(n12282), .A4(n12281), .ZN(
        n12285) );
  NAND2_X1 U15796 ( .A1(n12287), .A2(n12380), .ZN(n12288) );
  INV_X1 U15797 ( .A(n21172), .ZN(n12292) );
  NAND2_X1 U15798 ( .A1(n12294), .A2(n12380), .ZN(n12295) );
  NAND2_X1 U15799 ( .A1(n12213), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12303) );
  INV_X1 U15800 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21385) );
  NOR3_X1 U15801 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21389), .A3(
        n21468), .ZN(n21301) );
  NAND2_X1 U15802 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21301), .ZN(
        n21294) );
  NAND2_X1 U15803 ( .A1(n21385), .A2(n21294), .ZN(n12300) );
  NAND3_X1 U15804 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21587) );
  INV_X1 U15805 ( .A(n21587), .ZN(n12299) );
  NAND2_X1 U15806 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12299), .ZN(
        n21582) );
  AOI22_X1 U15807 ( .A1(n12301), .A2(n21328), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17524), .ZN(n12302) );
  INV_X1 U15808 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13433) );
  NAND2_X1 U15809 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12307) );
  NAND2_X1 U15810 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12306) );
  OAI211_X1 U15811 ( .C1(n13614), .C2(n13433), .A(n12307), .B(n12306), .ZN(
        n12308) );
  INV_X1 U15812 ( .A(n12308), .ZN(n12312) );
  AOI22_X1 U15813 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15814 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12310) );
  NAND2_X1 U15815 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12309) );
  NAND4_X1 U15816 ( .A1(n12312), .A2(n12311), .A3(n12310), .A4(n12309), .ZN(
        n12318) );
  AOI22_X1 U15817 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15818 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15819 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15820 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12313) );
  NAND4_X1 U15821 ( .A1(n12316), .A2(n12315), .A3(n12314), .A4(n12313), .ZN(
        n12317) );
  AOI22_X1 U15822 ( .A1(n12521), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12528), .B2(n12410), .ZN(n12319) );
  INV_X1 U15823 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13634) );
  OR2_X1 U15824 ( .A1(n12518), .A2(n13634), .ZN(n12335) );
  NAND2_X1 U15825 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12321) );
  NAND2_X1 U15826 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12320) );
  OAI211_X1 U15827 ( .C1(n13722), .C2(n12322), .A(n12321), .B(n12320), .ZN(
        n12323) );
  INV_X1 U15828 ( .A(n12323), .ZN(n12327) );
  AOI22_X1 U15829 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13647), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15830 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n9753), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U15831 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12324) );
  NAND4_X1 U15832 ( .A1(n12327), .A2(n12326), .A3(n12325), .A4(n12324), .ZN(
        n12333) );
  AOI22_X1 U15833 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13723), .B1(
        n12133), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15834 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n9746), .B1(
        n13724), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15835 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15836 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13646), .B1(
        n9777), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12328) );
  NAND4_X1 U15837 ( .A1(n12331), .A2(n12330), .A3(n12329), .A4(n12328), .ZN(
        n12332) );
  NAND2_X1 U15838 ( .A1(n12528), .A2(n12412), .ZN(n12334) );
  NAND2_X1 U15839 ( .A1(n12335), .A2(n12334), .ZN(n12409) );
  OR2_X1 U15840 ( .A1(n12518), .A2(n13348), .ZN(n12350) );
  NAND2_X1 U15841 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12337) );
  NAND2_X1 U15842 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12336) );
  OAI211_X1 U15843 ( .C1(n13614), .C2(n13348), .A(n12337), .B(n12336), .ZN(
        n12338) );
  INV_X1 U15844 ( .A(n12338), .ZN(n12342) );
  INV_X1 U15845 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n22019) );
  AOI22_X1 U15846 ( .A1(n9753), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15847 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U15848 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12339) );
  NAND4_X1 U15849 ( .A1(n12342), .A2(n12341), .A3(n12340), .A4(n12339), .ZN(
        n12348) );
  AOI22_X1 U15850 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15851 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15852 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15853 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12133), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12343) );
  NAND4_X1 U15854 ( .A1(n12346), .A2(n12345), .A3(n12344), .A4(n12343), .ZN(
        n12347) );
  NAND2_X1 U15855 ( .A1(n12528), .A2(n12434), .ZN(n12349) );
  NAND2_X1 U15856 ( .A1(n12350), .A2(n12349), .ZN(n12403) );
  OR2_X1 U15857 ( .A1(n12518), .A2(n13685), .ZN(n12365) );
  NAND2_X1 U15858 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12352) );
  NAND2_X1 U15859 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12351) );
  OAI211_X1 U15860 ( .C1(n13614), .C2(n13685), .A(n12352), .B(n12351), .ZN(
        n12353) );
  INV_X1 U15861 ( .A(n12353), .ZN(n12357) );
  AOI22_X1 U15862 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13725), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15863 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U15864 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12354) );
  NAND4_X1 U15865 ( .A1(n12357), .A2(n12356), .A3(n12355), .A4(n12354), .ZN(
        n12363) );
  AOI22_X1 U15866 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15867 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15868 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15869 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12358) );
  NAND4_X1 U15870 ( .A1(n12361), .A2(n12360), .A3(n12359), .A4(n12358), .ZN(
        n12362) );
  NAND2_X1 U15871 ( .A1(n12528), .A2(n12433), .ZN(n12364) );
  NOR2_X1 U15872 ( .A1(n13785), .A2(n12443), .ZN(n12366) );
  INV_X1 U15873 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15463) );
  NAND3_X1 U15874 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12367) );
  INV_X1 U15875 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15478) );
  INV_X1 U15876 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15456) );
  INV_X1 U15877 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12612) );
  OR2_X1 U15878 ( .A1(n15257), .A2(n12612), .ZN(n15214) );
  XNOR2_X1 U15879 ( .A(n15257), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15205) );
  NAND2_X1 U15880 ( .A1(n15257), .A2(n12612), .ZN(n15213) );
  NAND2_X1 U15881 ( .A1(n12386), .A2(n12380), .ZN(n12377) );
  NAND2_X1 U15882 ( .A1(n12377), .A2(n12376), .ZN(n12411) );
  INV_X1 U15883 ( .A(n12410), .ZN(n12370) );
  XNOR2_X1 U15884 ( .A(n12411), .B(n12370), .ZN(n12371) );
  NAND2_X1 U15885 ( .A1(n12371), .A2(n12438), .ZN(n12372) );
  NAND2_X1 U15886 ( .A1(n15293), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12402) );
  XNOR2_X1 U15887 ( .A(n12377), .B(n12376), .ZN(n12378) );
  AND2_X1 U15888 ( .A1(n9763), .A2(n12177), .ZN(n12387) );
  AOI21_X1 U15889 ( .B1(n12378), .B2(n12438), .A(n12387), .ZN(n12379) );
  AND2_X1 U15890 ( .A1(n12183), .A2(n12186), .ZN(n12384) );
  INV_X1 U15891 ( .A(n12380), .ZN(n12381) );
  XNOR2_X1 U15892 ( .A(n12381), .B(n12386), .ZN(n12382) );
  NAND2_X1 U15893 ( .A1(n12382), .A2(n12438), .ZN(n12383) );
  INV_X1 U15894 ( .A(n12385), .ZN(n12392) );
  INV_X1 U15895 ( .A(n12387), .ZN(n12388) );
  NAND2_X1 U15896 ( .A1(n12389), .A2(n12388), .ZN(n13786) );
  NOR2_X1 U15897 ( .A1(n13154), .A2(n13786), .ZN(n12391) );
  INV_X1 U15898 ( .A(n13785), .ZN(n12424) );
  OAI21_X1 U15899 ( .B1(n13786), .B2(n12424), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12390) );
  AOI21_X1 U15900 ( .B1(n12392), .B2(n12391), .A(n12390), .ZN(n12395) );
  OR2_X1 U15901 ( .A1(n12393), .A2(n13786), .ZN(n12394) );
  NAND2_X1 U15902 ( .A1(n12395), .A2(n12394), .ZN(n14291) );
  INV_X1 U15903 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21045) );
  OR2_X1 U15904 ( .A1(n14291), .A2(n21045), .ZN(n12396) );
  NAND2_X1 U15905 ( .A1(n14291), .A2(n21045), .ZN(n12397) );
  NAND2_X1 U15906 ( .A1(n12398), .A2(n12397), .ZN(n12399) );
  XNOR2_X1 U15907 ( .A(n12399), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14332) );
  INV_X1 U15908 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21034) );
  OR2_X1 U15909 ( .A1(n12399), .A2(n21034), .ZN(n12400) );
  INV_X1 U15910 ( .A(n15293), .ZN(n12401) );
  INV_X1 U15911 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21023) );
  XNOR2_X1 U15912 ( .A(n12404), .B(n12403), .ZN(n13188) );
  NAND2_X1 U15913 ( .A1(n13188), .A2(n12424), .ZN(n12408) );
  AND2_X1 U15914 ( .A1(n12410), .A2(n12412), .ZN(n12405) );
  NAND2_X1 U15915 ( .A1(n12411), .A2(n12405), .ZN(n12425) );
  XNOR2_X1 U15916 ( .A(n12425), .B(n12434), .ZN(n12406) );
  NAND2_X1 U15917 ( .A1(n12406), .A2(n12438), .ZN(n12407) );
  NAND2_X1 U15918 ( .A1(n12408), .A2(n12407), .ZN(n12420) );
  NAND2_X1 U15919 ( .A1(n13181), .A2(n12424), .ZN(n12416) );
  NAND2_X1 U15920 ( .A1(n12411), .A2(n12410), .ZN(n12413) );
  XNOR2_X1 U15921 ( .A(n12413), .B(n12412), .ZN(n12414) );
  NAND2_X1 U15922 ( .A1(n12414), .A2(n12438), .ZN(n12415) );
  OR2_X1 U15923 ( .A1(n20994), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12417) );
  NAND2_X1 U15924 ( .A1(n20994), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12419) );
  INV_X1 U15925 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17585) );
  AND2_X1 U15926 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12421) );
  INV_X1 U15927 ( .A(n12425), .ZN(n12436) );
  NAND2_X1 U15928 ( .A1(n12436), .A2(n12434), .ZN(n12426) );
  XNOR2_X1 U15929 ( .A(n12426), .B(n12433), .ZN(n12427) );
  NAND2_X1 U15930 ( .A1(n12427), .A2(n12438), .ZN(n12428) );
  NAND2_X1 U15931 ( .A1(n12429), .A2(n12428), .ZN(n17546) );
  OR2_X1 U15932 ( .A1(n17546), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12430) );
  NAND2_X1 U15933 ( .A1(n17546), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12431) );
  AOI22_X1 U15934 ( .A1(n12521), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12528), .B2(n12437), .ZN(n12432) );
  OR2_X1 U15935 ( .A1(n13249), .A2(n13785), .ZN(n12441) );
  AND2_X1 U15936 ( .A1(n12434), .A2(n12433), .ZN(n12435) );
  NAND2_X1 U15937 ( .A1(n12436), .A2(n12435), .ZN(n12442) );
  XNOR2_X1 U15938 ( .A(n12442), .B(n12437), .ZN(n12439) );
  NAND2_X1 U15939 ( .A1(n12439), .A2(n12438), .ZN(n12440) );
  NAND2_X1 U15940 ( .A1(n12441), .A2(n12440), .ZN(n12449) );
  OR2_X1 U15941 ( .A1(n12449), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17540) );
  INV_X1 U15942 ( .A(n12442), .ZN(n12445) );
  NAND2_X1 U15943 ( .A1(n12445), .A2(n12444), .ZN(n15254) );
  INV_X1 U15944 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17569) );
  OR2_X1 U15945 ( .A1(n15254), .A2(n17569), .ZN(n12446) );
  NAND2_X1 U15946 ( .A1(n15257), .A2(n12446), .ZN(n12448) );
  INV_X1 U15947 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15505) );
  NAND2_X1 U15948 ( .A1(n17569), .A2(n15505), .ZN(n12447) );
  NAND2_X1 U15949 ( .A1(n12448), .A2(n12447), .ZN(n12450) );
  NAND2_X1 U15950 ( .A1(n12449), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17539) );
  AOI21_X1 U15951 ( .B1(n15254), .B2(n17569), .A(n15505), .ZN(n15188) );
  NAND2_X1 U15952 ( .A1(n15188), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12452) );
  NAND2_X1 U15953 ( .A1(n15257), .A2(n12452), .ZN(n12453) );
  INV_X1 U15954 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15476) );
  INV_X1 U15955 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15266) );
  NAND2_X1 U15956 ( .A1(n15476), .A2(n15266), .ZN(n15236) );
  INV_X1 U15957 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12455) );
  INV_X1 U15958 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15430) );
  AND3_X1 U15959 ( .A1(n12455), .A2(n12612), .A3(n15430), .ZN(n12456) );
  NOR2_X1 U15960 ( .A1(n15257), .A2(n12456), .ZN(n12457) );
  AND2_X1 U15961 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12696) );
  NAND2_X1 U15962 ( .A1(n12696), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15378) );
  INV_X1 U15963 ( .A(n15378), .ZN(n12459) );
  INV_X1 U15964 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12633) );
  INV_X1 U15965 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15398) );
  NAND2_X1 U15966 ( .A1(n12633), .A2(n15398), .ZN(n12460) );
  NAND3_X1 U15967 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15338) );
  INV_X1 U15968 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12461) );
  INV_X1 U15969 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15128) );
  INV_X1 U15970 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15118) );
  INV_X1 U15971 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15099) );
  INV_X1 U15972 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15087) );
  NAND2_X1 U15973 ( .A1(n15099), .A2(n15087), .ZN(n15315) );
  INV_X1 U15974 ( .A(n15315), .ZN(n12462) );
  INV_X1 U15975 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15308) );
  AND2_X1 U15976 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15305) );
  NOR2_X1 U15977 ( .A1(n10812), .A2(n15308), .ZN(n12463) );
  NAND2_X1 U15978 ( .A1(n14500), .A2(n14501), .ZN(n12464) );
  XNOR2_X1 U15979 ( .A(n12464), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15075) );
  NOR2_X1 U15980 ( .A1(n12465), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n13862) );
  XNOR2_X1 U15981 ( .A(n12209), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12480) );
  INV_X1 U15982 ( .A(n12480), .ZN(n12467) );
  NAND2_X1 U15983 ( .A1(n21509), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12479) );
  INV_X1 U15984 ( .A(n12479), .ZN(n12466) );
  NAND2_X1 U15985 ( .A1(n12467), .A2(n12466), .ZN(n12481) );
  NAND2_X1 U15986 ( .A1(n21468), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12468) );
  NAND2_X1 U15987 ( .A1(n12481), .A2(n12468), .ZN(n12484) );
  XNOR2_X1 U15988 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12483) );
  NAND2_X1 U15989 ( .A1(n12484), .A2(n12483), .ZN(n12470) );
  NAND2_X1 U15990 ( .A1(n21389), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12469) );
  NOR2_X1 U15991 ( .A1(n12471), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12472) );
  INV_X1 U15992 ( .A(n12478), .ZN(n12474) );
  NOR2_X1 U15993 ( .A1(n17596), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12473) );
  INV_X1 U15994 ( .A(n12477), .ZN(n12475) );
  NAND2_X1 U15995 ( .A1(n12480), .A2(n12479), .ZN(n12482) );
  NAND2_X1 U15996 ( .A1(n12482), .A2(n12481), .ZN(n12503) );
  XNOR2_X1 U15997 ( .A(n12484), .B(n12483), .ZN(n12509) );
  XNOR2_X1 U15998 ( .A(n12486), .B(n12485), .ZN(n12516) );
  NAND2_X1 U15999 ( .A1(n12526), .A2(n12487), .ZN(n13869) );
  NOR2_X1 U16000 ( .A1(n13869), .A2(n21739), .ZN(n13744) );
  OAI21_X1 U16001 ( .B1(n12185), .B2(n13862), .A(n13744), .ZN(n12535) );
  XNOR2_X1 U16002 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12489) );
  NAND2_X1 U16003 ( .A1(n12528), .A2(n12489), .ZN(n12488) );
  NAND2_X1 U16004 ( .A1(n12524), .A2(n12488), .ZN(n12496) );
  INV_X1 U16005 ( .A(n12489), .ZN(n12492) );
  OAI211_X1 U16006 ( .C1(n12181), .C2(n12492), .A(n12490), .B(n12491), .ZN(
        n12494) );
  NAND2_X1 U16007 ( .A1(n14961), .A2(n12184), .ZN(n12493) );
  NAND2_X1 U16008 ( .A1(n12493), .A2(n12185), .ZN(n12511) );
  NAND2_X1 U16009 ( .A1(n12494), .A2(n12511), .ZN(n12495) );
  NAND2_X1 U16010 ( .A1(n12496), .A2(n12495), .ZN(n12504) );
  INV_X1 U16011 ( .A(n12504), .ZN(n12508) );
  INV_X1 U16012 ( .A(n12503), .ZN(n12497) );
  OR2_X1 U16013 ( .A1(n12518), .A2(n12497), .ZN(n12499) );
  NAND2_X1 U16014 ( .A1(n12528), .A2(n21060), .ZN(n12498) );
  OR2_X1 U16015 ( .A1(n12186), .A2(n21645), .ZN(n12500) );
  INV_X1 U16016 ( .A(n12505), .ZN(n12507) );
  INV_X1 U16017 ( .A(n12528), .ZN(n12502) );
  AND2_X1 U16018 ( .A1(n12500), .A2(n21060), .ZN(n12501) );
  NAND2_X1 U16019 ( .A1(n12502), .A2(n12501), .ZN(n12519) );
  OAI211_X1 U16020 ( .C1(n12505), .C2(n12504), .A(n12503), .B(n12519), .ZN(
        n12506) );
  OAI21_X1 U16021 ( .B1(n12508), .B2(n12507), .A(n12506), .ZN(n12515) );
  INV_X1 U16022 ( .A(n12509), .ZN(n12512) );
  NAND2_X1 U16023 ( .A1(n12528), .A2(n12512), .ZN(n12510) );
  OAI21_X1 U16024 ( .B1(n12518), .B2(n12512), .A(n12511), .ZN(n12513) );
  INV_X1 U16025 ( .A(n12513), .ZN(n12514) );
  INV_X1 U16026 ( .A(n12524), .ZN(n12517) );
  INV_X1 U16027 ( .A(n12519), .ZN(n12522) );
  NAND3_X1 U16028 ( .A1(n12522), .A2(n12521), .A3(n12520), .ZN(n12523) );
  NAND2_X1 U16029 ( .A1(n9762), .A2(n21653), .ZN(n14055) );
  NAND2_X1 U16030 ( .A1(n13862), .A2(n21653), .ZN(n14474) );
  NAND2_X1 U16031 ( .A1(n14055), .A2(n14474), .ZN(n14406) );
  NAND2_X1 U16032 ( .A1(n12531), .A2(n14406), .ZN(n12532) );
  NAND3_X1 U16033 ( .A1(n12532), .A2(n12184), .A3(n13749), .ZN(n12533) );
  NAND2_X1 U16034 ( .A1(n15557), .A2(n12533), .ZN(n12534) );
  NAND2_X1 U16035 ( .A1(n15582), .A2(n9763), .ZN(n12536) );
  INV_X1 U16036 ( .A(n12542), .ZN(n12541) );
  NAND2_X1 U16037 ( .A1(n12538), .A2(n21060), .ZN(n12679) );
  AND2_X1 U16038 ( .A1(n12679), .A2(n12184), .ZN(n12539) );
  AND2_X1 U16039 ( .A1(n12540), .A2(n12539), .ZN(n12662) );
  AOI21_X1 U16040 ( .B1(n12541), .B2(n12537), .A(n12662), .ZN(n14479) );
  INV_X1 U16041 ( .A(n12691), .ZN(n12548) );
  NOR2_X1 U16042 ( .A1(n12537), .A2(n21060), .ZN(n17593) );
  INV_X1 U16043 ( .A(n12199), .ZN(n13863) );
  NAND2_X1 U16044 ( .A1(n12542), .A2(n13863), .ZN(n15523) );
  NAND2_X1 U16045 ( .A1(n12542), .A2(n12176), .ZN(n17510) );
  NAND2_X1 U16046 ( .A1(n15523), .A2(n17510), .ZN(n13867) );
  OAI22_X1 U16047 ( .A1(n12543), .A2(n12185), .B1(n12181), .B2(n12544), .ZN(
        n12545) );
  OR2_X1 U16048 ( .A1(n13867), .A2(n12545), .ZN(n12546) );
  NOR2_X1 U16049 ( .A1(n17593), .A2(n12546), .ZN(n12547) );
  INV_X1 U16050 ( .A(n12562), .ZN(n12596) );
  NAND2_X1 U16051 ( .A1(n12560), .A2(n12549), .ZN(n12551) );
  AND2_X1 U16052 ( .A1(n12551), .A2(n12550), .ZN(n12552) );
  INV_X1 U16053 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12555) );
  NAND2_X1 U16054 ( .A1(n9783), .A2(n12555), .ZN(n12554) );
  XNOR2_X1 U16055 ( .A(n12557), .B(n14014), .ZN(n14186) );
  NAND2_X1 U16056 ( .A1(n14186), .A2(n13864), .ZN(n12559) );
  INV_X1 U16057 ( .A(n12557), .ZN(n12558) );
  NAND2_X1 U16058 ( .A1(n12559), .A2(n12558), .ZN(n14287) );
  INV_X1 U16059 ( .A(n9780), .ZN(n12636) );
  MUX2_X1 U16060 ( .A(n12636), .B(n12561), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12563) );
  NAND2_X1 U16061 ( .A1(n12563), .A2(n10809), .ZN(n14286) );
  INV_X1 U16062 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12567) );
  NAND2_X1 U16063 ( .A1(n12638), .A2(n12567), .ZN(n12571) );
  NAND2_X1 U16064 ( .A1(n12586), .A2(n21023), .ZN(n12569) );
  NAND2_X1 U16065 ( .A1(n13864), .A2(n12567), .ZN(n12568) );
  NAND3_X1 U16066 ( .A1(n12569), .A2(n12561), .A3(n12568), .ZN(n12570) );
  AND2_X1 U16067 ( .A1(n12571), .A2(n12570), .ZN(n14451) );
  INV_X1 U16068 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20977) );
  NAND2_X1 U16069 ( .A1(n9780), .A2(n20977), .ZN(n12574) );
  INV_X1 U16070 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21018) );
  NAND2_X1 U16071 ( .A1(n13864), .A2(n20977), .ZN(n12572) );
  OAI211_X1 U16072 ( .C1(n9783), .C2(n21018), .A(n12572), .B(n12586), .ZN(
        n12573) );
  AND2_X1 U16073 ( .A1(n12574), .A2(n12573), .ZN(n20935) );
  OAI21_X1 U16074 ( .B1(n9784), .B2(n17585), .A(n12586), .ZN(n12575) );
  OAI21_X1 U16075 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n14391), .A(n12575), .ZN(
        n12577) );
  INV_X1 U16076 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14960) );
  NAND2_X1 U16077 ( .A1(n12638), .A2(n14960), .ZN(n12576) );
  INV_X1 U16078 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20973) );
  NAND2_X1 U16079 ( .A1(n9780), .A2(n20973), .ZN(n12581) );
  INV_X1 U16080 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21843) );
  NAND2_X1 U16081 ( .A1(n13864), .A2(n20973), .ZN(n12579) );
  OAI211_X1 U16082 ( .C1(n9783), .C2(n21843), .A(n12579), .B(n12586), .ZN(
        n12580) );
  NAND2_X1 U16083 ( .A1(n12581), .A2(n12580), .ZN(n17577) );
  INV_X1 U16084 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17575) );
  OAI21_X1 U16085 ( .B1(n9783), .B2(n17575), .A(n12586), .ZN(n12583) );
  INV_X1 U16086 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14951) );
  NAND2_X1 U16087 ( .A1(n13864), .A2(n14951), .ZN(n12582) );
  NAND2_X1 U16088 ( .A1(n12583), .A2(n12582), .ZN(n12584) );
  OAI21_X1 U16089 ( .B1(n12656), .B2(P1_EBX_REG_7__SCAN_IN), .A(n12584), .ZN(
        n14949) );
  INV_X1 U16090 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U16091 ( .A1(n9780), .A2(n12585), .ZN(n12589) );
  NAND2_X1 U16092 ( .A1(n13864), .A2(n12585), .ZN(n12587) );
  OAI211_X1 U16093 ( .C1(n9784), .C2(n17569), .A(n12587), .B(n12586), .ZN(
        n12588) );
  AND2_X1 U16094 ( .A1(n12589), .A2(n12588), .ZN(n14880) );
  OAI21_X1 U16095 ( .B1(n9784), .B2(n15505), .A(n12586), .ZN(n12590) );
  OAI21_X1 U16096 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n14391), .A(n12590), .ZN(
        n12592) );
  INV_X1 U16097 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14942) );
  NAND2_X1 U16098 ( .A1(n12638), .A2(n14942), .ZN(n12591) );
  MUX2_X1 U16099 ( .A(n9780), .B(n9783), .S(P1_EBX_REG_10__SCAN_IN), .Z(n12595) );
  INV_X1 U16100 ( .A(n12595), .ZN(n12598) );
  NAND2_X1 U16101 ( .A1(n15266), .A2(n12596), .ZN(n12597) );
  NAND2_X1 U16102 ( .A1(n12598), .A2(n12597), .ZN(n14870) );
  INV_X1 U16103 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14933) );
  NAND2_X1 U16104 ( .A1(n12638), .A2(n14933), .ZN(n12602) );
  NAND2_X1 U16105 ( .A1(n12586), .A2(n15476), .ZN(n12600) );
  NAND2_X1 U16106 ( .A1(n13864), .A2(n14933), .ZN(n12599) );
  NAND3_X1 U16107 ( .A1(n12600), .A2(n12561), .A3(n12599), .ZN(n12601) );
  NAND2_X1 U16108 ( .A1(n12602), .A2(n12601), .ZN(n14852) );
  INV_X1 U16109 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14932) );
  NAND2_X1 U16110 ( .A1(n9780), .A2(n14932), .ZN(n12605) );
  NAND2_X1 U16111 ( .A1(n13864), .A2(n14932), .ZN(n12603) );
  OAI211_X1 U16112 ( .C1(n9783), .C2(n15478), .A(n12603), .B(n12586), .ZN(
        n12604) );
  AND2_X1 U16113 ( .A1(n12605), .A2(n12604), .ZN(n14839) );
  INV_X1 U16114 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n21859) );
  NAND2_X1 U16115 ( .A1(n12638), .A2(n21859), .ZN(n12608) );
  NAND2_X1 U16116 ( .A1(n12586), .A2(n15463), .ZN(n12606) );
  OAI211_X1 U16117 ( .C1(P1_EBX_REG_13__SCAN_IN), .C2(n14391), .A(n12606), .B(
        n12561), .ZN(n12607) );
  MUX2_X1 U16118 ( .A(n12636), .B(n12561), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12611) );
  OAI21_X1 U16119 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14392), .A(
        n12611), .ZN(n14794) );
  INV_X1 U16120 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14928) );
  NAND2_X1 U16121 ( .A1(n12638), .A2(n14928), .ZN(n12616) );
  NAND2_X1 U16122 ( .A1(n12586), .A2(n12612), .ZN(n12614) );
  NAND2_X1 U16123 ( .A1(n13864), .A2(n14928), .ZN(n12613) );
  NAND3_X1 U16124 ( .A1(n12614), .A2(n12561), .A3(n12613), .ZN(n12615) );
  NAND2_X1 U16125 ( .A1(n12616), .A2(n12615), .ZN(n14785) );
  MUX2_X1 U16126 ( .A(n12636), .B(n12561), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12617) );
  OAI21_X1 U16127 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n14392), .A(
        n12617), .ZN(n14767) );
  INV_X1 U16128 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14753) );
  NAND2_X1 U16129 ( .A1(n12638), .A2(n14753), .ZN(n12620) );
  NAND2_X1 U16130 ( .A1(n12586), .A2(n15430), .ZN(n12618) );
  OAI211_X1 U16131 ( .C1(P1_EBX_REG_17__SCAN_IN), .C2(n14391), .A(n12618), .B(
        n12561), .ZN(n12619) );
  OR2_X2 U16132 ( .A1(n14769), .A2(n14757), .ZN(n14759) );
  INV_X1 U16133 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n12621) );
  NAND2_X1 U16134 ( .A1(n9780), .A2(n12621), .ZN(n12624) );
  INV_X1 U16135 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21858) );
  NAND2_X1 U16136 ( .A1(n13864), .A2(n12621), .ZN(n12622) );
  OAI211_X1 U16137 ( .C1(n9783), .C2(n21858), .A(n12622), .B(n12586), .ZN(
        n12623) );
  NAND2_X1 U16138 ( .A1(n12624), .A2(n12623), .ZN(n14741) );
  NOR2_X4 U16139 ( .A1(n14759), .A2(n14741), .ZN(n14740) );
  INV_X1 U16140 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n22032) );
  OAI21_X1 U16141 ( .B1(n9784), .B2(n22032), .A(n12586), .ZN(n12625) );
  OAI21_X1 U16142 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(n14391), .A(n12625), .ZN(
        n12628) );
  INV_X1 U16143 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n12626) );
  NAND2_X1 U16144 ( .A1(n12638), .A2(n12626), .ZN(n12627) );
  INV_X1 U16145 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14921) );
  NAND2_X1 U16146 ( .A1(n9780), .A2(n14921), .ZN(n12631) );
  NAND2_X1 U16147 ( .A1(n13864), .A2(n14921), .ZN(n12629) );
  OAI211_X1 U16148 ( .C1(n9784), .C2(n15398), .A(n12629), .B(n12586), .ZN(
        n12630) );
  NAND2_X1 U16149 ( .A1(n12631), .A2(n12630), .ZN(n14702) );
  NOR2_X1 U16150 ( .A1(n14717), .A2(n14702), .ZN(n12632) );
  NAND2_X1 U16151 ( .A1(n12586), .A2(n12633), .ZN(n12634) );
  OAI211_X1 U16152 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n14391), .A(n12634), .B(
        n12561), .ZN(n12635) );
  OAI21_X1 U16153 ( .B1(n12656), .B2(P1_EBX_REG_21__SCAN_IN), .A(n12635), .ZN(
        n14693) );
  MUX2_X1 U16154 ( .A(n12636), .B(n12561), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12637) );
  OAI21_X1 U16155 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n14392), .A(
        n12637), .ZN(n14677) );
  INV_X1 U16156 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U16157 ( .A1(n12638), .A2(n14670), .ZN(n12641) );
  NAND2_X1 U16158 ( .A1(n12586), .A2(n12461), .ZN(n12639) );
  OAI211_X1 U16159 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n14391), .A(n12639), .B(
        n12561), .ZN(n12640) );
  MUX2_X1 U16160 ( .A(n9780), .B(n9784), .S(P1_EBX_REG_24__SCAN_IN), .Z(n12643) );
  NOR2_X1 U16161 ( .A1(n14392), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12642) );
  NOR2_X1 U16162 ( .A1(n12643), .A2(n12642), .ZN(n14654) );
  NAND2_X1 U16163 ( .A1(n12586), .A2(n15118), .ZN(n12644) );
  OAI211_X1 U16164 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n14391), .A(n12644), .B(
        n12561), .ZN(n12645) );
  OAI21_X1 U16165 ( .B1(n12656), .B2(P1_EBX_REG_25__SCAN_IN), .A(n12645), .ZN(
        n14641) );
  NAND2_X1 U16166 ( .A1(n14640), .A2(n14641), .ZN(n14617) );
  INV_X1 U16167 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21892) );
  NAND2_X1 U16168 ( .A1(n9780), .A2(n21892), .ZN(n12648) );
  INV_X1 U16169 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15335) );
  NAND2_X1 U16170 ( .A1(n13864), .A2(n21892), .ZN(n12646) );
  OAI211_X1 U16171 ( .C1(n9784), .C2(n15335), .A(n12646), .B(n12586), .ZN(
        n12647) );
  NAND2_X1 U16172 ( .A1(n12648), .A2(n12647), .ZN(n14618) );
  OR2_X2 U16173 ( .A1(n14617), .A2(n14618), .ZN(n14620) );
  MUX2_X1 U16174 ( .A(n9780), .B(n9783), .S(P1_EBX_REG_28__SCAN_IN), .Z(n12650) );
  NOR2_X1 U16175 ( .A1(n14392), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12649) );
  NOR2_X1 U16176 ( .A1(n12650), .A2(n12649), .ZN(n14594) );
  NAND2_X1 U16177 ( .A1(n12586), .A2(n15099), .ZN(n12651) );
  OAI211_X1 U16178 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n14391), .A(n12651), .B(
        n12561), .ZN(n12652) );
  OAI21_X1 U16179 ( .B1(n12656), .B2(P1_EBX_REG_27__SCAN_IN), .A(n12652), .ZN(
        n14591) );
  NAND2_X1 U16180 ( .A1(n14594), .A2(n14591), .ZN(n12653) );
  OR2_X1 U16181 ( .A1(n14392), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12655) );
  INV_X1 U16182 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U16183 ( .A1(n13864), .A2(n14907), .ZN(n12654) );
  NAND2_X1 U16184 ( .A1(n12655), .A2(n12654), .ZN(n12657) );
  OAI22_X1 U16185 ( .A1(n12657), .A2(n9783), .B1(P1_EBX_REG_29__SCAN_IN), .B2(
        n12656), .ZN(n14577) );
  NAND2_X1 U16186 ( .A1(n14578), .A2(n14577), .ZN(n14580) );
  INV_X1 U16187 ( .A(n14580), .ZN(n14390) );
  INV_X1 U16188 ( .A(n14578), .ZN(n14592) );
  OAI22_X1 U16189 ( .A1(n14390), .A2(n12561), .B1(n12657), .B2(n14592), .ZN(
        n12660) );
  NAND2_X1 U16190 ( .A1(n14392), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12659) );
  NAND2_X1 U16191 ( .A1(n14391), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12658) );
  NAND2_X1 U16192 ( .A1(n12659), .A2(n12658), .ZN(n14389) );
  XNOR2_X1 U16193 ( .A(n12660), .B(n14389), .ZN(n14904) );
  INV_X1 U16194 ( .A(n14904), .ZN(n14575) );
  INV_X1 U16195 ( .A(n12543), .ZN(n13861) );
  NAND2_X1 U16196 ( .A1(n13861), .A2(n12185), .ZN(n17522) );
  OAI21_X1 U16197 ( .B1(n12544), .B2(n12233), .A(n17522), .ZN(n12661) );
  INV_X1 U16198 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14513) );
  INV_X1 U16199 ( .A(n12537), .ZN(n13870) );
  NAND2_X1 U16200 ( .A1(n13870), .A2(n21060), .ZN(n17497) );
  INV_X1 U16201 ( .A(n17497), .ZN(n15542) );
  INV_X1 U16202 ( .A(n12662), .ZN(n12671) );
  NAND2_X1 U16203 ( .A1(n10386), .A2(n9783), .ZN(n12669) );
  AOI21_X1 U16204 ( .B1(n15538), .B2(n12176), .A(n12184), .ZN(n12666) );
  OAI21_X1 U16205 ( .B1(n12666), .B2(n12665), .A(n21060), .ZN(n12668) );
  AND4_X1 U16206 ( .A1(n12669), .A2(n12668), .A3(n10816), .A4(n12667), .ZN(
        n12670) );
  OAI211_X1 U16207 ( .C1(n12672), .C2(n12199), .A(n12671), .B(n12670), .ZN(
        n14492) );
  OAI21_X1 U16208 ( .B1(n14488), .B2(n12184), .A(n12673), .ZN(n12674) );
  OR2_X1 U16209 ( .A1(n14492), .A2(n12674), .ZN(n12675) );
  AND2_X2 U16210 ( .A1(n12691), .A2(n12675), .ZN(n15373) );
  OR2_X2 U16211 ( .A1(n15396), .A2(n15373), .ZN(n17559) );
  NOR2_X1 U16212 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15396), .ZN(
        n21040) );
  INV_X1 U16213 ( .A(n21040), .ZN(n12676) );
  AND3_X1 U16214 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15506) );
  AND2_X1 U16215 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12677) );
  NAND2_X1 U16216 ( .A1(n15506), .A2(n12677), .ZN(n15489) );
  NOR2_X1 U16217 ( .A1(n21018), .A2(n21023), .ZN(n21011) );
  NOR2_X1 U16218 ( .A1(n21034), .A2(n21045), .ZN(n15499) );
  NAND2_X1 U16219 ( .A1(n21011), .A2(n15499), .ZN(n17558) );
  NOR3_X1 U16220 ( .A1(n17585), .A2(n15489), .A3(n17558), .ZN(n15475) );
  NAND3_X1 U16221 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n15475), .ZN(n12693) );
  INV_X1 U16222 ( .A(n12693), .ZN(n15372) );
  AND2_X1 U16223 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15372), .ZN(
        n12678) );
  NAND2_X1 U16224 ( .A1(n21035), .A2(n12678), .ZN(n15355) );
  OR2_X1 U16225 ( .A1(n12680), .A2(n12679), .ZN(n15524) );
  INV_X1 U16226 ( .A(n15524), .ZN(n12681) );
  INV_X1 U16227 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15586) );
  OAI21_X1 U16228 ( .B1(n15586), .B2(n21045), .A(n21034), .ZN(n21007) );
  NAND3_X1 U16229 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21011), .A3(
        n21007), .ZN(n15472) );
  NAND2_X1 U16230 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12682) );
  OR2_X1 U16231 ( .A1(n15489), .A2(n12682), .ZN(n12683) );
  NOR2_X1 U16232 ( .A1(n15472), .A2(n12683), .ZN(n12695) );
  INV_X1 U16233 ( .A(n12695), .ZN(n12684) );
  NAND2_X1 U16234 ( .A1(n15355), .A2(n12685), .ZN(n15455) );
  NAND3_X1 U16235 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15420) );
  NAND2_X1 U16236 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12686) );
  NOR2_X1 U16237 ( .A1(n15420), .A2(n12686), .ZN(n12690) );
  INV_X1 U16238 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12687) );
  NOR2_X1 U16239 ( .A1(n15378), .A2(n12687), .ZN(n12688) );
  AND2_X1 U16240 ( .A1(n12690), .A2(n12688), .ZN(n12689) );
  NAND2_X1 U16241 ( .A1(n15455), .A2(n12689), .ZN(n15363) );
  NAND3_X1 U16242 ( .A1(n15316), .A2(n15305), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14514) );
  INV_X1 U16243 ( .A(n15305), .ZN(n15314) );
  INV_X1 U16244 ( .A(n21008), .ZN(n21028) );
  OR2_X2 U16245 ( .A1(n17559), .A2(n21028), .ZN(n17561) );
  NAND2_X1 U16246 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15334) );
  NAND2_X1 U16247 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12698) );
  NAND2_X1 U16248 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12690), .ZN(
        n15376) );
  NAND2_X1 U16249 ( .A1(n15373), .A2(n15586), .ZN(n12692) );
  NAND2_X1 U16250 ( .A1(n17559), .A2(n12693), .ZN(n12694) );
  OAI211_X1 U16251 ( .C1(n12695), .C2(n21008), .A(n21030), .B(n12694), .ZN(
        n15465) );
  AOI21_X2 U16252 ( .B1(n15376), .B2(n17559), .A(n15465), .ZN(n15394) );
  INV_X1 U16253 ( .A(n12696), .ZN(n15377) );
  NOR2_X1 U16254 ( .A1(n15377), .A2(n15376), .ZN(n12697) );
  INV_X1 U16255 ( .A(n17561), .ZN(n21041) );
  AND2_X1 U16256 ( .A1(n21041), .A2(n21030), .ZN(n15504) );
  OAI21_X1 U16257 ( .B1(n15335), .B2(n15118), .A(n17561), .ZN(n12699) );
  NAND2_X1 U16258 ( .A1(n15337), .A2(n12699), .ZN(n15327) );
  AOI21_X1 U16259 ( .B1(n15314), .B2(n17561), .A(n15327), .ZN(n15309) );
  INV_X1 U16260 ( .A(n15337), .ZN(n15347) );
  NOR2_X1 U16261 ( .A1(n15347), .A2(n17561), .ZN(n14510) );
  AOI21_X1 U16262 ( .B1(n15309), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14510), .ZN(n12700) );
  INV_X1 U16263 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21712) );
  NOR2_X1 U16264 ( .A1(n17570), .A2(n21712), .ZN(n15069) );
  OAI21_X1 U16265 ( .B1(n15075), .B2(n21012), .A(n12701), .ZN(P1_U3001) );
  NAND2_X1 U16266 ( .A1(n16646), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12703) );
  INV_X1 U16267 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12702) );
  NAND2_X1 U16268 ( .A1(n14433), .A2(n12704), .ZN(n12710) );
  INV_X1 U16269 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20781) );
  AOI22_X1 U16270 ( .A1(n12705), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12706) );
  OAI21_X1 U16271 ( .B1(n12707), .B2(n20781), .A(n12706), .ZN(n12708) );
  AOI21_X1 U16272 ( .B1(n9758), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12708), .ZN(n12709) );
  NAND2_X1 U16273 ( .A1(n13045), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13048) );
  INV_X1 U16274 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13052) );
  INV_X1 U16275 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13061) );
  INV_X1 U16276 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13065) );
  NAND2_X1 U16277 ( .A1(n13114), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12712) );
  NAND2_X1 U16278 ( .A1(n13006), .A2(n16924), .ZN(n12714) );
  NOR2_X1 U16279 ( .A1(n16877), .A2(n20781), .ZN(n12988) );
  AOI21_X1 U16280 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n12988), .ZN(n12713) );
  AND2_X1 U16281 ( .A1(n12714), .A2(n12713), .ZN(n12715) );
  INV_X1 U16282 ( .A(n12716), .ZN(n12730) );
  NAND2_X1 U16283 ( .A1(n12719), .A2(n12718), .ZN(n12723) );
  MUX2_X1 U16284 ( .A(n12726), .B(n12725), .S(n20166), .Z(n14562) );
  NAND2_X1 U16285 ( .A1(n14562), .A2(n11864), .ZN(n12727) );
  XOR2_X1 U16286 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12727), .Z(
        n12728) );
  NAND2_X1 U16287 ( .A1(n12995), .A2(n16899), .ZN(n12729) );
  AOI22_X1 U16288 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U16289 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U16290 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12732) );
  OAI21_X1 U16291 ( .B1(n12733), .B2(n21817), .A(n12732), .ZN(n12739) );
  AOI22_X1 U16292 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U16293 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U16294 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U16295 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12734) );
  NAND4_X1 U16296 ( .A1(n12737), .A2(n12736), .A3(n12735), .A4(n12734), .ZN(
        n12738) );
  AOI211_X1 U16297 ( .C1(n18334), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n12739), .B(n12738), .ZN(n12740) );
  NAND3_X1 U16298 ( .A1(n12742), .A2(n12741), .A3(n12740), .ZN(n12893) );
  AOI22_X1 U16299 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U16300 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12746) );
  AOI22_X1 U16301 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U16302 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12744) );
  NAND4_X1 U16303 ( .A1(n12747), .A2(n12746), .A3(n12745), .A4(n12744), .ZN(
        n12753) );
  AOI22_X1 U16304 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U16305 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12768), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U16306 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U16307 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17439), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12748) );
  NAND4_X1 U16308 ( .A1(n12751), .A2(n12750), .A3(n12749), .A4(n12748), .ZN(
        n12752) );
  AOI22_X1 U16309 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U16310 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12768), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U16311 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U16312 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12754) );
  NAND4_X1 U16313 ( .A1(n12757), .A2(n12756), .A3(n12755), .A4(n12754), .ZN(
        n12763) );
  AOI22_X1 U16314 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U16315 ( .A1(n18312), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18343), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U16316 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U16317 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12758) );
  NAND4_X1 U16318 ( .A1(n12761), .A2(n12760), .A3(n12759), .A4(n12758), .ZN(
        n12762) );
  AOI22_X1 U16319 ( .A1(n12808), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12819), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U16320 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n18212), .ZN(n12766) );
  AOI22_X1 U16321 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n9744), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n12816), .ZN(n12765) );
  AOI22_X1 U16322 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12818), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12764) );
  NAND4_X1 U16323 ( .A1(n12767), .A2(n12766), .A3(n12765), .A4(n12764), .ZN(
        n12774) );
  AOI22_X1 U16324 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12815), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n12768), .ZN(n12772) );
  AOI22_X1 U16325 ( .A1(n12731), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18343), .ZN(n12771) );
  AOI22_X1 U16326 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n12809), .ZN(n12769) );
  NAND4_X1 U16327 ( .A1(n12772), .A2(n12771), .A3(n12770), .A4(n12769), .ZN(
        n12773) );
  AOI22_X1 U16328 ( .A1(n12731), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9743), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12775) );
  OAI21_X1 U16329 ( .B1(n9732), .B2(n18381), .A(n12775), .ZN(n12780) );
  AOI22_X1 U16330 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12815), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U16331 ( .A1(n12818), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10901), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12777) );
  NAND3_X1 U16332 ( .A1(n12778), .A2(n12777), .A3(n12776), .ZN(n12779) );
  AOI22_X1 U16333 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18284), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U16334 ( .A1(n12808), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12809), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U16335 ( .A1(n12807), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12768), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12782) );
  AOI22_X1 U16336 ( .A1(n12819), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18343), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12781) );
  NAND2_X2 U16337 ( .A1(n12786), .A2(n12785), .ZN(n18532) );
  NAND2_X1 U16338 ( .A1(n18536), .A2(n18532), .ZN(n12829) );
  AOI22_X1 U16339 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U16340 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U16341 ( .A1(n18333), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12787) );
  OAI21_X1 U16342 ( .B1(n9732), .B2(n18370), .A(n12787), .ZN(n12793) );
  AOI22_X1 U16343 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12815), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U16344 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U16345 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U16346 ( .A1(n18312), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12810), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12788) );
  NAND4_X1 U16347 ( .A1(n12791), .A2(n12790), .A3(n12789), .A4(n12788), .ZN(
        n12792) );
  AOI211_X1 U16348 ( .C1(n18321), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n12793), .B(n12792), .ZN(n12794) );
  NAND3_X1 U16349 ( .A1(n12796), .A2(n12795), .A3(n12794), .ZN(n12892) );
  NAND2_X1 U16350 ( .A1(n12830), .A2(n12892), .ZN(n12833) );
  AOI22_X1 U16351 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U16352 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U16353 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12798) );
  AOI22_X1 U16354 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12797) );
  NAND4_X1 U16355 ( .A1(n12800), .A2(n12799), .A3(n12798), .A4(n12797), .ZN(
        n12806) );
  AOI22_X1 U16356 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U16357 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U16358 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U16359 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12801) );
  NAND4_X1 U16360 ( .A1(n12804), .A2(n12803), .A3(n12802), .A4(n12801), .ZN(
        n12805) );
  NOR2_X1 U16361 ( .A1(n18536), .A2(n10622), .ZN(n12826) );
  AOI22_X1 U16362 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12807), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U16363 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12808), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U16364 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12768), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U16365 ( .A1(n12810), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12809), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12811) );
  NAND4_X1 U16366 ( .A1(n12814), .A2(n12813), .A3(n12812), .A4(n12811), .ZN(
        n12825) );
  AOI22_X1 U16367 ( .A1(n12731), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12815), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U16368 ( .A1(n12817), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12816), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U16369 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12818), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U16370 ( .A1(n12819), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18343), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12820) );
  NAND4_X1 U16371 ( .A1(n12823), .A2(n12822), .A3(n12821), .A4(n12820), .ZN(
        n12824) );
  NAND2_X1 U16372 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n9733), .ZN(
        n19008) );
  NOR2_X1 U16373 ( .A1(n19303), .A2(n12827), .ZN(n12828) );
  XNOR2_X1 U16374 ( .A(n18524), .B(n12829), .ZN(n18976) );
  INV_X1 U16375 ( .A(n12892), .ZN(n18520) );
  XNOR2_X1 U16376 ( .A(n18520), .B(n12830), .ZN(n12831) );
  XNOR2_X1 U16377 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12831), .ZN(
        n18969) );
  AND2_X1 U16378 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12831), .ZN(
        n12832) );
  NOR2_X2 U16379 ( .A1(n18968), .A2(n12832), .ZN(n18953) );
  XNOR2_X1 U16380 ( .A(n18516), .B(n12833), .ZN(n18954) );
  NAND2_X1 U16381 ( .A1(n18953), .A2(n18954), .ZN(n18952) );
  XOR2_X1 U16382 ( .A(n18513), .B(n12834), .Z(n12835) );
  XNOR2_X1 U16383 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12835), .ZN(
        n18939) );
  NAND2_X1 U16384 ( .A1(n19207), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19181) );
  INV_X1 U16385 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19174) );
  NAND2_X1 U16386 ( .A1(n19134), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19120) );
  NAND2_X1 U16387 ( .A1(n19227), .A2(n18895), .ZN(n18891) );
  NOR4_X1 U16388 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n18891), .ZN(n12842) );
  NOR2_X1 U16389 ( .A1(n19136), .A2(n19127), .ZN(n19116) );
  NOR2_X1 U16390 ( .A1(n21877), .A2(n19070), .ZN(n18754) );
  INV_X1 U16391 ( .A(n18754), .ZN(n19091) );
  NOR2_X1 U16392 ( .A1(n21959), .A2(n19091), .ZN(n19076) );
  NAND2_X1 U16393 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n19076), .ZN(
        n18741) );
  NAND2_X1 U16394 ( .A1(n19077), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n19015) );
  INV_X1 U16395 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19014) );
  NOR2_X1 U16396 ( .A1(n19015), .A2(n19014), .ZN(n18714) );
  NAND2_X1 U16397 ( .A1(n18790), .A2(n21877), .ZN(n12845) );
  NAND2_X1 U16398 ( .A1(n18753), .A2(n21959), .ZN(n18740) );
  INV_X1 U16399 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19084) );
  NAND2_X1 U16400 ( .A1(n12848), .A2(n19116), .ZN(n18751) );
  INV_X1 U16401 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19042) );
  INV_X1 U16402 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12851) );
  NAND2_X1 U16403 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19018) );
  NAND2_X1 U16404 ( .A1(n18920), .A2(n19018), .ZN(n12849) );
  NAND2_X1 U16405 ( .A1(n18701), .A2(n12849), .ZN(n12850) );
  INV_X1 U16406 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18655) );
  NAND2_X1 U16407 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12919) );
  INV_X1 U16408 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17631) );
  NOR2_X1 U16409 ( .A1(n12919), .A2(n17631), .ZN(n13102) );
  INV_X1 U16410 ( .A(n13102), .ZN(n12932) );
  AOI21_X1 U16411 ( .B1(n13086), .B2(n9755), .A(n13089), .ZN(n12853) );
  INV_X1 U16412 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12943) );
  NOR2_X1 U16413 ( .A1(n10829), .A2(n13096), .ZN(n12931) );
  NOR2_X1 U16414 ( .A1(n19987), .A2(n12854), .ZN(n12863) );
  NAND2_X1 U16415 ( .A1(n12863), .A2(n18391), .ZN(n12858) );
  NOR2_X1 U16416 ( .A1(n12856), .A2(n12855), .ZN(n12857) );
  OAI211_X1 U16417 ( .C1(n19363), .C2(n19793), .A(n12885), .B(n12857), .ZN(
        n12866) );
  INV_X1 U16418 ( .A(n12858), .ZN(n12870) );
  OAI21_X1 U16419 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19797), .A(
        n12859), .ZN(n12872) );
  INV_X1 U16420 ( .A(n12872), .ZN(n12861) );
  OAI21_X1 U16421 ( .B1(n12861), .B2(n12860), .A(n12874), .ZN(n19817) );
  OAI21_X1 U16422 ( .B1(n19355), .B2(n18596), .A(n19986), .ZN(n12862) );
  OAI21_X1 U16423 ( .B1(n12863), .B2(n12862), .A(n19981), .ZN(n17732) );
  NOR3_X1 U16424 ( .A1(n12884), .A2(n17478), .A3(n17732), .ZN(n12869) );
  OAI21_X1 U16425 ( .B1(n12866), .B2(n12865), .A(n12864), .ZN(n12868) );
  NAND2_X1 U16426 ( .A1(n12868), .A2(n12867), .ZN(n17479) );
  NOR2_X1 U16427 ( .A1(n12872), .A2(n12871), .ZN(n12876) );
  INV_X1 U16428 ( .A(n12873), .ZN(n12875) );
  OAI21_X1 U16429 ( .B1(n12877), .B2(n14380), .A(n19816), .ZN(n12878) );
  NAND2_X1 U16430 ( .A1(n12931), .A2(n19239), .ZN(n12930) );
  NOR2_X1 U16431 ( .A1(n17635), .A2(n19297), .ZN(n19240) );
  INV_X1 U16432 ( .A(n19015), .ZN(n19029) );
  NAND3_X1 U16433 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18686) );
  NOR2_X1 U16434 ( .A1(n12851), .A2(n18686), .ZN(n12922) );
  NAND2_X1 U16435 ( .A1(n19029), .A2(n12922), .ZN(n19024) );
  INV_X1 U16436 ( .A(n19024), .ZN(n12886) );
  INV_X1 U16437 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19143) );
  NAND2_X1 U16438 ( .A1(n19134), .A2(n19177), .ZN(n18839) );
  NAND2_X1 U16439 ( .A1(n12886), .A2(n19141), .ZN(n19019) );
  NOR2_X1 U16440 ( .A1(n12919), .A2(n19019), .ZN(n17637) );
  OAI21_X1 U16441 ( .B1(n12885), .B2(n12883), .A(n12882), .ZN(n19778) );
  NOR2_X1 U16442 ( .A1(n19363), .A2(n18391), .ZN(n19780) );
  NAND3_X1 U16443 ( .A1(n12885), .A2(n12884), .A3(n19780), .ZN(n14382) );
  INV_X1 U16444 ( .A(n19812), .ZN(n19299) );
  INV_X1 U16445 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19255) );
  NAND3_X1 U16446 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19229) );
  NOR4_X1 U16447 ( .A1(n19251), .A2(n19255), .A3(n19233), .A4(n19229), .ZN(
        n19118) );
  INV_X1 U16448 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19964) );
  OAI21_X1 U16449 ( .B1(n19964), .B2(n10622), .A(n19303), .ZN(n19272) );
  NAND2_X1 U16450 ( .A1(n19118), .A2(n19272), .ZN(n19157) );
  OR2_X1 U16451 ( .A1(n19120), .A2(n19157), .ZN(n19112) );
  NOR2_X1 U16452 ( .A1(n19299), .A2(n19112), .ZN(n17645) );
  NOR2_X1 U16453 ( .A1(n19303), .A2(n10622), .ZN(n19271) );
  NAND2_X1 U16454 ( .A1(n19271), .A2(n19118), .ZN(n19178) );
  NOR2_X1 U16455 ( .A1(n19120), .A2(n19178), .ZN(n19068) );
  INV_X1 U16456 ( .A(n19068), .ZN(n19016) );
  NOR2_X1 U16457 ( .A1(n19964), .A2(n19016), .ZN(n19131) );
  OAI221_X1 U16458 ( .B1(n19792), .B2(n17645), .C1(n19131), .C2(n17645), .A(
        n12886), .ZN(n12887) );
  INV_X1 U16459 ( .A(n12887), .ZN(n12890) );
  NOR2_X1 U16460 ( .A1(n19024), .A2(n19016), .ZN(n12925) );
  OAI221_X1 U16461 ( .B1(n12890), .B2(n12925), .C1(n12890), .C2(n19326), .A(
        n19327), .ZN(n13105) );
  NAND2_X1 U16462 ( .A1(n19811), .A2(n19327), .ZN(n19288) );
  NOR2_X1 U16463 ( .A1(n12900), .A2(n18532), .ZN(n12898) );
  NOR2_X1 U16464 ( .A1(n12898), .A2(n18524), .ZN(n12907) );
  NAND2_X1 U16465 ( .A1(n12907), .A2(n12892), .ZN(n12896) );
  NOR2_X1 U16466 ( .A1(n18516), .A2(n12896), .ZN(n12895) );
  NAND2_X1 U16467 ( .A1(n12895), .A2(n12893), .ZN(n12894) );
  NOR2_X1 U16468 ( .A1(n18510), .A2(n12894), .ZN(n12916) );
  XNOR2_X1 U16469 ( .A(n12894), .B(n17635), .ZN(n18926) );
  XNOR2_X1 U16470 ( .A(n12895), .B(n18513), .ZN(n12910) );
  XOR2_X1 U16471 ( .A(n12896), .B(n18516), .Z(n12897) );
  NAND2_X1 U16472 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12897), .ZN(
        n12909) );
  INV_X1 U16473 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21839) );
  XNOR2_X1 U16474 ( .A(n21839), .B(n12897), .ZN(n18951) );
  XOR2_X1 U16475 ( .A(n18524), .B(n12898), .Z(n12899) );
  NAND2_X1 U16476 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12899), .ZN(
        n12905) );
  INV_X1 U16477 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19289) );
  XNOR2_X1 U16478 ( .A(n19289), .B(n12899), .ZN(n19286) );
  OR2_X1 U16479 ( .A1(n19303), .A2(n12901), .ZN(n12904) );
  XNOR2_X1 U16480 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12901), .ZN(
        n18992) );
  AOI21_X1 U16481 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18536), .A(
        n9733), .ZN(n12903) );
  NOR2_X1 U16482 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18536), .ZN(
        n12902) );
  AOI221_X1 U16483 ( .B1(n9733), .B2(n18536), .C1(n12903), .C2(n19964), .A(
        n12902), .ZN(n18991) );
  NAND2_X1 U16484 ( .A1(n18992), .A2(n18991), .ZN(n18990) );
  NAND2_X1 U16485 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12906), .ZN(
        n12908) );
  XNOR2_X1 U16486 ( .A(n12907), .B(n18520), .ZN(n18964) );
  NAND2_X1 U16487 ( .A1(n18951), .A2(n18950), .ZN(n18949) );
  NAND2_X1 U16488 ( .A1(n12909), .A2(n18949), .ZN(n12911) );
  NAND2_X1 U16489 ( .A1(n12910), .A2(n12911), .ZN(n12912) );
  XOR2_X1 U16490 ( .A(n12911), .B(n12910), .Z(n18943) );
  NAND2_X1 U16491 ( .A1(n18943), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18942) );
  NAND2_X1 U16492 ( .A1(n12916), .A2(n12913), .ZN(n12917) );
  NAND2_X1 U16493 ( .A1(n18926), .A2(n18927), .ZN(n18925) );
  NAND2_X1 U16494 ( .A1(n12916), .A2(n12915), .ZN(n12914) );
  OAI211_X1 U16495 ( .C1(n12916), .C2(n12915), .A(n18925), .B(n12914), .ZN(
        n18911) );
  INV_X1 U16496 ( .A(n12919), .ZN(n12918) );
  NAND2_X1 U16497 ( .A1(n18656), .A2(n12918), .ZN(n17641) );
  OAI22_X1 U16498 ( .A1(n13105), .A2(n12919), .B1(n19288), .B2(n17641), .ZN(
        n12920) );
  AOI21_X1 U16499 ( .B1(n19240), .B2(n17637), .A(n12920), .ZN(n17494) );
  NOR3_X1 U16500 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17494), .A3(
        n17631), .ZN(n12921) );
  NOR2_X1 U16501 ( .A1(n19328), .A2(n19921), .ZN(n12936) );
  NOR2_X1 U16502 ( .A1(n12932), .A2(n19019), .ZN(n13100) );
  INV_X1 U16503 ( .A(n13100), .ZN(n12942) );
  INV_X1 U16504 ( .A(n19288), .ZN(n19333) );
  NAND2_X1 U16505 ( .A1(n18656), .A2(n13102), .ZN(n12941) );
  AOI22_X1 U16506 ( .A1(n19240), .A2(n12942), .B1(n19333), .B2(n12941), .ZN(
        n17488) );
  OAI21_X1 U16507 ( .B1(n19024), .B2(n19112), .A(n19812), .ZN(n12924) );
  NAND2_X1 U16508 ( .A1(n19029), .A2(n19131), .ZN(n19074) );
  NAND2_X1 U16509 ( .A1(n12922), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17646) );
  OAI21_X1 U16510 ( .B1(n19074), .B2(n17646), .A(n19792), .ZN(n12923) );
  OAI211_X1 U16511 ( .C1(n19794), .C2(n12925), .A(n12924), .B(n12923), .ZN(
        n17486) );
  INV_X1 U16512 ( .A(n19270), .ZN(n19234) );
  OAI21_X1 U16513 ( .B1(n19234), .B2(n13102), .A(n19327), .ZN(n12926) );
  OAI21_X1 U16514 ( .B1(n17486), .B2(n12926), .A(n19328), .ZN(n13103) );
  AOI21_X1 U16515 ( .B1(n17488), .B2(n13103), .A(n12943), .ZN(n12927) );
  NAND2_X1 U16516 ( .A1(n12930), .A2(n12929), .ZN(P3_U2832) );
  NAND2_X1 U16517 ( .A1(n12931), .A2(n18921), .ZN(n12947) );
  NOR4_X1 U16518 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19024), .A3(
        n12932), .A4(n18819), .ZN(n12940) );
  INV_X1 U16519 ( .A(n20002), .ZN(n19949) );
  NAND2_X1 U16520 ( .A1(n20001), .A2(n19937), .ZN(n17730) );
  NAND2_X1 U16521 ( .A1(n19949), .A2(n17730), .ZN(n17470) );
  AOI21_X1 U16522 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19995), .ZN(n19845) );
  OAI21_X1 U16523 ( .B1(n19006), .B2(n18692), .A(n19369), .ZN(n18772) );
  INV_X1 U16524 ( .A(n18772), .ZN(n18846) );
  OR2_X1 U16525 ( .A1(n12933), .A2(n18846), .ZN(n13131) );
  NOR2_X1 U16526 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18692), .ZN(
        n17621) );
  INV_X1 U16527 ( .A(n18732), .ZN(n19848) );
  NAND2_X1 U16528 ( .A1(n19659), .A2(n12933), .ZN(n17625) );
  OAI211_X1 U16529 ( .C1(n12935), .C2(n19848), .A(n19009), .B(n17625), .ZN(
        n17620) );
  NOR2_X1 U16530 ( .A1(n17621), .A2(n17620), .ZN(n13129) );
  NAND2_X1 U16531 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18981) );
  NAND2_X2 U16532 ( .A1(n18981), .A2(n19009), .ZN(n18901) );
  AOI21_X1 U16533 ( .B1(n18865), .B2(n12968), .A(n12936), .ZN(n12937) );
  OAI221_X1 U16534 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n13131), .C1(
        n12938), .C2(n13129), .A(n12937), .ZN(n12939) );
  NAND2_X1 U16535 ( .A1(n18999), .A2(n12941), .ZN(n17619) );
  NAND2_X1 U16536 ( .A1(n18922), .A2(n12942), .ZN(n17632) );
  AOI21_X1 U16537 ( .B1(n17619), .B2(n17632), .A(n12943), .ZN(n12944) );
  NAND2_X1 U16538 ( .A1(n12947), .A2(n12946), .ZN(P3_U2800) );
  NAND2_X1 U16539 ( .A1(n12949), .A2(n12948), .ZN(n12950) );
  NAND2_X1 U16540 ( .A1(n15724), .A2(n12950), .ZN(n16591) );
  INV_X1 U16541 ( .A(n12957), .ZN(n17152) );
  AND2_X1 U16542 ( .A1(n17225), .A2(n17152), .ZN(n12951) );
  NAND2_X1 U16543 ( .A1(n12958), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12953) );
  NAND2_X1 U16544 ( .A1(n17225), .A2(n12953), .ZN(n12954) );
  NAND2_X1 U16545 ( .A1(n17143), .A2(n12954), .ZN(n17105) );
  AND2_X1 U16546 ( .A1(n17225), .A2(n12959), .ZN(n12956) );
  OR3_X1 U16547 ( .A1(n17105), .A2(n12956), .A3(n12955), .ZN(n17070) );
  AND2_X1 U16548 ( .A1(n17070), .A2(n12985), .ZN(n17057) );
  XNOR2_X1 U16549 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12960) );
  NOR2_X1 U16550 ( .A1(n17046), .A2(n16857), .ZN(n17164) );
  NAND2_X1 U16551 ( .A1(n17112), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17108) );
  NOR2_X1 U16552 ( .A1(n17108), .A2(n12959), .ZN(n17071) );
  NAND2_X1 U16553 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17071), .ZN(
        n17061) );
  NOR2_X1 U16554 ( .A1(n12960), .A2(n17061), .ZN(n12961) );
  AOI211_X1 U16555 ( .C1(n17057), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12962), .B(n12961), .ZN(n12963) );
  OAI21_X1 U16556 ( .B1(n16591), .B2(n17256), .A(n12963), .ZN(n12964) );
  OAI211_X1 U16557 ( .C1(n12966), .C2(n17266), .A(n12965), .B(n9875), .ZN(
        P2_U3026) );
  NAND2_X1 U16558 ( .A1(n18017), .A2(n18067), .ZN(n18077) );
  NOR3_X1 U16559 ( .A1(n12968), .A2(n12967), .A3(n18077), .ZN(n12981) );
  INV_X1 U16560 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n18103) );
  NAND2_X1 U16561 ( .A1(n12969), .A2(n18103), .ZN(n12979) );
  INV_X1 U16562 ( .A(n12970), .ZN(n12971) );
  INV_X1 U16563 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19919) );
  AOI21_X1 U16564 ( .B1(n17755), .B2(n12971), .A(n19919), .ZN(n12977) );
  NOR3_X1 U16565 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19921), .A3(n12972), 
        .ZN(n12973) );
  AOI21_X1 U16566 ( .B1(n18074), .B2(P3_EBX_REG_31__SCAN_IN), .A(n12973), .ZN(
        n12975) );
  INV_X1 U16567 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13128) );
  OR2_X1 U16568 ( .A1(n18076), .A2(n13128), .ZN(n12974) );
  NAND2_X1 U16569 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  NOR2_X1 U16570 ( .A1(n12977), .A2(n12976), .ZN(n12978) );
  NAND2_X1 U16571 ( .A1(n12979), .A2(n12978), .ZN(n12980) );
  AOI222_X1 U16572 ( .A1(n11647), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12982), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n11456), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n12983) );
  NAND3_X1 U16573 ( .A1(n12986), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12985), .ZN(n12992) );
  NOR2_X1 U16574 ( .A1(n12987), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12989) );
  AOI21_X1 U16575 ( .B1(n12990), .B2(n12989), .A(n12988), .ZN(n12991) );
  NOR2_X1 U16576 ( .A1(n16017), .A2(n17241), .ZN(n12996) );
  OAI211_X1 U16577 ( .C1(n12999), .C2(n17234), .A(n12998), .B(n12997), .ZN(
        P2_U3015) );
  OAI21_X1 U16578 ( .B1(n15623), .B2(n13000), .A(n14434), .ZN(n16964) );
  NAND2_X1 U16579 ( .A1(n20146), .A2(n20850), .ZN(n13001) );
  NAND2_X1 U16580 ( .A1(n13002), .A2(n13003), .ZN(n13004) );
  NAND2_X1 U16581 ( .A1(n14430), .A2(n13004), .ZN(n16963) );
  NAND2_X1 U16582 ( .A1(n13809), .A2(n20481), .ZN(n17367) );
  INV_X1 U16583 ( .A(n13007), .ZN(n13010) );
  INV_X1 U16584 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13008) );
  NAND2_X1 U16585 ( .A1(n15991), .A2(n13008), .ZN(n13009) );
  NAND2_X1 U16586 ( .A1(n13010), .A2(n13009), .ZN(n15976) );
  OAI21_X1 U16587 ( .B1(n13007), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13011), .ZN(n16932) );
  AND2_X1 U16588 ( .A1(n13011), .A2(n16920), .ZN(n13013) );
  NOR2_X1 U16589 ( .A1(n13012), .A2(n13013), .ZN(n16923) );
  NOR2_X1 U16590 ( .A1(n15950), .A2(n16923), .ZN(n15930) );
  OR2_X1 U16591 ( .A1(n13012), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13015) );
  NAND2_X1 U16592 ( .A1(n13014), .A2(n13015), .ZN(n16906) );
  NAND2_X1 U16593 ( .A1(n15930), .A2(n16906), .ZN(n20058) );
  NAND2_X1 U16594 ( .A1(n13014), .A2(n10665), .ZN(n13016) );
  AND2_X1 U16595 ( .A1(n13018), .A2(n13016), .ZN(n20061) );
  OR2_X1 U16596 ( .A1(n20058), .A2(n20061), .ZN(n15915) );
  AND2_X1 U16597 ( .A1(n13018), .A2(n16887), .ZN(n13019) );
  NOR2_X1 U16598 ( .A1(n13017), .A2(n13019), .ZN(n16889) );
  NOR2_X1 U16599 ( .A1(n15915), .A2(n16889), .ZN(n15898) );
  NOR2_X1 U16600 ( .A1(n13017), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13021) );
  OR2_X1 U16601 ( .A1(n13020), .A2(n13021), .ZN(n16878) );
  OR2_X1 U16602 ( .A1(n13020), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13023) );
  NAND2_X1 U16603 ( .A1(n13022), .A2(n13023), .ZN(n16861) );
  NAND2_X1 U16604 ( .A1(n13022), .A2(n16842), .ZN(n13025) );
  AND2_X1 U16605 ( .A1(n13024), .A2(n13025), .ZN(n16845) );
  NAND2_X1 U16606 ( .A1(n13024), .A2(n10659), .ZN(n13026) );
  AND2_X1 U16607 ( .A1(n13027), .A2(n13026), .ZN(n16833) );
  AND2_X1 U16608 ( .A1(n13027), .A2(n15851), .ZN(n13028) );
  OR2_X1 U16609 ( .A1(n13028), .A2(n13029), .ZN(n16819) );
  AND2_X1 U16610 ( .A1(n15845), .A2(n16819), .ZN(n15833) );
  OR2_X1 U16611 ( .A1(n13029), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13030) );
  NAND2_X1 U16612 ( .A1(n13032), .A2(n13030), .ZN(n16810) );
  NAND2_X1 U16613 ( .A1(n13032), .A2(n16800), .ZN(n13033) );
  AND2_X1 U16614 ( .A1(n13035), .A2(n13033), .ZN(n16798) );
  AND2_X1 U16615 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  OR2_X1 U16616 ( .A1(n13036), .A2(n13038), .ZN(n20045) );
  INV_X1 U16617 ( .A(n20045), .ZN(n20037) );
  NOR2_X1 U16618 ( .A1(n13038), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13039) );
  OR2_X1 U16619 ( .A1(n13037), .A2(n13039), .ZN(n16773) );
  XNOR2_X1 U16620 ( .A(n13037), .B(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16767) );
  NAND2_X1 U16621 ( .A1(n15788), .A2(n16767), .ZN(n15777) );
  NAND2_X1 U16622 ( .A1(n13037), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13040) );
  INV_X1 U16623 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16761) );
  NAND2_X1 U16624 ( .A1(n13040), .A2(n16761), .ZN(n13041) );
  AND2_X1 U16625 ( .A1(n13041), .A2(n13043), .ZN(n16759) );
  NAND2_X1 U16626 ( .A1(n13043), .A2(n13042), .ZN(n13044) );
  NAND2_X1 U16627 ( .A1(n12020), .A2(n13044), .ZN(n16747) );
  NAND2_X1 U16628 ( .A1(n15730), .A2(n20059), .ZN(n13047) );
  NOR2_X1 U16629 ( .A1(n12711), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13046) );
  OR2_X1 U16630 ( .A1(n13045), .A2(n13046), .ZN(n16738) );
  NAND2_X1 U16631 ( .A1(n13047), .A2(n16738), .ZN(n15715) );
  NAND2_X1 U16632 ( .A1(n15715), .A2(n20059), .ZN(n13050) );
  OR2_X1 U16633 ( .A1(n13045), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13049) );
  NAND2_X1 U16634 ( .A1(n13048), .A2(n13049), .ZN(n16719) );
  NAND2_X1 U16635 ( .A1(n13050), .A2(n16719), .ZN(n15699) );
  NAND2_X1 U16636 ( .A1(n13048), .A2(n15698), .ZN(n13051) );
  NAND2_X1 U16637 ( .A1(n13053), .A2(n13051), .ZN(n16708) );
  NAND2_X1 U16638 ( .A1(n13053), .A2(n13052), .ZN(n13054) );
  NAND2_X1 U16639 ( .A1(n13055), .A2(n13054), .ZN(n16703) );
  NAND2_X1 U16640 ( .A1(n15665), .A2(n20059), .ZN(n13057) );
  AND2_X1 U16641 ( .A1(n13055), .A2(n15664), .ZN(n13056) );
  OR2_X1 U16642 ( .A1(n13056), .A2(n13058), .ZN(n16690) );
  NAND2_X1 U16643 ( .A1(n13057), .A2(n16690), .ZN(n15643) );
  NAND2_X1 U16644 ( .A1(n15643), .A2(n20059), .ZN(n13060) );
  OR2_X1 U16645 ( .A1(n13058), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13059) );
  NAND2_X1 U16646 ( .A1(n9939), .A2(n13059), .ZN(n16678) );
  NAND2_X1 U16647 ( .A1(n13060), .A2(n16678), .ZN(n15629) );
  NAND2_X1 U16648 ( .A1(n15629), .A2(n20059), .ZN(n13063) );
  NAND2_X1 U16649 ( .A1(n9939), .A2(n13061), .ZN(n13062) );
  NAND2_X1 U16650 ( .A1(n9917), .A2(n13062), .ZN(n16667) );
  AND2_X1 U16651 ( .A1(n9917), .A2(n13065), .ZN(n13066) );
  NOR2_X1 U16652 ( .A1(n13064), .A2(n13066), .ZN(n16655) );
  NAND2_X1 U16653 ( .A1(n13067), .A2(n16655), .ZN(n13071) );
  INV_X1 U16654 ( .A(n13068), .ZN(n13070) );
  NOR2_X1 U16655 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13069) );
  NAND2_X1 U16656 ( .A1(n13070), .A2(n13069), .ZN(n20062) );
  AOI21_X1 U16657 ( .B1(n13071), .B2(n15999), .A(n20038), .ZN(n13072) );
  NOR2_X1 U16658 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20844), .ZN(n13073) );
  NOR2_X1 U16659 ( .A1(n13803), .A2(n13073), .ZN(n13078) );
  INV_X1 U16660 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13077) );
  NOR2_X1 U16661 ( .A1(n20854), .A2(n13077), .ZN(n13074) );
  INV_X1 U16662 ( .A(n16003), .ZN(n20053) );
  NAND2_X1 U16663 ( .A1(n13963), .A2(n17372), .ZN(n13075) );
  OR2_X1 U16664 ( .A1(n11426), .A2(n13075), .ZN(n16010) );
  NOR2_X1 U16665 ( .A1(n20814), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20552) );
  NAND3_X1 U16666 ( .A1(n17365), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20552), 
        .ZN(n17607) );
  AND3_X1 U16667 ( .A1(n20062), .A2(n16877), .A3(n17607), .ZN(n13076) );
  NAND2_X1 U16668 ( .A1(n14556), .A2(n17367), .ZN(n13080) );
  NAND2_X1 U16669 ( .A1(n13078), .A2(n13077), .ZN(n13079) );
  NAND2_X2 U16670 ( .A1(n13080), .A2(n13079), .ZN(n20032) );
  AOI22_X1 U16671 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_28__SCAN_IN), .ZN(n13082) );
  NAND2_X1 U16672 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13081) );
  OAI211_X1 U16673 ( .C1(n13083), .C2(n20053), .A(n13082), .B(n13081), .ZN(
        n13084) );
  INV_X1 U16674 ( .A(n13084), .ZN(n13085) );
  NAND4_X1 U16675 ( .A1(n10798), .A2(n9844), .A3(n10797), .A4(n13085), .ZN(
        P2_U2827) );
  INV_X1 U16676 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19945) );
  NAND2_X1 U16677 ( .A1(n19945), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13087) );
  NAND2_X1 U16678 ( .A1(n13088), .A2(n13087), .ZN(n13091) );
  NOR2_X1 U16679 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19945), .ZN(
        n13107) );
  AOI22_X1 U16680 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n9755), .B1(
        n18920), .B2(n19945), .ZN(n13093) );
  NAND2_X1 U16681 ( .A1(n13092), .A2(n13093), .ZN(n13098) );
  INV_X1 U16682 ( .A(n13093), .ZN(n13094) );
  OAI21_X1 U16683 ( .B1(n13096), .B2(n13095), .A(n13094), .ZN(n13097) );
  NAND2_X1 U16684 ( .A1(n13098), .A2(n13097), .ZN(n13127) );
  NAND2_X1 U16685 ( .A1(n13127), .A2(n19239), .ZN(n13113) );
  NAND3_X1 U16686 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n13102), .A3(
        n18656), .ZN(n13099) );
  XOR2_X1 U16687 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13099), .Z(
        n13135) );
  NAND2_X1 U16688 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n13100), .ZN(
        n13101) );
  XNOR2_X1 U16689 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13101), .ZN(
        n13134) );
  NOR2_X1 U16690 ( .A1(n19234), .A2(n19314), .ZN(n19321) );
  NOR2_X1 U16691 ( .A1(n19919), .A2(n19328), .ZN(n13133) );
  NAND3_X1 U16692 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n13102), .A3(
        n19945), .ZN(n13104) );
  OAI22_X1 U16693 ( .A1(n13105), .A2(n13104), .B1(n19945), .B2(n13103), .ZN(
        n13106) );
  AOI211_X1 U16694 ( .C1(n13107), .C2(n19321), .A(n13133), .B(n13106), .ZN(
        n13108) );
  OAI21_X1 U16695 ( .B1(n13135), .B2(n19288), .A(n13110), .ZN(n13111) );
  NAND2_X1 U16696 ( .A1(n13113), .A2(n13112), .ZN(P3_U2831) );
  NOR2_X1 U16697 ( .A1(n13064), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13115) );
  OR2_X1 U16698 ( .A1(n13114), .A2(n13115), .ZN(n16643) );
  INV_X1 U16699 ( .A(n14560), .ZN(n14436) );
  XNOR2_X1 U16700 ( .A(n13114), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14470) );
  NAND2_X1 U16701 ( .A1(n15975), .A2(n14470), .ZN(n14559) );
  INV_X1 U16702 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U16703 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_30__SCAN_IN), .ZN(n13116) );
  OAI21_X1 U16704 ( .B1(n20073), .B2(n13117), .A(n13116), .ZN(n13118) );
  AOI21_X1 U16705 ( .B1(n13119), .B2(n16003), .A(n13118), .ZN(n13120) );
  OAI21_X1 U16706 ( .B1(n14436), .B2(n14559), .A(n13120), .ZN(n13124) );
  INV_X1 U16707 ( .A(n14470), .ZN(n13121) );
  NAND3_X1 U16708 ( .A1(n10811), .A2(n13126), .A3(n13125), .ZN(P2_U2825) );
  NAND2_X1 U16709 ( .A1(n13127), .A2(n18921), .ZN(n13138) );
  XOR2_X1 U16710 ( .A(n13128), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n13130) );
  OAI22_X1 U16711 ( .A1(n13131), .A2(n13130), .B1(n13129), .B2(n13128), .ZN(
        n13132) );
  AOI211_X1 U16712 ( .C1(n18865), .C2(n18017), .A(n13133), .B(n13132), .ZN(
        n13137) );
  NAND2_X1 U16713 ( .A1(n13134), .A2(n18922), .ZN(n13136) );
  NAND2_X1 U16714 ( .A1(n13138), .A2(n10827), .ZN(P3_U2799) );
  INV_X1 U16715 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13139) );
  XNOR2_X1 U16716 ( .A(n13139), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20966) );
  NAND2_X1 U16717 ( .A1(n21647), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13256) );
  OAI21_X1 U16718 ( .B1(n20966), .B2(n14398), .A(n13256), .ZN(n13140) );
  AOI21_X1 U16719 ( .B1(n13627), .B2(P1_EAX_REG_2__SCAN_IN), .A(n13140), .ZN(
        n13141) );
  AND2_X1 U16720 ( .A1(n13142), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U16721 ( .A1(n13742), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13162) );
  NAND2_X1 U16722 ( .A1(n15564), .A2(n13335), .ZN(n13153) );
  NAND2_X1 U16723 ( .A1(n13173), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13151) );
  AOI22_X1 U16724 ( .A1(n13627), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21647), .ZN(n13150) );
  AND2_X1 U16725 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  NAND2_X1 U16726 ( .A1(n13153), .A2(n13152), .ZN(n14185) );
  NAND2_X1 U16727 ( .A1(n21139), .A2(n10026), .ZN(n13155) );
  NAND2_X1 U16728 ( .A1(n13155), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13781) );
  INV_X1 U16729 ( .A(n13173), .ZN(n13169) );
  NAND2_X1 U16730 ( .A1(n21647), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13158) );
  NAND2_X1 U16731 ( .A1(n13183), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13157) );
  OAI211_X1 U16732 ( .C1(n13169), .C2(n17498), .A(n13158), .B(n13157), .ZN(
        n13159) );
  AOI21_X1 U16733 ( .B1(n13156), .B2(n13335), .A(n13159), .ZN(n13780) );
  OR2_X1 U16734 ( .A1(n13781), .A2(n13780), .ZN(n13783) );
  INV_X1 U16735 ( .A(n13780), .ZN(n13160) );
  OR2_X1 U16736 ( .A1(n13160), .A2(n14398), .ZN(n13161) );
  NAND2_X1 U16737 ( .A1(n13783), .A2(n13161), .ZN(n14184) );
  NAND2_X1 U16738 ( .A1(n14185), .A2(n14184), .ZN(n14183) );
  INV_X1 U16739 ( .A(n14183), .ZN(n14282) );
  NAND2_X1 U16740 ( .A1(n14283), .A2(n14282), .ZN(n14281) );
  INV_X1 U16741 ( .A(n15573), .ZN(n13163) );
  NAND2_X1 U16742 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13164) );
  INV_X1 U16743 ( .A(n13164), .ZN(n13166) );
  NOR2_X2 U16744 ( .A1(n13164), .A2(n14460), .ZN(n13176) );
  INV_X1 U16745 ( .A(n13176), .ZN(n13165) );
  OAI21_X1 U16746 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13166), .A(
        n13165), .ZN(n15298) );
  AOI22_X1 U16747 ( .A1(n13740), .A2(n15298), .B1(n13742), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13168) );
  NAND2_X1 U16748 ( .A1(n13627), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n13167) );
  OAI211_X1 U16749 ( .C1(n13169), .C2(n12471), .A(n13168), .B(n13167), .ZN(
        n13170) );
  INV_X1 U16750 ( .A(n13170), .ZN(n13171) );
  NAND2_X1 U16751 ( .A1(n13172), .A2(n13171), .ZN(n14449) );
  NAND2_X1 U16752 ( .A1(n13173), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13179) );
  INV_X1 U16753 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13174) );
  AOI21_X1 U16754 ( .B1(n13174), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13175) );
  AOI21_X1 U16755 ( .B1(n13627), .B2(P1_EAX_REG_4__SCAN_IN), .A(n13175), .ZN(
        n13178) );
  NAND2_X1 U16756 ( .A1(n13176), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13184) );
  OAI21_X1 U16757 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13176), .A(
        n13184), .ZN(n21005) );
  NOR2_X1 U16758 ( .A1(n21005), .A2(n14398), .ZN(n13177) );
  AOI21_X1 U16759 ( .B1(n13179), .B2(n13178), .A(n13177), .ZN(n13180) );
  AOI21_X1 U16760 ( .B1(n13181), .B2(n13335), .A(n13180), .ZN(n15060) );
  INV_X1 U16761 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n15058) );
  INV_X1 U16762 ( .A(n13184), .ZN(n13185) );
  OAI21_X1 U16763 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13185), .A(
        n13190), .ZN(n20934) );
  AOI22_X1 U16764 ( .A1(n13740), .A2(n20934), .B1(n13742), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13186) );
  OAI21_X1 U16765 ( .B1(n13149), .B2(n15058), .A(n13186), .ZN(n13187) );
  NAND2_X1 U16766 ( .A1(n13189), .A2(n13335), .ZN(n13196) );
  INV_X1 U16767 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13193) );
  OAI21_X1 U16768 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13191), .A(
        n13251), .ZN(n20915) );
  NAND2_X1 U16769 ( .A1(n20915), .A2(n13740), .ZN(n13192) );
  OAI21_X1 U16770 ( .B1(n13193), .B2(n13256), .A(n13192), .ZN(n13194) );
  AOI21_X1 U16771 ( .B1(n13627), .B2(P1_EAX_REG_6__SCAN_IN), .A(n13194), .ZN(
        n13195) );
  AOI22_X1 U16772 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13200) );
  AOI22_X1 U16773 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U16774 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U16775 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13197) );
  NAND4_X1 U16776 ( .A1(n13200), .A2(n13199), .A3(n13198), .A4(n13197), .ZN(
        n13210) );
  NAND2_X1 U16777 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13202) );
  NAND2_X1 U16778 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13201) );
  OAI211_X1 U16779 ( .C1(n13722), .C2(n13203), .A(n13202), .B(n13201), .ZN(
        n13204) );
  INV_X1 U16780 ( .A(n13204), .ZN(n13208) );
  AOI22_X1 U16781 ( .A1(n9753), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U16782 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9777), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U16783 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13205) );
  NAND4_X1 U16784 ( .A1(n13208), .A2(n13207), .A3(n13206), .A4(n13205), .ZN(
        n13209) );
  NOR2_X1 U16785 ( .A1(n13210), .A2(n13209), .ZN(n13214) );
  OAI21_X1 U16786 ( .B1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n13211), .A(
        n13260), .ZN(n20894) );
  AOI22_X1 U16787 ( .A1(n13740), .A2(n20894), .B1(n13742), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13213) );
  NAND2_X1 U16788 ( .A1(n13627), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13212) );
  OAI211_X1 U16789 ( .C1(n13362), .C2(n13214), .A(n13213), .B(n13212), .ZN(
        n14938) );
  AOI22_X1 U16790 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13218) );
  AOI22_X1 U16791 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13217) );
  AOI22_X1 U16792 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13216) );
  AOI22_X1 U16793 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13215) );
  NAND4_X1 U16794 ( .A1(n13218), .A2(n13217), .A3(n13216), .A4(n13215), .ZN(
        n13227) );
  INV_X1 U16795 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13370) );
  NAND2_X1 U16796 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13220) );
  NAND2_X1 U16797 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13219) );
  OAI211_X1 U16798 ( .C1(n13614), .C2(n13370), .A(n13220), .B(n13219), .ZN(
        n13221) );
  INV_X1 U16799 ( .A(n13221), .ZN(n13225) );
  AOI22_X1 U16800 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13224) );
  AOI22_X1 U16801 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13223) );
  NAND2_X1 U16802 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13222) );
  NAND4_X1 U16803 ( .A1(n13225), .A2(n13224), .A3(n13223), .A4(n13222), .ZN(
        n13226) );
  NOR2_X1 U16804 ( .A1(n13227), .A2(n13226), .ZN(n13230) );
  XNOR2_X1 U16805 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n13252), .ZN(
        n15288) );
  AOI22_X1 U16806 ( .A1(n13740), .A2(n15288), .B1(n13742), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13229) );
  NAND2_X1 U16807 ( .A1(n13627), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13228) );
  OAI211_X1 U16808 ( .C1(n13362), .C2(n13230), .A(n13229), .B(n13228), .ZN(
        n14864) );
  AOI22_X1 U16809 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U16810 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13234) );
  INV_X2 U16811 ( .A(n13231), .ZN(n15537) );
  AOI22_X1 U16812 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13233) );
  AOI22_X1 U16813 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13232) );
  NAND4_X1 U16814 ( .A1(n13235), .A2(n13234), .A3(n13233), .A4(n13232), .ZN(
        n13245) );
  NAND2_X1 U16815 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13237) );
  NAND2_X1 U16816 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13236) );
  OAI211_X1 U16817 ( .C1(n13722), .C2(n13238), .A(n13237), .B(n13236), .ZN(
        n13239) );
  INV_X1 U16818 ( .A(n13239), .ZN(n13243) );
  AOI22_X1 U16819 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16820 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13241) );
  NAND2_X1 U16821 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13240) );
  NAND4_X1 U16822 ( .A1(n13243), .A2(n13242), .A3(n13241), .A4(n13240), .ZN(
        n13244) );
  NOR2_X1 U16823 ( .A1(n13245), .A2(n13244), .ZN(n13248) );
  INV_X1 U16824 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14872) );
  XNOR2_X1 U16825 ( .A(n13260), .B(n14872), .ZN(n15274) );
  AOI22_X1 U16826 ( .A1(n15274), .A2(n13740), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13742), .ZN(n13247) );
  NAND2_X1 U16827 ( .A1(n13627), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n13246) );
  OAI211_X1 U16828 ( .C1(n13362), .C2(n13248), .A(n13247), .B(n13246), .ZN(
        n14865) );
  INV_X1 U16829 ( .A(n13249), .ZN(n13250) );
  NAND2_X1 U16830 ( .A1(n13250), .A2(n13335), .ZN(n13259) );
  INV_X1 U16831 ( .A(n13251), .ZN(n13254) );
  INV_X1 U16832 ( .A(n13252), .ZN(n13253) );
  OAI21_X1 U16833 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13254), .A(
        n13253), .ZN(n20906) );
  NAND2_X1 U16834 ( .A1(n20906), .A2(n13740), .ZN(n13255) );
  OAI21_X1 U16835 ( .B1(n20900), .B2(n13256), .A(n13255), .ZN(n13257) );
  AOI21_X1 U16836 ( .B1(n13627), .B2(P1_EAX_REG_7__SCAN_IN), .A(n13257), .ZN(
        n13258) );
  AND3_X2 U16837 ( .A1(n14861), .A2(n9851), .A3(n14863), .ZN(n14762) );
  NAND2_X1 U16838 ( .A1(n13627), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n13267) );
  INV_X1 U16839 ( .A(n13356), .ZN(n13339) );
  INV_X1 U16840 ( .A(n13262), .ZN(n13264) );
  INV_X1 U16841 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13263) );
  NAND2_X1 U16842 ( .A1(n13264), .A2(n13263), .ZN(n13265) );
  NAND2_X1 U16843 ( .A1(n13339), .A2(n13265), .ZN(n15261) );
  AOI22_X1 U16844 ( .A1(n15261), .A2(n13740), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13742), .ZN(n13266) );
  NAND2_X1 U16845 ( .A1(n13267), .A2(n13266), .ZN(n14811) );
  INV_X1 U16846 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13270) );
  NAND2_X1 U16847 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13269) );
  NAND2_X1 U16848 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n13268) );
  OAI211_X1 U16849 ( .C1(n12104), .C2(n13270), .A(n13269), .B(n13268), .ZN(
        n13271) );
  INV_X1 U16850 ( .A(n13271), .ZN(n13275) );
  AOI22_X1 U16851 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13274) );
  AOI22_X1 U16852 ( .A1(n13697), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13273) );
  NAND2_X1 U16853 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13272) );
  NAND4_X1 U16854 ( .A1(n13275), .A2(n13274), .A3(n13273), .A4(n13272), .ZN(
        n13281) );
  AOI22_X1 U16855 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12133), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13279) );
  AOI22_X1 U16856 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U16857 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U16858 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13725), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13276) );
  NAND4_X1 U16859 ( .A1(n13279), .A2(n13278), .A3(n13277), .A4(n13276), .ZN(
        n13280) );
  OR2_X1 U16860 ( .A1(n13281), .A2(n13280), .ZN(n13282) );
  AOI22_X1 U16861 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13286) );
  AOI22_X1 U16862 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13285) );
  AOI22_X1 U16863 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13284) );
  AOI22_X1 U16864 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9753), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13283) );
  NAND4_X1 U16865 ( .A1(n13286), .A2(n13285), .A3(n13284), .A4(n13283), .ZN(
        n13296) );
  INV_X1 U16866 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13289) );
  NAND2_X1 U16867 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n13288) );
  NAND2_X1 U16868 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13287) );
  OAI211_X1 U16869 ( .C1(n12104), .C2(n13289), .A(n13288), .B(n13287), .ZN(
        n13290) );
  INV_X1 U16870 ( .A(n13290), .ZN(n13294) );
  AOI22_X1 U16871 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U16872 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13292) );
  NAND2_X1 U16873 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13291) );
  NAND4_X1 U16874 ( .A1(n13294), .A2(n13293), .A3(n13292), .A4(n13291), .ZN(
        n13295) );
  OAI21_X1 U16875 ( .B1(n13296), .B2(n13295), .A(n13335), .ZN(n13302) );
  NAND2_X1 U16876 ( .A1(n13627), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13301) );
  NAND2_X1 U16877 ( .A1(n13742), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13300) );
  INV_X1 U16878 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13298) );
  XNOR2_X1 U16879 ( .A(n13316), .B(n13298), .ZN(n15232) );
  NAND2_X1 U16880 ( .A1(n15232), .A2(n13740), .ZN(n13299) );
  NAND4_X1 U16881 ( .A1(n13302), .A2(n13301), .A3(n13300), .A4(n13299), .ZN(
        n14797) );
  AOI22_X1 U16882 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13306) );
  AOI22_X1 U16883 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13525), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U16884 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U16885 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9776), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13303) );
  NAND4_X1 U16886 ( .A1(n13306), .A2(n13305), .A3(n13304), .A4(n13303), .ZN(
        n13315) );
  INV_X1 U16887 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13712) );
  NAND2_X1 U16888 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n13308) );
  NAND2_X1 U16889 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13307) );
  OAI211_X1 U16890 ( .C1(n13614), .C2(n13712), .A(n13308), .B(n13307), .ZN(
        n13309) );
  INV_X1 U16891 ( .A(n13309), .ZN(n13313) );
  AOI22_X1 U16892 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13312) );
  AOI22_X1 U16893 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13311) );
  NAND2_X1 U16894 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13310) );
  NAND4_X1 U16895 ( .A1(n13313), .A2(n13312), .A3(n13311), .A4(n13310), .ZN(
        n13314) );
  OAI21_X1 U16896 ( .B1(n13315), .B2(n13314), .A(n13335), .ZN(n13321) );
  NAND2_X1 U16897 ( .A1(n13627), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13320) );
  INV_X1 U16898 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14784) );
  XNOR2_X1 U16899 ( .A(n13380), .B(n14784), .ZN(n15219) );
  NAND2_X1 U16900 ( .A1(n15219), .A2(n13740), .ZN(n13319) );
  NAND2_X1 U16901 ( .A1(n13742), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13318) );
  NAND4_X1 U16902 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n13318), .ZN(
        n14783) );
  OAI211_X1 U16903 ( .C1(n14811), .C2(n14848), .A(n14797), .B(n14783), .ZN(
        n13363) );
  INV_X1 U16904 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20983) );
  AOI22_X1 U16905 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13647), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13326) );
  AOI22_X1 U16906 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13724), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U16907 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U16908 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13323) );
  NAND4_X1 U16909 ( .A1(n13326), .A2(n13325), .A3(n13324), .A4(n13323), .ZN(
        n13337) );
  INV_X1 U16910 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13329) );
  NAND2_X1 U16911 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13328) );
  NAND2_X1 U16912 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13327) );
  OAI211_X1 U16913 ( .C1(n12104), .C2(n13329), .A(n13328), .B(n13327), .ZN(
        n13330) );
  INV_X1 U16914 ( .A(n13330), .ZN(n13334) );
  AOI22_X1 U16915 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13333) );
  AOI22_X1 U16916 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13332) );
  NAND2_X1 U16917 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13331) );
  NAND4_X1 U16918 ( .A1(n13334), .A2(n13333), .A3(n13332), .A4(n13331), .ZN(
        n13336) );
  OAI21_X1 U16919 ( .B1(n13337), .B2(n13336), .A(n13335), .ZN(n13341) );
  INV_X1 U16920 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13338) );
  XNOR2_X1 U16921 ( .A(n13339), .B(n13338), .ZN(n15246) );
  AOI22_X1 U16922 ( .A1(n15246), .A2(n13740), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13742), .ZN(n13340) );
  OAI211_X1 U16923 ( .C1(n13149), .C2(n20983), .A(n13341), .B(n13340), .ZN(
        n14835) );
  AOI22_X1 U16924 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13345) );
  AOI22_X1 U16925 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13344) );
  AOI22_X1 U16926 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U16927 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9753), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13342) );
  NAND4_X1 U16928 ( .A1(n13345), .A2(n13344), .A3(n13343), .A4(n13342), .ZN(
        n13355) );
  NAND2_X1 U16929 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13347) );
  NAND2_X1 U16930 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13346) );
  OAI211_X1 U16931 ( .C1(n13722), .C2(n13348), .A(n13347), .B(n13346), .ZN(
        n13349) );
  INV_X1 U16932 ( .A(n13349), .ZN(n13353) );
  AOI22_X1 U16933 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13352) );
  AOI22_X1 U16934 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9777), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U16935 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13350) );
  NAND4_X1 U16936 ( .A1(n13353), .A2(n13352), .A3(n13351), .A4(n13350), .ZN(
        n13354) );
  NOR2_X1 U16937 ( .A1(n13355), .A2(n13354), .ZN(n13361) );
  NAND2_X1 U16938 ( .A1(n13356), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13358) );
  INV_X1 U16939 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13357) );
  XNOR2_X1 U16940 ( .A(n13358), .B(n13357), .ZN(n15239) );
  AOI22_X1 U16941 ( .A1(n15239), .A2(n13740), .B1(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n13742), .ZN(n13360) );
  NAND2_X1 U16942 ( .A1(n13627), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13359) );
  OAI211_X1 U16943 ( .C1(n13362), .C2(n13361), .A(n13360), .B(n13359), .ZN(
        n14815) );
  NAND2_X1 U16944 ( .A1(n14835), .A2(n14815), .ZN(n14780) );
  NOR2_X1 U16945 ( .A1(n13363), .A2(n14780), .ZN(n14764) );
  AOI22_X1 U16946 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U16947 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U16948 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9781), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U16949 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13364) );
  NAND4_X1 U16950 ( .A1(n13367), .A2(n13366), .A3(n13365), .A4(n13364), .ZN(
        n13377) );
  NAND2_X1 U16951 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13369) );
  NAND2_X1 U16952 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13368) );
  OAI211_X1 U16953 ( .C1(n13722), .C2(n13370), .A(n13369), .B(n13368), .ZN(
        n13371) );
  INV_X1 U16954 ( .A(n13371), .ZN(n13375) );
  AOI22_X1 U16955 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U16956 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13373) );
  NAND2_X1 U16957 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13372) );
  NAND4_X1 U16958 ( .A1(n13375), .A2(n13374), .A3(n13373), .A4(n13372), .ZN(
        n13376) );
  NOR2_X1 U16959 ( .A1(n13377), .A2(n13376), .ZN(n13379) );
  AOI22_X1 U16960 ( .A1(n13627), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21647), .ZN(n13378) );
  OAI21_X1 U16961 ( .B1(n13737), .B2(n13379), .A(n13378), .ZN(n13386) );
  INV_X1 U16962 ( .A(n13382), .ZN(n13384) );
  INV_X1 U16963 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n13383) );
  NAND2_X1 U16964 ( .A1(n13384), .A2(n13383), .ZN(n13385) );
  NAND2_X1 U16965 ( .A1(n13425), .A2(n13385), .ZN(n15208) );
  MUX2_X1 U16966 ( .A(n13386), .B(n15208), .S(n13740), .Z(n14765) );
  AND2_X1 U16967 ( .A1(n14764), .A2(n14765), .ZN(n13387) );
  AOI22_X1 U16968 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13391) );
  AOI22_X1 U16969 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13390) );
  AOI22_X1 U16970 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9781), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13389) );
  AOI22_X1 U16971 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13388) );
  NAND4_X1 U16972 ( .A1(n13391), .A2(n13390), .A3(n13389), .A4(n13388), .ZN(
        n13401) );
  INV_X1 U16973 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13394) );
  NAND2_X1 U16974 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13393) );
  NAND2_X1 U16975 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13392) );
  OAI211_X1 U16976 ( .C1(n13722), .C2(n13394), .A(n13393), .B(n13392), .ZN(
        n13395) );
  INV_X1 U16977 ( .A(n13395), .ZN(n13399) );
  AOI22_X1 U16978 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U16979 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13397) );
  NAND2_X1 U16980 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13396) );
  NAND4_X1 U16981 ( .A1(n13399), .A2(n13398), .A3(n13397), .A4(n13396), .ZN(
        n13400) );
  NOR2_X1 U16982 ( .A1(n13401), .A2(n13400), .ZN(n13405) );
  AOI22_X1 U16983 ( .A1(n13627), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n13742), .ZN(n13404) );
  INV_X1 U16984 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13402) );
  XNOR2_X1 U16985 ( .A(n13425), .B(n13402), .ZN(n15198) );
  NAND2_X1 U16986 ( .A1(n15198), .A2(n13740), .ZN(n13403) );
  OAI211_X1 U16987 ( .C1(n13737), .C2(n13405), .A(n13404), .B(n13403), .ZN(
        n13406) );
  INV_X1 U16988 ( .A(n13406), .ZN(n14745) );
  AOI22_X1 U16989 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13410) );
  AOI22_X1 U16990 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9838), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13409) );
  AOI22_X1 U16991 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13408) );
  AOI22_X1 U16992 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13407) );
  NAND4_X1 U16993 ( .A1(n13410), .A2(n13409), .A3(n13408), .A4(n13407), .ZN(
        n13420) );
  INV_X1 U16994 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13413) );
  NAND2_X1 U16995 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13412) );
  NAND2_X1 U16996 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13411) );
  OAI211_X1 U16997 ( .C1(n13614), .C2(n13413), .A(n13412), .B(n13411), .ZN(
        n13414) );
  INV_X1 U16998 ( .A(n13414), .ZN(n13418) );
  AOI22_X1 U16999 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U17000 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13416) );
  NAND2_X1 U17001 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13415) );
  NAND4_X1 U17002 ( .A1(n13418), .A2(n13417), .A3(n13416), .A4(n13415), .ZN(
        n13419) );
  NOR2_X1 U17003 ( .A1(n13420), .A2(n13419), .ZN(n13424) );
  OAI21_X1 U17004 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21880), .A(
        n21647), .ZN(n13421) );
  INV_X1 U17005 ( .A(n13421), .ZN(n13422) );
  AOI21_X1 U17006 ( .B1(n13627), .B2(P1_EAX_REG_18__SCAN_IN), .A(n13422), .ZN(
        n13423) );
  OAI21_X1 U17007 ( .B1(n13737), .B2(n13424), .A(n13423), .ZN(n13432) );
  INV_X1 U17008 ( .A(n13427), .ZN(n13429) );
  INV_X1 U17009 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13428) );
  NAND2_X1 U17010 ( .A1(n13429), .A2(n13428), .ZN(n13430) );
  NAND2_X1 U17011 ( .A1(n13453), .A2(n13430), .ZN(n15181) );
  OR2_X1 U17012 ( .A1(n15181), .A2(n14398), .ZN(n13431) );
  XNOR2_X1 U17013 ( .A(n13453), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15177) );
  NAND2_X1 U17014 ( .A1(n15177), .A2(n13740), .ZN(n13452) );
  AOI22_X1 U17015 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13437) );
  AOI22_X1 U17016 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13436) );
  AOI22_X1 U17017 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U17018 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13434) );
  NAND4_X1 U17019 ( .A1(n13437), .A2(n13436), .A3(n13435), .A4(n13434), .ZN(
        n13447) );
  INV_X1 U17020 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13440) );
  NAND2_X1 U17021 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13439) );
  NAND2_X1 U17022 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13438) );
  OAI211_X1 U17023 ( .C1(n13614), .C2(n13440), .A(n13439), .B(n13438), .ZN(
        n13441) );
  INV_X1 U17024 ( .A(n13441), .ZN(n13445) );
  AOI22_X1 U17025 ( .A1(n9753), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9754), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13444) );
  AOI22_X1 U17026 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13443) );
  NAND2_X1 U17027 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13442) );
  NAND4_X1 U17028 ( .A1(n13445), .A2(n13444), .A3(n13443), .A4(n13442), .ZN(
        n13446) );
  NOR2_X1 U17029 ( .A1(n13447), .A2(n13446), .ZN(n13450) );
  AOI21_X1 U17030 ( .B1(n15172), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13448) );
  AOI21_X1 U17031 ( .B1(n13627), .B2(P1_EAX_REG_19__SCAN_IN), .A(n13448), .ZN(
        n13449) );
  OAI21_X1 U17032 ( .B1(n13737), .B2(n13450), .A(n13449), .ZN(n13451) );
  INV_X1 U17033 ( .A(n14706), .ZN(n13473) );
  OR2_X2 U17034 ( .A1(n13454), .A2(n14708), .ZN(n13510) );
  NAND2_X1 U17035 ( .A1(n13454), .A2(n14708), .ZN(n13455) );
  NAND2_X1 U17036 ( .A1(n13510), .A2(n13455), .ZN(n15166) );
  INV_X1 U17037 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13644) );
  NAND2_X1 U17038 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13457) );
  NAND2_X1 U17039 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13456) );
  OAI211_X1 U17040 ( .C1(n13614), .C2(n13644), .A(n13457), .B(n13456), .ZN(
        n13458) );
  INV_X1 U17041 ( .A(n13458), .ZN(n13462) );
  AOI22_X1 U17042 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13461) );
  AOI22_X1 U17043 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13522), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13460) );
  NAND2_X1 U17044 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13459) );
  NAND4_X1 U17045 ( .A1(n13462), .A2(n13461), .A3(n13460), .A4(n13459), .ZN(
        n13468) );
  AOI22_X1 U17046 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13466) );
  AOI22_X1 U17047 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9746), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U17048 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13725), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13464) );
  AOI22_X1 U17049 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13463) );
  NAND4_X1 U17050 ( .A1(n13466), .A2(n13465), .A3(n13464), .A4(n13463), .ZN(
        n13467) );
  NOR2_X1 U17051 ( .A1(n13468), .A2(n13467), .ZN(n13470) );
  AOI22_X1 U17052 ( .A1(n13627), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21647), .ZN(n13469) );
  OAI21_X1 U17053 ( .B1(n13737), .B2(n13470), .A(n13469), .ZN(n13471) );
  MUX2_X1 U17054 ( .A(n15166), .B(n13471), .S(n14398), .Z(n13472) );
  NAND2_X1 U17055 ( .A1(n13473), .A2(n13472), .ZN(n14688) );
  INV_X2 U17056 ( .A(n14688), .ZN(n13493) );
  XNOR2_X1 U17057 ( .A(n13510), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14694) );
  NAND2_X1 U17058 ( .A1(n14694), .A2(n13740), .ZN(n13491) );
  INV_X1 U17059 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n21940) );
  AOI22_X1 U17060 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13477) );
  AOI22_X1 U17061 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13476) );
  AOI22_X1 U17062 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12132), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13475) );
  AOI22_X1 U17063 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13474) );
  NAND4_X1 U17064 ( .A1(n13477), .A2(n13476), .A3(n13475), .A4(n13474), .ZN(
        n13486) );
  NAND2_X1 U17065 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13479) );
  NAND2_X1 U17066 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13478) );
  OAI211_X1 U17067 ( .C1(n13614), .C2(n9996), .A(n13479), .B(n13478), .ZN(
        n13480) );
  INV_X1 U17068 ( .A(n13480), .ZN(n13484) );
  AOI22_X1 U17069 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U17070 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13482) );
  NAND2_X1 U17071 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13481) );
  NAND4_X1 U17072 ( .A1(n13484), .A2(n13483), .A3(n13482), .A4(n13481), .ZN(
        n13485) );
  NOR2_X1 U17073 ( .A1(n13486), .A2(n13485), .ZN(n13489) );
  AOI21_X1 U17074 ( .B1(n14695), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13487) );
  AOI21_X1 U17075 ( .B1(n13627), .B2(P1_EAX_REG_21__SCAN_IN), .A(n13487), .ZN(
        n13488) );
  OAI21_X1 U17076 ( .B1(n13737), .B2(n13489), .A(n13488), .ZN(n13490) );
  NAND2_X1 U17077 ( .A1(n13491), .A2(n13490), .ZN(n14691) );
  AOI22_X1 U17078 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U17079 ( .A1(n9773), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13496) );
  AOI22_X1 U17080 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13495) );
  AOI22_X1 U17081 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13494) );
  NAND4_X1 U17082 ( .A1(n13497), .A2(n13496), .A3(n13495), .A4(n13494), .ZN(
        n13506) );
  INV_X1 U17083 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13696) );
  NAND2_X1 U17084 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13499) );
  NAND2_X1 U17085 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13498) );
  OAI211_X1 U17086 ( .C1(n13614), .C2(n13696), .A(n13499), .B(n13498), .ZN(
        n13500) );
  INV_X1 U17087 ( .A(n13500), .ZN(n13504) );
  AOI22_X1 U17088 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13503) );
  AOI22_X1 U17089 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9777), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13502) );
  NAND2_X1 U17090 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n13501) );
  NAND4_X1 U17091 ( .A1(n13504), .A2(n13503), .A3(n13502), .A4(n13501), .ZN(
        n13505) );
  NOR2_X1 U17092 ( .A1(n13506), .A2(n13505), .ZN(n13508) );
  AOI22_X1 U17093 ( .A1(n13627), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21647), .ZN(n13507) );
  OAI21_X1 U17094 ( .B1(n13737), .B2(n13508), .A(n13507), .ZN(n13509) );
  INV_X1 U17095 ( .A(n13509), .ZN(n13515) );
  INV_X1 U17096 ( .A(n13511), .ZN(n13513) );
  INV_X1 U17097 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13512) );
  NAND2_X1 U17098 ( .A1(n13513), .A2(n13512), .ZN(n13514) );
  AND2_X1 U17099 ( .A1(n13553), .A2(n13514), .ZN(n15145) );
  MUX2_X1 U17100 ( .A(n13515), .B(n15145), .S(n13740), .Z(n14673) );
  INV_X1 U17101 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13721) );
  INV_X1 U17102 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13517) );
  INV_X1 U17103 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13516) );
  OAI22_X1 U17104 ( .A1(n12097), .A2(n13517), .B1(n13711), .B2(n13516), .ZN(
        n13521) );
  INV_X1 U17105 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13519) );
  OAI22_X1 U17106 ( .A1(n13687), .A2(n13519), .B1(n12222), .B2(n13518), .ZN(
        n13520) );
  AOI211_X1 U17107 ( .C1(n13666), .C2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n13521), .B(n13520), .ZN(n13524) );
  AOI22_X1 U17108 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13523) );
  OAI211_X1 U17109 ( .C1(n12104), .C2(n13721), .A(n13524), .B(n13523), .ZN(
        n13531) );
  AOI22_X1 U17110 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13529) );
  AOI22_X1 U17111 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12132), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13528) );
  AOI22_X1 U17112 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U17113 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13526) );
  NAND4_X1 U17114 ( .A1(n13529), .A2(n13528), .A3(n13527), .A4(n13526), .ZN(
        n13530) );
  NOR2_X1 U17115 ( .A1(n13531), .A2(n13530), .ZN(n13558) );
  INV_X1 U17116 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13540) );
  INV_X1 U17117 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13533) );
  OAI22_X1 U17118 ( .A1(n13636), .A2(n13533), .B1(n12222), .B2(n13532), .ZN(
        n13537) );
  INV_X1 U17119 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13535) );
  INV_X1 U17120 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13534) );
  OAI22_X1 U17121 ( .A1(n13690), .A2(n13535), .B1(n13231), .B2(n13534), .ZN(
        n13536) );
  AOI211_X1 U17122 ( .C1(n13717), .C2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n13537), .B(n13536), .ZN(n13539) );
  AOI22_X1 U17123 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13538) );
  OAI211_X1 U17124 ( .C1(n13722), .C2(n13540), .A(n13539), .B(n13538), .ZN(
        n13547) );
  AOI22_X1 U17125 ( .A1(n13541), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13545) );
  AOI22_X1 U17126 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13544) );
  AOI22_X1 U17127 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13543) );
  AOI22_X1 U17128 ( .A1(n9753), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13542) );
  NAND4_X1 U17129 ( .A1(n13545), .A2(n13544), .A3(n13543), .A4(n13542), .ZN(
        n13546) );
  NOR2_X1 U17130 ( .A1(n13547), .A2(n13546), .ZN(n13559) );
  XOR2_X1 U17131 ( .A(n13558), .B(n13559), .Z(n13548) );
  NAND2_X1 U17132 ( .A1(n13548), .A2(n13706), .ZN(n13550) );
  AOI22_X1 U17133 ( .A1(n13627), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n21647), .ZN(n13549) );
  NAND2_X1 U17134 ( .A1(n13550), .A2(n13549), .ZN(n13552) );
  INV_X1 U17135 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13551) );
  XNOR2_X1 U17136 ( .A(n13553), .B(n13551), .ZN(n15138) );
  MUX2_X1 U17137 ( .A(n13552), .B(n15138), .S(n13740), .Z(n14660) );
  AND2_X2 U17138 ( .A1(n13554), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13555) );
  INV_X1 U17139 ( .A(n13555), .ZN(n13556) );
  INV_X1 U17140 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13575) );
  NAND2_X1 U17141 ( .A1(n13556), .A2(n13575), .ZN(n13557) );
  NAND2_X1 U17142 ( .A1(n13603), .A2(n13557), .ZN(n15131) );
  NOR2_X1 U17143 ( .A1(n13559), .A2(n13558), .ZN(n13582) );
  INV_X1 U17144 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13562) );
  NAND2_X1 U17145 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13561) );
  NAND2_X1 U17146 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13560) );
  OAI211_X1 U17147 ( .C1(n13614), .C2(n13562), .A(n13561), .B(n13560), .ZN(
        n13563) );
  INV_X1 U17148 ( .A(n13563), .ZN(n13568) );
  AOI22_X1 U17149 ( .A1(n9753), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U17150 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9777), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13566) );
  NAND2_X1 U17151 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13565) );
  NAND4_X1 U17152 ( .A1(n13568), .A2(n13567), .A3(n13566), .A4(n13565), .ZN(
        n13574) );
  AOI22_X1 U17153 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13572) );
  AOI22_X1 U17154 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13571) );
  AOI22_X1 U17155 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13570) );
  AOI22_X1 U17156 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13569) );
  NAND4_X1 U17157 ( .A1(n13572), .A2(n13571), .A3(n13570), .A4(n13569), .ZN(
        n13573) );
  OR2_X1 U17158 ( .A1(n13574), .A2(n13573), .ZN(n13581) );
  XNOR2_X1 U17159 ( .A(n13582), .B(n13581), .ZN(n13578) );
  AOI21_X1 U17160 ( .B1(n13575), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13576) );
  AOI21_X1 U17161 ( .B1(n13627), .B2(P1_EAX_REG_24__SCAN_IN), .A(n13576), .ZN(
        n13577) );
  OAI21_X1 U17162 ( .B1(n13578), .B2(n13737), .A(n13577), .ZN(n13579) );
  NAND2_X1 U17163 ( .A1(n13582), .A2(n13581), .ZN(n13608) );
  INV_X1 U17164 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13591) );
  INV_X1 U17165 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13584) );
  INV_X1 U17166 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13583) );
  OAI22_X1 U17167 ( .A1(n13231), .A2(n13584), .B1(n13711), .B2(n13583), .ZN(
        n13588) );
  INV_X1 U17168 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13586) );
  INV_X1 U17169 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13585) );
  OAI22_X1 U17170 ( .A1(n13690), .A2(n13586), .B1(n9772), .B2(n13585), .ZN(
        n13587) );
  AOI211_X1 U17171 ( .C1(n13666), .C2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n13588), .B(n13587), .ZN(n13590) );
  AOI22_X1 U17172 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13589) );
  OAI211_X1 U17173 ( .C1(n12104), .C2(n13591), .A(n13590), .B(n13589), .ZN(
        n13597) );
  AOI22_X1 U17174 ( .A1(n12132), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13595) );
  AOI22_X1 U17175 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U17176 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13725), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13593) );
  AOI22_X1 U17177 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9776), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13592) );
  NAND4_X1 U17178 ( .A1(n13595), .A2(n13594), .A3(n13593), .A4(n13592), .ZN(
        n13596) );
  NOR2_X1 U17179 ( .A1(n13597), .A2(n13596), .ZN(n13609) );
  XOR2_X1 U17180 ( .A(n13608), .B(n13609), .Z(n13598) );
  NAND2_X1 U17181 ( .A1(n13598), .A2(n13706), .ZN(n13600) );
  AOI22_X1 U17182 ( .A1(n13183), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n21647), .ZN(n13599) );
  NAND2_X1 U17183 ( .A1(n13600), .A2(n13599), .ZN(n13602) );
  INV_X1 U17184 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13601) );
  XNOR2_X1 U17185 ( .A(n13603), .B(n13601), .ZN(n15121) );
  MUX2_X1 U17186 ( .A(n13602), .B(n15121), .S(n13740), .Z(n14630) );
  AND2_X2 U17187 ( .A1(n13604), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13605) );
  INV_X1 U17188 ( .A(n13605), .ZN(n13606) );
  INV_X1 U17189 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14621) );
  NAND2_X1 U17190 ( .A1(n13606), .A2(n14621), .ZN(n13607) );
  NAND2_X1 U17191 ( .A1(n13658), .A2(n13607), .ZN(n15110) );
  NOR2_X1 U17192 ( .A1(n13609), .A2(n13608), .ZN(n13633) );
  INV_X1 U17193 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U17194 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13612) );
  NAND2_X1 U17195 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n13611) );
  OAI211_X1 U17196 ( .C1(n13614), .C2(n13613), .A(n13612), .B(n13611), .ZN(
        n13615) );
  INV_X1 U17197 ( .A(n13615), .ZN(n13619) );
  AOI22_X1 U17198 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U17199 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13564), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U17200 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13616) );
  NAND4_X1 U17201 ( .A1(n13619), .A2(n13618), .A3(n13617), .A4(n13616), .ZN(
        n13625) );
  AOI22_X1 U17202 ( .A1(n9782), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13623) );
  AOI22_X1 U17203 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13622) );
  AOI22_X1 U17204 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13621) );
  AOI22_X1 U17205 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13620) );
  NAND4_X1 U17206 ( .A1(n13623), .A2(n13622), .A3(n13621), .A4(n13620), .ZN(
        n13624) );
  OR2_X1 U17207 ( .A1(n13625), .A2(n13624), .ZN(n13632) );
  XNOR2_X1 U17208 ( .A(n13633), .B(n13632), .ZN(n13629) );
  AOI21_X1 U17209 ( .B1(n14621), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13626) );
  AOI21_X1 U17210 ( .B1(n13627), .B2(P1_EAX_REG_26__SCAN_IN), .A(n13626), .ZN(
        n13628) );
  OAI21_X1 U17211 ( .B1(n13629), .B2(n13737), .A(n13628), .ZN(n13630) );
  NAND2_X1 U17212 ( .A1(n13633), .A2(n13632), .ZN(n13660) );
  INV_X1 U17213 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13635) );
  OAI22_X1 U17214 ( .A1(n13636), .A2(n13635), .B1(n12222), .B2(n13634), .ZN(
        n13641) );
  INV_X1 U17215 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13638) );
  INV_X1 U17216 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13637) );
  OAI22_X1 U17217 ( .A1(n13639), .A2(n13638), .B1(n13231), .B2(n13637), .ZN(
        n13640) );
  AOI211_X1 U17218 ( .C1(n13717), .C2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n13641), .B(n13640), .ZN(n13643) );
  AOI22_X1 U17219 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n13693), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13642) );
  OAI211_X1 U17220 ( .C1(n13722), .C2(n13644), .A(n13643), .B(n13642), .ZN(
        n13653) );
  AOI22_X1 U17221 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13651) );
  AOI22_X1 U17222 ( .A1(n13525), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13650) );
  AOI22_X1 U17223 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13649) );
  AOI22_X1 U17224 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13725), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13648) );
  NAND4_X1 U17225 ( .A1(n13651), .A2(n13650), .A3(n13649), .A4(n13648), .ZN(
        n13652) );
  NOR2_X1 U17226 ( .A1(n13653), .A2(n13652), .ZN(n13661) );
  XOR2_X1 U17227 ( .A(n13660), .B(n13661), .Z(n13655) );
  INV_X1 U17228 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14979) );
  INV_X1 U17229 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14609) );
  OAI22_X1 U17230 ( .A1(n13149), .A2(n14979), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14609), .ZN(n13654) );
  AOI21_X1 U17231 ( .B1(n13655), .B2(n13706), .A(n13654), .ZN(n13656) );
  XNOR2_X1 U17232 ( .A(n13658), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14608) );
  MUX2_X1 U17233 ( .A(n13656), .B(n14608), .S(n13740), .Z(n14605) );
  INV_X1 U17234 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14597) );
  OAI21_X1 U17235 ( .B1(n13658), .B2(n14609), .A(n14597), .ZN(n13659) );
  NAND2_X1 U17236 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13657) );
  OR2_X2 U17237 ( .A1(n13658), .A2(n13657), .ZN(n13681) );
  NAND2_X1 U17238 ( .A1(n13659), .A2(n13681), .ZN(n15091) );
  NOR2_X1 U17239 ( .A1(n13661), .A2(n13660), .ZN(n13684) );
  NAND2_X1 U17240 ( .A1(n13662), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13664) );
  NAND2_X1 U17241 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n13663) );
  OAI211_X1 U17242 ( .C1(n12104), .C2(n9998), .A(n13664), .B(n13663), .ZN(
        n13665) );
  INV_X1 U17243 ( .A(n13665), .ZN(n13670) );
  AOI22_X1 U17244 ( .A1(n9753), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13669) );
  AOI22_X1 U17245 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9777), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13668) );
  NAND2_X1 U17246 ( .A1(n13666), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13667) );
  NAND4_X1 U17247 ( .A1(n13670), .A2(n13669), .A3(n13668), .A4(n13667), .ZN(
        n13676) );
  AOI22_X1 U17248 ( .A1(n9781), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U17249 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13723), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U17250 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13672) );
  AOI22_X1 U17251 ( .A1(n13724), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13671) );
  NAND4_X1 U17252 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13675) );
  OR2_X1 U17253 ( .A1(n13676), .A2(n13675), .ZN(n13683) );
  XNOR2_X1 U17254 ( .A(n13684), .B(n13683), .ZN(n13678) );
  AOI22_X1 U17255 ( .A1(n13183), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n21647), .ZN(n13677) );
  OAI21_X1 U17256 ( .B1(n13678), .B2(n13737), .A(n13677), .ZN(n13679) );
  MUX2_X1 U17257 ( .A(n15091), .B(n13679), .S(n14398), .Z(n14595) );
  INV_X1 U17258 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21867) );
  NAND2_X1 U17259 ( .A1(n13681), .A2(n21867), .ZN(n13682) );
  NAND2_X1 U17260 ( .A1(n13684), .A2(n13683), .ZN(n13732) );
  INV_X1 U17261 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13686) );
  OAI22_X1 U17262 ( .A1(n13687), .A2(n13686), .B1(n12222), .B2(n13685), .ZN(
        n13692) );
  INV_X1 U17263 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13689) );
  INV_X1 U17264 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13688) );
  OAI22_X1 U17265 ( .A1(n13690), .A2(n13689), .B1(n13231), .B2(n13688), .ZN(
        n13691) );
  AOI211_X1 U17266 ( .C1(n13717), .C2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n13692), .B(n13691), .ZN(n13695) );
  AOI22_X1 U17267 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13694) );
  OAI211_X1 U17268 ( .C1(n13722), .C2(n13696), .A(n13695), .B(n13694), .ZN(
        n13703) );
  AOI22_X1 U17269 ( .A1(n13522), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U17270 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13525), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U17271 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U17272 ( .A1(n13725), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13697), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13698) );
  NAND4_X1 U17273 ( .A1(n13701), .A2(n13700), .A3(n13699), .A4(n13698), .ZN(
        n13702) );
  NOR2_X1 U17274 ( .A1(n13703), .A2(n13702), .ZN(n13733) );
  XOR2_X1 U17275 ( .A(n13732), .B(n13733), .Z(n13707) );
  INV_X1 U17276 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14968) );
  OAI21_X1 U17277 ( .B1(n21880), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n21647), .ZN(n13704) );
  OAI21_X1 U17278 ( .B1(n13149), .B2(n14968), .A(n13704), .ZN(n13705) );
  AOI21_X1 U17279 ( .B1(n13707), .B2(n13706), .A(n13705), .ZN(n13708) );
  AOI21_X1 U17280 ( .B1(n14583), .B2(n13740), .A(n13708), .ZN(n14582) );
  INV_X1 U17281 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13710) );
  OAI22_X1 U17282 ( .A1(n13711), .A2(n13710), .B1(n12222), .B2(n13709), .ZN(
        n13716) );
  INV_X1 U17283 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13714) );
  OAI22_X1 U17284 ( .A1(n13231), .A2(n13714), .B1(n13713), .B2(n13712), .ZN(
        n13715) );
  AOI211_X1 U17285 ( .C1(n13717), .C2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n13716), .B(n13715), .ZN(n13720) );
  AOI22_X1 U17286 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13719) );
  OAI211_X1 U17287 ( .C1(n13722), .C2(n13721), .A(n13720), .B(n13719), .ZN(
        n13731) );
  AOI22_X1 U17288 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13522), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13729) );
  AOI22_X1 U17289 ( .A1(n13723), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13645), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13728) );
  AOI22_X1 U17290 ( .A1(n9838), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13724), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13727) );
  AOI22_X1 U17291 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9753), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13726) );
  NAND4_X1 U17292 ( .A1(n13729), .A2(n13728), .A3(n13727), .A4(n13726), .ZN(
        n13730) );
  NOR2_X1 U17293 ( .A1(n13731), .A2(n13730), .ZN(n13735) );
  NOR2_X1 U17294 ( .A1(n13733), .A2(n13732), .ZN(n13734) );
  XOR2_X1 U17295 ( .A(n13735), .B(n13734), .Z(n13738) );
  AOI22_X1 U17296 ( .A1(n13183), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21647), .ZN(n13736) );
  OAI21_X1 U17297 ( .B1(n13738), .B2(n13737), .A(n13736), .ZN(n13739) );
  INV_X1 U17298 ( .A(n13739), .ZN(n13741) );
  XNOR2_X1 U17299 ( .A(n14402), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15068) );
  MUX2_X1 U17300 ( .A(n13741), .B(n15068), .S(n13740), .Z(n14568) );
  AOI22_X1 U17301 ( .A1(n13183), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13742), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13743) );
  XNOR2_X1 U17302 ( .A(n14567), .B(n13743), .ZN(n14507) );
  OAI21_X1 U17303 ( .B1(n14055), .B2(n12543), .A(n15523), .ZN(n14476) );
  NAND2_X1 U17304 ( .A1(n15557), .A2(n14476), .ZN(n13747) );
  INV_X1 U17305 ( .A(n21106), .ZN(n14017) );
  NAND4_X1 U17306 ( .A1(n15522), .A2(n10378), .A3(n14017), .A4(n12182), .ZN(
        n14015) );
  NAND2_X1 U17307 ( .A1(n17593), .A2(n13744), .ZN(n14480) );
  OAI21_X1 U17308 ( .B1(n12199), .B2(n14015), .A(n14480), .ZN(n13745) );
  INV_X1 U17309 ( .A(n13745), .ZN(n13746) );
  NAND3_X1 U17310 ( .A1(n14507), .A2(n15066), .A3(n14017), .ZN(n13764) );
  NOR4_X1 U17311 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13753) );
  NOR4_X1 U17312 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13752) );
  NOR4_X1 U17313 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13751) );
  NOR4_X1 U17314 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13750) );
  AND4_X1 U17315 ( .A1(n13753), .A2(n13752), .A3(n13751), .A4(n13750), .ZN(
        n13758) );
  NOR4_X1 U17316 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n13756) );
  NOR4_X1 U17317 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .A3(P1_ADDRESS_REG_23__SCAN_IN), .A4(
        P1_ADDRESS_REG_22__SCAN_IN), .ZN(n13755) );
  NOR4_X1 U17318 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_28__SCAN_IN), .A3(P1_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_ADDRESS_REG_26__SCAN_IN), .ZN(n13754) );
  AND4_X1 U17319 ( .A1(n13756), .A2(n13755), .A3(n13754), .A4(n21666), .ZN(
        n13757) );
  NAND2_X1 U17320 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  INV_X1 U17321 ( .A(n15033), .ZN(n15039) );
  AOI22_X1 U17322 ( .A1(n15039), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15034), .ZN(n13762) );
  INV_X1 U17323 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n21103) );
  NAND2_X1 U17324 ( .A1(n15029), .A2(BUF1_REG_31__SCAN_IN), .ZN(n13761) );
  AND2_X1 U17325 ( .A1(n13762), .A2(n13761), .ZN(n13763) );
  NAND2_X1 U17326 ( .A1(n13764), .A2(n13763), .ZN(P1_U2873) );
  NOR2_X1 U17327 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13766) );
  NOR4_X1 U17328 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13765) );
  NAND4_X1 U17329 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13766), .A4(n13765), .ZN(n13779) );
  INV_X2 U17330 ( .A(n17721), .ZN(U215) );
  NOR3_X1 U17331 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21968), .ZN(n13768) );
  NOR4_X1 U17332 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13767) );
  NOR4_X1 U17333 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13772) );
  NOR4_X1 U17334 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_2__SCAN_IN), .A4(
        P2_ADDRESS_REG_1__SCAN_IN), .ZN(n13771) );
  NOR4_X1 U17335 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n13770) );
  NOR4_X1 U17336 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_20__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n13769) );
  AND4_X1 U17337 ( .A1(n13772), .A2(n13771), .A3(n13770), .A4(n13769), .ZN(
        n13777) );
  NOR4_X1 U17338 ( .A1(P2_ADDRESS_REG_9__SCAN_IN), .A2(
        P2_ADDRESS_REG_4__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13775) );
  NOR4_X1 U17339 ( .A1(P2_ADDRESS_REG_12__SCAN_IN), .A2(
        P2_ADDRESS_REG_11__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13774) );
  NOR4_X1 U17340 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n13773) );
  AND4_X1 U17341 ( .A1(n13775), .A2(n13774), .A3(n13773), .A4(n20775), .ZN(
        n13776) );
  NAND2_X1 U17342 ( .A1(n13777), .A2(n13776), .ZN(n13778) );
  NAND2_X1 U17343 ( .A1(n13781), .A2(n13780), .ZN(n13782) );
  NAND2_X1 U17344 ( .A1(n13783), .A2(n13782), .ZN(n14903) );
  AND2_X1 U17345 ( .A1(n21517), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15576) );
  NAND2_X1 U17346 ( .A1(n21645), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n17527) );
  INV_X1 U17347 ( .A(n17527), .ZN(n13784) );
  NOR2_X1 U17348 ( .A1(n14903), .A2(n15252), .ZN(n13797) );
  OR2_X1 U17349 ( .A1(n21139), .A2(n13785), .ZN(n13788) );
  NOR2_X1 U17350 ( .A1(n13786), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13787) );
  NAND2_X1 U17351 ( .A1(n13788), .A2(n13787), .ZN(n13789) );
  NAND2_X1 U17352 ( .A1(n13789), .A2(n14291), .ZN(n14040) );
  NOR2_X1 U17353 ( .A1(n14040), .A2(n20873), .ZN(n13796) );
  INV_X1 U17354 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13790) );
  NOR2_X1 U17355 ( .A1(n17570), .A2(n13790), .ZN(n14037) );
  NAND2_X1 U17356 ( .A1(n21579), .A2(n13791), .ZN(n21736) );
  NAND2_X1 U17357 ( .A1(n21736), .A2(n21645), .ZN(n13792) );
  NAND2_X1 U17358 ( .A1(n21645), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17525) );
  NAND2_X1 U17359 ( .A1(n21880), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13793) );
  AND2_X1 U17360 ( .A1(n17525), .A2(n13793), .ZN(n14290) );
  INV_X1 U17361 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13794) );
  AOI21_X1 U17362 ( .B1(n15173), .B2(n14290), .A(n13794), .ZN(n13795) );
  OR4_X1 U17363 ( .A1(n13797), .A2(n13796), .A3(n14037), .A4(n13795), .ZN(
        P1_U2999) );
  AOI22_X1 U17364 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n13799) );
  INV_X1 U17365 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21662) );
  INV_X1 U17366 ( .A(HOLD), .ZN(n20723) );
  NOR2_X1 U17367 ( .A1(n21662), .A2(n20723), .ZN(n13798) );
  INV_X1 U17368 ( .A(n13862), .ZN(n17521) );
  NAND2_X1 U17369 ( .A1(n21739), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21657) );
  OAI211_X1 U17370 ( .C1(n13799), .C2(n13798), .A(n17521), .B(n21657), .ZN(
        P1_U3195) );
  MUX2_X1 U17371 ( .A(P2_STATEBS16_REG_SCAN_IN), .B(n20850), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n13800) );
  AOI21_X1 U17372 ( .B1(n13800), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n13801) );
  NAND2_X1 U17373 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17270), .ZN(n17376) );
  INV_X1 U17374 ( .A(n17376), .ZN(n17610) );
  NOR2_X1 U17375 ( .A1(n13801), .A2(n17610), .ZN(P2_U3178) );
  INV_X1 U17376 ( .A(n16010), .ZN(n13805) );
  INV_X1 U17377 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13804) );
  AND2_X1 U17378 ( .A1(n20800), .A2(n17365), .ZN(n20009) );
  INV_X1 U17379 ( .A(n20009), .ZN(n13802) );
  OAI211_X1 U17380 ( .C1(n13805), .C2(n13804), .A(n13803), .B(n13802), .ZN(
        P2_U2814) );
  OAI21_X1 U17381 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n20009), .A(n20847), 
        .ZN(n13806) );
  OAI21_X1 U17382 ( .B1(n13807), .B2(n20847), .A(n13806), .ZN(P2_U3612) );
  NOR3_X1 U17383 ( .A1(n13962), .A2(n13809), .A3(n17348), .ZN(n13810) );
  NAND2_X1 U17384 ( .A1(n17349), .A2(n13810), .ZN(n17357) );
  AND2_X1 U17385 ( .A1(n17357), .A2(n17372), .ZN(n20842) );
  OAI21_X1 U17386 ( .B1(n20842), .B2(n17273), .A(n13811), .ZN(P2_U2819) );
  INV_X1 U17387 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13815) );
  NAND2_X1 U17388 ( .A1(n17307), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13813) );
  NAND2_X1 U17389 ( .A1(n17305), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13812) );
  AND2_X1 U17390 ( .A1(n13813), .A2(n13812), .ZN(n20163) );
  NOR2_X1 U17391 ( .A1(n13857), .A2(n20163), .ZN(n13853) );
  AOI21_X1 U17392 ( .B1(n14556), .B2(P2_EAX_REG_4__SCAN_IN), .A(n13853), .ZN(
        n13814) );
  OAI21_X1 U17393 ( .B1(n13907), .B2(n13815), .A(n13814), .ZN(P2_U2971) );
  INV_X1 U17394 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n13819) );
  INV_X1 U17395 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n13817) );
  NAND2_X1 U17396 ( .A1(n17305), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13816) );
  OAI21_X1 U17397 ( .B1(n17305), .B2(n13817), .A(n13816), .ZN(n16535) );
  NAND2_X1 U17398 ( .A1(n13942), .A2(n16535), .ZN(n13938) );
  NAND2_X1 U17399 ( .A1(n14556), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n13818) );
  OAI211_X1 U17400 ( .C1(n13907), .C2(n13819), .A(n13938), .B(n13818), .ZN(
        P2_U2978) );
  INV_X1 U17401 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n13823) );
  INV_X1 U17402 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n13821) );
  NAND2_X1 U17403 ( .A1(n17305), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13820) );
  OAI21_X1 U17404 ( .B1(n17305), .B2(n13821), .A(n13820), .ZN(n16550) );
  NAND2_X1 U17405 ( .A1(n13942), .A2(n16550), .ZN(n13945) );
  NAND2_X1 U17406 ( .A1(n14556), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n13822) );
  OAI211_X1 U17407 ( .C1(n13907), .C2(n13823), .A(n13945), .B(n13822), .ZN(
        P2_U2976) );
  INV_X1 U17408 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n13827) );
  INV_X1 U17409 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n13825) );
  NAND2_X1 U17410 ( .A1(n17305), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13824) );
  OAI21_X1 U17411 ( .B1(n17305), .B2(n13825), .A(n13824), .ZN(n16557) );
  NAND2_X1 U17412 ( .A1(n13942), .A2(n16557), .ZN(n13947) );
  NAND2_X1 U17413 ( .A1(n14556), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n13826) );
  OAI211_X1 U17414 ( .C1(n13907), .C2(n13827), .A(n13947), .B(n13826), .ZN(
        P2_U2975) );
  INV_X1 U17415 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13831) );
  INV_X1 U17416 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n13829) );
  NAND2_X1 U17417 ( .A1(n17305), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13828) );
  OAI21_X1 U17418 ( .B1(n17305), .B2(n13829), .A(n13828), .ZN(n20168) );
  NAND2_X1 U17419 ( .A1(n13942), .A2(n20168), .ZN(n13916) );
  NAND2_X1 U17420 ( .A1(n14556), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n13830) );
  OAI211_X1 U17421 ( .C1(n13907), .C2(n13831), .A(n13916), .B(n13830), .ZN(
        P2_U2972) );
  INV_X1 U17422 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n13835) );
  INV_X1 U17423 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n13833) );
  NAND2_X1 U17424 ( .A1(n17305), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13832) );
  OAI21_X1 U17425 ( .B1(n17305), .B2(n13833), .A(n13832), .ZN(n16521) );
  NAND2_X1 U17426 ( .A1(n13942), .A2(n16521), .ZN(n13932) );
  NAND2_X1 U17427 ( .A1(n14556), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n13834) );
  OAI211_X1 U17428 ( .C1(n13907), .C2(n13835), .A(n13932), .B(n13834), .ZN(
        P2_U2980) );
  INV_X1 U17429 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13889) );
  INV_X1 U17430 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19354) );
  NAND2_X1 U17431 ( .A1(n17305), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13836) );
  OAI21_X1 U17432 ( .B1(n17305), .B2(n19354), .A(n13836), .ZN(n16601) );
  INV_X1 U17433 ( .A(n16601), .ZN(n20153) );
  NOR2_X1 U17434 ( .A1(n13857), .A2(n20153), .ZN(n13846) );
  AOI21_X1 U17435 ( .B1(n14556), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13846), .ZN(
        n13837) );
  OAI21_X1 U17436 ( .B1(n13889), .B2(n13907), .A(n13837), .ZN(P2_U2954) );
  INV_X1 U17437 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13841) );
  INV_X1 U17438 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n13839) );
  INV_X1 U17439 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13838) );
  MUX2_X1 U17440 ( .A(n13839), .B(n13838), .S(n17305), .Z(n17309) );
  NOR2_X1 U17441 ( .A1(n13857), .A2(n17309), .ZN(n13849) );
  AOI21_X1 U17442 ( .B1(n14556), .B2(P2_EAX_REG_6__SCAN_IN), .A(n13849), .ZN(
        n13840) );
  OAI21_X1 U17443 ( .B1(n13841), .B2(n13907), .A(n13840), .ZN(P2_U2973) );
  INV_X1 U17444 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13845) );
  NAND2_X1 U17445 ( .A1(n17307), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13843) );
  NAND2_X1 U17446 ( .A1(n17305), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13842) );
  NOR2_X1 U17447 ( .A1(n13857), .A2(n22063), .ZN(n13851) );
  AOI21_X1 U17448 ( .B1(n14556), .B2(P2_EAX_REG_3__SCAN_IN), .A(n13851), .ZN(
        n13844) );
  OAI21_X1 U17449 ( .B1(n13845), .B2(n13907), .A(n13844), .ZN(P2_U2970) );
  INV_X1 U17450 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13848) );
  AOI21_X1 U17451 ( .B1(n14556), .B2(P2_EAX_REG_2__SCAN_IN), .A(n13846), .ZN(
        n13847) );
  OAI21_X1 U17452 ( .B1(n13848), .B2(n13907), .A(n13847), .ZN(P2_U2969) );
  INV_X1 U17453 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13900) );
  AOI21_X1 U17454 ( .B1(n14556), .B2(P2_EAX_REG_22__SCAN_IN), .A(n13849), .ZN(
        n13850) );
  OAI21_X1 U17455 ( .B1(n13900), .B2(n13907), .A(n13850), .ZN(P2_U2958) );
  INV_X1 U17456 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13903) );
  AOI21_X1 U17457 ( .B1(n14556), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13851), .ZN(
        n13852) );
  OAI21_X1 U17458 ( .B1(n13903), .B2(n13907), .A(n13852), .ZN(P2_U2955) );
  INV_X1 U17459 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13893) );
  AOI21_X1 U17460 ( .B1(n14556), .B2(P2_EAX_REG_20__SCAN_IN), .A(n13853), .ZN(
        n13854) );
  OAI21_X1 U17461 ( .B1(n13893), .B2(n13907), .A(n13854), .ZN(P2_U2956) );
  INV_X1 U17462 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13858) );
  INV_X1 U17463 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n13855) );
  INV_X1 U17464 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14162) );
  MUX2_X1 U17465 ( .A(n13855), .B(n14162), .S(n17305), .Z(n16627) );
  INV_X1 U17466 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13856) );
  OAI222_X1 U17467 ( .A1(n13858), .A2(n13907), .B1(n13857), .B2(n16627), .C1(
        n13856), .C2(n13958), .ZN(P2_U2982) );
  NOR2_X1 U17468 ( .A1(n12537), .A2(n13869), .ZN(n13860) );
  NAND2_X1 U17469 ( .A1(n13860), .A2(n14486), .ZN(n14396) );
  NAND2_X1 U17470 ( .A1(n21517), .A2(n21644), .ZN(n20869) );
  INV_X1 U17471 ( .A(n20869), .ZN(n14719) );
  AOI21_X1 U17472 ( .B1(n14396), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14719), 
        .ZN(n13859) );
  NAND2_X1 U17473 ( .A1(n14056), .A2(n13859), .ZN(P1_U2801) );
  OAI22_X1 U17474 ( .A1(n15557), .A2(n13863), .B1(n13861), .B2(n13860), .ZN(
        n20867) );
  NOR3_X1 U17475 ( .A1(n13864), .A2(n13863), .A3(n13862), .ZN(n13865) );
  NOR2_X1 U17476 ( .A1(n13865), .A2(n21739), .ZN(n21740) );
  NOR2_X1 U17477 ( .A1(n20867), .A2(n21740), .ZN(n17514) );
  NOR2_X1 U17478 ( .A1(n17514), .A2(n20866), .ZN(n20875) );
  INV_X1 U17479 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13874) );
  NOR2_X1 U17480 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  MUX2_X1 U17481 ( .A(n13868), .B(n15524), .S(n15557), .Z(n13872) );
  NAND2_X1 U17482 ( .A1(n13870), .A2(n13869), .ZN(n13871) );
  AOI21_X1 U17483 ( .B1(n13872), .B2(n13871), .A(n14017), .ZN(n17511) );
  NAND2_X1 U17484 ( .A1(n20875), .A2(n17511), .ZN(n13873) );
  OAI21_X1 U17485 ( .B1(n20875), .B2(n13874), .A(n13873), .ZN(P1_U3484) );
  OR2_X1 U17486 ( .A1(n11426), .A2(n17617), .ZN(n13875) );
  INV_X1 U17487 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n17720) );
  INV_X1 U17488 ( .A(n20132), .ZN(n13879) );
  INV_X1 U17489 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13911) );
  INV_X1 U17490 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n21946) );
  OAI222_X1 U17491 ( .A1(n20101), .A2(n17720), .B1(n13977), .B2(n13911), .C1(
        n20845), .C2(n21946), .ZN(P2_U2921) );
  OAI21_X1 U17492 ( .B1(n13881), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13880), .ZN(n14045) );
  INV_X1 U17493 ( .A(n14045), .ZN(n13887) );
  NOR2_X1 U17494 ( .A1(n20051), .A2(n16008), .ZN(n14048) );
  INV_X1 U17495 ( .A(n13882), .ZN(n16004) );
  OAI21_X1 U17496 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16004), .A(
        n13883), .ZN(n14046) );
  OAI21_X1 U17497 ( .B1(n16930), .B2(n13884), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13885) );
  OAI21_X1 U17498 ( .B1(n16942), .B2(n14046), .A(n13885), .ZN(n13886) );
  AOI211_X1 U17499 ( .C1(n16939), .C2(n13887), .A(n14048), .B(n13886), .ZN(
        n13888) );
  OAI21_X1 U17500 ( .B1(n14052), .B2(n17306), .A(n13888), .ZN(P2_U3014) );
  INV_X1 U17501 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n13891) );
  INV_X1 U17502 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13890) );
  OAI222_X1 U17503 ( .A1(n13891), .A2(n20101), .B1(n13977), .B2(n13890), .C1(
        n20845), .C2(n13889), .ZN(P2_U2933) );
  INV_X1 U17504 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n13892) );
  INV_X1 U17505 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n20083) );
  OAI222_X1 U17506 ( .A1(n13892), .A2(n20101), .B1(n20845), .B2(n13815), .C1(
        n20083), .C2(n20132), .ZN(P2_U2947) );
  INV_X1 U17507 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13895) );
  INV_X1 U17508 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13894) );
  OAI222_X1 U17509 ( .A1(n13895), .A2(n20101), .B1(n13977), .B2(n13894), .C1(
        n20845), .C2(n13893), .ZN(P2_U2931) );
  INV_X1 U17510 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13897) );
  INV_X1 U17511 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13937) );
  INV_X1 U17512 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n13896) );
  OAI222_X1 U17513 ( .A1(n13897), .A2(n20101), .B1(n13977), .B2(n13937), .C1(
        n20845), .C2(n13896), .ZN(P2_U2923) );
  INV_X1 U17514 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13899) );
  INV_X1 U17515 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13944) );
  INV_X1 U17516 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n13898) );
  OAI222_X1 U17517 ( .A1(n13899), .A2(n20101), .B1(n13977), .B2(n13944), .C1(
        n20845), .C2(n13898), .ZN(P2_U2925) );
  INV_X1 U17518 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n13902) );
  INV_X1 U17519 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13901) );
  OAI222_X1 U17520 ( .A1(n13902), .A2(n20101), .B1(n13977), .B2(n13901), .C1(
        n20845), .C2(n13900), .ZN(P2_U2929) );
  INV_X1 U17521 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n13904) );
  INV_X1 U17522 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16592) );
  OAI222_X1 U17523 ( .A1(n13904), .A2(n20101), .B1(n13977), .B2(n16592), .C1(
        n20845), .C2(n13903), .ZN(P2_U2932) );
  INV_X1 U17524 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n13906) );
  INV_X1 U17525 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13931) );
  INV_X1 U17526 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13905) );
  OAI222_X1 U17527 ( .A1(n13906), .A2(n20101), .B1(n13977), .B2(n13931), .C1(
        n20845), .C2(n13905), .ZN(P2_U2935) );
  INV_X1 U17528 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13918) );
  INV_X1 U17529 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n17713) );
  INV_X1 U17530 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n21865) );
  OAI222_X1 U17531 ( .A1(n13977), .A2(n13918), .B1(n20101), .B2(n17713), .C1(
        n20845), .C2(n21865), .ZN(P2_U2930) );
  NAND2_X1 U17532 ( .A1(n13955), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13910) );
  INV_X1 U17533 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n13909) );
  NAND2_X1 U17534 ( .A1(n17305), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13908) );
  OAI21_X1 U17535 ( .B1(n17305), .B2(n13909), .A(n13908), .ZN(n16507) );
  NAND2_X1 U17536 ( .A1(n13942), .A2(n16507), .ZN(n13914) );
  OAI211_X1 U17537 ( .C1(n13911), .C2(n13958), .A(n13910), .B(n13914), .ZN(
        P2_U2966) );
  INV_X1 U17538 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20108) );
  NAND2_X1 U17539 ( .A1(n13955), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13913) );
  INV_X1 U17540 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18642) );
  NAND2_X1 U17541 ( .A1(n17305), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13912) );
  OAI21_X1 U17542 ( .B1(n17305), .B2(n18642), .A(n13912), .ZN(n16527) );
  NAND2_X1 U17543 ( .A1(n13942), .A2(n16527), .ZN(n13935) );
  OAI211_X1 U17544 ( .C1(n20108), .C2(n13958), .A(n13913), .B(n13935), .ZN(
        P2_U2979) );
  INV_X1 U17545 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20104) );
  NAND2_X1 U17546 ( .A1(n13955), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13915) );
  OAI211_X1 U17547 ( .C1(n20104), .C2(n13958), .A(n13915), .B(n13914), .ZN(
        P2_U2981) );
  NAND2_X1 U17548 ( .A1(n13955), .A2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13917) );
  OAI211_X1 U17549 ( .C1(n13958), .C2(n13918), .A(n13917), .B(n13916), .ZN(
        P2_U2957) );
  INV_X1 U17550 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20118) );
  NAND2_X1 U17551 ( .A1(n13955), .A2(P2_LWORD_REG_7__SCAN_IN), .ZN(n13921) );
  INV_X1 U17552 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n13920) );
  NAND2_X1 U17553 ( .A1(n17305), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13919) );
  OAI21_X1 U17554 ( .B1(n17305), .B2(n13920), .A(n13919), .ZN(n16565) );
  NAND2_X1 U17555 ( .A1(n13942), .A2(n16565), .ZN(n13950) );
  OAI211_X1 U17556 ( .C1(n13958), .C2(n20118), .A(n13921), .B(n13950), .ZN(
        P2_U2974) );
  INV_X1 U17557 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13924) );
  NAND2_X1 U17558 ( .A1(n13955), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n13923) );
  INV_X1 U17559 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19345) );
  NAND2_X1 U17560 ( .A1(n17305), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13922) );
  OAI21_X1 U17561 ( .B1(n17305), .B2(n19345), .A(n13922), .ZN(n16617) );
  NAND2_X1 U17562 ( .A1(n13942), .A2(n16617), .ZN(n13929) );
  OAI211_X1 U17563 ( .C1(n13958), .C2(n13924), .A(n13923), .B(n13929), .ZN(
        P2_U2967) );
  INV_X1 U17564 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13928) );
  NAND2_X1 U17565 ( .A1(n13955), .A2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13927) );
  NAND2_X1 U17566 ( .A1(n17307), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13926) );
  NAND2_X1 U17567 ( .A1(n17305), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13925) );
  AND2_X1 U17568 ( .A1(n13926), .A2(n13925), .ZN(n20148) );
  INV_X1 U17569 ( .A(n20148), .ZN(n16608) );
  NAND2_X1 U17570 ( .A1(n13942), .A2(n16608), .ZN(n13956) );
  OAI211_X1 U17571 ( .C1(n13958), .C2(n13928), .A(n13927), .B(n13956), .ZN(
        P2_U2953) );
  NAND2_X1 U17572 ( .A1(n13955), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13930) );
  OAI211_X1 U17573 ( .C1(n13931), .C2(n13958), .A(n13930), .B(n13929), .ZN(
        P2_U2952) );
  INV_X1 U17574 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13934) );
  NAND2_X1 U17575 ( .A1(n13955), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13933) );
  OAI211_X1 U17576 ( .C1(n13958), .C2(n13934), .A(n13933), .B(n13932), .ZN(
        P2_U2965) );
  NAND2_X1 U17577 ( .A1(n13955), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13936) );
  OAI211_X1 U17578 ( .C1(n13937), .C2(n13958), .A(n13936), .B(n13935), .ZN(
        P2_U2964) );
  INV_X1 U17579 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13940) );
  NAND2_X1 U17580 ( .A1(n13955), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13939) );
  OAI211_X1 U17581 ( .C1(n13958), .C2(n13940), .A(n13939), .B(n13938), .ZN(
        P2_U2963) );
  NAND2_X1 U17582 ( .A1(n13955), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13943) );
  INV_X1 U17583 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18639) );
  NAND2_X1 U17584 ( .A1(n17305), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13941) );
  OAI21_X1 U17585 ( .B1(n17305), .B2(n18639), .A(n13941), .ZN(n16543) );
  NAND2_X1 U17586 ( .A1(n13942), .A2(n16543), .ZN(n13953) );
  OAI211_X1 U17587 ( .C1(n13944), .C2(n13958), .A(n13943), .B(n13953), .ZN(
        P2_U2962) );
  INV_X1 U17588 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n21823) );
  NAND2_X1 U17589 ( .A1(n13955), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13946) );
  OAI211_X1 U17590 ( .C1(n13958), .C2(n21823), .A(n13946), .B(n13945), .ZN(
        P2_U2961) );
  INV_X1 U17591 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13949) );
  NAND2_X1 U17592 ( .A1(n13955), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13948) );
  OAI211_X1 U17593 ( .C1(n13958), .C2(n13949), .A(n13948), .B(n13947), .ZN(
        P2_U2960) );
  INV_X1 U17594 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13952) );
  NAND2_X1 U17595 ( .A1(n13955), .A2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13951) );
  OAI211_X1 U17596 ( .C1(n13958), .C2(n13952), .A(n13951), .B(n13950), .ZN(
        P2_U2959) );
  INV_X1 U17597 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20112) );
  NAND2_X1 U17598 ( .A1(n13955), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13954) );
  OAI211_X1 U17599 ( .C1(n20112), .C2(n13958), .A(n13954), .B(n13953), .ZN(
        P2_U2977) );
  INV_X1 U17600 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n20128) );
  NAND2_X1 U17601 ( .A1(n13955), .A2(P2_LWORD_REG_1__SCAN_IN), .ZN(n13957) );
  OAI211_X1 U17602 ( .C1(n13958), .C2(n20128), .A(n13957), .B(n13956), .ZN(
        P2_U2968) );
  NAND2_X1 U17603 ( .A1(n13959), .A2(n11078), .ZN(n13960) );
  NAND2_X1 U17604 ( .A1(n13961), .A2(n13960), .ZN(n13967) );
  NAND3_X1 U17605 ( .A1(n17349), .A2(n13963), .A3(n13962), .ZN(n13964) );
  INV_X1 U17606 ( .A(n17347), .ZN(n13966) );
  NAND2_X1 U17607 ( .A1(n17345), .A2(n13966), .ZN(n13994) );
  NAND2_X1 U17608 ( .A1(n17361), .A2(n17372), .ZN(n13970) );
  NOR2_X1 U17609 ( .A1(n17376), .A2(n17273), .ZN(n13968) );
  NOR2_X1 U17610 ( .A1(n17375), .A2(n13968), .ZN(n13969) );
  AND2_X1 U17611 ( .A1(n13970), .A2(n13969), .ZN(n20798) );
  INV_X1 U17612 ( .A(n20798), .ZN(n17298) );
  INV_X1 U17613 ( .A(n13971), .ZN(n20803) );
  INV_X1 U17614 ( .A(n13972), .ZN(n13973) );
  AND2_X1 U17615 ( .A1(n13974), .A2(n13973), .ZN(n13975) );
  OR3_X1 U17616 ( .A1(n20798), .A2(n20803), .A3(n17355), .ZN(n13976) );
  OAI21_X1 U17617 ( .B1(n17298), .B2(n17362), .A(n13976), .ZN(P2_U3595) );
  INV_X1 U17618 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13979) );
  INV_X1 U17619 ( .A(n20845), .ZN(n20129) );
  AOI22_X1 U17620 ( .A1(n14053), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n20129), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13978) );
  OAI21_X1 U17621 ( .B1(n20101), .B2(n13979), .A(n13978), .ZN(P2_U2928) );
  INV_X1 U17622 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13981) );
  AOI22_X1 U17623 ( .A1(n14053), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n20129), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13980) );
  OAI21_X1 U17624 ( .B1(n20101), .B2(n13981), .A(n13980), .ZN(P2_U2924) );
  INV_X1 U17625 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13983) );
  AOI22_X1 U17626 ( .A1(n14053), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n20129), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13982) );
  OAI21_X1 U17627 ( .B1(n20101), .B2(n13983), .A(n13982), .ZN(P2_U2922) );
  INV_X1 U17628 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n13985) );
  AOI22_X1 U17629 ( .A1(n14053), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n20129), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13984) );
  OAI21_X1 U17630 ( .B1(n20101), .B2(n13985), .A(n13984), .ZN(P2_U2934) );
  INV_X1 U17631 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13987) );
  AOI22_X1 U17632 ( .A1(n14053), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n20129), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13986) );
  OAI21_X1 U17633 ( .B1(n20101), .B2(n13987), .A(n13986), .ZN(P2_U2927) );
  INV_X1 U17634 ( .A(n14206), .ZN(n13988) );
  AOI22_X1 U17635 ( .A1(n14204), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20800), .B2(n17269), .ZN(n13990) );
  INV_X1 U17636 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16041) );
  NOR2_X1 U17637 ( .A1(n10286), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13991) );
  OAI211_X1 U17638 ( .C1(n20854), .C2(n16041), .A(n13989), .B(n13991), .ZN(
        n13992) );
  INV_X1 U17639 ( .A(n13992), .ZN(n13993) );
  NAND2_X1 U17640 ( .A1(n13994), .A2(n9919), .ZN(n13995) );
  MUX2_X1 U17641 ( .A(n14052), .B(n13996), .S(n16503), .Z(n13997) );
  OAI21_X1 U17642 ( .B1(n20133), .B2(n20076), .A(n13997), .ZN(P2_U2887) );
  INV_X1 U17643 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15991) );
  AOI21_X1 U17644 ( .B1(n13999), .B2(n21897), .A(n13998), .ZN(n14021) );
  NAND2_X1 U17645 ( .A1(n14001), .A2(n14000), .ZN(n14002) );
  XNOR2_X1 U17646 ( .A(n14002), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14022) );
  AOI22_X1 U17647 ( .A1(n16939), .A2(n14021), .B1(n16899), .B2(n14022), .ZN(
        n14003) );
  OR2_X1 U17648 ( .A1(n16877), .A2(n20732), .ZN(n14023) );
  OAI211_X1 U17649 ( .C1(n16921), .C2(n15991), .A(n14003), .B(n14023), .ZN(
        n14004) );
  AOI21_X1 U17650 ( .B1(n16924), .B2(n15991), .A(n14004), .ZN(n14005) );
  OAI21_X1 U17651 ( .B1(n15994), .B2(n17306), .A(n14005), .ZN(P2_U3013) );
  NAND2_X1 U17652 ( .A1(n17269), .A2(n20831), .ZN(n20416) );
  NAND2_X1 U17653 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20253) );
  AND2_X1 U17654 ( .A1(n20296), .A2(n20800), .ZN(n20358) );
  AOI21_X1 U17655 ( .B1(n14204), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n20358), .ZN(n14006) );
  NAND2_X1 U17656 ( .A1(n14009), .A2(n14008), .ZN(n14010) );
  NOR2_X1 U17657 ( .A1(n15994), .A2(n16503), .ZN(n14011) );
  AOI21_X1 U17658 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n16503), .A(n14011), .ZN(
        n14012) );
  OAI21_X1 U17659 ( .B1(n20134), .B2(n20076), .A(n14012), .ZN(P2_U2886) );
  NOR2_X1 U17660 ( .A1(n14392), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14013) );
  OR2_X1 U17661 ( .A1(n14014), .A2(n14013), .ZN(n14896) );
  OAI22_X1 U17662 ( .A1(n15557), .A2(n15524), .B1(n14015), .B2(n14391), .ZN(
        n14016) );
  INV_X2 U17663 ( .A(n20975), .ZN(n14927) );
  OAI222_X1 U17664 ( .A1(n14896), .A2(n14959), .B1(n12555), .B2(n20978), .C1(
        n14903), .C2(n14927), .ZN(P1_U2872) );
  INV_X1 U17665 ( .A(n14018), .ZN(n14019) );
  AOI211_X1 U17666 ( .C1(n21897), .C2(n14020), .A(n14019), .B(n14049), .ZN(
        n14033) );
  INV_X1 U17667 ( .A(n14021), .ZN(n14025) );
  NAND2_X1 U17668 ( .A1(n17221), .A2(n14022), .ZN(n14024) );
  OAI211_X1 U17669 ( .C1(n17234), .C2(n14025), .A(n14024), .B(n14023), .ZN(
        n14032) );
  OR2_X1 U17670 ( .A1(n14027), .A2(n14026), .ZN(n14028) );
  NAND2_X1 U17671 ( .A1(n14029), .A2(n14028), .ZN(n20828) );
  INV_X1 U17672 ( .A(n20828), .ZN(n14030) );
  OAI22_X1 U17673 ( .A1(n14030), .A2(n17256), .B1(n14525), .B2(n21897), .ZN(
        n14031) );
  NOR3_X1 U17674 ( .A1(n14033), .A2(n14032), .A3(n14031), .ZN(n14034) );
  OAI21_X1 U17675 ( .B1(n15994), .B2(n17241), .A(n14034), .ZN(P2_U3045) );
  INV_X1 U17676 ( .A(n14896), .ZN(n14038) );
  INV_X1 U17677 ( .A(n15396), .ZN(n14035) );
  AOI21_X1 U17678 ( .B1(n14035), .B2(n21047), .A(n15586), .ZN(n14036) );
  AOI211_X1 U17679 ( .C1(n14038), .C2(n21027), .A(n14037), .B(n14036), .ZN(
        n14039) );
  OAI21_X1 U17680 ( .B1(n21028), .B2(n15373), .A(n15586), .ZN(n21046) );
  OAI211_X1 U17681 ( .C1(n14040), .C2(n21012), .A(n14039), .B(n21046), .ZN(
        P1_U3031) );
  OR2_X1 U17682 ( .A1(n14042), .A2(n14041), .ZN(n14044) );
  AND2_X1 U17683 ( .A1(n14044), .A2(n14043), .ZN(n16005) );
  OAI22_X1 U17684 ( .A1(n17266), .A2(n14046), .B1(n17234), .B2(n14045), .ZN(
        n14047) );
  AOI211_X1 U17685 ( .C1(n16005), .C2(n12994), .A(n14048), .B(n14047), .ZN(
        n14051) );
  MUX2_X1 U17686 ( .A(n14049), .B(n14525), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n14050) );
  OAI211_X1 U17687 ( .C1(n17241), .C2(n14052), .A(n14051), .B(n14050), .ZN(
        P2_U3046) );
  AOI222_X1 U17688 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n14053), .B1(n20130), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .C1(n20129), .C2(
        P2_UWORD_REG_9__SCAN_IN), .ZN(n14054) );
  INV_X1 U17689 ( .A(n14054), .ZN(P2_U2926) );
  INV_X1 U17690 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14102) );
  OR2_X2 U17691 ( .A1(n20988), .A2(n9762), .ZN(n14215) );
  NAND2_X1 U17692 ( .A1(n15614), .A2(DATAI_5_), .ZN(n14058) );
  NAND2_X1 U17693 ( .A1(n15615), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14057) );
  AND2_X1 U17694 ( .A1(n14058), .A2(n14057), .ZN(n21092) );
  NOR2_X1 U17695 ( .A1(n14242), .A2(n21092), .ZN(n14218) );
  AOI21_X1 U17696 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n20988), .A(n14218), 
        .ZN(n14059) );
  OAI21_X1 U17697 ( .B1(n14102), .B2(n14215), .A(n14059), .ZN(P1_U2942) );
  INV_X1 U17698 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U17699 ( .A1(n15614), .A2(DATAI_7_), .ZN(n14061) );
  NAND2_X1 U17700 ( .A1(n15615), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14060) );
  NOR2_X1 U17701 ( .A1(n14242), .A2(n21108), .ZN(n14072) );
  AOI21_X1 U17702 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n20988), .A(n14072), 
        .ZN(n14062) );
  OAI21_X1 U17703 ( .B1(n14139), .B2(n14215), .A(n14062), .ZN(P1_U2959) );
  INV_X1 U17704 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n14142) );
  NAND2_X1 U17705 ( .A1(n15614), .A2(DATAI_6_), .ZN(n14064) );
  NAND2_X1 U17706 ( .A1(n15615), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14063) );
  AND2_X1 U17707 ( .A1(n14064), .A2(n14063), .ZN(n21097) );
  NOR2_X1 U17708 ( .A1(n14242), .A2(n21097), .ZN(n14237) );
  AOI21_X1 U17709 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n20988), .A(n14237), 
        .ZN(n14065) );
  OAI21_X1 U17710 ( .B1(n14142), .B2(n14215), .A(n14065), .ZN(P1_U2958) );
  INV_X1 U17711 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14110) );
  INV_X1 U17712 ( .A(DATAI_3_), .ZN(n14067) );
  NAND2_X1 U17713 ( .A1(n15615), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14066) );
  OAI21_X1 U17714 ( .B1(n15615), .B2(n14067), .A(n14066), .ZN(n21078) );
  INV_X1 U17715 ( .A(n21078), .ZN(n15063) );
  NOR2_X1 U17716 ( .A1(n14242), .A2(n15063), .ZN(n14235) );
  AOI21_X1 U17717 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n20988), .A(n14235), 
        .ZN(n14068) );
  OAI21_X1 U17718 ( .B1(n14110), .B2(n14215), .A(n14068), .ZN(P1_U2940) );
  INV_X1 U17719 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14107) );
  NAND2_X1 U17720 ( .A1(n15614), .A2(DATAI_1_), .ZN(n14070) );
  NAND2_X1 U17721 ( .A1(n15615), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14069) );
  AND2_X1 U17722 ( .A1(n14070), .A2(n14069), .ZN(n21062) );
  NOR2_X1 U17723 ( .A1(n14242), .A2(n21062), .ZN(n14216) );
  AOI21_X1 U17724 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n20988), .A(n14216), 
        .ZN(n14071) );
  OAI21_X1 U17725 ( .B1(n14107), .B2(n14215), .A(n14071), .ZN(P1_U2938) );
  INV_X1 U17726 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14119) );
  AOI21_X1 U17727 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n20988), .A(n14072), 
        .ZN(n14073) );
  OAI21_X1 U17728 ( .B1(n14119), .B2(n14215), .A(n14073), .ZN(P1_U2944) );
  INV_X1 U17729 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21797) );
  INV_X1 U17730 ( .A(DATAI_9_), .ZN(n14075) );
  INV_X1 U17731 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14074) );
  MUX2_X1 U17732 ( .A(n14075), .B(n14074), .S(n15615), .Z(n15053) );
  NOR2_X1 U17733 ( .A1(n14242), .A2(n15053), .ZN(n14226) );
  AOI21_X1 U17734 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n20988), .A(n14226), 
        .ZN(n14076) );
  OAI21_X1 U17735 ( .B1(n21797), .B2(n14215), .A(n14076), .ZN(P1_U2946) );
  INV_X1 U17736 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n21910) );
  NAND2_X1 U17737 ( .A1(n15614), .A2(DATAI_4_), .ZN(n14078) );
  NAND2_X1 U17738 ( .A1(n15615), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14077) );
  AND2_X1 U17739 ( .A1(n14078), .A2(n14077), .ZN(n21084) );
  NOR2_X1 U17740 ( .A1(n14242), .A2(n21084), .ZN(n14232) );
  AOI21_X1 U17741 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n20988), .A(n14232), 
        .ZN(n14079) );
  OAI21_X1 U17742 ( .B1(n21910), .B2(n14215), .A(n14079), .ZN(P1_U2941) );
  INV_X1 U17743 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14984) );
  INV_X1 U17744 ( .A(DATAI_10_), .ZN(n14080) );
  INV_X1 U17745 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17675) );
  MUX2_X1 U17746 ( .A(n14080), .B(n17675), .S(n15615), .Z(n15051) );
  NOR2_X1 U17747 ( .A1(n14242), .A2(n15051), .ZN(n14229) );
  AOI21_X1 U17748 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n20988), .A(n14229), 
        .ZN(n14081) );
  OAI21_X1 U17749 ( .B1(n14984), .B2(n14215), .A(n14081), .ZN(P1_U2947) );
  INV_X1 U17750 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n22013) );
  NAND2_X1 U17751 ( .A1(n15614), .A2(DATAI_2_), .ZN(n14083) );
  NAND2_X1 U17752 ( .A1(n15615), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14082) );
  NOR2_X1 U17753 ( .A1(n14242), .A2(n21072), .ZN(n14249) );
  AOI21_X1 U17754 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n20988), .A(n14249), 
        .ZN(n14084) );
  OAI21_X1 U17755 ( .B1(n22013), .B2(n14215), .A(n14084), .ZN(P1_U2939) );
  AND2_X1 U17756 ( .A1(n17497), .A2(n12543), .ZN(n14085) );
  AND2_X1 U17757 ( .A1(n12537), .A2(n21060), .ZN(n14087) );
  NOR2_X1 U17758 ( .A1(n21647), .A2(n21644), .ZN(n15558) );
  INV_X1 U17759 ( .A(n15558), .ZN(n17600) );
  INV_X1 U17760 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n21830) );
  INV_X1 U17761 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21955) );
  INV_X1 U17762 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n14088) );
  OAI222_X1 U17763 ( .A1(n20985), .A2(n21830), .B1(n20982), .B2(n21955), .C1(
        n14088), .C2(n14160), .ZN(P1_U2936) );
  INV_X1 U17764 ( .A(n14242), .ZN(n14095) );
  INV_X1 U17765 ( .A(DATAI_13_), .ZN(n14090) );
  INV_X1 U17766 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14089) );
  MUX2_X1 U17767 ( .A(n14090), .B(n14089), .S(n15615), .Z(n15045) );
  INV_X1 U17768 ( .A(n15045), .ZN(n14091) );
  NAND2_X1 U17769 ( .A1(n14095), .A2(n14091), .ZN(n20990) );
  NAND2_X1 U17770 ( .A1(n20988), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n14092) );
  OAI211_X1 U17771 ( .C1(n14215), .C2(n14968), .A(n20990), .B(n14092), .ZN(
        P1_U2950) );
  INV_X1 U17772 ( .A(DATAI_0_), .ZN(n14094) );
  NAND2_X1 U17773 ( .A1(n15615), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14093) );
  OAI21_X1 U17774 ( .B1(n15615), .B2(n14094), .A(n14093), .ZN(n15607) );
  NAND2_X1 U17775 ( .A1(n14095), .A2(n15607), .ZN(n14098) );
  NAND2_X1 U17776 ( .A1(n20988), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n14096) );
  OAI211_X1 U17777 ( .C1(n14215), .C2(n21955), .A(n14098), .B(n14096), .ZN(
        P1_U2952) );
  INV_X1 U17778 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14126) );
  NAND2_X1 U17779 ( .A1(n20988), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14097) );
  OAI211_X1 U17780 ( .C1(n14215), .C2(n14126), .A(n14098), .B(n14097), .ZN(
        P1_U2937) );
  INV_X1 U17781 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n14100) );
  INV_X1 U17782 ( .A(n20982), .ZN(n20980) );
  INV_X1 U17783 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14099) );
  OAI222_X1 U17784 ( .A1(n14100), .A2(n14160), .B1(n14153), .B2(n14968), .C1(
        n20985), .C2(n14099), .ZN(P1_U2907) );
  INV_X1 U17785 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n14103) );
  INV_X1 U17786 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n14101) );
  OAI222_X1 U17787 ( .A1(n14103), .A2(n14160), .B1(n14153), .B2(n14102), .C1(
        n20985), .C2(n14101), .ZN(P1_U2915) );
  INV_X1 U17788 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n14105) );
  INV_X1 U17789 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n14104) );
  OAI222_X1 U17790 ( .A1(n14105), .A2(n14160), .B1(n14153), .B2(n21910), .C1(
        n20985), .C2(n14104), .ZN(P1_U2916) );
  INV_X1 U17791 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n14108) );
  INV_X1 U17792 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n14106) );
  OAI222_X1 U17793 ( .A1(n14108), .A2(n14160), .B1(n14153), .B2(n14107), .C1(
        n20985), .C2(n14106), .ZN(P1_U2919) );
  INV_X1 U17794 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n14111) );
  INV_X1 U17795 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n14109) );
  OAI222_X1 U17796 ( .A1(n14111), .A2(n14160), .B1(n14153), .B2(n14110), .C1(
        n20985), .C2(n14109), .ZN(P1_U2917) );
  INV_X1 U17797 ( .A(P1_UWORD_REG_9__SCAN_IN), .ZN(n14113) );
  INV_X1 U17798 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14112) );
  OAI222_X1 U17799 ( .A1(n14113), .A2(n14160), .B1(n14153), .B2(n21797), .C1(
        n20985), .C2(n14112), .ZN(P1_U2911) );
  INV_X1 U17800 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n14115) );
  INV_X1 U17801 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14239) );
  INV_X1 U17802 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n14114) );
  OAI222_X1 U17803 ( .A1(n14115), .A2(n14160), .B1(n14153), .B2(n14239), .C1(
        n20985), .C2(n14114), .ZN(P1_U2914) );
  INV_X1 U17804 ( .A(P1_UWORD_REG_14__SCAN_IN), .ZN(n14117) );
  INV_X1 U17805 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14116) );
  OAI222_X1 U17806 ( .A1(n14117), .A2(n14160), .B1(n14153), .B2(n14963), .C1(
        n20985), .C2(n14116), .ZN(P1_U2906) );
  INV_X1 U17807 ( .A(P1_UWORD_REG_7__SCAN_IN), .ZN(n14120) );
  INV_X1 U17808 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n14118) );
  OAI222_X1 U17809 ( .A1(n14120), .A2(n14160), .B1(n14153), .B2(n14119), .C1(
        n20985), .C2(n14118), .ZN(P1_U2913) );
  INV_X1 U17810 ( .A(P1_UWORD_REG_11__SCAN_IN), .ZN(n14122) );
  INV_X1 U17811 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14121) );
  OAI222_X1 U17812 ( .A1(n14122), .A2(n14160), .B1(n14153), .B2(n14979), .C1(
        n20985), .C2(n14121), .ZN(P1_U2909) );
  INV_X1 U17813 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n14124) );
  INV_X1 U17814 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14256) );
  INV_X1 U17815 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14123) );
  OAI222_X1 U17816 ( .A1(n14124), .A2(n14160), .B1(n14153), .B2(n14256), .C1(
        n20985), .C2(n14123), .ZN(P1_U2908) );
  INV_X1 U17817 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n14127) );
  INV_X1 U17818 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n14125) );
  OAI222_X1 U17819 ( .A1(n14127), .A2(n14160), .B1(n14153), .B2(n14126), .C1(
        n20985), .C2(n14125), .ZN(P1_U2920) );
  INV_X1 U17820 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n14129) );
  INV_X1 U17821 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14253) );
  INV_X1 U17822 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n14128) );
  OAI222_X1 U17823 ( .A1(n14129), .A2(n14160), .B1(n20982), .B2(n14253), .C1(
        n20985), .C2(n14128), .ZN(P1_U2925) );
  INV_X1 U17824 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n14131) );
  INV_X1 U17825 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14223) );
  INV_X1 U17826 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n14130) );
  OAI222_X1 U17827 ( .A1(n14131), .A2(n14160), .B1(n20982), .B2(n14223), .C1(
        n20985), .C2(n14130), .ZN(P1_U2922) );
  INV_X1 U17828 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n14133) );
  INV_X1 U17829 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14231) );
  INV_X1 U17830 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n14132) );
  OAI222_X1 U17831 ( .A1(n14133), .A2(n14160), .B1(n20982), .B2(n14231), .C1(
        n20985), .C2(n14132), .ZN(P1_U2926) );
  INV_X1 U17832 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n14135) );
  INV_X1 U17833 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14228) );
  INV_X1 U17834 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n14134) );
  OAI222_X1 U17835 ( .A1(n14135), .A2(n14160), .B1(n20982), .B2(n14228), .C1(
        n20985), .C2(n14134), .ZN(P1_U2927) );
  INV_X1 U17836 ( .A(P1_LWORD_REG_8__SCAN_IN), .ZN(n14137) );
  INV_X1 U17837 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14244) );
  INV_X1 U17838 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n14136) );
  OAI222_X1 U17839 ( .A1(n14137), .A2(n14160), .B1(n20982), .B2(n14244), .C1(
        n20985), .C2(n14136), .ZN(P1_U2928) );
  INV_X1 U17840 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n14140) );
  INV_X1 U17841 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n14138) );
  OAI222_X1 U17842 ( .A1(n14140), .A2(n14160), .B1(n20982), .B2(n14139), .C1(
        n20985), .C2(n14138), .ZN(P1_U2929) );
  INV_X1 U17843 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n14143) );
  INV_X1 U17844 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n14141) );
  OAI222_X1 U17845 ( .A1(n14143), .A2(n14160), .B1(n20982), .B2(n14142), .C1(
        n20985), .C2(n14141), .ZN(P1_U2930) );
  INV_X1 U17846 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n14145) );
  INV_X1 U17847 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n14144) );
  OAI222_X1 U17848 ( .A1(n14145), .A2(n14160), .B1(n20982), .B2(n15058), .C1(
        n20985), .C2(n14144), .ZN(P1_U2931) );
  INV_X1 U17849 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n15061) );
  INV_X1 U17850 ( .A(P1_LWORD_REG_4__SCAN_IN), .ZN(n14146) );
  INV_X1 U17851 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n21879) );
  OAI222_X1 U17852 ( .A1(n20982), .A2(n15061), .B1(n14160), .B2(n14146), .C1(
        n20985), .C2(n21879), .ZN(P1_U2932) );
  INV_X1 U17853 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n14289) );
  INV_X1 U17854 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n22038) );
  INV_X1 U17855 ( .A(P1_LWORD_REG_2__SCAN_IN), .ZN(n14147) );
  OAI222_X1 U17856 ( .A1(n20982), .A2(n14289), .B1(n20985), .B2(n22038), .C1(
        n14147), .C2(n14160), .ZN(P1_U2934) );
  INV_X1 U17857 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n14149) );
  INV_X1 U17858 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n14148) );
  OAI222_X1 U17859 ( .A1(n14149), .A2(n14160), .B1(n14153), .B2(n22013), .C1(
        n14148), .C2(n20985), .ZN(P1_U2918) );
  INV_X1 U17860 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n14151) );
  INV_X1 U17861 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14994) );
  INV_X1 U17862 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n14150) );
  OAI222_X1 U17863 ( .A1(n14151), .A2(n14160), .B1(n14153), .B2(n14994), .C1(
        n14150), .C2(n20985), .ZN(P1_U2912) );
  INV_X1 U17864 ( .A(P1_UWORD_REG_10__SCAN_IN), .ZN(n14154) );
  INV_X1 U17865 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14152) );
  OAI222_X1 U17866 ( .A1(n14154), .A2(n14160), .B1(n14153), .B2(n14984), .C1(
        n14152), .C2(n20985), .ZN(P1_U2910) );
  INV_X1 U17867 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n14156) );
  INV_X1 U17868 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21990) );
  INV_X1 U17869 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n14155) );
  OAI222_X1 U17870 ( .A1(n14156), .A2(n14160), .B1(n20982), .B2(n21990), .C1(
        n14155), .C2(n20985), .ZN(P1_U2935) );
  INV_X1 U17871 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14158) );
  INV_X1 U17872 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n15042) );
  INV_X1 U17873 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n14157) );
  OAI222_X1 U17874 ( .A1(n14158), .A2(n14160), .B1(n20982), .B2(n15042), .C1(
        n14157), .C2(n20985), .ZN(P1_U2921) );
  INV_X1 U17875 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n14161) );
  INV_X1 U17876 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n15065) );
  INV_X1 U17877 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n14159) );
  OAI222_X1 U17878 ( .A1(n14161), .A2(n14160), .B1(n20982), .B2(n15065), .C1(
        n14159), .C2(n20985), .ZN(P1_U2933) );
  INV_X1 U17879 ( .A(DATAI_15_), .ZN(n14163) );
  MUX2_X1 U17880 ( .A(n14163), .B(n14162), .S(n15615), .Z(n15041) );
  OAI222_X1 U17881 ( .A1(n14215), .A2(n15042), .B1(n14242), .B2(n15041), .C1(
        n14164), .C2(n14158), .ZN(P1_U2967) );
  INV_X1 U17882 ( .A(n14165), .ZN(n14166) );
  INV_X1 U17883 ( .A(n15064), .ZN(n14167) );
  AOI22_X1 U17884 ( .A1(n14167), .A2(n15607), .B1(P1_EAX_REG_0__SCAN_IN), .B2(
        n15034), .ZN(n14168) );
  OAI21_X1 U17885 ( .B1(n14903), .B2(n15067), .A(n14168), .ZN(P1_U2904) );
  NAND2_X1 U17886 ( .A1(n20253), .A2(n20821), .ZN(n14169) );
  NOR2_X1 U17887 ( .A1(n20821), .A2(n20831), .ZN(n20609) );
  NAND2_X1 U17888 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20609), .ZN(
        n14200) );
  AND2_X1 U17889 ( .A1(n20548), .A2(n20800), .ZN(n20295) );
  AOI21_X1 U17890 ( .B1(n14204), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n20295), .ZN(n14170) );
  NAND2_X1 U17891 ( .A1(n14172), .A2(n14173), .ZN(n14176) );
  OR2_X1 U17892 ( .A1(n17283), .A2(n14177), .ZN(n14178) );
  NAND2_X2 U17893 ( .A1(n14179), .A2(n14180), .ZN(n14198) );
  MUX2_X1 U17894 ( .A(n14181), .B(n17320), .S(n20082), .Z(n14182) );
  OAI21_X1 U17895 ( .B1(n20817), .B2(n20076), .A(n14182), .ZN(P2_U2885) );
  OAI21_X1 U17896 ( .B1(n14185), .B2(n14184), .A(n14183), .ZN(n14895) );
  OAI222_X1 U17897 ( .A1(n14895), .A2(n15067), .B1(n15066), .B2(n21990), .C1(
        n15064), .C2(n21062), .ZN(P1_U2903) );
  XNOR2_X1 U17898 ( .A(n14186), .B(n14391), .ZN(n21055) );
  OAI222_X1 U17899 ( .A1(n21055), .A2(n14959), .B1(n12549), .B2(n20978), .C1(
        n14895), .C2(n14927), .ZN(P1_U2871) );
  INV_X2 U17900 ( .A(n20084), .ZN(n20093) );
  INV_X1 U17901 ( .A(n14191), .ZN(n14192) );
  NAND2_X1 U17902 ( .A1(n11073), .A2(n20181), .ZN(n14193) );
  INV_X1 U17903 ( .A(n16617), .ZN(n20139) );
  NAND2_X1 U17904 ( .A1(n20198), .A2(n16005), .ZN(n20095) );
  OAI211_X1 U17905 ( .C1(n20198), .C2(n16005), .A(n20095), .B(n22058), .ZN(
        n14196) );
  INV_X1 U17906 ( .A(n20085), .ZN(n22053) );
  AOI22_X1 U17907 ( .A1(n22053), .A2(n16005), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n20093), .ZN(n14195) );
  OAI211_X1 U17908 ( .C1(n22062), .C2(n20139), .A(n14196), .B(n14195), .ZN(
        P2_U2919) );
  BUF_X2 U17909 ( .A(n14199), .Z(n14213) );
  INV_X1 U17910 ( .A(n14200), .ZN(n14201) );
  NAND2_X1 U17911 ( .A1(n14201), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20657) );
  OAI211_X1 U17912 ( .C1(n14201), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n20657), .B(n20800), .ZN(n14202) );
  INV_X1 U17913 ( .A(n14202), .ZN(n14203) );
  AOI21_X1 U17914 ( .B1(n14204), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14203), .ZN(n14205) );
  OAI21_X2 U17915 ( .B1(n14213), .B2(n14206), .A(n14205), .ZN(n14305) );
  INV_X1 U17916 ( .A(n14305), .ZN(n14207) );
  NAND2_X1 U17917 ( .A1(n14207), .A2(n14208), .ZN(n14210) );
  INV_X1 U17918 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n21842) );
  MUX2_X1 U17919 ( .A(n21842), .B(n14213), .S(n20082), .Z(n14214) );
  OAI21_X1 U17920 ( .B1(n20199), .B2(n20076), .A(n14214), .ZN(P2_U2884) );
  AOI21_X1 U17921 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n20988), .A(n14216), 
        .ZN(n14217) );
  OAI21_X1 U17922 ( .B1(n21990), .B2(n14215), .A(n14217), .ZN(P1_U2953) );
  AOI21_X1 U17923 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n20988), .A(n14218), 
        .ZN(n14219) );
  OAI21_X1 U17924 ( .B1(n15058), .B2(n14215), .A(n14219), .ZN(P1_U2957) );
  INV_X1 U17925 ( .A(DATAI_14_), .ZN(n14221) );
  INV_X1 U17926 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14220) );
  MUX2_X1 U17927 ( .A(n14221), .B(n14220), .S(n15615), .Z(n15043) );
  NOR2_X1 U17928 ( .A1(n14242), .A2(n15043), .ZN(n14245) );
  AOI21_X1 U17929 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n20988), .A(n14245), 
        .ZN(n14222) );
  OAI21_X1 U17930 ( .B1(n14223), .B2(n14215), .A(n14222), .ZN(P1_U2966) );
  INV_X1 U17931 ( .A(DATAI_12_), .ZN(n14224) );
  INV_X1 U17932 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17671) );
  MUX2_X1 U17933 ( .A(n14224), .B(n17671), .S(n15615), .Z(n15048) );
  NOR2_X1 U17934 ( .A1(n14242), .A2(n15048), .ZN(n14254) );
  AOI21_X1 U17935 ( .B1(n20988), .B2(P1_LWORD_REG_12__SCAN_IN), .A(n14254), 
        .ZN(n14225) );
  OAI21_X1 U17936 ( .B1(n20983), .B2(n14215), .A(n14225), .ZN(P1_U2964) );
  AOI21_X1 U17937 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n20988), .A(n14226), 
        .ZN(n14227) );
  OAI21_X1 U17938 ( .B1(n14228), .B2(n14215), .A(n14227), .ZN(P1_U2961) );
  AOI21_X1 U17939 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n20988), .A(n14229), 
        .ZN(n14230) );
  OAI21_X1 U17940 ( .B1(n14231), .B2(n14215), .A(n14230), .ZN(P1_U2962) );
  AOI21_X1 U17941 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n20988), .A(n14232), 
        .ZN(n14233) );
  OAI21_X1 U17942 ( .B1(n15061), .B2(n14215), .A(n14233), .ZN(P1_U2956) );
  INV_X1 U17943 ( .A(DATAI_11_), .ZN(n21757) );
  INV_X1 U17944 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n17673) );
  MUX2_X1 U17945 ( .A(n21757), .B(n17673), .S(n15615), .Z(n15049) );
  NOR2_X1 U17946 ( .A1(n14242), .A2(n15049), .ZN(n14251) );
  AOI21_X1 U17947 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n20988), .A(n14251), 
        .ZN(n14234) );
  OAI21_X1 U17948 ( .B1(n14979), .B2(n14215), .A(n14234), .ZN(P1_U2948) );
  AOI21_X1 U17949 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n20988), .A(n14235), 
        .ZN(n14236) );
  OAI21_X1 U17950 ( .B1(n15065), .B2(n14215), .A(n14236), .ZN(P1_U2955) );
  AOI21_X1 U17951 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n20988), .A(n14237), 
        .ZN(n14238) );
  OAI21_X1 U17952 ( .B1(n14239), .B2(n14215), .A(n14238), .ZN(P1_U2943) );
  INV_X1 U17953 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n14240) );
  NOR2_X1 U17954 ( .A1(n15614), .A2(n14240), .ZN(n14241) );
  AOI21_X1 U17955 ( .B1(DATAI_8_), .B2(n15614), .A(n14241), .ZN(n15054) );
  NOR2_X1 U17956 ( .A1(n14242), .A2(n15054), .ZN(n14247) );
  AOI21_X1 U17957 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n20988), .A(n14247), 
        .ZN(n14243) );
  OAI21_X1 U17958 ( .B1(n14244), .B2(n14215), .A(n14243), .ZN(P1_U2960) );
  AOI21_X1 U17959 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n20988), .A(n14245), 
        .ZN(n14246) );
  OAI21_X1 U17960 ( .B1(n14963), .B2(n14215), .A(n14246), .ZN(P1_U2951) );
  AOI21_X1 U17961 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n20988), .A(n14247), 
        .ZN(n14248) );
  OAI21_X1 U17962 ( .B1(n14994), .B2(n14215), .A(n14248), .ZN(P1_U2945) );
  AOI21_X1 U17963 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n20988), .A(n14249), 
        .ZN(n14250) );
  OAI21_X1 U17964 ( .B1(n14289), .B2(n14215), .A(n14250), .ZN(P1_U2954) );
  AOI21_X1 U17965 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n20988), .A(n14251), 
        .ZN(n14252) );
  OAI21_X1 U17966 ( .B1(n14253), .B2(n14215), .A(n14252), .ZN(P1_U2963) );
  AOI21_X1 U17967 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n20988), .A(n14254), 
        .ZN(n14255) );
  OAI21_X1 U17968 ( .B1(n14256), .B2(n14215), .A(n14255), .ZN(P1_U2949) );
  AND2_X1 U17969 ( .A1(n14273), .A2(n14257), .ZN(n14258) );
  NOR2_X1 U17970 ( .A1(n14279), .A2(n14258), .ZN(n17171) );
  INV_X1 U17971 ( .A(n17171), .ZN(n14260) );
  AOI22_X1 U17972 ( .A1(n16634), .A2(n16543), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n20093), .ZN(n14259) );
  OAI21_X1 U17973 ( .B1(n14260), .B2(n16637), .A(n14259), .ZN(P2_U2909) );
  OR2_X1 U17974 ( .A1(n14264), .A2(n14263), .ZN(n14265) );
  AND2_X1 U17975 ( .A1(n14262), .A2(n14265), .ZN(n17206) );
  INV_X1 U17976 ( .A(n17206), .ZN(n14266) );
  INV_X1 U17977 ( .A(n16565), .ZN(n20184) );
  OAI222_X1 U17978 ( .A1(n20118), .A2(n20084), .B1(n14266), .B2(n16637), .C1(
        n22062), .C2(n20184), .ZN(P2_U2912) );
  NAND2_X1 U17979 ( .A1(n14262), .A2(n14268), .ZN(n14269) );
  NAND2_X1 U17980 ( .A1(n14267), .A2(n14269), .ZN(n17195) );
  INV_X1 U17981 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20116) );
  INV_X1 U17982 ( .A(n16557), .ZN(n14270) );
  OAI222_X1 U17983 ( .A1(n17195), .A2(n16637), .B1(n20084), .B2(n20116), .C1(
        n22062), .C2(n14270), .ZN(P2_U2911) );
  NAND2_X1 U17984 ( .A1(n14267), .A2(n14271), .ZN(n14272) );
  NAND2_X1 U17985 ( .A1(n14273), .A2(n14272), .ZN(n17181) );
  INV_X1 U17986 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20114) );
  INV_X1 U17987 ( .A(n16550), .ZN(n14274) );
  OAI222_X1 U17988 ( .A1(n17181), .A2(n16637), .B1(n20084), .B2(n20114), .C1(
        n22062), .C2(n14274), .ZN(P2_U2910) );
  INV_X1 U17989 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20120) );
  XNOR2_X1 U17990 ( .A(n14275), .B(n9938), .ZN(n17218) );
  INV_X1 U17991 ( .A(n17218), .ZN(n20064) );
  OAI222_X1 U17992 ( .A1(n20120), .A2(n20084), .B1(n20064), .B2(n16637), .C1(
        n22062), .C2(n17309), .ZN(P2_U2913) );
  OAI21_X1 U17993 ( .B1(n14279), .B2(n14278), .A(n14277), .ZN(n17151) );
  INV_X1 U17994 ( .A(n16535), .ZN(n14280) );
  INV_X1 U17995 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20110) );
  OAI222_X1 U17996 ( .A1(n17151), .A2(n16637), .B1(n14280), .B2(n22062), .C1(
        n20110), .C2(n20084), .ZN(P2_U2908) );
  OAI21_X1 U17997 ( .B1(n14283), .B2(n14282), .A(n14281), .ZN(n20963) );
  INV_X1 U17998 ( .A(n14284), .ZN(n14285) );
  AOI21_X1 U17999 ( .B1(n14287), .B2(n14286), .A(n14285), .ZN(n21026) );
  AOI22_X1 U18000 ( .A1(n20974), .A2(n21026), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14943), .ZN(n14288) );
  OAI21_X1 U18001 ( .B1(n20963), .B2(n14927), .A(n14288), .ZN(P1_U2870) );
  OAI222_X1 U18002 ( .A1(n20963), .A2(n15067), .B1(n15066), .B2(n14289), .C1(
        n15064), .C2(n21072), .ZN(P1_U2902) );
  INV_X2 U18003 ( .A(n15173), .ZN(n20992) );
  INV_X1 U18004 ( .A(n14291), .ZN(n14292) );
  XNOR2_X1 U18005 ( .A(n14293), .B(n14292), .ZN(n14294) );
  NAND2_X1 U18006 ( .A1(n14294), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n21044) );
  INV_X1 U18007 ( .A(n14294), .ZN(n14295) );
  NAND2_X1 U18008 ( .A1(n14295), .A2(n21045), .ZN(n21043) );
  NAND3_X1 U18009 ( .A1(n21044), .A2(n21043), .A3(n21001), .ZN(n14297) );
  AOI22_X1 U18010 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n21051), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14296) );
  OAI211_X1 U18011 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n21006), .A(
        n14297), .B(n14296), .ZN(n14298) );
  INV_X1 U18012 ( .A(n14298), .ZN(n14299) );
  OAI21_X1 U18013 ( .B1(n14895), .B2(n15252), .A(n14299), .ZN(P1_U2998) );
  INV_X1 U18014 ( .A(n14277), .ZN(n14302) );
  OAI21_X1 U18015 ( .B1(n14302), .B2(n10821), .A(n14301), .ZN(n17139) );
  AOI22_X1 U18016 ( .A1(n16634), .A2(n16527), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n20093), .ZN(n14303) );
  OAI21_X1 U18017 ( .B1(n17139), .B2(n16637), .A(n14303), .ZN(P2_U2907) );
  NAND2_X1 U18018 ( .A1(n11073), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14304) );
  NAND2_X1 U18019 ( .A1(n16020), .A2(n14304), .ZN(n14310) );
  NAND2_X1 U18020 ( .A1(n14305), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n16019) );
  NOR2_X1 U18021 ( .A1(n14349), .A2(n16133), .ZN(n14306) );
  NAND2_X1 U18022 ( .A1(n14346), .A2(n14306), .ZN(n14361) );
  INV_X1 U18023 ( .A(n14306), .ZN(n14307) );
  NAND2_X1 U18024 ( .A1(n14308), .A2(n14307), .ZN(n14309) );
  OR2_X1 U18025 ( .A1(n14310), .A2(n14309), .ZN(n14311) );
  NAND2_X1 U18026 ( .A1(n14361), .A2(n14311), .ZN(n20088) );
  INV_X1 U18027 ( .A(n14313), .ZN(n14314) );
  NOR2_X1 U18028 ( .A1(n14312), .A2(n14314), .ZN(n14318) );
  OAI21_X1 U18029 ( .B1(n14318), .B2(n14317), .A(n14316), .ZN(n17242) );
  NOR2_X1 U18030 ( .A1(n17242), .A2(n16503), .ZN(n14319) );
  AOI21_X1 U18031 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n16503), .A(n14319), .ZN(
        n14320) );
  OAI21_X1 U18032 ( .B1(n20088), .B2(n20076), .A(n14320), .ZN(P2_U2883) );
  OR2_X1 U18033 ( .A1(n14322), .A2(n14321), .ZN(n14323) );
  NAND2_X1 U18034 ( .A1(n14324), .A2(n14323), .ZN(n16630) );
  INV_X1 U18035 ( .A(n16630), .ZN(n20815) );
  XNOR2_X1 U18036 ( .A(n20817), .B(n16630), .ZN(n14328) );
  NOR2_X1 U18037 ( .A1(n20824), .A2(n20828), .ZN(n14325) );
  AOI21_X1 U18038 ( .B1(n20824), .B2(n20828), .A(n14325), .ZN(n20096) );
  NAND2_X1 U18039 ( .A1(n20096), .A2(n20095), .ZN(n20094) );
  INV_X1 U18040 ( .A(n14325), .ZN(n14326) );
  NAND2_X1 U18041 ( .A1(n20094), .A2(n14326), .ZN(n14327) );
  NAND2_X1 U18042 ( .A1(n14328), .A2(n14327), .ZN(n16629) );
  OAI21_X1 U18043 ( .B1(n14328), .B2(n14327), .A(n16629), .ZN(n14329) );
  NAND2_X1 U18044 ( .A1(n14329), .A2(n22058), .ZN(n14331) );
  AOI22_X1 U18045 ( .A1(n16634), .A2(n16601), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n20093), .ZN(n14330) );
  OAI211_X1 U18046 ( .C1(n20815), .C2(n20085), .A(n14331), .B(n14330), .ZN(
        P2_U2917) );
  OR2_X1 U18047 ( .A1(n14333), .A2(n14332), .ZN(n14334) );
  AND2_X1 U18048 ( .A1(n14335), .A2(n14334), .ZN(n21033) );
  INV_X1 U18049 ( .A(n20966), .ZN(n14337) );
  AOI22_X1 U18050 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21051), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14336) );
  OAI21_X1 U18051 ( .B1(n21006), .B2(n14337), .A(n14336), .ZN(n14338) );
  AOI21_X1 U18052 ( .B1(n21033), .B2(n21001), .A(n14338), .ZN(n14339) );
  OAI21_X1 U18053 ( .B1(n20963), .B2(n15252), .A(n14339), .ZN(P1_U2997) );
  XNOR2_X1 U18054 ( .A(n16493), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U18055 ( .A1(n14341), .A2(n14342), .ZN(n14343) );
  NAND2_X1 U18056 ( .A1(n14340), .A2(n14343), .ZN(n20067) );
  INV_X1 U18057 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n21970) );
  MUX2_X1 U18058 ( .A(n20067), .B(n21970), .S(n16503), .Z(n14344) );
  OAI21_X1 U18059 ( .B1(n14345), .B2(n20076), .A(n14344), .ZN(P2_U2881) );
  INV_X1 U18060 ( .A(n14346), .ZN(n14350) );
  AND4_X1 U18061 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__5__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14347) );
  NAND2_X1 U18062 ( .A1(n16498), .A2(n14347), .ZN(n14348) );
  OR2_X1 U18063 ( .A1(n14349), .A2(n14348), .ZN(n16024) );
  NAND2_X1 U18064 ( .A1(n16495), .A2(n16021), .ZN(n20077) );
  OAI211_X1 U18065 ( .C1(n16495), .C2(n16021), .A(n20077), .B(n16497), .ZN(
        n14356) );
  NAND2_X1 U18066 ( .A1(n14352), .A2(n14353), .ZN(n14354) );
  NAND2_X1 U18067 ( .A1(n17183), .A2(n20082), .ZN(n14355) );
  OAI211_X1 U18068 ( .C1(n20082), .C2(n11772), .A(n14356), .B(n14355), .ZN(
        P2_U2878) );
  AOI21_X1 U18069 ( .B1(n14358), .B2(n14301), .A(n14357), .ZN(n17129) );
  INV_X1 U18070 ( .A(n17129), .ZN(n14360) );
  INV_X1 U18071 ( .A(n16521), .ZN(n14359) );
  INV_X1 U18072 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20106) );
  OAI222_X1 U18073 ( .A1(n14360), .A2(n16637), .B1(n14359), .B2(n22062), .C1(
        n20106), .C2(n20084), .ZN(P2_U2906) );
  AOI211_X1 U18074 ( .C1(n16156), .C2(n14361), .A(n20076), .B(n16493), .ZN(
        n14365) );
  NAND2_X1 U18075 ( .A1(n14316), .A2(n14362), .ZN(n14363) );
  AND2_X1 U18076 ( .A1(n14341), .A2(n14363), .ZN(n17238) );
  MUX2_X1 U18077 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n17238), .S(n20082), .Z(
        n14364) );
  OR2_X1 U18078 ( .A1(n14365), .A2(n14364), .ZN(P2_U2882) );
  INV_X1 U18079 ( .A(n14366), .ZN(n14367) );
  OAI21_X1 U18080 ( .B1(n14357), .B2(n14368), .A(n14367), .ZN(n17111) );
  AOI22_X1 U18081 ( .A1(n16634), .A2(n16507), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n20093), .ZN(n14369) );
  OAI21_X1 U18082 ( .B1(n17111), .B2(n16637), .A(n14369), .ZN(P2_U2905) );
  AOI22_X1 U18083 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14373) );
  AOI22_X1 U18084 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U18085 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14371) );
  AOI22_X1 U18086 ( .A1(n18315), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14370) );
  NAND4_X1 U18087 ( .A1(n14373), .A2(n14372), .A3(n14371), .A4(n14370), .ZN(
        n14379) );
  AOI22_X1 U18088 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18312), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U18089 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U18090 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14375) );
  AOI22_X1 U18091 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14374) );
  NAND4_X1 U18092 ( .A1(n14377), .A2(n14376), .A3(n14375), .A4(n14374), .ZN(
        n14378) );
  NOR2_X1 U18093 ( .A1(n14379), .A2(n14378), .ZN(n18492) );
  INV_X1 U18094 ( .A(n18492), .ZN(n14388) );
  INV_X1 U18095 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n18058) );
  NAND2_X1 U18096 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18376) );
  NOR2_X1 U18097 ( .A1(n18058), .A2(n18376), .ZN(n18367) );
  INV_X1 U18098 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n14384) );
  NAND3_X1 U18099 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n18352) );
  NOR2_X1 U18100 ( .A1(n14384), .A2(n18352), .ZN(n17464) );
  NAND3_X1 U18101 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .ZN(n17466) );
  INV_X1 U18102 ( .A(n18354), .ZN(n18330) );
  AND2_X1 U18103 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .ZN(n14385) );
  AOI21_X1 U18104 ( .B1(n18330), .B2(n14385), .A(P3_EBX_REG_11__SCAN_IN), .ZN(
        n14386) );
  NOR2_X1 U18105 ( .A1(n9936), .A2(n14386), .ZN(n14387) );
  MUX2_X1 U18106 ( .A(n14388), .B(n14387), .S(n18379), .Z(P3_U2692) );
  NAND2_X1 U18107 ( .A1(n14390), .A2(n14389), .ZN(n14394) );
  AOI22_X1 U18108 ( .A1(n14392), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14391), .ZN(n14393) );
  INV_X1 U18109 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14421) );
  OAI22_X1 U18110 ( .A1(n14509), .A2(n14959), .B1(n20978), .B2(n14421), .ZN(
        P1_U2841) );
  NAND2_X1 U18111 ( .A1(n21647), .A2(n21644), .ZN(n17529) );
  NOR2_X1 U18112 ( .A1(n21474), .A2(n17529), .ZN(n17601) );
  NAND2_X1 U18113 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17601), .ZN(n17532) );
  INV_X1 U18114 ( .A(n17532), .ZN(n14400) );
  OAI21_X1 U18115 ( .B1(n17527), .B2(n14398), .A(n17570), .ZN(n14399) );
  OR2_X1 U18116 ( .A1(n14456), .A2(n9763), .ZN(n14419) );
  NAND2_X1 U18117 ( .A1(n21653), .A2(n21880), .ZN(n17520) );
  NAND3_X1 U18118 ( .A1(n9762), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n17520), .ZN(
        n14401) );
  OR2_X2 U18119 ( .A1(n14419), .A2(n14401), .ZN(n20927) );
  INV_X1 U18120 ( .A(n14402), .ZN(n14403) );
  NAND2_X1 U18121 ( .A1(n14403), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14404) );
  INV_X1 U18122 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14420) );
  NAND2_X1 U18123 ( .A1(n14507), .A2(n20914), .ZN(n14428) );
  NAND2_X1 U18124 ( .A1(n14406), .A2(n21880), .ZN(n14417) );
  INV_X1 U18125 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21702) );
  INV_X1 U18126 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21698) );
  INV_X1 U18127 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21694) );
  INV_X1 U18128 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21686) );
  NAND3_X1 U18129 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n14801) );
  NOR2_X1 U18130 ( .A1(n21686), .A2(n14801), .ZN(n14747) );
  AND3_X1 U18131 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14407) );
  AND2_X1 U18132 ( .A1(n14747), .A2(n14407), .ZN(n14722) );
  INV_X1 U18133 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21667) );
  NAND3_X1 U18134 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20939) );
  NOR2_X1 U18135 ( .A1(n21667), .A2(n20939), .ZN(n20940) );
  INV_X1 U18136 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21674) );
  NAND2_X1 U18137 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20905) );
  NOR2_X1 U18138 ( .A1(n21674), .A2(n20905), .ZN(n14887) );
  NAND3_X1 U18139 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20940), .A3(n14887), 
        .ZN(n20889) );
  INV_X1 U18140 ( .A(n20889), .ZN(n14408) );
  NAND4_X1 U18141 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .A4(n14408), .ZN(n14410) );
  NAND2_X1 U18142 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14409) );
  NOR2_X1 U18143 ( .A1(n14410), .A2(n14409), .ZN(n14411) );
  NAND2_X1 U18144 ( .A1(n14722), .A2(n14411), .ZN(n14696) );
  NOR2_X1 U18145 ( .A1(n21694), .A2(n14696), .ZN(n14681) );
  NAND2_X1 U18146 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n14681), .ZN(n14664) );
  NOR2_X1 U18147 ( .A1(n21698), .A2(n14664), .ZN(n14648) );
  NAND2_X1 U18148 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14648), .ZN(n14634) );
  NOR2_X1 U18149 ( .A1(n21702), .A2(n14634), .ZN(n14623) );
  NAND2_X1 U18150 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n14623), .ZN(n14422) );
  INV_X1 U18151 ( .A(n14422), .ZN(n14412) );
  OAI21_X1 U18152 ( .B1(n20938), .B2(n14412), .A(n20904), .ZN(n14622) );
  NAND2_X1 U18153 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14585) );
  INV_X1 U18154 ( .A(n14585), .ZN(n14423) );
  NOR2_X1 U18155 ( .A1(n20938), .A2(n14423), .ZN(n14413) );
  OR2_X1 U18156 ( .A1(n14622), .A2(n14413), .ZN(n14599) );
  INV_X1 U18157 ( .A(n14599), .ZN(n14415) );
  INV_X1 U18158 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21708) );
  OAI21_X1 U18159 ( .B1(n21708), .B2(n21712), .A(n20959), .ZN(n14414) );
  NAND2_X1 U18160 ( .A1(n14415), .A2(n14414), .ZN(n14570) );
  NAND2_X1 U18161 ( .A1(n9762), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14416) );
  NAND2_X1 U18162 ( .A1(n14417), .A2(n14416), .ZN(n14418) );
  OAI22_X1 U18163 ( .A1(n20948), .A2(n14421), .B1(n20901), .B2(n14420), .ZN(
        n14426) );
  NOR2_X1 U18164 ( .A1(n20938), .A2(n14422), .ZN(n14584) );
  AND2_X1 U18165 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n14423), .ZN(n14424) );
  NAND2_X1 U18166 ( .A1(n14584), .A2(n14424), .ZN(n14569) );
  NOR3_X1 U18167 ( .A1(n14569), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21712), 
        .ZN(n14425) );
  AOI211_X1 U18168 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14570), .A(n14426), 
        .B(n14425), .ZN(n14427) );
  OAI211_X1 U18169 ( .C1(n14509), .C2(n20927), .A(n14428), .B(n14427), .ZN(
        P1_U2809) );
  AND2_X1 U18170 ( .A1(n14430), .A2(n14429), .ZN(n14432) );
  AOI21_X1 U18171 ( .B1(n14435), .B2(n14434), .A(n14433), .ZN(n16952) );
  NAND2_X1 U18172 ( .A1(n16952), .A2(n20041), .ZN(n14446) );
  OAI21_X1 U18173 ( .B1(n14437), .B2(n16643), .A(n15999), .ZN(n14438) );
  INV_X1 U18174 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21894) );
  AOI22_X1 U18175 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_29__SCAN_IN), .ZN(n14439) );
  OAI21_X1 U18176 ( .B1(n20073), .B2(n21894), .A(n14439), .ZN(n14440) );
  AOI21_X1 U18177 ( .B1(n14441), .B2(n16003), .A(n14440), .ZN(n14442) );
  INV_X1 U18178 ( .A(n14442), .ZN(n14443) );
  OAI211_X1 U18179 ( .C1(n20065), .C2(n16950), .A(n14446), .B(n14445), .ZN(
        P2_U2826) );
  OAI21_X1 U18180 ( .B1(n14447), .B2(n14449), .A(n14448), .ZN(n15296) );
  AND2_X1 U18181 ( .A1(n14284), .A2(n14451), .ZN(n14452) );
  NOR2_X1 U18182 ( .A1(n14450), .A2(n14452), .ZN(n21020) );
  AOI22_X1 U18183 ( .A1(n20974), .A2(n21020), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14943), .ZN(n14453) );
  OAI21_X1 U18184 ( .B1(n15296), .B2(n14927), .A(n14453), .ZN(P1_U2869) );
  NOR2_X1 U18185 ( .A1(n14456), .A2(n12199), .ZN(n14454) );
  NAND2_X1 U18186 ( .A1(n9763), .A2(n21060), .ZN(n14481) );
  NOR2_X1 U18187 ( .A1(n14456), .A2(n14481), .ZN(n20958) );
  INV_X1 U18188 ( .A(n21020), .ZN(n14464) );
  INV_X1 U18189 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21989) );
  NAND4_X1 U18190 ( .A1(n20959), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .A4(n21989), .ZN(n14459) );
  OAI221_X1 U18191 ( .B1(n20938), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n20938), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n20904), .ZN(n14457) );
  NAND2_X1 U18192 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n14457), .ZN(n14458) );
  OAI211_X1 U18193 ( .C1(n20901), .C2(n14460), .A(n14459), .B(n14458), .ZN(
        n14462) );
  AND3_X2 U18194 ( .A1(n20904), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n14505), 
        .ZN(n20965) );
  NOR2_X1 U18195 ( .A1(n20952), .A2(n15298), .ZN(n14461) );
  AOI211_X1 U18196 ( .C1(P1_EBX_REG_3__SCAN_IN), .C2(n20955), .A(n14462), .B(
        n14461), .ZN(n14463) );
  OAI21_X1 U18197 ( .B1(n20927), .B2(n14464), .A(n14463), .ZN(n14465) );
  AOI21_X1 U18198 ( .B1(n20958), .B2(n21327), .A(n14465), .ZN(n14466) );
  OAI21_X1 U18199 ( .B1(n15296), .B2(n20962), .A(n14466), .ZN(P1_U2837) );
  NOR2_X1 U18200 ( .A1(n16388), .A2(n17306), .ZN(n14472) );
  NAND2_X1 U18201 ( .A1(n16930), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14468) );
  OAI211_X1 U18202 ( .C1(n14470), .C2(n16933), .A(n14469), .B(n14468), .ZN(
        n14471) );
  OAI21_X1 U18203 ( .B1(n16911), .B2(n14473), .A(n10830), .ZN(P2_U2984) );
  INV_X1 U18204 ( .A(n14474), .ZN(n14477) );
  INV_X1 U18205 ( .A(n12531), .ZN(n14490) );
  NAND3_X1 U18206 ( .A1(n17497), .A2(n14490), .A3(n15523), .ZN(n14475) );
  OAI21_X1 U18207 ( .B1(n14477), .B2(n14476), .A(n14475), .ZN(n14478) );
  MUX2_X1 U18208 ( .A(n15524), .B(n14478), .S(n15557), .Z(n14484) );
  OAI211_X1 U18209 ( .C1(n10013), .C2(n14481), .A(n14480), .B(n14479), .ZN(
        n14482) );
  INV_X1 U18210 ( .A(n14482), .ZN(n14483) );
  NAND2_X1 U18211 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15558), .ZN(n17604) );
  INV_X1 U18212 ( .A(n17604), .ZN(n14485) );
  AOI22_X1 U18213 ( .A1(n15552), .A2(n14486), .B1(n14485), .B2(
        P1_FLUSH_REG_SCAN_IN), .ZN(n17591) );
  INV_X1 U18214 ( .A(n17597), .ZN(n14498) );
  AOI21_X1 U18215 ( .B1(n15542), .B2(n17592), .A(n14498), .ZN(n14499) );
  INV_X1 U18216 ( .A(n13156), .ZN(n15561) );
  INV_X1 U18217 ( .A(n14487), .ZN(n14489) );
  NAND3_X1 U18218 ( .A1(n14490), .A2(n14489), .A3(n14488), .ZN(n14491) );
  NOR2_X1 U18219 ( .A1(n14492), .A2(n14491), .ZN(n14494) );
  INV_X1 U18220 ( .A(n17593), .ZN(n14493) );
  NAND2_X1 U18221 ( .A1(n14494), .A2(n14493), .ZN(n15585) );
  INV_X1 U18222 ( .A(n15585), .ZN(n14495) );
  OAI22_X1 U18223 ( .A1(n15561), .A2(n14495), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15582), .ZN(n17495) );
  NAND2_X1 U18224 ( .A1(n15557), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15599) );
  OAI22_X1 U18225 ( .A1(n15599), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21644), .ZN(n14496) );
  AOI21_X1 U18226 ( .B1(n17592), .B2(n17495), .A(n14496), .ZN(n14497) );
  OAI22_X1 U18227 ( .A1(n14499), .A2(n17498), .B1(n14498), .B2(n14497), .ZN(
        P1_U3474) );
  INV_X1 U18228 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21710) );
  NOR2_X1 U18229 ( .A1(n17570), .A2(n21710), .ZN(n14512) );
  AOI21_X1 U18230 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14512), .ZN(n14504) );
  OAI21_X1 U18231 ( .B1(n21006), .B2(n14505), .A(n14504), .ZN(n14506) );
  AOI21_X1 U18232 ( .B1(n14507), .B2(n21000), .A(n14506), .ZN(n14508) );
  OAI21_X1 U18233 ( .B1(n14519), .B2(n20873), .A(n14508), .ZN(P1_U2968) );
  INV_X1 U18234 ( .A(n14509), .ZN(n14517) );
  INV_X1 U18235 ( .A(n14512), .ZN(n14515) );
  NAND3_X1 U18236 ( .A1(n10796), .A2(n14515), .A3(n10810), .ZN(n14516) );
  AOI21_X1 U18237 ( .B1(n14517), .B2(n21027), .A(n14516), .ZN(n14518) );
  OAI21_X1 U18238 ( .B1(n14519), .B2(n21012), .A(n14518), .ZN(P1_U3000) );
  XOR2_X1 U18239 ( .A(n14521), .B(n14520), .Z(n14539) );
  NAND2_X1 U18240 ( .A1(n14523), .A2(n14522), .ZN(n14528) );
  OAI22_X1 U18241 ( .A1(n17082), .A2(n14528), .B1(n14525), .B2(n14524), .ZN(
        n14532) );
  XNOR2_X1 U18242 ( .A(n14527), .B(n14526), .ZN(n14534) );
  NOR2_X1 U18243 ( .A1(n20051), .A2(n20734), .ZN(n14535) );
  AOI21_X1 U18244 ( .B1(n17080), .B2(n14528), .A(n14535), .ZN(n14530) );
  NAND2_X1 U18245 ( .A1(n12994), .A2(n16630), .ZN(n14529) );
  OAI211_X1 U18246 ( .C1(n17266), .C2(n14534), .A(n14530), .B(n14529), .ZN(
        n14531) );
  AOI211_X1 U18247 ( .C1(n17262), .C2(n14539), .A(n14532), .B(n14531), .ZN(
        n14533) );
  OAI21_X1 U18248 ( .B1(n17320), .B2(n17241), .A(n14533), .ZN(P2_U3044) );
  NOR2_X1 U18249 ( .A1(n14534), .A2(n16942), .ZN(n14538) );
  AOI21_X1 U18250 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14535), .ZN(n14536) );
  OAI21_X1 U18251 ( .B1(n16933), .B2(n15976), .A(n14536), .ZN(n14537) );
  AOI211_X1 U18252 ( .C1(n14539), .C2(n16939), .A(n14538), .B(n14537), .ZN(
        n14540) );
  OAI21_X1 U18253 ( .B1(n17320), .B2(n17306), .A(n14540), .ZN(P2_U3012) );
  MUX2_X1 U18254 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n16002), .S(
        n20059), .Z(n17282) );
  NAND2_X1 U18255 ( .A1(n17282), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20795) );
  AND2_X1 U18256 ( .A1(n14541), .A2(n16002), .ZN(n14542) );
  NOR2_X1 U18257 ( .A1(n15973), .A2(n14542), .ZN(n14543) );
  NAND2_X1 U18258 ( .A1(n20059), .A2(n14543), .ZN(n15989) );
  OAI21_X1 U18259 ( .B1(n20059), .B2(n21897), .A(n15989), .ZN(n20793) );
  NOR2_X1 U18260 ( .A1(n20795), .A2(n20793), .ZN(n14549) );
  AND2_X1 U18261 ( .A1(n10510), .A2(n14544), .ZN(n17277) );
  NOR3_X1 U18262 ( .A1(n17277), .A2(n11169), .A3(n14545), .ZN(n14547) );
  INV_X1 U18263 ( .A(n17280), .ZN(n17319) );
  NOR2_X1 U18264 ( .A1(n15994), .A2(n17319), .ZN(n14546) );
  AOI211_X1 U18265 ( .C1(n21769), .C2(n17327), .A(n14547), .B(n14546), .ZN(
        n17315) );
  OR2_X1 U18266 ( .A1(n17345), .A2(n20814), .ZN(n20797) );
  OAI22_X1 U18267 ( .A1(n17315), .A2(n20803), .B1(n20134), .B2(n20797), .ZN(
        n14548) );
  OAI21_X1 U18268 ( .B1(n14549), .B2(n14548), .A(n17298), .ZN(n14550) );
  OAI21_X1 U18269 ( .B1(n17298), .B2(n21769), .A(n14550), .ZN(P2_U3600) );
  AOI22_X1 U18270 ( .A1(n16616), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n20093), .ZN(n14554) );
  NAND2_X1 U18271 ( .A1(n16615), .A2(BUF1_REG_31__SCAN_IN), .ZN(n14553) );
  OAI211_X1 U18272 ( .C1(n14551), .C2(n20085), .A(n14554), .B(n14553), .ZN(
        P2_U2888) );
  INV_X1 U18273 ( .A(n16017), .ZN(n14555) );
  NAND2_X1 U18274 ( .A1(n14555), .A2(n20041), .ZN(n14563) );
  NAND2_X1 U18275 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14558) );
  NAND3_X1 U18276 ( .A1(n14556), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n17367), 
        .ZN(n14557) );
  OAI211_X1 U18277 ( .C1(n16009), .C2(n20781), .A(n14558), .B(n14557), .ZN(
        n14561) );
  OR2_X1 U18278 ( .A1(n14719), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14565) );
  NAND2_X1 U18279 ( .A1(n12561), .A2(n12199), .ZN(n14564) );
  MUX2_X1 U18280 ( .A(n14565), .B(n14564), .S(n21735), .Z(P1_U3487) );
  AOI21_X2 U18281 ( .B1(n14568), .B2(n14566), .A(n14567), .ZN(n15073) );
  INV_X1 U18282 ( .A(n15073), .ZN(n14906) );
  INV_X1 U18283 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14905) );
  INV_X1 U18284 ( .A(n14569), .ZN(n14571) );
  OAI21_X1 U18285 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14571), .A(n14570), 
        .ZN(n14573) );
  AOI22_X1 U18286 ( .A1(n20965), .A2(n15068), .B1(n20956), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14572) );
  OAI211_X1 U18287 ( .C1(n20948), .C2(n14905), .A(n14573), .B(n14572), .ZN(
        n14574) );
  OAI21_X1 U18288 ( .B1(n14906), .B2(n20907), .A(n14576), .ZN(P1_U2810) );
  OR2_X1 U18289 ( .A1(n14578), .A2(n14577), .ZN(n14579) );
  NAND2_X1 U18290 ( .A1(n14580), .A2(n14579), .ZN(n15303) );
  OAI21_X1 U18291 ( .B1(n14581), .B2(n14582), .A(n14566), .ZN(n14908) );
  INV_X1 U18292 ( .A(n14908), .ZN(n15079) );
  NAND2_X1 U18293 ( .A1(n15079), .A2(n20914), .ZN(n14590) );
  INV_X1 U18294 ( .A(n14583), .ZN(n15077) );
  OAI22_X1 U18295 ( .A1(n20952), .A2(n15077), .B1(n20901), .B2(n21867), .ZN(
        n14588) );
  INV_X1 U18296 ( .A(n14584), .ZN(n14612) );
  NOR2_X1 U18297 ( .A1(n14612), .A2(n14585), .ZN(n14586) );
  MUX2_X1 U18298 ( .A(n14586), .B(n14599), .S(P1_REIP_REG_29__SCAN_IN), .Z(
        n14587) );
  AOI211_X1 U18299 ( .C1(P1_EBX_REG_29__SCAN_IN), .C2(n20955), .A(n14588), .B(
        n14587), .ZN(n14589) );
  OAI211_X1 U18300 ( .C1(n20927), .C2(n15303), .A(n14590), .B(n14589), .ZN(
        P1_U2811) );
  INV_X1 U18301 ( .A(n14591), .ZN(n14613) );
  NOR2_X1 U18302 ( .A1(n14620), .A2(n14613), .ZN(n14593) );
  OAI21_X1 U18303 ( .B1(n14594), .B2(n14593), .A(n14592), .ZN(n15319) );
  NAND2_X1 U18304 ( .A1(n15093), .A2(n20914), .ZN(n14603) );
  OAI22_X1 U18305 ( .A1(n20952), .A2(n15091), .B1(n20901), .B2(n14597), .ZN(
        n14601) );
  INV_X1 U18306 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n22020) );
  NOR2_X1 U18307 ( .A1(n14612), .A2(n22020), .ZN(n14598) );
  INV_X1 U18308 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15089) );
  MUX2_X1 U18309 ( .A(n14599), .B(n14598), .S(n15089), .Z(n14600) );
  AOI211_X1 U18310 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n20955), .A(n14601), .B(
        n14600), .ZN(n14602) );
  OAI211_X1 U18311 ( .C1(n15319), .C2(n20927), .A(n14603), .B(n14602), .ZN(
        P1_U2812) );
  INV_X1 U18312 ( .A(n14604), .ZN(n14607) );
  OAI21_X2 U18313 ( .B1(n14607), .B2(n10773), .A(n14606), .ZN(n14978) );
  INV_X1 U18314 ( .A(n14608), .ZN(n15101) );
  OAI22_X1 U18315 ( .A1(n20952), .A2(n15101), .B1(n20901), .B2(n14609), .ZN(
        n14610) );
  AOI21_X1 U18316 ( .B1(n20955), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14610), .ZN(
        n14611) );
  OAI21_X1 U18317 ( .B1(n14612), .B2(P1_REIP_REG_27__SCAN_IN), .A(n14611), 
        .ZN(n14615) );
  XNOR2_X1 U18318 ( .A(n14620), .B(n14613), .ZN(n15328) );
  NOR2_X1 U18319 ( .A1(n15328), .A2(n20927), .ZN(n14614) );
  AOI211_X1 U18320 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14622), .A(n14615), 
        .B(n14614), .ZN(n14616) );
  OAI21_X1 U18321 ( .B1(n14978), .B2(n20907), .A(n14616), .ZN(P1_U2813) );
  NAND2_X1 U18322 ( .A1(n14617), .A2(n14618), .ZN(n14619) );
  NAND2_X1 U18323 ( .A1(n14620), .A2(n14619), .ZN(n15333) );
  OAI21_X1 U18324 ( .B1(n9834), .B2(n9871), .A(n14604), .ZN(n14911) );
  INV_X1 U18325 ( .A(n14911), .ZN(n15112) );
  NAND2_X1 U18326 ( .A1(n15112), .A2(n20914), .ZN(n14629) );
  OAI22_X1 U18327 ( .A1(n20952), .A2(n15110), .B1(n20901), .B2(n14621), .ZN(
        n14627) );
  INV_X1 U18328 ( .A(n14622), .ZN(n14625) );
  AOI21_X1 U18329 ( .B1(n20959), .B2(n14623), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14624) );
  NOR2_X1 U18330 ( .A1(n14625), .A2(n14624), .ZN(n14626) );
  AOI211_X1 U18331 ( .C1(n20955), .C2(P1_EBX_REG_26__SCAN_IN), .A(n14627), .B(
        n14626), .ZN(n14628) );
  OAI211_X1 U18332 ( .C1(n15333), .C2(n20927), .A(n14629), .B(n14628), .ZN(
        P1_U2814) );
  INV_X1 U18333 ( .A(n14630), .ZN(n14633) );
  INV_X1 U18334 ( .A(n14631), .ZN(n14632) );
  AOI21_X1 U18335 ( .B1(n14633), .B2(n14632), .A(n9834), .ZN(n15123) );
  INV_X1 U18336 ( .A(n15123), .ZN(n14913) );
  OAI21_X1 U18337 ( .B1(n20938), .B2(n14648), .A(n20904), .ZN(n14665) );
  INV_X1 U18338 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14912) );
  INV_X1 U18339 ( .A(n14634), .ZN(n14636) );
  NAND2_X1 U18340 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14635) );
  OAI211_X1 U18341 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14636), .A(n20959), 
        .B(n14635), .ZN(n14639) );
  INV_X1 U18342 ( .A(n15121), .ZN(n14637) );
  AOI22_X1 U18343 ( .A1(n20965), .A2(n14637), .B1(n20956), .B2(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14638) );
  OAI211_X1 U18344 ( .C1(n14912), .C2(n20948), .A(n14639), .B(n14638), .ZN(
        n14644) );
  OR2_X1 U18345 ( .A1(n14640), .A2(n14641), .ZN(n14642) );
  NAND2_X1 U18346 ( .A1(n14617), .A2(n14642), .ZN(n15348) );
  NOR2_X1 U18347 ( .A1(n15348), .A2(n20927), .ZN(n14643) );
  AOI211_X1 U18348 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14665), .A(n14644), 
        .B(n14643), .ZN(n14645) );
  OAI21_X1 U18349 ( .B1(n14913), .B2(n20907), .A(n14645), .ZN(P1_U2815) );
  INV_X1 U18350 ( .A(n14646), .ZN(n14647) );
  AOI21_X1 U18351 ( .B1(n14647), .B2(n9831), .A(n14631), .ZN(n15133) );
  INV_X1 U18352 ( .A(n15133), .ZN(n14998) );
  INV_X1 U18353 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14652) );
  INV_X1 U18354 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21700) );
  NAND3_X1 U18355 ( .A1(n20959), .A2(n14648), .A3(n21700), .ZN(n14651) );
  INV_X1 U18356 ( .A(n15131), .ZN(n14649) );
  AOI22_X1 U18357 ( .A1(n20965), .A2(n14649), .B1(n20956), .B2(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14650) );
  OAI211_X1 U18358 ( .C1(n14652), .C2(n20948), .A(n14651), .B(n14650), .ZN(
        n14653) );
  AOI21_X1 U18359 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n14665), .A(n14653), 
        .ZN(n14658) );
  INV_X1 U18360 ( .A(n14654), .ZN(n14656) );
  INV_X1 U18361 ( .A(n14663), .ZN(n14655) );
  AOI21_X1 U18362 ( .B1(n14656), .B2(n14655), .A(n14640), .ZN(n15359) );
  NAND2_X1 U18363 ( .A1(n15359), .A2(n20954), .ZN(n14657) );
  OAI211_X1 U18364 ( .C1(n14998), .C2(n20907), .A(n14658), .B(n14657), .ZN(
        P1_U2816) );
  OAI21_X1 U18365 ( .B1(n14659), .B2(n14660), .A(n9831), .ZN(n14999) );
  AND2_X1 U18366 ( .A1(n14675), .A2(n14661), .ZN(n14662) );
  NOR2_X1 U18367 ( .A1(n14663), .A2(n14662), .ZN(n15369) );
  NOR2_X1 U18368 ( .A1(n20938), .A2(n14664), .ZN(n14666) );
  OAI21_X1 U18369 ( .B1(n14666), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14665), 
        .ZN(n14669) );
  INV_X1 U18370 ( .A(n15138), .ZN(n14667) );
  AOI22_X1 U18371 ( .A1(n20965), .A2(n14667), .B1(n20956), .B2(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14668) );
  OAI211_X1 U18372 ( .C1(n14670), .C2(n20948), .A(n14669), .B(n14668), .ZN(
        n14671) );
  AOI21_X1 U18373 ( .B1(n15369), .B2(n20954), .A(n14671), .ZN(n14672) );
  OAI21_X1 U18374 ( .B1(n14999), .B2(n20907), .A(n14672), .ZN(P1_U2817) );
  AOI21_X1 U18375 ( .B1(n14673), .B2(n14689), .A(n14659), .ZN(n15149) );
  INV_X1 U18376 ( .A(n15149), .ZN(n14917) );
  INV_X1 U18377 ( .A(n14675), .ZN(n14676) );
  AOI21_X1 U18378 ( .B1(n14677), .B2(n14674), .A(n14676), .ZN(n15382) );
  NAND2_X1 U18379 ( .A1(n20938), .A2(n20904), .ZN(n14901) );
  INV_X1 U18380 ( .A(n14696), .ZN(n14678) );
  NAND2_X1 U18381 ( .A1(n20904), .A2(n14678), .ZN(n14679) );
  NAND2_X1 U18382 ( .A1(n14901), .A2(n14679), .ZN(n14710) );
  INV_X1 U18383 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21696) );
  NOR2_X1 U18384 ( .A1(n14710), .A2(n21696), .ZN(n14686) );
  INV_X1 U18385 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14684) );
  NAND2_X1 U18386 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14680) );
  OAI211_X1 U18387 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14681), .A(n20959), 
        .B(n14680), .ZN(n14683) );
  AOI22_X1 U18388 ( .A1(n20965), .A2(n15145), .B1(n20956), .B2(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14682) );
  OAI211_X1 U18389 ( .C1(n14684), .C2(n20948), .A(n14683), .B(n14682), .ZN(
        n14685) );
  AOI211_X1 U18390 ( .C1(n15382), .C2(n20954), .A(n14686), .B(n14685), .ZN(
        n14687) );
  OAI21_X1 U18391 ( .B1(n14917), .B2(n20907), .A(n14687), .ZN(P1_U2818) );
  INV_X1 U18392 ( .A(n14689), .ZN(n14690) );
  AOI21_X1 U18393 ( .B1(n14691), .B2(n14688), .A(n14690), .ZN(n15157) );
  INV_X1 U18394 ( .A(n15157), .ZN(n14920) );
  OAI21_X1 U18395 ( .B1(n14692), .B2(n14693), .A(n14674), .ZN(n14918) );
  INV_X1 U18396 ( .A(n14918), .ZN(n15389) );
  INV_X1 U18397 ( .A(n14694), .ZN(n15155) );
  OAI22_X1 U18398 ( .A1(n20952), .A2(n15155), .B1(n20901), .B2(n14695), .ZN(
        n14698) );
  NOR3_X1 U18399 ( .A1(n20938), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14696), 
        .ZN(n14697) );
  AOI211_X1 U18400 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n20955), .A(n14698), .B(
        n14697), .ZN(n14699) );
  OAI21_X1 U18401 ( .B1(n21694), .B2(n14710), .A(n14699), .ZN(n14700) );
  AOI21_X1 U18402 ( .B1(n15389), .B2(n20954), .A(n14700), .ZN(n14701) );
  OAI21_X1 U18403 ( .B1(n14920), .B2(n20907), .A(n14701), .ZN(P1_U2819) );
  INV_X1 U18404 ( .A(n14717), .ZN(n14704) );
  INV_X1 U18405 ( .A(n14702), .ZN(n14703) );
  AOI21_X1 U18406 ( .B1(n14740), .B2(n14704), .A(n14703), .ZN(n14705) );
  OR2_X1 U18407 ( .A1(n14692), .A2(n14705), .ZN(n15393) );
  AOI21_X1 U18408 ( .B1(n14707), .B2(n14706), .A(n13493), .ZN(n15168) );
  NAND2_X1 U18409 ( .A1(n15168), .A2(n20914), .ZN(n14715) );
  OAI22_X1 U18410 ( .A1(n20952), .A2(n15166), .B1(n20901), .B2(n14708), .ZN(
        n14713) );
  NAND2_X1 U18411 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14709) );
  NOR2_X1 U18412 ( .A1(n20889), .A2(n14709), .ZN(n14724) );
  NAND2_X1 U18413 ( .A1(n20959), .A2(n14724), .ZN(n14855) );
  INV_X1 U18414 ( .A(n14722), .ZN(n14726) );
  INV_X1 U18415 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21690) );
  NOR3_X1 U18416 ( .A1(n14855), .A2(n14726), .A3(n21690), .ZN(n14718) );
  AOI21_X1 U18417 ( .B1(n14718), .B2(P1_REIP_REG_19__SCAN_IN), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n14711) );
  NOR2_X1 U18418 ( .A1(n14711), .A2(n14710), .ZN(n14712) );
  AOI211_X1 U18419 ( .C1(P1_EBX_REG_20__SCAN_IN), .C2(n20955), .A(n14713), .B(
        n14712), .ZN(n14714) );
  OAI211_X1 U18420 ( .C1(n15393), .C2(n20927), .A(n14715), .B(n14714), .ZN(
        P1_U2820) );
  OAI21_X1 U18421 ( .B1(n9786), .B2(n14716), .A(n14706), .ZN(n15174) );
  XNOR2_X1 U18422 ( .A(n14740), .B(n14717), .ZN(n15412) );
  INV_X1 U18423 ( .A(n14718), .ZN(n14730) );
  NAND2_X1 U18424 ( .A1(n20904), .A2(n14719), .ZN(n20925) );
  NAND2_X1 U18425 ( .A1(n20965), .A2(n15177), .ZN(n14720) );
  OAI211_X1 U18426 ( .C1(n20901), .C2(n15172), .A(n20925), .B(n14720), .ZN(
        n14721) );
  AOI21_X1 U18427 ( .B1(n20955), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14721), .ZN(
        n14729) );
  NAND2_X1 U18428 ( .A1(n14722), .A2(n21690), .ZN(n14723) );
  NOR2_X1 U18429 ( .A1(n14855), .A2(n14723), .ZN(n14738) );
  NAND2_X1 U18430 ( .A1(n20904), .A2(n14724), .ZN(n14725) );
  NAND2_X1 U18431 ( .A1(n14901), .A2(n14725), .ZN(n14850) );
  NAND2_X1 U18432 ( .A1(n14901), .A2(n14726), .ZN(n14727) );
  NAND2_X1 U18433 ( .A1(n14850), .A2(n14727), .ZN(n14755) );
  OAI21_X1 U18434 ( .B1(n14738), .B2(n14755), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14728) );
  OAI211_X1 U18435 ( .C1(n14730), .C2(P1_REIP_REG_19__SCAN_IN), .A(n14729), 
        .B(n14728), .ZN(n14731) );
  AOI21_X1 U18436 ( .B1(n15412), .B2(n20954), .A(n14731), .ZN(n14732) );
  OAI21_X1 U18437 ( .B1(n15174), .B2(n20907), .A(n14732), .ZN(P1_U2821) );
  INV_X1 U18438 ( .A(n14733), .ZN(n14735) );
  AOI21_X1 U18439 ( .B1(n14735), .B2(n10766), .A(n9786), .ZN(n15186) );
  INV_X1 U18440 ( .A(n15186), .ZN(n14925) );
  NAND2_X1 U18441 ( .A1(n20955), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14737) );
  AOI21_X1 U18442 ( .B1(n20956), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20945), .ZN(n14736) );
  OAI211_X1 U18443 ( .C1(n20952), .C2(n15181), .A(n14737), .B(n14736), .ZN(
        n14739) );
  AOI211_X1 U18444 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n14755), .A(n14739), 
        .B(n14738), .ZN(n14743) );
  AOI21_X1 U18445 ( .B1(n14741), .B2(n14759), .A(n14740), .ZN(n15415) );
  NAND2_X1 U18446 ( .A1(n15415), .A2(n20954), .ZN(n14742) );
  OAI211_X1 U18447 ( .C1(n14925), .C2(n20907), .A(n14743), .B(n14742), .ZN(
        P1_U2822) );
  AND2_X1 U18448 ( .A1(n14744), .A2(n14745), .ZN(n14746) );
  OR2_X1 U18449 ( .A1(n14746), .A2(n14734), .ZN(n15025) );
  INV_X1 U18450 ( .A(n14747), .ZN(n14774) );
  OR2_X1 U18451 ( .A1(n14855), .A2(n14774), .ZN(n14773) );
  NAND2_X1 U18452 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14748) );
  INV_X1 U18453 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21799) );
  OAI21_X1 U18454 ( .B1(n14773), .B2(n14748), .A(n21799), .ZN(n14756) );
  NAND2_X1 U18455 ( .A1(n20956), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14749) );
  AND2_X1 U18456 ( .A1(n14749), .A2(n20925), .ZN(n14752) );
  INV_X1 U18457 ( .A(n15198), .ZN(n14750) );
  NAND2_X1 U18458 ( .A1(n20965), .A2(n14750), .ZN(n14751) );
  OAI211_X1 U18459 ( .C1(n20948), .C2(n14753), .A(n14752), .B(n14751), .ZN(
        n14754) );
  AOI21_X1 U18460 ( .B1(n14756), .B2(n14755), .A(n14754), .ZN(n14761) );
  NAND2_X1 U18461 ( .A1(n14769), .A2(n14757), .ZN(n14758) );
  AND2_X1 U18462 ( .A1(n14759), .A2(n14758), .ZN(n15433) );
  NAND2_X1 U18463 ( .A1(n15433), .A2(n20954), .ZN(n14760) );
  OAI211_X1 U18464 ( .C1(n15025), .C2(n20907), .A(n14761), .B(n14760), .ZN(
        P1_U2823) );
  NAND2_X1 U18465 ( .A1(n14763), .A2(n14764), .ZN(n14782) );
  INV_X1 U18466 ( .A(n14782), .ZN(n14766) );
  OAI21_X1 U18467 ( .B1(n14766), .B2(n14765), .A(n14744), .ZN(n15212) );
  NAND2_X1 U18468 ( .A1(n14787), .A2(n14767), .ZN(n14768) );
  NAND2_X1 U18469 ( .A1(n14769), .A2(n14768), .ZN(n15442) );
  AOI21_X1 U18470 ( .B1(n20956), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20945), .ZN(n14770) );
  OAI21_X1 U18471 ( .B1(n15208), .B2(n20952), .A(n14770), .ZN(n14772) );
  INV_X1 U18472 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21993) );
  NOR3_X1 U18473 ( .A1(n14773), .A2(P1_REIP_REG_16__SCAN_IN), .A3(n21993), 
        .ZN(n14771) );
  AOI211_X1 U18474 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n20955), .A(n14772), .B(
        n14771), .ZN(n14777) );
  NOR2_X1 U18475 ( .A1(n14773), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14791) );
  NAND2_X1 U18476 ( .A1(n14901), .A2(n14774), .ZN(n14775) );
  NAND2_X1 U18477 ( .A1(n14850), .A2(n14775), .ZN(n14807) );
  OAI21_X1 U18478 ( .B1(n14791), .B2(n14807), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14776) );
  OAI211_X1 U18479 ( .C1(n15442), .C2(n20927), .A(n14777), .B(n14776), .ZN(
        n14778) );
  INV_X1 U18480 ( .A(n14778), .ZN(n14779) );
  OAI21_X1 U18481 ( .B1(n15212), .B2(n20907), .A(n14779), .ZN(P1_U2824) );
  NAND2_X1 U18482 ( .A1(n14763), .A2(n14811), .ZN(n14813) );
  NAND2_X1 U18483 ( .A1(n14763), .A2(n14848), .ZN(n14781) );
  AOI21_X1 U18484 ( .B1(n14813), .B2(n14781), .A(n14780), .ZN(n14816) );
  AND2_X1 U18485 ( .A1(n14816), .A2(n14797), .ZN(n14798) );
  OAI22_X1 U18486 ( .A1(n14784), .A2(n20901), .B1(n14928), .B2(n20948), .ZN(
        n14789) );
  OR2_X1 U18487 ( .A1(n14795), .A2(n14785), .ZN(n14786) );
  NAND2_X1 U18488 ( .A1(n14787), .A2(n14786), .ZN(n15450) );
  NOR2_X1 U18489 ( .A1(n20927), .A2(n15450), .ZN(n14788) );
  NOR3_X1 U18490 ( .A1(n20945), .A2(n14789), .A3(n14788), .ZN(n14790) );
  OAI21_X1 U18491 ( .B1(n15219), .B2(n20952), .A(n14790), .ZN(n14792) );
  AOI211_X1 U18492 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n14807), .A(n14792), 
        .B(n14791), .ZN(n14793) );
  OAI21_X1 U18493 ( .B1(n15223), .B2(n20907), .A(n14793), .ZN(P1_U2825) );
  AND2_X1 U18494 ( .A1(n14820), .A2(n14794), .ZN(n14796) );
  OR2_X1 U18495 ( .A1(n14796), .A2(n14795), .ZN(n15451) );
  INV_X1 U18496 ( .A(n14797), .ZN(n14800) );
  INV_X1 U18497 ( .A(n14816), .ZN(n14799) );
  AOI21_X1 U18498 ( .B1(n14800), .B2(n14799), .A(n14798), .ZN(n15234) );
  NAND2_X1 U18499 ( .A1(n15234), .A2(n20914), .ZN(n14810) );
  OAI21_X1 U18500 ( .B1(n14855), .B2(n14801), .A(n21686), .ZN(n14808) );
  INV_X1 U18501 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14931) );
  NAND2_X1 U18502 ( .A1(n20956), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14802) );
  AND2_X1 U18503 ( .A1(n14802), .A2(n20925), .ZN(n14805) );
  INV_X1 U18504 ( .A(n15232), .ZN(n14803) );
  NAND2_X1 U18505 ( .A1(n20965), .A2(n14803), .ZN(n14804) );
  OAI211_X1 U18506 ( .C1(n20948), .C2(n14931), .A(n14805), .B(n14804), .ZN(
        n14806) );
  AOI21_X1 U18507 ( .B1(n14808), .B2(n14807), .A(n14806), .ZN(n14809) );
  OAI211_X1 U18508 ( .C1(n15451), .C2(n20927), .A(n14810), .B(n14809), .ZN(
        P1_U2826) );
  OR2_X1 U18509 ( .A1(n14763), .A2(n14811), .ZN(n14812) );
  NAND2_X1 U18510 ( .A1(n14813), .A2(n14812), .ZN(n14849) );
  INV_X1 U18511 ( .A(n14848), .ZN(n14814) );
  OAI21_X1 U18512 ( .B1(n14849), .B2(n14814), .A(n14813), .ZN(n14836) );
  NAND2_X1 U18513 ( .A1(n14836), .A2(n14835), .ZN(n14834) );
  INV_X1 U18514 ( .A(n14815), .ZN(n14817) );
  AOI21_X1 U18515 ( .B1(n14834), .B2(n14817), .A(n14816), .ZN(n15241) );
  NAND2_X1 U18516 ( .A1(n14841), .A2(n14818), .ZN(n14819) );
  NAND2_X1 U18517 ( .A1(n14820), .A2(n14819), .ZN(n15468) );
  NOR2_X1 U18518 ( .A1(n15468), .A2(n20927), .ZN(n14832) );
  NAND2_X1 U18519 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n14822) );
  INV_X1 U18520 ( .A(n14822), .ZN(n14821) );
  INV_X1 U18521 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21685) );
  NAND2_X1 U18522 ( .A1(n14821), .A2(n21685), .ZN(n14830) );
  NAND2_X1 U18523 ( .A1(n14901), .A2(n14822), .ZN(n14823) );
  NAND2_X1 U18524 ( .A1(n14850), .A2(n14823), .ZN(n14844) );
  NAND2_X1 U18525 ( .A1(n14844), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n14829) );
  INV_X1 U18526 ( .A(n15239), .ZN(n14824) );
  NAND2_X1 U18527 ( .A1(n20965), .A2(n14824), .ZN(n14826) );
  NAND2_X1 U18528 ( .A1(n20956), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14825) );
  NAND3_X1 U18529 ( .A1(n14826), .A2(n20925), .A3(n14825), .ZN(n14827) );
  AOI21_X1 U18530 ( .B1(n20955), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14827), .ZN(
        n14828) );
  OAI211_X1 U18531 ( .C1(n14855), .C2(n14830), .A(n14829), .B(n14828), .ZN(
        n14831) );
  AOI211_X1 U18532 ( .C1(n15241), .C2(n20914), .A(n14832), .B(n14831), .ZN(
        n14833) );
  INV_X1 U18533 ( .A(n14833), .ZN(P1_U2827) );
  OAI21_X1 U18534 ( .B1(n14836), .B2(n14835), .A(n14834), .ZN(n15251) );
  AOI21_X1 U18535 ( .B1(n20956), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20945), .ZN(n14837) );
  OAI21_X1 U18536 ( .B1(n15246), .B2(n20952), .A(n14837), .ZN(n14843) );
  OR2_X1 U18537 ( .A1(n14838), .A2(n14839), .ZN(n14840) );
  NAND2_X1 U18538 ( .A1(n14841), .A2(n14840), .ZN(n15482) );
  NOR2_X1 U18539 ( .A1(n15482), .A2(n20927), .ZN(n14842) );
  AOI211_X1 U18540 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n20955), .A(n14843), .B(
        n14842), .ZN(n14847) );
  INV_X1 U18541 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21682) );
  NOR2_X1 U18542 ( .A1(n14855), .A2(n21682), .ZN(n14845) );
  OAI21_X1 U18543 ( .B1(n14845), .B2(P1_REIP_REG_12__SCAN_IN), .A(n14844), 
        .ZN(n14846) );
  OAI211_X1 U18544 ( .C1(n15251), .C2(n20907), .A(n14847), .B(n14846), .ZN(
        P1_U2828) );
  XNOR2_X1 U18545 ( .A(n14849), .B(n14848), .ZN(n15263) );
  INV_X1 U18546 ( .A(n15263), .ZN(n15050) );
  INV_X1 U18547 ( .A(n14850), .ZN(n14875) );
  NOR2_X1 U18548 ( .A1(n14851), .A2(n14852), .ZN(n14853) );
  OR2_X1 U18549 ( .A1(n14838), .A2(n14853), .ZN(n15488) );
  AOI21_X1 U18550 ( .B1(n20956), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20945), .ZN(n14854) );
  OAI21_X1 U18551 ( .B1(n15261), .B2(n20952), .A(n14854), .ZN(n14857) );
  NOR2_X1 U18552 ( .A1(n14855), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n14856) );
  AOI211_X1 U18553 ( .C1(n20955), .C2(P1_EBX_REG_11__SCAN_IN), .A(n14857), .B(
        n14856), .ZN(n14858) );
  OAI21_X1 U18554 ( .B1(n20927), .B2(n15488), .A(n14858), .ZN(n14859) );
  AOI21_X1 U18555 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n14875), .A(n14859), 
        .ZN(n14860) );
  OAI21_X1 U18556 ( .B1(n15050), .B2(n20907), .A(n14860), .ZN(P1_U2829) );
  NAND2_X1 U18557 ( .A1(n14861), .A2(n14862), .ZN(n14946) );
  INV_X1 U18558 ( .A(n14863), .ZN(n14945) );
  INV_X1 U18559 ( .A(n14864), .ZN(n14877) );
  NAND2_X1 U18560 ( .A1(n14939), .A2(n14938), .ZN(n14937) );
  INV_X1 U18561 ( .A(n14865), .ZN(n14866) );
  AOI21_X1 U18562 ( .B1(n14937), .B2(n14866), .A(n14763), .ZN(n15276) );
  INV_X1 U18563 ( .A(n15276), .ZN(n15052) );
  INV_X1 U18564 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21678) );
  NOR2_X1 U18565 ( .A1(n20889), .A2(n21678), .ZN(n14867) );
  INV_X1 U18566 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21680) );
  NAND3_X1 U18567 ( .A1(n20959), .A2(n14867), .A3(n21680), .ZN(n14868) );
  OAI21_X1 U18568 ( .B1(n20952), .B2(n15274), .A(n14868), .ZN(n14874) );
  AOI21_X1 U18569 ( .B1(n14870), .B2(n14869), .A(n14851), .ZN(n15498) );
  AOI22_X1 U18570 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n20955), .B1(n20954), 
        .B2(n15498), .ZN(n14871) );
  OAI211_X1 U18571 ( .C1(n20901), .C2(n14872), .A(n14871), .B(n20925), .ZN(
        n14873) );
  AOI211_X1 U18572 ( .C1(n14875), .C2(P1_REIP_REG_10__SCAN_IN), .A(n14874), 
        .B(n14873), .ZN(n14876) );
  OAI21_X1 U18573 ( .B1(n15052), .B2(n20907), .A(n14876), .ZN(P1_U2830) );
  AOI21_X1 U18574 ( .B1(n14877), .B2(n14948), .A(n14939), .ZN(n15290) );
  INV_X1 U18575 ( .A(n15290), .ZN(n15055) );
  NAND2_X1 U18576 ( .A1(n20959), .A2(n20940), .ZN(n20923) );
  NOR2_X1 U18577 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20923), .ZN(n14886) );
  OR2_X1 U18578 ( .A1(n14879), .A2(n14880), .ZN(n14881) );
  AND2_X1 U18579 ( .A1(n14878), .A2(n14881), .ZN(n17562) );
  INV_X1 U18580 ( .A(n17562), .ZN(n14882) );
  OAI22_X1 U18581 ( .A1(n20927), .A2(n14882), .B1(n20952), .B2(n15288), .ZN(
        n14885) );
  INV_X1 U18582 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21675) );
  INV_X1 U18583 ( .A(n20904), .ZN(n20953) );
  AOI21_X1 U18584 ( .B1(n20959), .B2(n20889), .A(n20953), .ZN(n20891) );
  AOI22_X1 U18585 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20956), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(n20955), .ZN(n14883) );
  OAI211_X1 U18586 ( .C1(n21675), .C2(n20891), .A(n14883), .B(n20925), .ZN(
        n14884) );
  AOI211_X1 U18587 ( .C1(n14887), .C2(n14886), .A(n14885), .B(n14884), .ZN(
        n14888) );
  OAI21_X1 U18588 ( .B1(n15055), .B2(n20907), .A(n14888), .ZN(P1_U2832) );
  AOI22_X1 U18589 ( .A1(n20956), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20953), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14890) );
  NAND2_X1 U18590 ( .A1(n20958), .A2(n21540), .ZN(n14889) );
  OAI211_X1 U18591 ( .C1(n20952), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14890), .B(n14889), .ZN(n14893) );
  INV_X1 U18592 ( .A(n14186), .ZN(n14891) );
  OAI22_X1 U18593 ( .A1(n14891), .A2(n20927), .B1(n20938), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14892) );
  AOI211_X1 U18594 ( .C1(n20955), .C2(P1_EBX_REG_1__SCAN_IN), .A(n14893), .B(
        n14892), .ZN(n14894) );
  OAI21_X1 U18595 ( .B1(n20962), .B2(n14895), .A(n14894), .ZN(P1_U2839) );
  NOR2_X1 U18596 ( .A1(n20927), .A2(n14896), .ZN(n14900) );
  OAI21_X1 U18597 ( .B1(n20965), .B2(n20956), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14898) );
  NAND2_X1 U18598 ( .A1(n20958), .A2(n13156), .ZN(n14897) );
  OAI211_X1 U18599 ( .C1(n20948), .C2(n12555), .A(n14898), .B(n14897), .ZN(
        n14899) );
  AOI211_X1 U18600 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n14901), .A(n14900), .B(
        n14899), .ZN(n14902) );
  OAI21_X1 U18601 ( .B1(n20962), .B2(n14903), .A(n14902), .ZN(P1_U2840) );
  OAI222_X1 U18602 ( .A1(n14927), .A2(n14906), .B1(n14905), .B2(n20978), .C1(
        n14904), .C2(n14959), .ZN(P1_U2842) );
  OAI222_X1 U18603 ( .A1(n14927), .A2(n14908), .B1(n14907), .B2(n20978), .C1(
        n15303), .C2(n14959), .ZN(P1_U2843) );
  INV_X1 U18604 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14909) );
  OAI222_X1 U18605 ( .A1(n14927), .A2(n14910), .B1(n14909), .B2(n20978), .C1(
        n15319), .C2(n14959), .ZN(P1_U2844) );
  INV_X1 U18606 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n21956) );
  OAI222_X1 U18607 ( .A1(n14978), .A2(n14927), .B1(n21956), .B2(n20978), .C1(
        n14959), .C2(n15328), .ZN(P1_U2845) );
  OAI222_X1 U18608 ( .A1(n14911), .A2(n14927), .B1(n21892), .B2(n20978), .C1(
        n15333), .C2(n14959), .ZN(P1_U2846) );
  OAI222_X1 U18609 ( .A1(n14927), .A2(n14913), .B1(n14912), .B2(n20978), .C1(
        n15348), .C2(n14959), .ZN(P1_U2847) );
  AOI22_X1 U18610 ( .A1(n15359), .A2(n20974), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14943), .ZN(n14914) );
  OAI21_X1 U18611 ( .B1(n14998), .B2(n14927), .A(n14914), .ZN(P1_U2848) );
  AOI22_X1 U18612 ( .A1(n15369), .A2(n20974), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14943), .ZN(n14915) );
  OAI21_X1 U18613 ( .B1(n14999), .B2(n14927), .A(n14915), .ZN(P1_U2849) );
  AOI22_X1 U18614 ( .A1(n15382), .A2(n20974), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14943), .ZN(n14916) );
  OAI21_X1 U18615 ( .B1(n14917), .B2(n14927), .A(n14916), .ZN(P1_U2850) );
  INV_X1 U18616 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14919) );
  OAI222_X1 U18617 ( .A1(n14920), .A2(n14927), .B1(n14919), .B2(n20978), .C1(
        n14918), .C2(n14959), .ZN(P1_U2851) );
  INV_X1 U18618 ( .A(n15168), .ZN(n14922) );
  OAI222_X1 U18619 ( .A1(n14922), .A2(n14927), .B1(n14921), .B2(n20978), .C1(
        n15393), .C2(n14959), .ZN(P1_U2852) );
  AOI22_X1 U18620 ( .A1(n15412), .A2(n20974), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14943), .ZN(n14923) );
  OAI21_X1 U18621 ( .B1(n15174), .B2(n14927), .A(n14923), .ZN(P1_U2853) );
  AOI22_X1 U18622 ( .A1(n15415), .A2(n20974), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n14943), .ZN(n14924) );
  OAI21_X1 U18623 ( .B1(n14925), .B2(n14927), .A(n14924), .ZN(P1_U2854) );
  AOI22_X1 U18624 ( .A1(n15433), .A2(n20974), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14943), .ZN(n14926) );
  OAI21_X1 U18625 ( .B1(n15025), .B2(n14927), .A(n14926), .ZN(P1_U2855) );
  INV_X1 U18626 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21929) );
  OAI222_X1 U18627 ( .A1(n15212), .A2(n14927), .B1(n21929), .B2(n20978), .C1(
        n15442), .C2(n14959), .ZN(P1_U2856) );
  OAI22_X1 U18628 ( .A1(n15450), .A2(n14959), .B1(n14928), .B2(n20978), .ZN(
        n14929) );
  INV_X1 U18629 ( .A(n14929), .ZN(n14930) );
  OAI21_X1 U18630 ( .B1(n15223), .B2(n14927), .A(n14930), .ZN(P1_U2857) );
  INV_X1 U18631 ( .A(n15234), .ZN(n15044) );
  OAI222_X1 U18632 ( .A1(n15044), .A2(n14927), .B1(n14931), .B2(n20978), .C1(
        n15451), .C2(n14959), .ZN(P1_U2858) );
  INV_X1 U18633 ( .A(n15241), .ZN(n15047) );
  OAI222_X1 U18634 ( .A1(n15047), .A2(n14927), .B1(n21859), .B2(n20978), .C1(
        n15468), .C2(n14959), .ZN(P1_U2859) );
  OAI222_X1 U18635 ( .A1(n15251), .A2(n14927), .B1(n14932), .B2(n20978), .C1(
        n15482), .C2(n14959), .ZN(P1_U2860) );
  OAI22_X1 U18636 ( .A1(n15488), .A2(n14959), .B1(n14933), .B2(n20978), .ZN(
        n14934) );
  AOI21_X1 U18637 ( .B1(n15263), .B2(n20975), .A(n14934), .ZN(n14935) );
  INV_X1 U18638 ( .A(n14935), .ZN(P1_U2861) );
  AOI22_X1 U18639 ( .A1(n15498), .A2(n20974), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14943), .ZN(n14936) );
  OAI21_X1 U18640 ( .B1(n15052), .B2(n14927), .A(n14936), .ZN(P1_U2862) );
  OAI21_X1 U18641 ( .B1(n14939), .B2(n14938), .A(n14937), .ZN(n15280) );
  NAND2_X1 U18642 ( .A1(n14878), .A2(n14940), .ZN(n14941) );
  NAND2_X1 U18643 ( .A1(n14869), .A2(n14941), .ZN(n20892) );
  OAI222_X1 U18644 ( .A1(n15280), .A2(n14927), .B1(n14942), .B2(n20978), .C1(
        n14959), .C2(n20892), .ZN(P1_U2863) );
  AOI22_X1 U18645 ( .A1(n17562), .A2(n20974), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14943), .ZN(n14944) );
  OAI21_X1 U18646 ( .B1(n15055), .B2(n14927), .A(n14944), .ZN(P1_U2864) );
  NAND2_X1 U18647 ( .A1(n14946), .A2(n14945), .ZN(n14947) );
  NAND2_X1 U18648 ( .A1(n14948), .A2(n14947), .ZN(n20908) );
  NOR2_X1 U18649 ( .A1(n9926), .A2(n14949), .ZN(n14950) );
  OR2_X1 U18650 ( .A1(n14879), .A2(n14950), .ZN(n20912) );
  OAI222_X1 U18651 ( .A1(n20908), .A2(n14927), .B1(n14951), .B2(n20978), .C1(
        n14959), .C2(n20912), .ZN(P1_U2865) );
  AND2_X1 U18652 ( .A1(n14953), .A2(n14952), .ZN(n14954) );
  NOR2_X1 U18653 ( .A1(n14861), .A2(n14954), .ZN(n20931) );
  INV_X1 U18654 ( .A(n20931), .ZN(n15059) );
  NAND2_X1 U18655 ( .A1(n14956), .A2(n14957), .ZN(n14958) );
  NAND2_X1 U18656 ( .A1(n14955), .A2(n14958), .ZN(n20926) );
  OAI222_X1 U18657 ( .A1(n15059), .A2(n14927), .B1(n14960), .B2(n20978), .C1(
        n14959), .C2(n20926), .ZN(P1_U2867) );
  INV_X1 U18658 ( .A(DATAI_30_), .ZN(n14967) );
  NAND2_X1 U18659 ( .A1(n15073), .A2(n15026), .ZN(n14966) );
  AND2_X1 U18660 ( .A1(n14961), .A2(n21106), .ZN(n14962) );
  INV_X1 U18661 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14963) );
  OAI22_X1 U18662 ( .A1(n15027), .A2(n15043), .B1(n15066), .B2(n14963), .ZN(
        n14964) );
  AOI21_X1 U18663 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n15029), .A(n14964), .ZN(
        n14965) );
  OAI211_X1 U18664 ( .C1(n15033), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        P1_U2874) );
  INV_X1 U18665 ( .A(DATAI_29_), .ZN(n14972) );
  NAND2_X1 U18666 ( .A1(n15079), .A2(n15026), .ZN(n14971) );
  OAI22_X1 U18667 ( .A1(n15027), .A2(n15045), .B1(n15066), .B2(n14968), .ZN(
        n14969) );
  AOI21_X1 U18668 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n15029), .A(n14969), .ZN(
        n14970) );
  OAI211_X1 U18669 ( .C1(n15033), .C2(n14972), .A(n14971), .B(n14970), .ZN(
        P1_U2875) );
  INV_X1 U18670 ( .A(DATAI_28_), .ZN(n14977) );
  NAND2_X1 U18671 ( .A1(n15093), .A2(n15026), .ZN(n14976) );
  INV_X1 U18672 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n21082) );
  NOR2_X1 U18673 ( .A1(n15037), .A2(n21082), .ZN(n14974) );
  OAI22_X1 U18674 ( .A1(n15027), .A2(n15048), .B1(n15066), .B2(n14256), .ZN(
        n14973) );
  NOR2_X1 U18675 ( .A1(n14974), .A2(n14973), .ZN(n14975) );
  OAI211_X1 U18676 ( .C1(n15033), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        P1_U2876) );
  INV_X1 U18677 ( .A(DATAI_27_), .ZN(n14983) );
  INV_X1 U18678 ( .A(n14978), .ZN(n15103) );
  NAND2_X1 U18679 ( .A1(n15103), .A2(n15026), .ZN(n14982) );
  OAI22_X1 U18680 ( .A1(n15027), .A2(n15049), .B1(n15066), .B2(n14979), .ZN(
        n14980) );
  AOI21_X1 U18681 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n15029), .A(n14980), .ZN(
        n14981) );
  OAI211_X1 U18682 ( .C1(n15033), .C2(n14983), .A(n14982), .B(n14981), .ZN(
        P1_U2877) );
  INV_X1 U18683 ( .A(DATAI_26_), .ZN(n14989) );
  NAND2_X1 U18684 ( .A1(n15112), .A2(n15026), .ZN(n14988) );
  INV_X1 U18685 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n21068) );
  NOR2_X1 U18686 ( .A1(n15037), .A2(n21068), .ZN(n14986) );
  OAI22_X1 U18687 ( .A1(n15027), .A2(n15051), .B1(n15066), .B2(n14984), .ZN(
        n14985) );
  NOR2_X1 U18688 ( .A1(n14986), .A2(n14985), .ZN(n14987) );
  OAI211_X1 U18689 ( .C1(n15033), .C2(n14989), .A(n14988), .B(n14987), .ZN(
        P1_U2878) );
  INV_X1 U18690 ( .A(DATAI_25_), .ZN(n14993) );
  NAND2_X1 U18691 ( .A1(n15123), .A2(n15026), .ZN(n14992) );
  OAI22_X1 U18692 ( .A1(n15027), .A2(n15053), .B1(n15066), .B2(n21797), .ZN(
        n14990) );
  AOI21_X1 U18693 ( .B1(n15029), .B2(BUF1_REG_25__SCAN_IN), .A(n14990), .ZN(
        n14991) );
  OAI211_X1 U18694 ( .C1(n15033), .C2(n14993), .A(n14992), .B(n14991), .ZN(
        P1_U2879) );
  OAI22_X1 U18695 ( .A1(n15027), .A2(n15054), .B1(n15066), .B2(n14994), .ZN(
        n14995) );
  AOI21_X1 U18696 ( .B1(n15029), .B2(BUF1_REG_24__SCAN_IN), .A(n14995), .ZN(
        n14997) );
  NAND2_X1 U18697 ( .A1(n15039), .A2(DATAI_24_), .ZN(n14996) );
  OAI211_X1 U18698 ( .C1(n14998), .C2(n15067), .A(n14997), .B(n14996), .ZN(
        P1_U2880) );
  INV_X1 U18699 ( .A(DATAI_23_), .ZN(n15003) );
  INV_X1 U18700 ( .A(n14999), .ZN(n15140) );
  NAND2_X1 U18701 ( .A1(n15140), .A2(n15026), .ZN(n15002) );
  OAI22_X1 U18702 ( .A1(n15027), .A2(n21108), .B1(n15066), .B2(n14119), .ZN(
        n15000) );
  AOI21_X1 U18703 ( .B1(n15029), .B2(BUF1_REG_23__SCAN_IN), .A(n15000), .ZN(
        n15001) );
  OAI211_X1 U18704 ( .C1(n15033), .C2(n15003), .A(n15002), .B(n15001), .ZN(
        P1_U2881) );
  INV_X1 U18705 ( .A(DATAI_22_), .ZN(n15007) );
  NAND2_X1 U18706 ( .A1(n15149), .A2(n15026), .ZN(n15006) );
  OAI22_X1 U18707 ( .A1(n15027), .A2(n21097), .B1(n15066), .B2(n14239), .ZN(
        n15004) );
  AOI21_X1 U18708 ( .B1(n15029), .B2(BUF1_REG_22__SCAN_IN), .A(n15004), .ZN(
        n15005) );
  OAI211_X1 U18709 ( .C1(n15033), .C2(n15007), .A(n15006), .B(n15005), .ZN(
        P1_U2882) );
  INV_X1 U18710 ( .A(DATAI_21_), .ZN(n15011) );
  NAND2_X1 U18711 ( .A1(n15157), .A2(n15026), .ZN(n15010) );
  OAI22_X1 U18712 ( .A1(n15027), .A2(n21092), .B1(n15066), .B2(n14102), .ZN(
        n15008) );
  AOI21_X1 U18713 ( .B1(n15029), .B2(BUF1_REG_21__SCAN_IN), .A(n15008), .ZN(
        n15009) );
  OAI211_X1 U18714 ( .C1(n15033), .C2(n15011), .A(n15010), .B(n15009), .ZN(
        P1_U2883) );
  INV_X1 U18715 ( .A(DATAI_20_), .ZN(n15016) );
  NAND2_X1 U18716 ( .A1(n15168), .A2(n15026), .ZN(n15015) );
  INV_X1 U18717 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n21081) );
  NOR2_X1 U18718 ( .A1(n15037), .A2(n21081), .ZN(n15013) );
  OAI22_X1 U18719 ( .A1(n15027), .A2(n21084), .B1(n15066), .B2(n21910), .ZN(
        n15012) );
  NOR2_X1 U18720 ( .A1(n15013), .A2(n15012), .ZN(n15014) );
  OAI211_X1 U18721 ( .C1(n15033), .C2(n15016), .A(n15015), .B(n15014), .ZN(
        P1_U2884) );
  INV_X1 U18722 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16594) );
  INV_X1 U18723 ( .A(n15027), .ZN(n15035) );
  AOI22_X1 U18724 ( .A1(n15035), .A2(n21078), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15034), .ZN(n15017) );
  OAI21_X1 U18725 ( .B1(n15037), .B2(n16594), .A(n15017), .ZN(n15018) );
  AOI21_X1 U18726 ( .B1(n15039), .B2(DATAI_19_), .A(n15018), .ZN(n15019) );
  OAI21_X1 U18727 ( .B1(n15174), .B2(n15067), .A(n15019), .ZN(P1_U2885) );
  INV_X1 U18728 ( .A(DATAI_18_), .ZN(n15024) );
  NAND2_X1 U18729 ( .A1(n15186), .A2(n15026), .ZN(n15023) );
  INV_X1 U18730 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n21067) );
  NOR2_X1 U18731 ( .A1(n15037), .A2(n21067), .ZN(n15021) );
  OAI22_X1 U18732 ( .A1(n15027), .A2(n21072), .B1(n15066), .B2(n22013), .ZN(
        n15020) );
  NOR2_X1 U18733 ( .A1(n15021), .A2(n15020), .ZN(n15022) );
  OAI211_X1 U18734 ( .C1(n15033), .C2(n15024), .A(n15023), .B(n15022), .ZN(
        P1_U2886) );
  INV_X1 U18735 ( .A(DATAI_17_), .ZN(n15032) );
  INV_X1 U18736 ( .A(n15025), .ZN(n15200) );
  NAND2_X1 U18737 ( .A1(n15200), .A2(n15026), .ZN(n15031) );
  OAI22_X1 U18738 ( .A1(n15027), .A2(n21062), .B1(n15066), .B2(n14107), .ZN(
        n15028) );
  AOI21_X1 U18739 ( .B1(n15029), .B2(BUF1_REG_17__SCAN_IN), .A(n15028), .ZN(
        n15030) );
  OAI211_X1 U18740 ( .C1(n15033), .C2(n15032), .A(n15031), .B(n15030), .ZN(
        P1_U2887) );
  INV_X1 U18741 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n22004) );
  AOI22_X1 U18742 ( .A1(n15035), .A2(n15607), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15034), .ZN(n15036) );
  OAI21_X1 U18743 ( .B1(n15037), .B2(n22004), .A(n15036), .ZN(n15038) );
  AOI21_X1 U18744 ( .B1(n15039), .B2(DATAI_16_), .A(n15038), .ZN(n15040) );
  OAI21_X1 U18745 ( .B1(n15212), .B2(n15067), .A(n15040), .ZN(P1_U2888) );
  OAI222_X1 U18746 ( .A1(n15223), .A2(n15067), .B1(n15066), .B2(n15042), .C1(
        n15064), .C2(n15041), .ZN(P1_U2889) );
  OAI222_X1 U18747 ( .A1(n15044), .A2(n15067), .B1(n14223), .B2(n15066), .C1(
        n15064), .C2(n15043), .ZN(P1_U2890) );
  INV_X1 U18748 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15046) );
  OAI222_X1 U18749 ( .A1(n15047), .A2(n15067), .B1(n15046), .B2(n15066), .C1(
        n15064), .C2(n15045), .ZN(P1_U2891) );
  OAI222_X1 U18750 ( .A1(n15251), .A2(n15067), .B1(n20983), .B2(n15066), .C1(
        n15064), .C2(n15048), .ZN(P1_U2892) );
  OAI222_X1 U18751 ( .A1(n15050), .A2(n15067), .B1(n14253), .B2(n15066), .C1(
        n15064), .C2(n15049), .ZN(P1_U2893) );
  OAI222_X1 U18752 ( .A1(n15052), .A2(n15067), .B1(n14231), .B2(n15066), .C1(
        n15064), .C2(n15051), .ZN(P1_U2894) );
  OAI222_X1 U18753 ( .A1(n15280), .A2(n15067), .B1(n14228), .B2(n15066), .C1(
        n15064), .C2(n15053), .ZN(P1_U2895) );
  OAI222_X1 U18754 ( .A1(n15055), .A2(n15067), .B1(n14244), .B2(n15066), .C1(
        n15064), .C2(n15054), .ZN(P1_U2896) );
  OAI222_X1 U18755 ( .A1(n20908), .A2(n15067), .B1(n14139), .B2(n15066), .C1(
        n15064), .C2(n21108), .ZN(P1_U2897) );
  INV_X1 U18756 ( .A(n14862), .ZN(n15056) );
  XNOR2_X1 U18757 ( .A(n14861), .B(n15056), .ZN(n20971) );
  INV_X1 U18758 ( .A(n20971), .ZN(n15057) );
  OAI222_X1 U18759 ( .A1(n15064), .A2(n21097), .B1(n15067), .B2(n15057), .C1(
        n14142), .C2(n15066), .ZN(P1_U2898) );
  OAI222_X1 U18760 ( .A1(n15059), .A2(n15067), .B1(n15058), .B2(n15066), .C1(
        n15064), .C2(n21092), .ZN(P1_U2899) );
  XOR2_X1 U18761 ( .A(n14448), .B(n15060), .Z(n20999) );
  INV_X1 U18762 ( .A(n20999), .ZN(n15062) );
  OAI222_X1 U18763 ( .A1(n15064), .A2(n21084), .B1(n15067), .B2(n15062), .C1(
        n15061), .C2(n15066), .ZN(P1_U2900) );
  OAI222_X1 U18764 ( .A1(n15296), .A2(n15067), .B1(n15066), .B2(n15065), .C1(
        n15064), .C2(n15063), .ZN(P1_U2901) );
  INV_X1 U18765 ( .A(n15068), .ZN(n15071) );
  AOI21_X1 U18766 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15069), .ZN(n15070) );
  OAI21_X1 U18767 ( .B1(n21006), .B2(n15071), .A(n15070), .ZN(n15072) );
  AOI21_X1 U18768 ( .B1(n15073), .B2(n21000), .A(n15072), .ZN(n15074) );
  OAI21_X1 U18769 ( .B1(n15075), .B2(n20873), .A(n15074), .ZN(P1_U2969) );
  NOR2_X1 U18770 ( .A1(n17570), .A2(n21708), .ZN(n15304) );
  AOI21_X1 U18771 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15304), .ZN(n15076) );
  OAI21_X1 U18772 ( .B1(n21006), .B2(n15077), .A(n15076), .ZN(n15078) );
  AOI21_X1 U18773 ( .B1(n15079), .B2(n21000), .A(n15078), .ZN(n15080) );
  OAI21_X1 U18774 ( .B1(n15313), .B2(n20873), .A(n15080), .ZN(P1_U2970) );
  NAND2_X1 U18775 ( .A1(n15257), .A2(n15338), .ZN(n15081) );
  NAND2_X1 U18776 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15082) );
  AND3_X1 U18777 ( .A1(n15118), .A2(n15335), .A3(n15099), .ZN(n15083) );
  NAND4_X1 U18778 ( .A1(n15084), .A2(n15083), .A3(n12461), .A4(n15128), .ZN(
        n15085) );
  MUX2_X1 U18779 ( .A(n15086), .B(n15085), .S(n10812), .Z(n15088) );
  XNOR2_X1 U18780 ( .A(n15088), .B(n15087), .ZN(n15323) );
  NOR2_X1 U18781 ( .A1(n17570), .A2(n15089), .ZN(n15318) );
  AOI21_X1 U18782 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15318), .ZN(n15090) );
  OAI21_X1 U18783 ( .B1(n21006), .B2(n15091), .A(n15090), .ZN(n15092) );
  AOI21_X1 U18784 ( .B1(n15093), .B2(n21000), .A(n15092), .ZN(n15094) );
  OR2_X1 U18785 ( .A1(n15096), .A2(n15095), .ZN(n15098) );
  NOR2_X1 U18786 ( .A1(n17570), .A2(n22020), .ZN(n15326) );
  AOI21_X1 U18787 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15326), .ZN(n15100) );
  OAI21_X1 U18788 ( .B1(n21006), .B2(n15101), .A(n15100), .ZN(n15102) );
  AOI21_X1 U18789 ( .B1(n15103), .B2(n21000), .A(n15102), .ZN(n15104) );
  INV_X1 U18790 ( .A(n15136), .ZN(n15125) );
  OAI21_X1 U18791 ( .B1(n15125), .B2(n15338), .A(n15257), .ZN(n15106) );
  NAND2_X1 U18792 ( .A1(n15105), .A2(n15106), .ZN(n15107) );
  XNOR2_X1 U18793 ( .A(n15107), .B(n15335), .ZN(n15344) );
  INV_X1 U18794 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15108) );
  NOR2_X1 U18795 ( .A1(n17570), .A2(n15108), .ZN(n15340) );
  AOI21_X1 U18796 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15340), .ZN(n15109) );
  OAI21_X1 U18797 ( .B1(n21006), .B2(n15110), .A(n15109), .ZN(n15111) );
  AOI21_X1 U18798 ( .B1(n15112), .B2(n21000), .A(n15111), .ZN(n15113) );
  OAI21_X1 U18799 ( .B1(n20873), .B2(n15344), .A(n15113), .ZN(P1_U2973) );
  INV_X1 U18800 ( .A(n15114), .ZN(n15115) );
  MUX2_X1 U18801 ( .A(n15115), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .S(
        n15257), .Z(n15117) );
  NAND2_X1 U18802 ( .A1(n15126), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15116) );
  NAND2_X1 U18803 ( .A1(n15117), .A2(n15116), .ZN(n15119) );
  XNOR2_X1 U18804 ( .A(n15119), .B(n15118), .ZN(n15352) );
  NOR2_X1 U18805 ( .A1(n17570), .A2(n21702), .ZN(n15346) );
  AOI21_X1 U18806 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15346), .ZN(n15120) );
  OAI21_X1 U18807 ( .B1(n21006), .B2(n15121), .A(n15120), .ZN(n15122) );
  AOI21_X1 U18808 ( .B1(n15123), .B2(n21000), .A(n15122), .ZN(n15124) );
  OAI21_X1 U18809 ( .B1(n20873), .B2(n15352), .A(n15124), .ZN(P1_U2974) );
  NAND2_X1 U18810 ( .A1(n15126), .A2(n15125), .ZN(n15127) );
  MUX2_X1 U18811 ( .A(n15127), .B(n15126), .S(n15257), .Z(n15129) );
  XNOR2_X1 U18812 ( .A(n15129), .B(n15128), .ZN(n15362) );
  NOR2_X1 U18813 ( .A1(n17570), .A2(n21700), .ZN(n15357) );
  AOI21_X1 U18814 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15357), .ZN(n15130) );
  OAI21_X1 U18815 ( .B1(n21006), .B2(n15131), .A(n15130), .ZN(n15132) );
  AOI21_X1 U18816 ( .B1(n15133), .B2(n21000), .A(n15132), .ZN(n15134) );
  XNOR2_X1 U18817 ( .A(n15257), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15135) );
  XNOR2_X1 U18818 ( .A(n15136), .B(n15135), .ZN(n15371) );
  NOR2_X1 U18819 ( .A1(n17570), .A2(n21698), .ZN(n15364) );
  AOI21_X1 U18820 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15364), .ZN(n15137) );
  OAI21_X1 U18821 ( .B1(n21006), .B2(n15138), .A(n15137), .ZN(n15139) );
  AOI21_X1 U18822 ( .B1(n15140), .B2(n21000), .A(n15139), .ZN(n15141) );
  OAI21_X1 U18823 ( .B1(n15371), .B2(n20873), .A(n15141), .ZN(P1_U2976) );
  NAND2_X1 U18824 ( .A1(n15143), .A2(n15142), .ZN(n15144) );
  XOR2_X1 U18825 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15144), .Z(
        n15385) );
  INV_X1 U18826 ( .A(n15145), .ZN(n15147) );
  NOR2_X1 U18827 ( .A1(n17570), .A2(n21696), .ZN(n15380) );
  AOI21_X1 U18828 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15380), .ZN(n15146) );
  OAI21_X1 U18829 ( .B1(n21006), .B2(n15147), .A(n15146), .ZN(n15148) );
  AOI21_X1 U18830 ( .B1(n15149), .B2(n21000), .A(n15148), .ZN(n15150) );
  OAI21_X1 U18831 ( .B1(n20873), .B2(n15385), .A(n15150), .ZN(P1_U2977) );
  INV_X1 U18832 ( .A(n15151), .ZN(n15416) );
  NAND3_X1 U18833 ( .A1(n15416), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15257), .ZN(n15162) );
  NOR2_X1 U18834 ( .A1(n15152), .A2(n15257), .ZN(n15159) );
  NAND2_X1 U18835 ( .A1(n15159), .A2(n15398), .ZN(n15160) );
  OAI21_X1 U18836 ( .B1(n15162), .B2(n15398), .A(n15160), .ZN(n15153) );
  XNOR2_X1 U18837 ( .A(n15153), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15392) );
  NOR2_X1 U18838 ( .A1(n17570), .A2(n21694), .ZN(n15387) );
  AOI21_X1 U18839 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15387), .ZN(n15154) );
  OAI21_X1 U18840 ( .B1(n21006), .B2(n15155), .A(n15154), .ZN(n15156) );
  AOI21_X1 U18841 ( .B1(n15157), .B2(n21000), .A(n15156), .ZN(n15158) );
  OAI21_X1 U18842 ( .B1(n15392), .B2(n20873), .A(n15158), .ZN(P1_U2978) );
  NOR2_X1 U18843 ( .A1(n15159), .A2(n15398), .ZN(n15163) );
  OAI21_X1 U18844 ( .B1(n15162), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15160), .ZN(n15161) );
  AOI21_X1 U18845 ( .B1(n15163), .B2(n15162), .A(n15161), .ZN(n15406) );
  INV_X1 U18846 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15164) );
  NOR2_X1 U18847 ( .A1(n17570), .A2(n15164), .ZN(n15402) );
  AOI21_X1 U18848 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15402), .ZN(n15165) );
  OAI21_X1 U18849 ( .B1(n21006), .B2(n15166), .A(n15165), .ZN(n15167) );
  AOI21_X1 U18850 ( .B1(n15168), .B2(n21000), .A(n15167), .ZN(n15169) );
  OAI21_X1 U18851 ( .B1(n15406), .B2(n20873), .A(n15169), .ZN(P1_U2979) );
  NOR2_X1 U18852 ( .A1(n15257), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15170) );
  MUX2_X1 U18853 ( .A(n15257), .B(n15170), .S(n15151), .Z(n15171) );
  XNOR2_X1 U18854 ( .A(n15171), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15414) );
  NAND2_X1 U18855 ( .A1(n21051), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15408) );
  OAI21_X1 U18856 ( .B1(n15173), .B2(n15172), .A(n15408), .ZN(n15176) );
  NOR2_X1 U18857 ( .A1(n15174), .A2(n15252), .ZN(n15175) );
  AOI211_X1 U18858 ( .C1(n15178), .C2(n15177), .A(n15176), .B(n15175), .ZN(
        n15179) );
  OAI21_X1 U18859 ( .B1(n20873), .B2(n15414), .A(n15179), .ZN(P1_U2980) );
  NOR2_X1 U18860 ( .A1(n17570), .A2(n21690), .ZN(n15422) );
  AOI21_X1 U18861 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15422), .ZN(n15180) );
  OAI21_X1 U18862 ( .B1(n21006), .B2(n15181), .A(n15180), .ZN(n15185) );
  NOR2_X1 U18863 ( .A1(n15182), .A2(n15183), .ZN(n15417) );
  NOR3_X1 U18864 ( .A1(n15417), .A2(n15416), .A3(n20873), .ZN(n15184) );
  AOI211_X1 U18865 ( .C1(n21000), .C2(n15186), .A(n15185), .B(n15184), .ZN(
        n15187) );
  INV_X1 U18866 ( .A(n15187), .ZN(P1_U2981) );
  NOR2_X1 U18867 ( .A1(n15257), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15195) );
  INV_X1 U18868 ( .A(n15188), .ZN(n15189) );
  NAND2_X1 U18869 ( .A1(n15257), .A2(n15189), .ZN(n15190) );
  NOR2_X1 U18870 ( .A1(n15265), .A2(n15192), .ZN(n15228) );
  AOI21_X1 U18871 ( .B1(n15228), .B2(n15193), .A(n9879), .ZN(n15194) );
  MUX2_X1 U18872 ( .A(n15195), .B(n15257), .S(n15194), .Z(n15196) );
  XNOR2_X1 U18873 ( .A(n15196), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15435) );
  NOR2_X1 U18874 ( .A1(n17570), .A2(n21799), .ZN(n15432) );
  AOI21_X1 U18875 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15432), .ZN(n15197) );
  OAI21_X1 U18876 ( .B1(n21006), .B2(n15198), .A(n15197), .ZN(n15199) );
  AOI21_X1 U18877 ( .B1(n15200), .B2(n21000), .A(n15199), .ZN(n15201) );
  OAI21_X1 U18878 ( .B1(n15435), .B2(n20873), .A(n15201), .ZN(P1_U2982) );
  INV_X1 U18879 ( .A(n15202), .ZN(n15204) );
  AOI21_X1 U18880 ( .B1(n15265), .B2(n15204), .A(n15203), .ZN(n15216) );
  NAND2_X1 U18881 ( .A1(n15216), .A2(n15214), .ZN(n15218) );
  NAND2_X1 U18882 ( .A1(n15218), .A2(n15213), .ZN(n15206) );
  XNOR2_X1 U18883 ( .A(n15206), .B(n15205), .ZN(n15436) );
  NAND2_X1 U18884 ( .A1(n15436), .A2(n21001), .ZN(n15211) );
  INV_X1 U18885 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15207) );
  NOR2_X1 U18886 ( .A1(n17570), .A2(n15207), .ZN(n15439) );
  NOR2_X1 U18887 ( .A1(n21006), .A2(n15208), .ZN(n15209) );
  AOI211_X1 U18888 ( .C1(n20992), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15439), .B(n15209), .ZN(n15210) );
  OAI211_X1 U18889 ( .C1(n15252), .C2(n15212), .A(n15211), .B(n15210), .ZN(
        P1_U2983) );
  INV_X1 U18890 ( .A(n15213), .ZN(n15217) );
  AND2_X1 U18891 ( .A1(n15214), .A2(n15213), .ZN(n15215) );
  OAI22_X1 U18892 ( .A1(n15218), .A2(n15217), .B1(n15216), .B2(n15215), .ZN(
        n15443) );
  NAND2_X1 U18893 ( .A1(n15443), .A2(n21001), .ZN(n15222) );
  NOR2_X1 U18894 ( .A1(n17570), .A2(n21993), .ZN(n15446) );
  NOR2_X1 U18895 ( .A1(n21006), .A2(n15219), .ZN(n15220) );
  AOI211_X1 U18896 ( .C1(n20992), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15446), .B(n15220), .ZN(n15221) );
  OAI211_X1 U18897 ( .C1(n15252), .C2(n15223), .A(n15222), .B(n15221), .ZN(
        P1_U2984) );
  NAND2_X1 U18898 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15225) );
  NAND2_X1 U18899 ( .A1(n15257), .A2(n15225), .ZN(n15237) );
  OAI21_X1 U18900 ( .B1(n15228), .B2(n15227), .A(n15226), .ZN(n15230) );
  XNOR2_X1 U18901 ( .A(n15257), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15229) );
  XNOR2_X1 U18902 ( .A(n15230), .B(n15229), .ZN(n15458) );
  AND2_X1 U18903 ( .A1(n21051), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15454) );
  AOI21_X1 U18904 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15454), .ZN(n15231) );
  OAI21_X1 U18905 ( .B1(n21006), .B2(n15232), .A(n15231), .ZN(n15233) );
  AOI21_X1 U18906 ( .B1(n15234), .B2(n21000), .A(n15233), .ZN(n15235) );
  OAI21_X1 U18907 ( .B1(n15458), .B2(n20873), .A(n15235), .ZN(P1_U2985) );
  AOI22_X1 U18908 ( .A1(n15265), .A2(n15237), .B1(n10812), .B2(n15236), .ZN(
        n15245) );
  AND2_X1 U18909 ( .A1(n15245), .A2(n9884), .ZN(n15243) );
  XOR2_X1 U18910 ( .A(n15224), .B(n9892), .Z(n15471) );
  NOR2_X1 U18911 ( .A1(n17570), .A2(n21685), .ZN(n15462) );
  AOI21_X1 U18912 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15462), .ZN(n15238) );
  OAI21_X1 U18913 ( .B1(n21006), .B2(n15239), .A(n15238), .ZN(n15240) );
  AOI21_X1 U18914 ( .B1(n15241), .B2(n21000), .A(n15240), .ZN(n15242) );
  OAI21_X1 U18915 ( .B1(n15471), .B2(n20873), .A(n15242), .ZN(P1_U2986) );
  INV_X1 U18916 ( .A(n15243), .ZN(n15244) );
  OAI21_X1 U18917 ( .B1(n9884), .B2(n15245), .A(n15244), .ZN(n15485) );
  NAND2_X1 U18918 ( .A1(n15485), .A2(n21001), .ZN(n15250) );
  NAND2_X1 U18919 ( .A1(n21051), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15481) );
  INV_X1 U18920 ( .A(n15481), .ZN(n15248) );
  NOR2_X1 U18921 ( .A1(n21006), .A2(n15246), .ZN(n15247) );
  AOI211_X1 U18922 ( .C1(n20992), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15248), .B(n15247), .ZN(n15249) );
  OAI211_X1 U18923 ( .C1(n15252), .C2(n15251), .A(n15250), .B(n15249), .ZN(
        P1_U2987) );
  NAND2_X1 U18924 ( .A1(n15253), .A2(n17539), .ZN(n15286) );
  INV_X1 U18925 ( .A(n15286), .ZN(n15256) );
  NAND2_X1 U18926 ( .A1(n15257), .A2(n15254), .ZN(n15284) );
  OAI21_X1 U18927 ( .B1(n15286), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n15284), .ZN(n15255) );
  OAI21_X1 U18928 ( .B1(n15256), .B2(n17569), .A(n15255), .ZN(n15279) );
  NOR2_X1 U18929 ( .A1(n15279), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15267) );
  NAND3_X1 U18930 ( .A1(n15267), .A2(n10812), .A3(n15266), .ZN(n15270) );
  NAND3_X1 U18931 ( .A1(n15265), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15257), .ZN(n15258) );
  NAND2_X1 U18932 ( .A1(n15270), .A2(n15258), .ZN(n15259) );
  XNOR2_X1 U18933 ( .A(n15259), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15494) );
  OR2_X1 U18934 ( .A1(n17570), .A2(n21682), .ZN(n15487) );
  NAND2_X1 U18935 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15260) );
  OAI211_X1 U18936 ( .C1(n21006), .C2(n15261), .A(n15487), .B(n15260), .ZN(
        n15262) );
  AOI21_X1 U18937 ( .B1(n15263), .B2(n21000), .A(n15262), .ZN(n15264) );
  OAI21_X1 U18938 ( .B1(n15494), .B2(n20873), .A(n15264), .ZN(P1_U2988) );
  XNOR2_X1 U18939 ( .A(n15265), .B(n15266), .ZN(n15269) );
  NOR2_X1 U18940 ( .A1(n15267), .A2(n15266), .ZN(n15268) );
  MUX2_X1 U18941 ( .A(n15269), .B(n15268), .S(n10812), .Z(n15272) );
  INV_X1 U18942 ( .A(n15270), .ZN(n15271) );
  NOR2_X1 U18943 ( .A1(n15272), .A2(n15271), .ZN(n15510) );
  NOR2_X1 U18944 ( .A1(n17570), .A2(n21680), .ZN(n15497) );
  AOI21_X1 U18945 ( .B1(n20992), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15497), .ZN(n15273) );
  OAI21_X1 U18946 ( .B1(n21006), .B2(n15274), .A(n15273), .ZN(n15275) );
  AOI21_X1 U18947 ( .B1(n15276), .B2(n21000), .A(n15275), .ZN(n15277) );
  OAI21_X1 U18948 ( .B1(n15510), .B2(n20873), .A(n15277), .ZN(P1_U2989) );
  XNOR2_X1 U18949 ( .A(n15257), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15278) );
  XNOR2_X1 U18950 ( .A(n15279), .B(n15278), .ZN(n15519) );
  INV_X1 U18951 ( .A(n15280), .ZN(n20896) );
  NAND2_X1 U18952 ( .A1(n21051), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15512) );
  NAND2_X1 U18953 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15281) );
  OAI211_X1 U18954 ( .C1(n21006), .C2(n20894), .A(n15512), .B(n15281), .ZN(
        n15282) );
  AOI21_X1 U18955 ( .B1(n20896), .B2(n21000), .A(n15282), .ZN(n15283) );
  OAI21_X1 U18956 ( .B1(n15519), .B2(n20873), .A(n15283), .ZN(P1_U2990) );
  XNOR2_X1 U18957 ( .A(n15284), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15285) );
  XNOR2_X1 U18958 ( .A(n15286), .B(n15285), .ZN(n17564) );
  INV_X1 U18959 ( .A(n17564), .ZN(n15292) );
  AOI22_X1 U18960 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n21051), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15287) );
  OAI21_X1 U18961 ( .B1(n21006), .B2(n15288), .A(n15287), .ZN(n15289) );
  AOI21_X1 U18962 ( .B1(n15290), .B2(n21000), .A(n15289), .ZN(n15291) );
  OAI21_X1 U18963 ( .B1(n20873), .B2(n15292), .A(n15291), .ZN(P1_U2991) );
  XNOR2_X1 U18964 ( .A(n15293), .B(n21023), .ZN(n15295) );
  XNOR2_X1 U18965 ( .A(n15295), .B(n15294), .ZN(n21019) );
  INV_X1 U18966 ( .A(n21019), .ZN(n15302) );
  INV_X1 U18967 ( .A(n15296), .ZN(n15300) );
  AOI22_X1 U18968 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n21051), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n15297) );
  OAI21_X1 U18969 ( .B1(n21006), .B2(n15298), .A(n15297), .ZN(n15299) );
  AOI21_X1 U18970 ( .B1(n15300), .B2(n21000), .A(n15299), .ZN(n15301) );
  OAI21_X1 U18971 ( .B1(n20873), .B2(n15302), .A(n15301), .ZN(P1_U2996) );
  INV_X1 U18972 ( .A(n15303), .ZN(n15311) );
  INV_X1 U18973 ( .A(n15304), .ZN(n15307) );
  NAND3_X1 U18974 ( .A1(n15316), .A2(n15305), .A3(n15308), .ZN(n15306) );
  OAI211_X1 U18975 ( .C1(n15309), .C2(n15308), .A(n15307), .B(n15306), .ZN(
        n15310) );
  AOI21_X1 U18976 ( .B1(n15311), .B2(n21027), .A(n15310), .ZN(n15312) );
  OAI21_X1 U18977 ( .B1(n15313), .B2(n21012), .A(n15312), .ZN(P1_U3002) );
  AND3_X1 U18978 ( .A1(n15316), .A2(n15315), .A3(n15314), .ZN(n15317) );
  AOI211_X1 U18979 ( .C1(n15327), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15318), .B(n15317), .ZN(n15322) );
  INV_X1 U18980 ( .A(n15319), .ZN(n15320) );
  NAND2_X1 U18981 ( .A1(n15320), .A2(n21027), .ZN(n15321) );
  OAI211_X1 U18982 ( .C1(n15323), .C2(n21012), .A(n15322), .B(n15321), .ZN(
        P1_U3003) );
  NOR2_X1 U18983 ( .A1(n15324), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15325) );
  AOI211_X1 U18984 ( .C1(n15327), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15326), .B(n15325), .ZN(n15331) );
  INV_X1 U18985 ( .A(n15328), .ZN(n15329) );
  NAND2_X1 U18986 ( .A1(n15329), .A2(n21027), .ZN(n15330) );
  OAI211_X1 U18987 ( .C1(n15332), .C2(n21012), .A(n15331), .B(n15330), .ZN(
        P1_U3004) );
  NOR2_X1 U18988 ( .A1(n15333), .A2(n21054), .ZN(n15342) );
  NOR3_X1 U18989 ( .A1(n15363), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15334), .ZN(n15345) );
  INV_X1 U18990 ( .A(n15345), .ZN(n15336) );
  AOI21_X1 U18991 ( .B1(n15337), .B2(n15336), .A(n15335), .ZN(n15341) );
  NOR3_X1 U18992 ( .A1(n15363), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15338), .ZN(n15339) );
  NOR4_X1 U18993 ( .A1(n15342), .A2(n15341), .A3(n15340), .A4(n15339), .ZN(
        n15343) );
  OAI21_X1 U18994 ( .B1(n15344), .B2(n21012), .A(n15343), .ZN(P1_U3005) );
  AOI211_X1 U18995 ( .C1(n15347), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15346), .B(n15345), .ZN(n15351) );
  INV_X1 U18996 ( .A(n15348), .ZN(n15349) );
  NAND2_X1 U18997 ( .A1(n15349), .A2(n21027), .ZN(n15350) );
  OAI211_X1 U18998 ( .C1(n15352), .C2(n21012), .A(n15351), .B(n15350), .ZN(
        P1_U3006) );
  INV_X1 U18999 ( .A(n15353), .ZN(n15354) );
  OAI21_X1 U19000 ( .B1(n15355), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15354), .ZN(n15358) );
  NOR3_X1 U19001 ( .A1(n15363), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n12461), .ZN(n15356) );
  AOI211_X1 U19002 ( .C1(n15358), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15357), .B(n15356), .ZN(n15361) );
  NAND2_X1 U19003 ( .A1(n15359), .A2(n21027), .ZN(n15360) );
  OAI211_X1 U19004 ( .C1(n15362), .C2(n21012), .A(n15361), .B(n15360), .ZN(
        P1_U3007) );
  INV_X1 U19005 ( .A(n15363), .ZN(n15365) );
  AOI21_X1 U19006 ( .B1(n15365), .B2(n12461), .A(n15364), .ZN(n15366) );
  OAI21_X1 U19007 ( .B1(n15367), .B2(n12461), .A(n15366), .ZN(n15368) );
  AOI21_X1 U19008 ( .B1(n15369), .B2(n21027), .A(n15368), .ZN(n15370) );
  OAI21_X1 U19009 ( .B1(n15371), .B2(n21012), .A(n15370), .ZN(P1_U3008) );
  AND2_X1 U19010 ( .A1(n15396), .A2(n15372), .ZN(n15459) );
  INV_X1 U19011 ( .A(n15376), .ZN(n15395) );
  NAND3_X1 U19012 ( .A1(n15373), .A2(n15372), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15375) );
  NOR2_X1 U19013 ( .A1(n15460), .A2(n15376), .ZN(n15397) );
  AOI21_X1 U19014 ( .B1(n15459), .B2(n15395), .A(n15397), .ZN(n15410) );
  NOR3_X1 U19015 ( .A1(n15410), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15377), .ZN(n15386) );
  OR2_X1 U19016 ( .A1(n15386), .A2(n15388), .ZN(n15381) );
  NOR3_X1 U19017 ( .A1(n15410), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n15378), .ZN(n15379) );
  AOI211_X1 U19018 ( .C1(n15381), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15380), .B(n15379), .ZN(n15384) );
  NAND2_X1 U19019 ( .A1(n15382), .A2(n21027), .ZN(n15383) );
  OAI211_X1 U19020 ( .C1(n15385), .C2(n21012), .A(n15384), .B(n15383), .ZN(
        P1_U3009) );
  AOI211_X1 U19021 ( .C1(n15388), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15387), .B(n15386), .ZN(n15391) );
  NAND2_X1 U19022 ( .A1(n15389), .A2(n21027), .ZN(n15390) );
  OAI211_X1 U19023 ( .C1(n15392), .C2(n21012), .A(n15391), .B(n15390), .ZN(
        P1_U3010) );
  NOR2_X1 U19024 ( .A1(n15393), .A2(n21054), .ZN(n15404) );
  OAI21_X1 U19025 ( .B1(n21008), .B2(n15395), .A(n15394), .ZN(n15407) );
  INV_X1 U19026 ( .A(n15407), .ZN(n15400) );
  OAI21_X1 U19027 ( .B1(n15397), .B2(n15396), .A(n22032), .ZN(n15399) );
  AOI21_X1 U19028 ( .B1(n15400), .B2(n15399), .A(n15398), .ZN(n15403) );
  NOR3_X1 U19029 ( .A1(n15410), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n22032), .ZN(n15401) );
  NOR4_X1 U19030 ( .A1(n15404), .A2(n15403), .A3(n15402), .A4(n15401), .ZN(
        n15405) );
  OAI21_X1 U19031 ( .B1(n15406), .B2(n21012), .A(n15405), .ZN(P1_U3011) );
  NAND2_X1 U19032 ( .A1(n15407), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15409) );
  OAI211_X1 U19033 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15410), .A(
        n15409), .B(n15408), .ZN(n15411) );
  AOI21_X1 U19034 ( .B1(n15412), .B2(n21027), .A(n15411), .ZN(n15413) );
  OAI21_X1 U19035 ( .B1(n15414), .B2(n21012), .A(n15413), .ZN(P1_U3012) );
  INV_X1 U19036 ( .A(n15415), .ZN(n15426) );
  OR3_X1 U19037 ( .A1(n15417), .A2(n15416), .A3(n21012), .ZN(n15425) );
  NOR2_X1 U19038 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15460), .ZN(
        n15418) );
  AOI211_X1 U19039 ( .C1(n15463), .C2(n17559), .A(n15418), .B(n15465), .ZN(
        n15452) );
  OAI21_X1 U19040 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21041), .A(
        n15452), .ZN(n15447) );
  AOI21_X1 U19041 ( .B1(n17561), .B2(n15420), .A(n15447), .ZN(n15428) );
  INV_X1 U19042 ( .A(n15428), .ZN(n15423) );
  INV_X1 U19043 ( .A(n15455), .ZN(n15419) );
  NOR2_X1 U19044 ( .A1(n15419), .A2(n15456), .ZN(n15427) );
  INV_X1 U19045 ( .A(n15427), .ZN(n15444) );
  NOR3_X1 U19046 ( .A1(n15444), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15420), .ZN(n15421) );
  AOI211_X1 U19047 ( .C1(n15423), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15422), .B(n15421), .ZN(n15424) );
  OAI211_X1 U19048 ( .C1(n21054), .C2(n15426), .A(n15425), .B(n15424), .ZN(
        P1_U3013) );
  NAND3_X1 U19049 ( .A1(n15427), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15429) );
  AOI21_X1 U19050 ( .B1(n15430), .B2(n15429), .A(n15428), .ZN(n15431) );
  AOI211_X1 U19051 ( .C1(n15433), .C2(n21027), .A(n15432), .B(n15431), .ZN(
        n15434) );
  OAI21_X1 U19052 ( .B1(n15435), .B2(n21012), .A(n15434), .ZN(P1_U3014) );
  NAND2_X1 U19053 ( .A1(n15436), .A2(n21042), .ZN(n15441) );
  XNOR2_X1 U19054 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15437) );
  NOR2_X1 U19055 ( .A1(n15444), .A2(n15437), .ZN(n15438) );
  AOI211_X1 U19056 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15447), .A(
        n15439), .B(n15438), .ZN(n15440) );
  OAI211_X1 U19057 ( .C1(n21054), .C2(n15442), .A(n15441), .B(n15440), .ZN(
        P1_U3015) );
  NAND2_X1 U19058 ( .A1(n15443), .A2(n21042), .ZN(n15449) );
  NOR2_X1 U19059 ( .A1(n15444), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15445) );
  AOI211_X1 U19060 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15447), .A(
        n15446), .B(n15445), .ZN(n15448) );
  OAI211_X1 U19061 ( .C1(n21054), .C2(n15450), .A(n15449), .B(n15448), .ZN(
        P1_U3016) );
  OAI22_X1 U19062 ( .A1(n15452), .A2(n15456), .B1(n21054), .B2(n15451), .ZN(
        n15453) );
  AOI211_X1 U19063 ( .C1(n15456), .C2(n15455), .A(n15454), .B(n15453), .ZN(
        n15457) );
  OAI21_X1 U19064 ( .B1(n15458), .B2(n21012), .A(n15457), .ZN(P1_U3017) );
  INV_X1 U19065 ( .A(n15459), .ZN(n15461) );
  NAND2_X1 U19066 ( .A1(n15461), .A2(n15460), .ZN(n15464) );
  AOI21_X1 U19067 ( .B1(n15464), .B2(n15463), .A(n15462), .ZN(n15467) );
  NAND2_X1 U19068 ( .A1(n15465), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15466) );
  OAI211_X1 U19069 ( .C1(n15468), .C2(n21054), .A(n15467), .B(n15466), .ZN(
        n15469) );
  INV_X1 U19070 ( .A(n15469), .ZN(n15470) );
  OAI21_X1 U19071 ( .B1(n15471), .B2(n21012), .A(n15470), .ZN(P1_U3018) );
  INV_X1 U19072 ( .A(n17559), .ZN(n21031) );
  INV_X1 U19073 ( .A(n15472), .ZN(n17556) );
  INV_X1 U19074 ( .A(n15489), .ZN(n15479) );
  NAND3_X1 U19075 ( .A1(n17556), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15479), .ZN(n15473) );
  NAND2_X1 U19076 ( .A1(n21028), .A2(n15473), .ZN(n15474) );
  OAI211_X1 U19077 ( .C1(n21031), .C2(n15475), .A(n21030), .B(n15474), .ZN(
        n15492) );
  AOI21_X1 U19078 ( .B1(n21035), .B2(n15476), .A(n15492), .ZN(n15477) );
  NOR2_X1 U19079 ( .A1(n15477), .A2(n15478), .ZN(n15484) );
  NAND2_X1 U19080 ( .A1(n15499), .A2(n21035), .ZN(n17560) );
  NAND2_X1 U19081 ( .A1(n21008), .A2(n17560), .ZN(n17583) );
  NAND4_X1 U19082 ( .A1(n17563), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15479), .A4(n15478), .ZN(n15480) );
  OAI211_X1 U19083 ( .C1(n15482), .C2(n21054), .A(n15481), .B(n15480), .ZN(
        n15483) );
  AOI211_X1 U19084 ( .C1(n15485), .C2(n21042), .A(n15484), .B(n15483), .ZN(
        n15486) );
  INV_X1 U19085 ( .A(n15486), .ZN(P1_U3019) );
  OAI21_X1 U19086 ( .B1(n15488), .B2(n21054), .A(n15487), .ZN(n15491) );
  INV_X1 U19087 ( .A(n17563), .ZN(n17582) );
  NOR3_X1 U19088 ( .A1(n17582), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15489), .ZN(n15490) );
  AOI211_X1 U19089 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15492), .A(
        n15491), .B(n15490), .ZN(n15493) );
  OAI21_X1 U19090 ( .B1(n15494), .B2(n21012), .A(n15493), .ZN(P1_U3020) );
  INV_X1 U19091 ( .A(n15506), .ZN(n15495) );
  NOR4_X1 U19092 ( .A1(n17582), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15505), .A4(n15495), .ZN(n15496) );
  AOI211_X1 U19093 ( .C1(n21027), .C2(n15498), .A(n15497), .B(n15496), .ZN(
        n15509) );
  INV_X1 U19094 ( .A(n15499), .ZN(n15500) );
  NAND2_X1 U19095 ( .A1(n17559), .A2(n15500), .ZN(n15501) );
  NAND2_X1 U19096 ( .A1(n21030), .A2(n15501), .ZN(n21009) );
  NAND2_X1 U19097 ( .A1(n17556), .A2(n15506), .ZN(n15502) );
  NOR2_X1 U19098 ( .A1(n21009), .A2(n15502), .ZN(n15503) );
  NOR2_X1 U19099 ( .A1(n15504), .A2(n15503), .ZN(n15516) );
  AND2_X1 U19100 ( .A1(n15506), .A2(n15505), .ZN(n15507) );
  AND2_X1 U19101 ( .A1(n17563), .A2(n15507), .ZN(n15515) );
  OAI21_X1 U19102 ( .B1(n15516), .B2(n15515), .A(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15508) );
  OAI211_X1 U19103 ( .C1(n15510), .C2(n21012), .A(n15509), .B(n15508), .ZN(
        P1_U3021) );
  INV_X1 U19104 ( .A(n20892), .ZN(n15511) );
  NAND2_X1 U19105 ( .A1(n15511), .A2(n21027), .ZN(n15513) );
  NAND2_X1 U19106 ( .A1(n15513), .A2(n15512), .ZN(n15514) );
  NOR2_X1 U19107 ( .A1(n15515), .A2(n15514), .ZN(n15518) );
  NAND2_X1 U19108 ( .A1(n15516), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15517) );
  OAI211_X1 U19109 ( .C1(n15519), .C2(n21012), .A(n15518), .B(n15517), .ZN(
        P1_U3022) );
  NOR2_X1 U19110 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21644), .ZN(n15553) );
  INV_X1 U19111 ( .A(n15520), .ZN(n20957) );
  XNOR2_X1 U19112 ( .A(n15521), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15525) );
  INV_X1 U19113 ( .A(n15525), .ZN(n15593) );
  NAND2_X1 U19114 ( .A1(n15522), .A2(n15593), .ZN(n15529) );
  NAND2_X1 U19115 ( .A1(n15524), .A2(n15523), .ZN(n15535) );
  NAND2_X1 U19116 ( .A1(n15535), .A2(n15525), .ZN(n15528) );
  XNOR2_X1 U19117 ( .A(n12209), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15526) );
  NAND2_X1 U19118 ( .A1(n15542), .A2(n15526), .ZN(n15527) );
  OAI211_X1 U19119 ( .C1(n15585), .C2(n15529), .A(n15528), .B(n15527), .ZN(
        n15530) );
  AOI21_X1 U19120 ( .B1(n20957), .B2(n15585), .A(n15530), .ZN(n15596) );
  INV_X1 U19121 ( .A(n15596), .ZN(n15531) );
  MUX2_X1 U19122 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15531), .S(
        n15552), .Z(n17504) );
  AOI22_X1 U19123 ( .A1(n15553), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n17504), .B2(n21644), .ZN(n15548) );
  NAND2_X1 U19124 ( .A1(n21327), .A2(n15585), .ZN(n15546) );
  NOR2_X1 U19125 ( .A1(n15533), .A2(n15532), .ZN(n15534) );
  NAND2_X1 U19126 ( .A1(n15535), .A2(n15534), .ZN(n15545) );
  AOI21_X1 U19127 ( .B1(n15521), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12471), .ZN(n15536) );
  NOR2_X1 U19128 ( .A1(n9782), .A2(n15536), .ZN(n15600) );
  OR3_X1 U19129 ( .A1(n15585), .A2(n15600), .A3(n15538), .ZN(n15544) );
  NAND2_X1 U19130 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15539) );
  NAND2_X1 U19131 ( .A1(n12471), .A2(n15539), .ZN(n15540) );
  NAND3_X1 U19132 ( .A1(n15542), .A2(n15541), .A3(n15540), .ZN(n15543) );
  NAND4_X1 U19133 ( .A1(n15546), .A2(n15545), .A3(n15544), .A4(n15543), .ZN(
        n15598) );
  MUX2_X1 U19134 ( .A(n15598), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17500), .Z(n17507) );
  AOI22_X1 U19135 ( .A1(n15553), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21644), .B2(n17507), .ZN(n15547) );
  NOR2_X1 U19136 ( .A1(n15548), .A2(n15547), .ZN(n17519) );
  INV_X1 U19137 ( .A(n17519), .ZN(n15549) );
  NOR2_X1 U19138 ( .A1(n15549), .A2(n12042), .ZN(n15560) );
  OR2_X1 U19139 ( .A1(n15550), .A2(n10611), .ZN(n15551) );
  XNOR2_X1 U19140 ( .A(n15551), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20942) );
  AOI21_X1 U19141 ( .B1(n17593), .B2(n20942), .A(n17500), .ZN(n15556) );
  OAI21_X1 U19142 ( .B1(n15552), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n21644), .ZN(n15555) );
  INV_X1 U19143 ( .A(n15553), .ZN(n15554) );
  OAI22_X1 U19144 ( .A1(n15556), .A2(n15555), .B1(n15554), .B2(n17596), .ZN(
        n17518) );
  NOR3_X1 U19145 ( .A1(n15560), .A2(n17518), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n15559) );
  NAND2_X1 U19146 ( .A1(n21645), .A2(n17529), .ZN(n21742) );
  INV_X1 U19147 ( .A(n21114), .ZN(n21206) );
  NOR3_X1 U19148 ( .A1(n15560), .A2(n17518), .A3(n17600), .ZN(n17528) );
  NAND2_X1 U19149 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21474), .ZN(n15578) );
  INV_X1 U19150 ( .A(n15578), .ZN(n15569) );
  OAI22_X1 U19151 ( .A1(n21139), .A2(n21579), .B1(n15561), .B2(n15569), .ZN(
        n15562) );
  OAI21_X1 U19152 ( .B1(n17528), .B2(n15562), .A(n21056), .ZN(n15563) );
  OAI21_X1 U19153 ( .B1(n21056), .B2(n21509), .A(n15563), .ZN(P1_U3478) );
  NAND2_X1 U19154 ( .A1(n9770), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15568) );
  NAND2_X1 U19155 ( .A1(n15568), .A2(n21517), .ZN(n15567) );
  NOR2_X1 U19156 ( .A1(n9770), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15565) );
  OAI22_X1 U19157 ( .A1(n15567), .A2(n15565), .B1(n21384), .B2(n15569), .ZN(
        n15566) );
  MUX2_X1 U19158 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15566), .S(
        n21056), .Z(P1_U3477) );
  NOR2_X1 U19159 ( .A1(n15574), .A2(n21579), .ZN(n21228) );
  NOR2_X1 U19160 ( .A1(n21228), .A2(n21430), .ZN(n21297) );
  AOI21_X1 U19161 ( .B1(n13145), .B2(n15568), .A(n21297), .ZN(n15571) );
  NOR2_X1 U19162 ( .A1(n15520), .A2(n15569), .ZN(n15570) );
  OAI21_X1 U19163 ( .B1(n15571), .B2(n15570), .A(n21056), .ZN(n15572) );
  OAI21_X1 U19164 ( .B1(n21056), .B2(n21389), .A(n15572), .ZN(P1_U3476) );
  NAND2_X1 U19165 ( .A1(n21517), .A2(n21880), .ZN(n21464) );
  MUX2_X1 U19166 ( .A(n21539), .B(n21303), .S(n9770), .Z(n15577) );
  OAI21_X1 U19167 ( .B1(n21381), .B2(n15577), .A(n15576), .ZN(n15580) );
  NAND2_X1 U19168 ( .A1(n21327), .A2(n15578), .ZN(n15579) );
  OAI211_X1 U19169 ( .C1(n15573), .C2(n21464), .A(n15580), .B(n15579), .ZN(
        n15581) );
  MUX2_X1 U19170 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15581), .S(
        n21056), .Z(P1_U3475) );
  NOR2_X1 U19171 ( .A1(n12042), .A2(n15521), .ZN(n15588) );
  INV_X1 U19172 ( .A(n15588), .ZN(n15583) );
  OAI22_X1 U19173 ( .A1(n17497), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n15583), .B2(n15582), .ZN(n15584) );
  AOI21_X1 U19174 ( .B1(n21540), .B2(n15585), .A(n15584), .ZN(n17499) );
  INV_X1 U19175 ( .A(n15599), .ZN(n15594) );
  NOR2_X1 U19176 ( .A1(n21644), .A2(n15586), .ZN(n15592) );
  AOI22_X1 U19177 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n21045), .B2(n14503), .ZN(
        n15591) );
  INV_X1 U19178 ( .A(n15591), .ZN(n15587) );
  AOI22_X1 U19179 ( .A1(n15594), .A2(n15588), .B1(n15592), .B2(n15587), .ZN(
        n15589) );
  OAI21_X1 U19180 ( .B1(n17499), .B2(n15601), .A(n15589), .ZN(n15590) );
  MUX2_X1 U19181 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15590), .S(
        n17597), .Z(P1_U3473) );
  AOI22_X1 U19182 ( .A1(n15594), .A2(n15593), .B1(n15592), .B2(n15591), .ZN(
        n15595) );
  OAI21_X1 U19183 ( .B1(n15596), .B2(n15601), .A(n15595), .ZN(n15597) );
  MUX2_X1 U19184 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15597), .S(
        n17597), .Z(P1_U3472) );
  INV_X1 U19185 ( .A(n15598), .ZN(n15602) );
  OAI22_X1 U19186 ( .A1(n15602), .A2(n15601), .B1(n15600), .B2(n15599), .ZN(
        n15603) );
  MUX2_X1 U19187 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15603), .S(
        n17597), .Z(P1_U3469) );
  INV_X1 U19188 ( .A(n21139), .ZN(n15604) );
  OAI21_X1 U19189 ( .B1(n21135), .B2(n21638), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15605) );
  NAND2_X1 U19190 ( .A1(n15605), .A2(n21517), .ZN(n15613) );
  OR2_X1 U19191 ( .A1(n21327), .A2(n20957), .ZN(n21142) );
  NAND2_X1 U19192 ( .A1(n21173), .A2(n21384), .ZN(n15608) );
  NOR2_X1 U19193 ( .A1(n15609), .A2(n21647), .ZN(n21388) );
  INV_X1 U19194 ( .A(n21388), .ZN(n21329) );
  INV_X1 U19195 ( .A(n21328), .ZN(n15606) );
  NAND2_X1 U19196 ( .A1(n15606), .A2(n21386), .ZN(n21203) );
  INV_X1 U19197 ( .A(n21110), .ZN(n15620) );
  INV_X1 U19198 ( .A(n21584), .ZN(n21477) );
  INV_X1 U19199 ( .A(n15608), .ZN(n15612) );
  NAND3_X1 U19200 ( .A1(n21385), .A2(n21389), .A3(n21468), .ZN(n21113) );
  NOR2_X1 U19201 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21113), .ZN(
        n21107) );
  INV_X1 U19202 ( .A(n21107), .ZN(n21090) );
  NAND2_X1 U19203 ( .A1(n15609), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21541) );
  NAND2_X1 U19204 ( .A1(n21114), .A2(n21541), .ZN(n21330) );
  AOI21_X1 U19205 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21090), .A(n21330), 
        .ZN(n15611) );
  NAND2_X1 U19206 ( .A1(n21203), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15610) );
  OAI211_X1 U19207 ( .C1(n15613), .C2(n15612), .A(n15611), .B(n15610), .ZN(
        n21058) );
  INV_X1 U19208 ( .A(DATAI_16_), .ZN(n15616) );
  OAI22_X1 U19209 ( .A1(n15616), .A2(n21104), .B1(n22004), .B2(n21102), .ZN(
        n21591) );
  INV_X1 U19210 ( .A(n21591), .ZN(n21552) );
  INV_X1 U19211 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17660) );
  INV_X1 U19212 ( .A(DATAI_24_), .ZN(n21904) );
  OAI22_X2 U19213 ( .A1(n17660), .A2(n21102), .B1(n21904), .B2(n21104), .ZN(
        n21549) );
  AOI22_X1 U19214 ( .A1(n21638), .A2(n21549), .B1(n21583), .B2(n21107), .ZN(
        n15617) );
  OAI21_X1 U19215 ( .B1(n21132), .B2(n21552), .A(n15617), .ZN(n15618) );
  AOI21_X1 U19216 ( .B1(n21058), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n15618), .ZN(n15619) );
  OAI21_X1 U19217 ( .B1(n15620), .B2(n21477), .A(n15619), .ZN(P1_U3033) );
  NOR2_X1 U19218 ( .A1(n15637), .A2(n15621), .ZN(n15622) );
  OAI21_X1 U19219 ( .B1(n15624), .B2(n15625), .A(n13002), .ZN(n16970) );
  INV_X1 U19220 ( .A(n16970), .ZN(n15635) );
  AOI22_X1 U19221 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_27__SCAN_IN), .ZN(n15627) );
  NAND2_X1 U19222 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15626) );
  OAI211_X1 U19223 ( .C1(n15628), .C2(n20053), .A(n15627), .B(n15626), .ZN(
        n15634) );
  INV_X1 U19224 ( .A(n15629), .ZN(n15630) );
  OAI21_X1 U19225 ( .B1(n15630), .B2(n16667), .A(n15999), .ZN(n15632) );
  INV_X1 U19226 ( .A(n13067), .ZN(n15631) );
  AOI21_X1 U19227 ( .B1(n15740), .B2(n15632), .A(n15631), .ZN(n15633) );
  AOI211_X1 U19228 ( .C1(n20040), .C2(n15635), .A(n15634), .B(n15633), .ZN(
        n15636) );
  OAI21_X1 U19229 ( .B1(n16665), .B2(n20066), .A(n15636), .ZN(P2_U2828) );
  AOI21_X1 U19230 ( .B1(n15638), .B2(n15659), .A(n15637), .ZN(n16984) );
  INV_X1 U19231 ( .A(n16984), .ZN(n16681) );
  NOR2_X1 U19232 ( .A1(n15640), .A2(n15641), .ZN(n15642) );
  OR2_X1 U19233 ( .A1(n15624), .A2(n15642), .ZN(n16991) );
  INV_X1 U19234 ( .A(n16991), .ZN(n15652) );
  INV_X1 U19235 ( .A(n16678), .ZN(n15644) );
  AOI21_X1 U19236 ( .B1(n15643), .B2(n15644), .A(n20062), .ZN(n15645) );
  OAI21_X1 U19237 ( .B1(n15645), .B2(n20038), .A(n15629), .ZN(n15650) );
  AOI22_X1 U19238 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_26__SCAN_IN), .ZN(n15649) );
  NAND2_X1 U19239 ( .A1(n15646), .A2(n16003), .ZN(n15648) );
  NAND2_X1 U19240 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15647) );
  NAND4_X1 U19241 ( .A1(n15650), .A2(n15649), .A3(n15648), .A4(n15647), .ZN(
        n15651) );
  AOI21_X1 U19242 ( .B1(n15652), .B2(n20040), .A(n15651), .ZN(n15653) );
  OAI21_X1 U19243 ( .B1(n16681), .B2(n20066), .A(n15653), .ZN(P2_U2829) );
  AND2_X1 U19244 ( .A1(n15654), .A2(n15655), .ZN(n15656) );
  OR2_X1 U19245 ( .A1(n15656), .A2(n15640), .ZN(n17003) );
  INV_X1 U19246 ( .A(n15659), .ZN(n15660) );
  AOI21_X1 U19247 ( .B1(n15661), .B2(n15658), .A(n15660), .ZN(n16995) );
  NAND2_X1 U19248 ( .A1(n16995), .A2(n20041), .ZN(n15673) );
  XOR2_X1 U19249 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n15662), .Z(n15671) );
  AOI22_X1 U19250 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_25__SCAN_IN), .ZN(n15663) );
  OAI21_X1 U19251 ( .B1(n20073), .B2(n15664), .A(n15663), .ZN(n15670) );
  INV_X1 U19252 ( .A(n15665), .ZN(n15666) );
  OAI21_X1 U19253 ( .B1(n15666), .B2(n16690), .A(n15999), .ZN(n15668) );
  INV_X1 U19254 ( .A(n15643), .ZN(n15667) );
  AOI21_X1 U19255 ( .B1(n15740), .B2(n15668), .A(n15667), .ZN(n15669) );
  AOI211_X1 U19256 ( .C1(n16003), .C2(n15671), .A(n15670), .B(n15669), .ZN(
        n15672) );
  OAI211_X1 U19257 ( .C1(n20065), .C2(n17003), .A(n15673), .B(n15672), .ZN(
        P2_U2830) );
  INV_X1 U19258 ( .A(n15658), .ZN(n15675) );
  AOI21_X1 U19259 ( .B1(n15676), .B2(n15674), .A(n15675), .ZN(n17008) );
  NAND2_X1 U19260 ( .A1(n15677), .A2(n15678), .ZN(n15679) );
  NAND2_X1 U19261 ( .A1(n15654), .A2(n15679), .ZN(n17014) );
  AOI22_X1 U19262 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_24__SCAN_IN), .ZN(n15681) );
  NAND2_X1 U19263 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15680) );
  OAI211_X1 U19264 ( .C1(n15682), .C2(n20053), .A(n15681), .B(n15680), .ZN(
        n15683) );
  INV_X1 U19265 ( .A(n15683), .ZN(n15688) );
  INV_X1 U19266 ( .A(n16703), .ZN(n15685) );
  AOI21_X1 U19267 ( .B1(n15684), .B2(n15685), .A(n20062), .ZN(n15686) );
  OAI21_X1 U19268 ( .B1(n15686), .B2(n20038), .A(n15665), .ZN(n15687) );
  OAI211_X1 U19269 ( .C1(n17014), .C2(n20065), .A(n15688), .B(n15687), .ZN(
        n15689) );
  AOI21_X1 U19270 ( .B1(n17008), .B2(n20041), .A(n15689), .ZN(n15690) );
  INV_X1 U19271 ( .A(n15690), .ZN(P2_U2831) );
  OR2_X1 U19272 ( .A1(n15691), .A2(n15692), .ZN(n15693) );
  NAND2_X1 U19273 ( .A1(n15677), .A2(n15693), .ZN(n17023) );
  OR2_X1 U19274 ( .A1(n15694), .A2(n15695), .ZN(n15696) );
  AND2_X1 U19275 ( .A1(n15674), .A2(n15696), .ZN(n17028) );
  NAND2_X1 U19276 ( .A1(n17028), .A2(n20041), .ZN(n15706) );
  AOI22_X1 U19277 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_23__SCAN_IN), .ZN(n15697) );
  OAI21_X1 U19278 ( .B1(n20073), .B2(n15698), .A(n15697), .ZN(n15703) );
  INV_X1 U19279 ( .A(n15699), .ZN(n15716) );
  OAI21_X1 U19280 ( .B1(n15716), .B2(n16708), .A(n15999), .ZN(n15701) );
  INV_X1 U19281 ( .A(n15684), .ZN(n15700) );
  AOI21_X1 U19282 ( .B1(n15740), .B2(n15701), .A(n15700), .ZN(n15702) );
  AOI211_X1 U19283 ( .C1(n16003), .C2(n15704), .A(n15703), .B(n15702), .ZN(
        n15705) );
  OAI211_X1 U19284 ( .C1(n20065), .C2(n17023), .A(n15706), .B(n15705), .ZN(
        P2_U2832) );
  NOR2_X1 U19285 ( .A1(n15707), .A2(n15708), .ZN(n15709) );
  OR2_X1 U19286 ( .A1(n15694), .A2(n15709), .ZN(n16716) );
  NOR2_X1 U19287 ( .A1(n15722), .A2(n15710), .ZN(n15711) );
  OR2_X1 U19288 ( .A1(n15691), .A2(n15711), .ZN(n17036) );
  INV_X1 U19289 ( .A(n17036), .ZN(n15720) );
  AOI22_X1 U19290 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_22__SCAN_IN), .ZN(n15713) );
  NAND2_X1 U19291 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15712) );
  OAI211_X1 U19292 ( .C1(n15714), .C2(n20053), .A(n15713), .B(n15712), .ZN(
        n15719) );
  INV_X1 U19293 ( .A(n15715), .ZN(n15731) );
  OAI21_X1 U19294 ( .B1(n15731), .B2(n16719), .A(n15999), .ZN(n15717) );
  AOI21_X1 U19295 ( .B1(n15740), .B2(n15717), .A(n15716), .ZN(n15718) );
  AOI211_X1 U19296 ( .C1(n15720), .C2(n20040), .A(n15719), .B(n15718), .ZN(
        n15721) );
  OAI21_X1 U19297 ( .B1(n16716), .B2(n20066), .A(n15721), .ZN(P2_U2833) );
  INV_X1 U19298 ( .A(n15722), .ZN(n15726) );
  NAND2_X1 U19299 ( .A1(n15724), .A2(n15723), .ZN(n15725) );
  NAND2_X1 U19300 ( .A1(n15726), .A2(n15725), .ZN(n17052) );
  AOI21_X1 U19301 ( .B1(n15727), .B2(n12011), .A(n15707), .ZN(n17043) );
  NAND2_X1 U19302 ( .A1(n17043), .A2(n20041), .ZN(n15737) );
  INV_X1 U19303 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15729) );
  AOI22_X1 U19304 ( .A1(P2_REIP_REG_21__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_21__SCAN_IN), .ZN(n15728) );
  OAI21_X1 U19305 ( .B1(n20073), .B2(n15729), .A(n15728), .ZN(n15734) );
  INV_X1 U19306 ( .A(n15730), .ZN(n15744) );
  OAI21_X1 U19307 ( .B1(n15744), .B2(n16738), .A(n15999), .ZN(n15732) );
  AOI21_X1 U19308 ( .B1(n15740), .B2(n15732), .A(n15731), .ZN(n15733) );
  AOI211_X1 U19309 ( .C1(n16003), .C2(n15735), .A(n15734), .B(n15733), .ZN(
        n15736) );
  OAI211_X1 U19310 ( .C1(n20065), .C2(n17052), .A(n15737), .B(n15736), .ZN(
        P2_U2834) );
  NAND2_X1 U19311 ( .A1(n16438), .A2(n20041), .ZN(n15750) );
  AOI22_X1 U19312 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_20__SCAN_IN), .ZN(n15738) );
  OAI21_X1 U19313 ( .B1(n20073), .B2(n15739), .A(n15738), .ZN(n15747) );
  INV_X1 U19314 ( .A(n15741), .ZN(n15743) );
  OAI21_X1 U19315 ( .B1(n15743), .B2(n15742), .A(n15999), .ZN(n15745) );
  AOI21_X1 U19316 ( .B1(n15740), .B2(n15745), .A(n15744), .ZN(n15746) );
  AOI211_X1 U19317 ( .C1(n16003), .C2(n15748), .A(n15747), .B(n15746), .ZN(
        n15749) );
  OAI211_X1 U19318 ( .C1(n20065), .C2(n16591), .A(n15750), .B(n15749), .ZN(
        P2_U2835) );
  OR2_X1 U19319 ( .A1(n15751), .A2(n15752), .ZN(n15753) );
  NAND2_X1 U19320 ( .A1(n12010), .A2(n15753), .ZN(n17065) );
  INV_X1 U19321 ( .A(n15756), .ZN(n15757) );
  XNOR2_X1 U19322 ( .A(n15755), .B(n15757), .ZN(n17063) );
  AOI21_X1 U19323 ( .B1(n15758), .B2(n10655), .A(n20062), .ZN(n15759) );
  OAI21_X1 U19324 ( .B1(n20038), .B2(n15759), .A(n15741), .ZN(n15763) );
  AOI21_X1 U19325 ( .B1(n20032), .B2(P2_EBX_REG_19__SCAN_IN), .A(n20033), .ZN(
        n15760) );
  OAI21_X1 U19326 ( .B1(n20760), .B2(n16009), .A(n15760), .ZN(n15761) );
  AOI21_X1 U19327 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20031), .A(
        n15761), .ZN(n15762) );
  OAI211_X1 U19328 ( .C1(n20053), .C2(n15764), .A(n15763), .B(n15762), .ZN(
        n15765) );
  AOI21_X1 U19329 ( .B1(n17063), .B2(n20040), .A(n15765), .ZN(n15766) );
  OAI21_X1 U19330 ( .B1(n17065), .B2(n20066), .A(n15766), .ZN(P2_U2836) );
  AOI21_X1 U19331 ( .B1(n15768), .B2(n15767), .A(n15751), .ZN(n17076) );
  INV_X1 U19332 ( .A(n17076), .ZN(n16455) );
  AOI21_X1 U19333 ( .B1(n15770), .B2(n15769), .A(n15755), .ZN(n16600) );
  AOI21_X1 U19334 ( .B1(n20032), .B2(P2_EBX_REG_18__SCAN_IN), .A(n20033), .ZN(
        n15771) );
  OAI21_X1 U19335 ( .B1(n15772), .B2(n16009), .A(n15771), .ZN(n15773) );
  AOI21_X1 U19336 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20031), .A(
        n15773), .ZN(n15774) );
  OAI21_X1 U19337 ( .B1(n15775), .B2(n20053), .A(n15774), .ZN(n15780) );
  INV_X1 U19338 ( .A(n15777), .ZN(n15776) );
  NOR2_X1 U19339 ( .A1(n16015), .A2(n15776), .ZN(n15787) );
  OAI21_X1 U19340 ( .B1(n20062), .B2(n15777), .A(n15740), .ZN(n15778) );
  MUX2_X1 U19341 ( .A(n15787), .B(n15778), .S(n16759), .Z(n15779) );
  AOI211_X1 U19342 ( .C1(n16600), .C2(n20040), .A(n15780), .B(n15779), .ZN(
        n15781) );
  OAI21_X1 U19343 ( .B1(n16455), .B2(n20066), .A(n15781), .ZN(P2_U2837) );
  INV_X1 U19344 ( .A(n15767), .ZN(n15783) );
  AOI21_X1 U19345 ( .B1(n15784), .B2(n15782), .A(n15783), .ZN(n17083) );
  OAI21_X1 U19346 ( .B1(n15786), .B2(n10805), .A(n15769), .ZN(n17085) );
  INV_X1 U19347 ( .A(n17085), .ZN(n15796) );
  OAI21_X1 U19348 ( .B1(n15788), .B2(n16767), .A(n15787), .ZN(n15794) );
  NAND2_X1 U19349 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15790) );
  AOI21_X1 U19350 ( .B1(n20032), .B2(P2_EBX_REG_17__SCAN_IN), .A(n20033), .ZN(
        n15789) );
  OAI211_X1 U19351 ( .C1(n16009), .C2(n20757), .A(n15790), .B(n15789), .ZN(
        n15791) );
  AOI21_X1 U19352 ( .B1(n15792), .B2(n16003), .A(n15791), .ZN(n15793) );
  OAI211_X1 U19353 ( .C1(n15740), .C2(n16767), .A(n15794), .B(n15793), .ZN(
        n15795) );
  AOI21_X1 U19354 ( .B1(n15796), .B2(n20040), .A(n15795), .ZN(n15797) );
  OAI21_X1 U19355 ( .B1(n17089), .B2(n20066), .A(n15797), .ZN(P2_U2838) );
  OR2_X1 U19356 ( .A1(n15798), .A2(n15799), .ZN(n15800) );
  NAND2_X1 U19357 ( .A1(n15782), .A2(n15800), .ZN(n17101) );
  INV_X1 U19358 ( .A(n15801), .ZN(n15808) );
  NAND2_X1 U19359 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15803) );
  AOI21_X1 U19360 ( .B1(n20032), .B2(P2_EBX_REG_16__SCAN_IN), .A(n20033), .ZN(
        n15802) );
  OAI211_X1 U19361 ( .C1(n16009), .C2(n20755), .A(n15803), .B(n15802), .ZN(
        n15807) );
  OAI21_X1 U19362 ( .B1(n20062), .B2(n10274), .A(n15740), .ZN(n15805) );
  NOR2_X1 U19363 ( .A1(n16015), .A2(n15804), .ZN(n20044) );
  MUX2_X1 U19364 ( .A(n15805), .B(n20044), .S(n16773), .Z(n15806) );
  AOI211_X1 U19365 ( .C1(n16003), .C2(n15808), .A(n15807), .B(n15806), .ZN(
        n15812) );
  AOI21_X1 U19366 ( .B1(n15810), .B2(n15809), .A(n15786), .ZN(n17099) );
  NAND2_X1 U19367 ( .A1(n17099), .A2(n20040), .ZN(n15811) );
  OAI211_X1 U19368 ( .C1(n20066), .C2(n17101), .A(n15812), .B(n15811), .ZN(
        P2_U2839) );
  NOR2_X1 U19369 ( .A1(n16009), .A2(n15813), .ZN(n15814) );
  AOI211_X1 U19370 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n20032), .A(n20033), .B(
        n15814), .ZN(n15815) );
  OAI21_X1 U19371 ( .B1(n16800), .B2(n20073), .A(n15815), .ZN(n15820) );
  INV_X1 U19372 ( .A(n15817), .ZN(n15816) );
  NOR2_X1 U19373 ( .A1(n16015), .A2(n15816), .ZN(n15832) );
  OAI21_X1 U19374 ( .B1(n20062), .B2(n15817), .A(n15740), .ZN(n15818) );
  MUX2_X1 U19375 ( .A(n15832), .B(n15818), .S(n16798), .Z(n15819) );
  AOI211_X1 U19376 ( .C1(n16003), .C2(n15821), .A(n15820), .B(n15819), .ZN(
        n15828) );
  INV_X1 U19377 ( .A(n15824), .ZN(n15825) );
  AOI21_X1 U19378 ( .B1(n15826), .B2(n15822), .A(n15825), .ZN(n17119) );
  NAND2_X1 U19379 ( .A1(n17119), .A2(n20041), .ZN(n15827) );
  OAI211_X1 U19380 ( .C1(n20065), .C2(n17111), .A(n15828), .B(n15827), .ZN(
        P2_U2841) );
  NAND2_X1 U19381 ( .A1(n15829), .A2(n15830), .ZN(n15831) );
  NAND2_X1 U19382 ( .A1(n15822), .A2(n15831), .ZN(n17132) );
  OAI21_X1 U19383 ( .B1(n15833), .B2(n16810), .A(n15832), .ZN(n15839) );
  NAND2_X1 U19384 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15835) );
  AOI21_X1 U19385 ( .B1(n20032), .B2(P2_EBX_REG_13__SCAN_IN), .A(n20033), .ZN(
        n15834) );
  OAI211_X1 U19386 ( .C1(n16809), .C2(n16009), .A(n15835), .B(n15834), .ZN(
        n15836) );
  AOI21_X1 U19387 ( .B1(n15837), .B2(n16003), .A(n15836), .ZN(n15838) );
  OAI211_X1 U19388 ( .C1(n15740), .C2(n16810), .A(n15839), .B(n15838), .ZN(
        n15840) );
  AOI21_X1 U19389 ( .B1(n17129), .B2(n20040), .A(n15840), .ZN(n15841) );
  OAI21_X1 U19390 ( .B1(n17132), .B2(n20066), .A(n15841), .ZN(P2_U2842) );
  OR2_X1 U19391 ( .A1(n15842), .A2(n15843), .ZN(n15844) );
  AND2_X1 U19392 ( .A1(n15829), .A2(n15844), .ZN(n17146) );
  INV_X1 U19393 ( .A(n17146), .ZN(n16486) );
  AOI21_X1 U19394 ( .B1(n15999), .B2(n15845), .A(n20038), .ZN(n15848) );
  INV_X1 U19395 ( .A(n15845), .ZN(n15846) );
  NAND2_X1 U19396 ( .A1(n15975), .A2(n15846), .ZN(n15847) );
  MUX2_X1 U19397 ( .A(n15848), .B(n15847), .S(n16819), .Z(n15856) );
  INV_X1 U19398 ( .A(n20032), .ZN(n20052) );
  OAI21_X1 U19399 ( .B1(n20052), .B2(n16485), .A(n20051), .ZN(n15849) );
  AOI21_X1 U19400 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n20057), .A(n15849), 
        .ZN(n15850) );
  OAI21_X1 U19401 ( .B1(n15851), .B2(n20073), .A(n15850), .ZN(n15853) );
  NOR2_X1 U19402 ( .A1(n17139), .A2(n20065), .ZN(n15852) );
  AOI211_X1 U19403 ( .C1(n16003), .C2(n15854), .A(n15853), .B(n15852), .ZN(
        n15855) );
  OAI211_X1 U19404 ( .C1(n20066), .C2(n16486), .A(n15856), .B(n15855), .ZN(
        P2_U2843) );
  NOR2_X1 U19405 ( .A1(n15857), .A2(n15858), .ZN(n15859) );
  OR2_X1 U19406 ( .A1(n15842), .A2(n15859), .ZN(n17150) );
  NAND2_X1 U19407 ( .A1(n15975), .A2(n15860), .ZN(n15863) );
  INV_X1 U19408 ( .A(n15860), .ZN(n15861) );
  AOI21_X1 U19409 ( .B1(n15999), .B2(n15861), .A(n20038), .ZN(n15862) );
  MUX2_X1 U19410 ( .A(n15863), .B(n15862), .S(n16833), .Z(n15870) );
  OAI21_X1 U19411 ( .B1(n20052), .B2(n11774), .A(n20051), .ZN(n15864) );
  AOI21_X1 U19412 ( .B1(P2_REIP_REG_11__SCAN_IN), .B2(n20057), .A(n15864), 
        .ZN(n15865) );
  OAI21_X1 U19413 ( .B1(n10659), .B2(n20073), .A(n15865), .ZN(n15867) );
  NOR2_X1 U19414 ( .A1(n17151), .A2(n20065), .ZN(n15866) );
  AOI211_X1 U19415 ( .C1(n16003), .C2(n15868), .A(n15867), .B(n15866), .ZN(
        n15869) );
  OAI211_X1 U19416 ( .C1(n20066), .C2(n17150), .A(n15870), .B(n15869), .ZN(
        P2_U2844) );
  NAND2_X1 U19417 ( .A1(n15975), .A2(n15871), .ZN(n15874) );
  OR2_X1 U19418 ( .A1(n15871), .A2(n20062), .ZN(n15872) );
  AND2_X1 U19419 ( .A1(n15740), .A2(n15872), .ZN(n15873) );
  MUX2_X1 U19420 ( .A(n15874), .B(n15873), .S(n16845), .Z(n15886) );
  AND2_X1 U19421 ( .A1(n14351), .A2(n15875), .ZN(n15876) );
  OR2_X1 U19422 ( .A1(n15876), .A2(n15857), .ZN(n20074) );
  INV_X1 U19423 ( .A(n15877), .ZN(n15881) );
  NAND2_X1 U19424 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15879) );
  AOI21_X1 U19425 ( .B1(n20032), .B2(P2_EBX_REG_10__SCAN_IN), .A(n20033), .ZN(
        n15878) );
  OAI211_X1 U19426 ( .C1(n16009), .C2(n16841), .A(n15879), .B(n15878), .ZN(
        n15880) );
  AOI21_X1 U19427 ( .B1(n15881), .B2(n16003), .A(n15880), .ZN(n15883) );
  NAND2_X1 U19428 ( .A1(n17171), .A2(n20040), .ZN(n15882) );
  OAI211_X1 U19429 ( .C1(n20074), .C2(n20066), .A(n15883), .B(n15882), .ZN(
        n15884) );
  INV_X1 U19430 ( .A(n15884), .ZN(n15885) );
  NAND2_X1 U19431 ( .A1(n15886), .A2(n15885), .ZN(P2_U2845) );
  NOR2_X1 U19432 ( .A1(n10279), .A2(n15887), .ZN(n15888) );
  XOR2_X1 U19433 ( .A(n16861), .B(n15888), .Z(n15896) );
  NAND2_X1 U19434 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15890) );
  AOI21_X1 U19435 ( .B1(n20032), .B2(P2_EBX_REG_9__SCAN_IN), .A(n20033), .ZN(
        n15889) );
  OAI211_X1 U19436 ( .C1(n16009), .C2(n20745), .A(n15890), .B(n15889), .ZN(
        n15891) );
  AOI21_X1 U19437 ( .B1(n15892), .B2(n16003), .A(n15891), .ZN(n15893) );
  OAI21_X1 U19438 ( .B1(n17181), .B2(n20065), .A(n15893), .ZN(n15894) );
  AOI21_X1 U19439 ( .B1(n17183), .B2(n20041), .A(n15894), .ZN(n15895) );
  OAI21_X1 U19440 ( .B1(n15896), .B2(n20062), .A(n15895), .ZN(P2_U2846) );
  NAND2_X1 U19441 ( .A1(n15898), .A2(n15999), .ZN(n15897) );
  AND2_X1 U19442 ( .A1(n15740), .A2(n15897), .ZN(n15901) );
  INV_X1 U19443 ( .A(n15898), .ZN(n15899) );
  NAND2_X1 U19444 ( .A1(n15975), .A2(n15899), .ZN(n15900) );
  MUX2_X1 U19445 ( .A(n15901), .B(n15900), .S(n16878), .Z(n15914) );
  OR2_X1 U19446 ( .A1(n15902), .A2(n15903), .ZN(n15904) );
  NAND2_X1 U19447 ( .A1(n14352), .A2(n15904), .ZN(n17187) );
  INV_X1 U19448 ( .A(n17187), .ZN(n15912) );
  INV_X1 U19449 ( .A(n15905), .ZN(n15909) );
  INV_X1 U19450 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21984) );
  NAND2_X1 U19451 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15907) );
  AOI21_X1 U19452 ( .B1(n20032), .B2(P2_EBX_REG_8__SCAN_IN), .A(n20033), .ZN(
        n15906) );
  OAI211_X1 U19453 ( .C1(n16009), .C2(n20743), .A(n15907), .B(n15906), .ZN(
        n15908) );
  AOI21_X1 U19454 ( .B1(n15909), .B2(n16003), .A(n15908), .ZN(n15910) );
  OAI21_X1 U19455 ( .B1(n17195), .B2(n20065), .A(n15910), .ZN(n15911) );
  AOI21_X1 U19456 ( .B1(n15912), .B2(n20041), .A(n15911), .ZN(n15913) );
  NAND2_X1 U19457 ( .A1(n15914), .A2(n15913), .ZN(P2_U2847) );
  NAND2_X1 U19458 ( .A1(n15975), .A2(n15915), .ZN(n15918) );
  INV_X1 U19459 ( .A(n15915), .ZN(n20063) );
  NAND2_X1 U19460 ( .A1(n20063), .A2(n15999), .ZN(n15916) );
  AND2_X1 U19461 ( .A1(n15740), .A2(n15916), .ZN(n15917) );
  MUX2_X1 U19462 ( .A(n15918), .B(n15917), .S(n16889), .Z(n15929) );
  AND2_X1 U19463 ( .A1(n14340), .A2(n15919), .ZN(n15920) );
  OR2_X1 U19464 ( .A1(n15920), .A2(n15902), .ZN(n17208) );
  NAND2_X1 U19465 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15922) );
  AOI21_X1 U19466 ( .B1(n20032), .B2(P2_EBX_REG_7__SCAN_IN), .A(n20033), .ZN(
        n15921) );
  OAI211_X1 U19467 ( .C1(n16009), .C2(n20741), .A(n15922), .B(n15921), .ZN(
        n15923) );
  AOI21_X1 U19468 ( .B1(n15924), .B2(n16003), .A(n15923), .ZN(n15926) );
  NAND2_X1 U19469 ( .A1(n17206), .A2(n20040), .ZN(n15925) );
  OAI211_X1 U19470 ( .C1(n17208), .C2(n20066), .A(n15926), .B(n15925), .ZN(
        n15927) );
  INV_X1 U19471 ( .A(n15927), .ZN(n15928) );
  NAND2_X1 U19472 ( .A1(n15929), .A2(n15928), .ZN(P2_U2848) );
  NOR2_X1 U19473 ( .A1(n10279), .A2(n15930), .ZN(n15931) );
  XOR2_X1 U19474 ( .A(n16906), .B(n15931), .Z(n15941) );
  XNOR2_X1 U19475 ( .A(n15932), .B(n15933), .ZN(n17233) );
  NAND2_X1 U19476 ( .A1(n20032), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n15934) );
  OAI211_X1 U19477 ( .C1(n16904), .C2(n16009), .A(n15934), .B(n20051), .ZN(
        n15937) );
  NOR2_X1 U19478 ( .A1(n15935), .A2(n20053), .ZN(n15936) );
  AOI211_X1 U19479 ( .C1(n20031), .C2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n15937), .B(n15936), .ZN(n15938) );
  OAI21_X1 U19480 ( .B1(n17233), .B2(n20065), .A(n15938), .ZN(n15939) );
  AOI21_X1 U19481 ( .B1(n17238), .B2(n20041), .A(n15939), .ZN(n15940) );
  OAI21_X1 U19482 ( .B1(n15941), .B2(n20062), .A(n15940), .ZN(P2_U2850) );
  INV_X1 U19483 ( .A(n17242), .ZN(n15955) );
  NAND2_X1 U19484 ( .A1(n15961), .A2(n15943), .ZN(n15944) );
  NAND2_X1 U19485 ( .A1(n15932), .A2(n15944), .ZN(n20086) );
  NOR2_X1 U19486 ( .A1(n16916), .A2(n20053), .ZN(n15947) );
  INV_X1 U19487 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20738) );
  NAND2_X1 U19488 ( .A1(n20032), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n15945) );
  OAI211_X1 U19489 ( .C1(n20738), .C2(n16009), .A(n15945), .B(n20051), .ZN(
        n15946) );
  AOI211_X1 U19490 ( .C1(n20031), .C2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n15947), .B(n15946), .ZN(n15948) );
  OAI21_X1 U19491 ( .B1(n20086), .B2(n20065), .A(n15948), .ZN(n15954) );
  INV_X1 U19492 ( .A(n15950), .ZN(n15949) );
  NOR2_X1 U19493 ( .A1(n16015), .A2(n15949), .ZN(n15952) );
  OAI21_X1 U19494 ( .B1(n20062), .B2(n15950), .A(n15740), .ZN(n15951) );
  MUX2_X1 U19495 ( .A(n15952), .B(n15951), .S(n16923), .Z(n15953) );
  AOI211_X1 U19496 ( .C1(n15955), .C2(n20041), .A(n15954), .B(n15953), .ZN(
        n15956) );
  OAI21_X1 U19497 ( .B1(n16010), .B2(n20088), .A(n15956), .ZN(P2_U2851) );
  INV_X1 U19498 ( .A(n14213), .ZN(n15957) );
  NAND2_X1 U19499 ( .A1(n15959), .A2(n15958), .ZN(n15960) );
  NAND2_X1 U19500 ( .A1(n15961), .A2(n15960), .ZN(n17257) );
  NOR2_X1 U19501 ( .A1(n20053), .A2(n15962), .ZN(n15964) );
  INV_X1 U19502 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20736) );
  OAI22_X1 U19503 ( .A1(n20052), .A2(n21842), .B1(n20736), .B2(n16009), .ZN(
        n15963) );
  AOI211_X1 U19504 ( .C1(n20031), .C2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15964), .B(n15963), .ZN(n15965) );
  OAI21_X1 U19505 ( .B1(n17257), .B2(n20065), .A(n15965), .ZN(n15970) );
  OAI21_X1 U19506 ( .B1(n20062), .B2(n15966), .A(n15740), .ZN(n15968) );
  NOR2_X1 U19507 ( .A1(n16015), .A2(n10281), .ZN(n15967) );
  MUX2_X1 U19508 ( .A(n15968), .B(n15967), .S(n16932), .Z(n15969) );
  AOI211_X1 U19509 ( .C1(n20041), .C2(n15957), .A(n15970), .B(n15969), .ZN(
        n15971) );
  OAI21_X1 U19510 ( .B1(n16010), .B2(n20199), .A(n15971), .ZN(P2_U2852) );
  NAND2_X1 U19511 ( .A1(n15973), .A2(n15999), .ZN(n15972) );
  AND2_X1 U19512 ( .A1(n15740), .A2(n15972), .ZN(n15978) );
  INV_X1 U19513 ( .A(n15973), .ZN(n15974) );
  NAND2_X1 U19514 ( .A1(n15975), .A2(n15974), .ZN(n15977) );
  MUX2_X1 U19515 ( .A(n15978), .B(n15977), .S(n15976), .Z(n15988) );
  NAND2_X1 U19516 ( .A1(n16630), .A2(n20040), .ZN(n15984) );
  AOI22_X1 U19517 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n20057), .B1(n20032), 
        .B2(P2_EBX_REG_2__SCAN_IN), .ZN(n15983) );
  NAND2_X1 U19518 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15982) );
  INV_X1 U19519 ( .A(n15979), .ZN(n15980) );
  NAND2_X1 U19520 ( .A1(n16003), .A2(n15980), .ZN(n15981) );
  NAND4_X1 U19521 ( .A1(n15984), .A2(n15983), .A3(n15982), .A4(n15981), .ZN(
        n15985) );
  AOI21_X1 U19522 ( .B1(n15986), .B2(n20041), .A(n15985), .ZN(n15987) );
  OAI211_X1 U19523 ( .C1(n20817), .C2(n16010), .A(n15988), .B(n15987), .ZN(
        P2_U2853) );
  INV_X1 U19524 ( .A(n15989), .ZN(n16000) );
  AOI22_X1 U19525 ( .A1(n20032), .A2(P2_EBX_REG_1__SCAN_IN), .B1(n15990), .B2(
        n16003), .ZN(n15993) );
  NAND2_X1 U19526 ( .A1(n20031), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15992) );
  OAI211_X1 U19527 ( .C1(n16009), .C2(n20732), .A(n15993), .B(n15992), .ZN(
        n15996) );
  NOR2_X1 U19528 ( .A1(n15994), .A2(n20066), .ZN(n15995) );
  AOI211_X1 U19529 ( .C1(n20040), .C2(n20828), .A(n15996), .B(n15995), .ZN(
        n15997) );
  OAI21_X1 U19530 ( .B1(n20134), .B2(n16010), .A(n15997), .ZN(n15998) );
  AOI21_X1 U19531 ( .B1(n16000), .B2(n15999), .A(n15998), .ZN(n16001) );
  OAI21_X1 U19532 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n15740), .A(
        n16001), .ZN(P2_U2854) );
  INV_X1 U19533 ( .A(n16002), .ZN(n16016) );
  OAI21_X1 U19534 ( .B1(n20038), .B2(n20031), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16014) );
  AOI22_X1 U19535 ( .A1(n20040), .A2(n16005), .B1(n16004), .B2(n16003), .ZN(
        n16007) );
  NAND2_X1 U19536 ( .A1(n20032), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n16006) );
  OAI211_X1 U19537 ( .C1(n16009), .C2(n16008), .A(n16007), .B(n16006), .ZN(
        n16012) );
  NOR2_X1 U19538 ( .A1(n20133), .A2(n16010), .ZN(n16011) );
  AOI211_X1 U19539 ( .C1(n20041), .C2(n17281), .A(n16012), .B(n16011), .ZN(
        n16013) );
  OAI211_X1 U19540 ( .C1(n16016), .C2(n16015), .A(n16014), .B(n16013), .ZN(
        P2_U2855) );
  NAND2_X1 U19541 ( .A1(n16503), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n16018) );
  OAI21_X1 U19542 ( .B1(n16017), .B2(n16503), .A(n16018), .ZN(P2_U2856) );
  AND2_X1 U19543 ( .A1(n16484), .A2(n16479), .ZN(n16022) );
  NAND4_X1 U19544 ( .A1(n16022), .A2(n16489), .A3(n16477), .A4(n16021), .ZN(
        n16023) );
  NOR2_X1 U19545 ( .A1(n16024), .A2(n16023), .ZN(n16025) );
  OAI22_X1 U19546 ( .A1(n16225), .A2(n16028), .B1(n16229), .B2(n16027), .ZN(
        n16032) );
  OAI22_X1 U19547 ( .A1(n16221), .A2(n16030), .B1(n16228), .B2(n16029), .ZN(
        n16031) );
  NOR2_X1 U19548 ( .A1(n16032), .A2(n16031), .ZN(n16049) );
  AOI22_X1 U19549 ( .A1(n16203), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16036) );
  AOI22_X1 U19550 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16035) );
  NAND2_X1 U19551 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n16034) );
  NAND2_X1 U19552 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n16033) );
  NAND4_X1 U19553 ( .A1(n16036), .A2(n16035), .A3(n16034), .A4(n16033), .ZN(
        n16040) );
  INV_X1 U19554 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16037) );
  OAI22_X1 U19555 ( .A1(n16153), .A2(n16038), .B1(n11252), .B2(n16037), .ZN(
        n16039) );
  NOR2_X1 U19556 ( .A1(n16040), .A2(n16039), .ZN(n16048) );
  OAI22_X1 U19557 ( .A1(n16217), .A2(n16042), .B1(n16109), .B2(n16041), .ZN(
        n16046) );
  INV_X1 U19558 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16043) );
  OAI22_X1 U19559 ( .A1(n16215), .A2(n16044), .B1(n16219), .B2(n16043), .ZN(
        n16045) );
  NOR2_X1 U19560 ( .A1(n16046), .A2(n16045), .ZN(n16047) );
  NAND3_X1 U19561 ( .A1(n16049), .A2(n16048), .A3(n16047), .ZN(n16462) );
  OAI22_X1 U19562 ( .A1(n16225), .A2(n16051), .B1(n16229), .B2(n16050), .ZN(
        n16055) );
  OAI22_X1 U19563 ( .A1(n16221), .A2(n16053), .B1(n16228), .B2(n16052), .ZN(
        n16054) );
  NOR2_X1 U19564 ( .A1(n16055), .A2(n16054), .ZN(n16071) );
  AOI22_X1 U19565 ( .A1(n16203), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16059) );
  AOI22_X1 U19566 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16058) );
  NAND2_X1 U19567 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n16057) );
  NAND2_X1 U19568 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n16056) );
  NAND4_X1 U19569 ( .A1(n16059), .A2(n16058), .A3(n16057), .A4(n16056), .ZN(
        n16063) );
  OAI22_X1 U19570 ( .A1(n16153), .A2(n16061), .B1(n11252), .B2(n16060), .ZN(
        n16062) );
  NOR2_X1 U19571 ( .A1(n16063), .A2(n16062), .ZN(n16070) );
  OAI22_X1 U19572 ( .A1(n16217), .A2(n16064), .B1(n16109), .B2(n21861), .ZN(
        n16068) );
  OAI22_X1 U19573 ( .A1(n16215), .A2(n16066), .B1(n16219), .B2(n16065), .ZN(
        n16067) );
  NOR2_X1 U19574 ( .A1(n16068), .A2(n16067), .ZN(n16069) );
  NAND3_X1 U19575 ( .A1(n16071), .A2(n16070), .A3(n16069), .ZN(n16457) );
  NAND4_X1 U19576 ( .A1(n16462), .A2(n16456), .A3(n16457), .A4(n16472), .ZN(
        n16440) );
  OAI22_X1 U19577 ( .A1(n16072), .A2(n16229), .B1(n16225), .B2(n11545), .ZN(
        n16076) );
  OAI22_X1 U19578 ( .A1(n16074), .A2(n16228), .B1(n16221), .B2(n16073), .ZN(
        n16075) );
  NOR2_X1 U19579 ( .A1(n16076), .A2(n16075), .ZN(n16093) );
  AOI22_X1 U19580 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n16203), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16080) );
  AOI22_X1 U19581 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n16205), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U19582 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n16078) );
  NAND2_X1 U19583 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n16077) );
  NAND4_X1 U19584 ( .A1(n16080), .A2(n16079), .A3(n16078), .A4(n16077), .ZN(
        n16084) );
  OAI22_X1 U19585 ( .A1(n16082), .A2(n16153), .B1(n11252), .B2(n16081), .ZN(
        n16083) );
  NOR2_X1 U19586 ( .A1(n16084), .A2(n16083), .ZN(n16092) );
  OAI22_X1 U19587 ( .A1(n16086), .A2(n16109), .B1(n16217), .B2(n16085), .ZN(
        n16090) );
  INV_X1 U19588 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16088) );
  INV_X1 U19589 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16087) );
  OAI22_X1 U19590 ( .A1(n16088), .A2(n16215), .B1(n16219), .B2(n16087), .ZN(
        n16089) );
  NOR2_X1 U19591 ( .A1(n16090), .A2(n16089), .ZN(n16091) );
  NAND3_X1 U19592 ( .A1(n16093), .A2(n16092), .A3(n16091), .ZN(n16447) );
  OAI22_X1 U19593 ( .A1(n16095), .A2(n16229), .B1(n16225), .B2(n16094), .ZN(
        n16099) );
  OAI22_X1 U19594 ( .A1(n16097), .A2(n16228), .B1(n16221), .B2(n16096), .ZN(
        n16098) );
  NOR2_X1 U19595 ( .A1(n16099), .A2(n16098), .ZN(n16117) );
  AOI22_X1 U19596 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n16203), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16103) );
  AOI22_X1 U19597 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n16205), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16102) );
  NAND2_X1 U19598 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n16101) );
  NAND2_X1 U19599 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n16100) );
  NAND4_X1 U19600 ( .A1(n16103), .A2(n16102), .A3(n16101), .A4(n16100), .ZN(
        n16107) );
  OAI22_X1 U19601 ( .A1(n16105), .A2(n16153), .B1(n11252), .B2(n16104), .ZN(
        n16106) );
  NOR2_X1 U19602 ( .A1(n16107), .A2(n16106), .ZN(n16116) );
  OAI22_X1 U19603 ( .A1(n16110), .A2(n16109), .B1(n16217), .B2(n16108), .ZN(
        n16114) );
  INV_X1 U19604 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16112) );
  INV_X1 U19605 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16111) );
  OAI22_X1 U19606 ( .A1(n16112), .A2(n16215), .B1(n16219), .B2(n16111), .ZN(
        n16113) );
  NOR2_X1 U19607 ( .A1(n16114), .A2(n16113), .ZN(n16115) );
  NAND3_X1 U19608 ( .A1(n16117), .A2(n16116), .A3(n16115), .ZN(n16450) );
  OAI22_X1 U19609 ( .A1(n16119), .A2(n16229), .B1(n16225), .B2(n16118), .ZN(
        n16123) );
  OAI22_X1 U19610 ( .A1(n16121), .A2(n16228), .B1(n16221), .B2(n16120), .ZN(
        n16122) );
  NOR2_X1 U19611 ( .A1(n16123), .A2(n16122), .ZN(n16139) );
  AOI22_X1 U19612 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n16203), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16127) );
  AOI22_X1 U19613 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n16205), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16126) );
  NAND2_X1 U19614 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n16125) );
  NAND2_X1 U19615 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n16124) );
  NAND4_X1 U19616 ( .A1(n16127), .A2(n16126), .A3(n16125), .A4(n16124), .ZN(
        n16131) );
  OAI22_X1 U19617 ( .A1(n16129), .A2(n16153), .B1(n11252), .B2(n16128), .ZN(
        n16130) );
  NOR2_X1 U19618 ( .A1(n16131), .A2(n16130), .ZN(n16138) );
  OAI22_X1 U19619 ( .A1(n16133), .A2(n16109), .B1(n16217), .B2(n16132), .ZN(
        n16136) );
  INV_X1 U19620 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16134) );
  OAI22_X1 U19621 ( .A1(n16134), .A2(n16215), .B1(n16219), .B2(n21882), .ZN(
        n16135) );
  NOR2_X1 U19622 ( .A1(n16136), .A2(n16135), .ZN(n16137) );
  NAND3_X1 U19623 ( .A1(n16139), .A2(n16138), .A3(n16137), .ZN(n16441) );
  NAND3_X1 U19624 ( .A1(n16447), .A2(n16450), .A3(n16441), .ZN(n16140) );
  OAI22_X1 U19625 ( .A1(n16225), .A2(n16142), .B1(n16229), .B2(n16141), .ZN(
        n16146) );
  OAI22_X1 U19626 ( .A1(n16221), .A2(n16144), .B1(n16228), .B2(n16143), .ZN(
        n16145) );
  NOR2_X1 U19627 ( .A1(n16146), .A2(n16145), .ZN(n16164) );
  AOI22_X1 U19628 ( .A1(n16203), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16150) );
  AOI22_X1 U19629 ( .A1(n16205), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16149) );
  NAND2_X1 U19630 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n16148) );
  NAND2_X1 U19631 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n16147) );
  NAND4_X1 U19632 ( .A1(n16150), .A2(n16149), .A3(n16148), .A4(n16147), .ZN(
        n16155) );
  OAI22_X1 U19633 ( .A1(n16153), .A2(n16152), .B1(n11252), .B2(n16151), .ZN(
        n16154) );
  NOR2_X1 U19634 ( .A1(n16155), .A2(n16154), .ZN(n16163) );
  OAI22_X1 U19635 ( .A1(n16217), .A2(n16157), .B1(n16109), .B2(n16156), .ZN(
        n16161) );
  INV_X1 U19636 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16158) );
  OAI22_X1 U19637 ( .A1(n16215), .A2(n16159), .B1(n16219), .B2(n16158), .ZN(
        n16160) );
  NOR2_X1 U19638 ( .A1(n16161), .A2(n16160), .ZN(n16162) );
  OAI22_X1 U19639 ( .A1(n16351), .A2(n16229), .B1(n16225), .B2(n16165), .ZN(
        n16167) );
  OAI22_X1 U19640 ( .A1(n16342), .A2(n9764), .B1(n16221), .B2(n17312), .ZN(
        n16166) );
  NOR2_X1 U19641 ( .A1(n16167), .A2(n16166), .ZN(n16181) );
  AOI22_X1 U19642 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n16203), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16171) );
  AOI22_X1 U19643 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n16205), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16170) );
  NAND2_X1 U19644 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n16169) );
  NAND2_X1 U19645 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n16168) );
  NAND4_X1 U19646 ( .A1(n16171), .A2(n16170), .A3(n16169), .A4(n16168), .ZN(
        n16173) );
  OAI22_X1 U19647 ( .A1(n21796), .A2(n11252), .B1(n16153), .B2(n16341), .ZN(
        n16172) );
  NOR2_X1 U19648 ( .A1(n16173), .A2(n16172), .ZN(n16180) );
  OAI22_X1 U19649 ( .A1(n16339), .A2(n16217), .B1(n16109), .B2(n16174), .ZN(
        n16178) );
  INV_X1 U19650 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16175) );
  OAI22_X1 U19651 ( .A1(n16215), .A2(n16176), .B1(n16219), .B2(n16175), .ZN(
        n16177) );
  NOR2_X1 U19652 ( .A1(n16178), .A2(n16177), .ZN(n16179) );
  NAND3_X1 U19653 ( .A1(n16181), .A2(n16180), .A3(n16179), .ZN(n16428) );
  INV_X1 U19654 ( .A(n16182), .ZN(n16373) );
  AOI22_X1 U19655 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16193) );
  AOI22_X1 U19656 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16192) );
  AOI22_X1 U19657 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16191) );
  INV_X1 U19658 ( .A(n16184), .ZN(n16187) );
  INV_X1 U19659 ( .A(n16185), .ZN(n16186) );
  NAND2_X1 U19660 ( .A1(n16187), .A2(n16186), .ZN(n16368) );
  INV_X1 U19661 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n21972) );
  NAND2_X1 U19662 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n16189) );
  NAND2_X1 U19663 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n16188) );
  AND3_X1 U19664 ( .A1(n16368), .A2(n16189), .A3(n16188), .ZN(n16190) );
  NAND4_X1 U19665 ( .A1(n16193), .A2(n16192), .A3(n16191), .A4(n16190), .ZN(
        n16201) );
  AOI22_X1 U19666 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16199) );
  AOI22_X1 U19667 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9768), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16198) );
  AOI22_X1 U19668 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16197) );
  INV_X1 U19669 ( .A(n16368), .ZN(n16381) );
  NAND2_X1 U19670 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n16195) );
  NAND2_X1 U19671 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n16194) );
  AND3_X1 U19672 ( .A1(n16381), .A2(n16195), .A3(n16194), .ZN(n16196) );
  NAND4_X1 U19673 ( .A1(n16199), .A2(n16198), .A3(n16197), .A4(n16196), .ZN(
        n16200) );
  NAND2_X1 U19674 ( .A1(n16201), .A2(n16200), .ZN(n16255) );
  NOR2_X1 U19675 ( .A1(n20854), .A2(n16255), .ZN(n16253) );
  AOI22_X1 U19676 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n16203), .B1(
        n16202), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16210) );
  AOI22_X1 U19677 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n16205), .B1(
        n16204), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16209) );
  NAND2_X1 U19678 ( .A1(n11189), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n16208) );
  NAND2_X1 U19679 ( .A1(n16206), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n16207) );
  NAND4_X1 U19680 ( .A1(n16210), .A2(n16209), .A3(n16208), .A4(n16207), .ZN(
        n16213) );
  OAI22_X1 U19681 ( .A1(n16211), .A2(n11252), .B1(n16153), .B2(n21759), .ZN(
        n16212) );
  NOR2_X1 U19682 ( .A1(n16213), .A2(n16212), .ZN(n16235) );
  INV_X1 U19683 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16214) );
  OAI22_X1 U19684 ( .A1(n16217), .A2(n16216), .B1(n16215), .B2(n16214), .ZN(
        n16223) );
  INV_X1 U19685 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16218) );
  OAI22_X1 U19686 ( .A1(n16221), .A2(n16220), .B1(n16219), .B2(n16218), .ZN(
        n16222) );
  NOR2_X1 U19687 ( .A1(n16223), .A2(n16222), .ZN(n16234) );
  OAI22_X1 U19688 ( .A1(n16494), .A2(n16109), .B1(n16225), .B2(n16224), .ZN(
        n16226) );
  INV_X1 U19689 ( .A(n16226), .ZN(n16233) );
  OAI22_X1 U19690 ( .A1(n16230), .A2(n16229), .B1(n16228), .B2(n16227), .ZN(
        n16231) );
  INV_X1 U19691 ( .A(n16231), .ZN(n16232) );
  NAND4_X1 U19692 ( .A1(n16235), .A2(n16234), .A3(n16233), .A4(n16232), .ZN(
        n16256) );
  NOR2_X1 U19693 ( .A1(n20146), .A2(n16255), .ZN(n16423) );
  AOI22_X1 U19694 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16243) );
  AOI22_X1 U19695 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16242) );
  AOI22_X1 U19696 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16241) );
  NAND2_X1 U19697 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n16239) );
  NAND2_X1 U19698 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n16238) );
  AND3_X1 U19699 ( .A1(n16368), .A2(n16239), .A3(n16238), .ZN(n16240) );
  NAND4_X1 U19700 ( .A1(n16243), .A2(n16242), .A3(n16241), .A4(n16240), .ZN(
        n16252) );
  AOI22_X1 U19701 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16372), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16250) );
  AOI22_X1 U19702 ( .A1(n16377), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9768), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16249) );
  AOI22_X1 U19703 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9765), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16248) );
  NAND2_X1 U19704 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n16246) );
  NAND2_X1 U19705 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n16245) );
  AND3_X1 U19706 ( .A1(n16381), .A2(n16246), .A3(n16245), .ZN(n16247) );
  NAND4_X1 U19707 ( .A1(n16250), .A2(n16249), .A3(n16248), .A4(n16247), .ZN(
        n16251) );
  AND2_X1 U19708 ( .A1(n16252), .A2(n16251), .ZN(n16254) );
  AOI21_X1 U19709 ( .B1(n16253), .B2(n16256), .A(n16254), .ZN(n16259) );
  INV_X1 U19710 ( .A(n16254), .ZN(n16258) );
  NOR2_X1 U19711 ( .A1(n16258), .A2(n16255), .ZN(n16257) );
  AND2_X1 U19712 ( .A1(n16257), .A2(n16256), .ZN(n16277) );
  OAI22_X1 U19713 ( .A1(n16259), .A2(n16277), .B1(n16258), .B2(n20146), .ZN(
        n16417) );
  AOI22_X1 U19714 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16265) );
  AOI22_X1 U19715 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16264) );
  AOI22_X1 U19716 ( .A1(n16340), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16263) );
  NAND2_X1 U19717 ( .A1(n9765), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n16261) );
  NAND2_X1 U19718 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n16260) );
  AND3_X1 U19719 ( .A1(n16368), .A2(n16261), .A3(n16260), .ZN(n16262) );
  NAND4_X1 U19720 ( .A1(n16265), .A2(n16264), .A3(n16263), .A4(n16262), .ZN(
        n16275) );
  AOI22_X1 U19721 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16266), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16273) );
  AOI22_X1 U19722 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9768), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16272) );
  AOI22_X1 U19723 ( .A1(n16374), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16271) );
  NAND2_X1 U19724 ( .A1(n9765), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n16269) );
  NAND2_X1 U19725 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n16268) );
  AND3_X1 U19726 ( .A1(n16381), .A2(n16269), .A3(n16268), .ZN(n16270) );
  NAND4_X1 U19727 ( .A1(n16273), .A2(n16272), .A3(n16271), .A4(n16270), .ZN(
        n16274) );
  NAND2_X1 U19728 ( .A1(n16275), .A2(n16274), .ZN(n16280) );
  INV_X1 U19729 ( .A(n16280), .ZN(n16278) );
  INV_X1 U19730 ( .A(n16277), .ZN(n16276) );
  OAI211_X1 U19731 ( .C1(n16278), .C2(n16277), .A(n16319), .B(n16314), .ZN(
        n16281) );
  INV_X1 U19732 ( .A(n16281), .ZN(n16279) );
  NOR2_X1 U19733 ( .A1(n20146), .A2(n16280), .ZN(n16412) );
  NAND2_X2 U19734 ( .A1(n16411), .A2(n10813), .ZN(n16299) );
  AOI22_X1 U19735 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16377), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16288) );
  AOI22_X1 U19736 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16287) );
  AOI22_X1 U19737 ( .A1(n16374), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16286) );
  NAND2_X1 U19738 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n16284) );
  NAND2_X1 U19739 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n16283) );
  AND3_X1 U19740 ( .A1(n16368), .A2(n16284), .A3(n16283), .ZN(n16285) );
  NAND4_X1 U19741 ( .A1(n16288), .A2(n16287), .A3(n16286), .A4(n16285), .ZN(
        n16297) );
  AOI22_X1 U19742 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16377), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16295) );
  AOI22_X1 U19743 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16294) );
  AOI22_X1 U19744 ( .A1(n16374), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16293) );
  NAND2_X1 U19745 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n16291) );
  NAND2_X1 U19746 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n16290) );
  AND3_X1 U19747 ( .A1(n16381), .A2(n16291), .A3(n16290), .ZN(n16292) );
  NAND4_X1 U19748 ( .A1(n16295), .A2(n16294), .A3(n16293), .A4(n16292), .ZN(
        n16296) );
  XNOR2_X1 U19749 ( .A(n16314), .B(n16315), .ZN(n16298) );
  NAND2_X1 U19750 ( .A1(n20854), .A2(n16315), .ZN(n16407) );
  AOI22_X1 U19751 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16377), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16305) );
  AOI22_X1 U19752 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16304) );
  AOI22_X1 U19753 ( .A1(n16374), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16303) );
  NAND2_X1 U19754 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n16301) );
  NAND2_X1 U19755 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n16300) );
  AND3_X1 U19756 ( .A1(n16368), .A2(n16301), .A3(n16300), .ZN(n16302) );
  NAND4_X1 U19757 ( .A1(n16305), .A2(n16304), .A3(n16303), .A4(n16302), .ZN(
        n16313) );
  AOI22_X1 U19758 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16377), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16311) );
  AOI22_X1 U19759 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16310) );
  AOI22_X1 U19760 ( .A1(n16374), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16309) );
  NAND2_X1 U19761 ( .A1(n9765), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n16307) );
  NAND2_X1 U19762 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n16306) );
  AND3_X1 U19763 ( .A1(n16381), .A2(n16307), .A3(n16306), .ZN(n16308) );
  NAND4_X1 U19764 ( .A1(n16311), .A2(n16310), .A3(n16309), .A4(n16308), .ZN(
        n16312) );
  NAND2_X1 U19765 ( .A1(n16313), .A2(n16312), .ZN(n16317) );
  INV_X1 U19766 ( .A(n16317), .ZN(n16323) );
  INV_X1 U19767 ( .A(n16314), .ZN(n16316) );
  NAND2_X1 U19768 ( .A1(n16316), .A2(n16315), .ZN(n16318) );
  INV_X1 U19769 ( .A(n16318), .ZN(n16320) );
  OR2_X1 U19770 ( .A1(n16318), .A2(n16317), .ZN(n16395) );
  OAI211_X1 U19771 ( .C1(n16323), .C2(n16320), .A(n16395), .B(n16319), .ZN(
        n16321) );
  INV_X1 U19772 ( .A(n16321), .ZN(n16322) );
  NAND2_X1 U19773 ( .A1(n20854), .A2(n16323), .ZN(n16402) );
  AOI22_X1 U19774 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16377), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16329) );
  AOI22_X1 U19775 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9768), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16328) );
  AOI22_X1 U19776 ( .A1(n16374), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16327) );
  NAND2_X1 U19777 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n16325) );
  NAND2_X1 U19778 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n16324) );
  AND3_X1 U19779 ( .A1(n16368), .A2(n16325), .A3(n16324), .ZN(n16326) );
  NAND4_X1 U19780 ( .A1(n16329), .A2(n16328), .A3(n16327), .A4(n16326), .ZN(
        n16337) );
  AOI22_X1 U19781 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16377), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16335) );
  AOI22_X1 U19782 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16334) );
  AOI22_X1 U19783 ( .A1(n16374), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16333) );
  NAND2_X1 U19784 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n16331) );
  NAND2_X1 U19785 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n16330) );
  AND3_X1 U19786 ( .A1(n16381), .A2(n16331), .A3(n16330), .ZN(n16332) );
  NAND4_X1 U19787 ( .A1(n16335), .A2(n16334), .A3(n16333), .A4(n16332), .ZN(
        n16336) );
  AND2_X1 U19788 ( .A1(n16337), .A2(n16336), .ZN(n16397) );
  INV_X1 U19789 ( .A(n16397), .ZN(n16338) );
  NOR3_X1 U19790 ( .A1(n16395), .A2(n20854), .A3(n16338), .ZN(n16363) );
  INV_X1 U19791 ( .A(n16377), .ZN(n16353) );
  OAI22_X1 U19792 ( .A1(n16182), .A2(n21796), .B1(n16353), .B2(n16339), .ZN(
        n16348) );
  OAI22_X1 U19793 ( .A1(n11164), .A2(n16342), .B1(n16183), .B2(n16341), .ZN(
        n16347) );
  AOI22_X1 U19794 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16345) );
  NAND2_X1 U19795 ( .A1(n9765), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n16344) );
  NAND2_X1 U19796 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n16343) );
  NAND4_X1 U19797 ( .A1(n16345), .A2(n16344), .A3(n16381), .A4(n16343), .ZN(
        n16346) );
  NOR3_X1 U19798 ( .A1(n16348), .A2(n16347), .A3(n16346), .ZN(n16361) );
  AOI22_X1 U19799 ( .A1(n16372), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16350) );
  NAND2_X1 U19800 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n16349) );
  OAI211_X1 U19801 ( .C1(n16174), .C2(n11164), .A(n16350), .B(n16349), .ZN(
        n16359) );
  OAI22_X1 U19802 ( .A1(n16353), .A2(n16175), .B1(n9736), .B2(n16351), .ZN(
        n16358) );
  NAND2_X1 U19803 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n16354) );
  OAI211_X1 U19804 ( .C1(n16356), .C2(n16355), .A(n16354), .B(n16368), .ZN(
        n16357) );
  NOR3_X1 U19805 ( .A1(n16359), .A2(n16358), .A3(n16357), .ZN(n16360) );
  NOR2_X1 U19806 ( .A1(n16361), .A2(n16360), .ZN(n16362) );
  NAND2_X1 U19807 ( .A1(n16363), .A2(n16362), .ZN(n16364) );
  OAI21_X1 U19808 ( .B1(n16363), .B2(n16362), .A(n16364), .ZN(n16391) );
  INV_X1 U19809 ( .A(n16364), .ZN(n16365) );
  AOI22_X1 U19810 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16372), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U19811 ( .A1(n16374), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9767), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16366) );
  NAND2_X1 U19812 ( .A1(n16367), .A2(n16366), .ZN(n16386) );
  AOI22_X1 U19813 ( .A1(n16377), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16371) );
  NAND2_X1 U19814 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n16370) );
  NAND2_X1 U19815 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n16369) );
  NAND4_X1 U19816 ( .A1(n16371), .A2(n16370), .A3(n16369), .A4(n16368), .ZN(
        n16385) );
  AOI22_X1 U19817 ( .A1(n16373), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16372), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16376) );
  AOI22_X1 U19818 ( .A1(n16374), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9768), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16375) );
  NAND2_X1 U19819 ( .A1(n16376), .A2(n16375), .ZN(n16384) );
  AOI22_X1 U19820 ( .A1(n16377), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16382) );
  NAND2_X1 U19821 ( .A1(n16378), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n16380) );
  NAND2_X1 U19822 ( .A1(n16244), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n16379) );
  NAND4_X1 U19823 ( .A1(n16382), .A2(n16381), .A3(n16380), .A4(n16379), .ZN(
        n16383) );
  OAI22_X1 U19824 ( .A1(n16386), .A2(n16385), .B1(n16384), .B2(n16383), .ZN(
        n16387) );
  NOR2_X1 U19825 ( .A1(n16388), .A2(n16503), .ZN(n16389) );
  OAI21_X1 U19826 ( .B1(n16518), .B2(n20076), .A(n16390), .ZN(P2_U2857) );
  INV_X1 U19827 ( .A(n16952), .ZN(n16394) );
  NAND2_X1 U19828 ( .A1(n16503), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16392) );
  OAI211_X1 U19829 ( .C1(n16503), .C2(n16394), .A(n16393), .B(n16392), .ZN(
        P2_U2858) );
  NAND2_X1 U19830 ( .A1(n16396), .A2(n16395), .ZN(n16398) );
  XNOR2_X1 U19831 ( .A(n16398), .B(n16397), .ZN(n16533) );
  NOR2_X1 U19832 ( .A1(n16964), .A2(n16503), .ZN(n16399) );
  AOI21_X1 U19833 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16503), .A(n16399), .ZN(
        n16400) );
  OAI21_X1 U19834 ( .B1(n16533), .B2(n20076), .A(n16400), .ZN(P2_U2859) );
  AOI21_X1 U19835 ( .B1(n16403), .B2(n16402), .A(n16401), .ZN(n16534) );
  NAND2_X1 U19836 ( .A1(n16534), .A2(n16497), .ZN(n16405) );
  NAND2_X1 U19837 ( .A1(n16503), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16404) );
  OAI211_X1 U19838 ( .C1(n16503), .C2(n16665), .A(n16405), .B(n16404), .ZN(
        P2_U2860) );
  AOI21_X1 U19839 ( .B1(n16408), .B2(n16407), .A(n16406), .ZN(n16542) );
  NAND2_X1 U19840 ( .A1(n16542), .A2(n16497), .ZN(n16410) );
  NAND2_X1 U19841 ( .A1(n16503), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16409) );
  OAI211_X1 U19842 ( .C1(n16681), .C2(n16503), .A(n16410), .B(n16409), .ZN(
        P2_U2861) );
  OAI21_X1 U19843 ( .B1(n16413), .B2(n16412), .A(n16411), .ZN(n16556) );
  NAND2_X1 U19844 ( .A1(n16995), .A2(n20082), .ZN(n16415) );
  NAND2_X1 U19845 ( .A1(n16503), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16414) );
  OAI211_X1 U19846 ( .C1(n16556), .C2(n20076), .A(n16415), .B(n16414), .ZN(
        P2_U2862) );
  NAND2_X1 U19847 ( .A1(n17008), .A2(n20082), .ZN(n16420) );
  OR2_X1 U19848 ( .A1(n16418), .A2(n16417), .ZN(n16562) );
  NAND3_X1 U19849 ( .A1(n16416), .A2(n16562), .A3(n16497), .ZN(n16419) );
  OAI211_X1 U19850 ( .C1(n20082), .C2(n16421), .A(n16420), .B(n16419), .ZN(
        P2_U2863) );
  INV_X1 U19851 ( .A(n17028), .ZN(n16427) );
  OAI21_X1 U19852 ( .B1(n16424), .B2(n16423), .A(n16422), .ZN(n16571) );
  INV_X1 U19853 ( .A(n16571), .ZN(n16425) );
  AOI22_X1 U19854 ( .A1(n16425), .A2(n16497), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n16503), .ZN(n16426) );
  OAI21_X1 U19855 ( .B1(n16427), .B2(n16503), .A(n16426), .ZN(P2_U2864) );
  INV_X1 U19856 ( .A(n16428), .ZN(n16431) );
  INV_X1 U19857 ( .A(n16434), .ZN(n16430) );
  AOI21_X1 U19858 ( .B1(n16431), .B2(n16430), .A(n16429), .ZN(n16577) );
  AOI22_X1 U19859 ( .A1(n16577), .A2(n16497), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n16503), .ZN(n16432) );
  OAI21_X1 U19860 ( .B1(n16716), .B2(n16503), .A(n16432), .ZN(P2_U2865) );
  INV_X1 U19861 ( .A(n17043), .ZN(n16437) );
  AOI21_X1 U19862 ( .B1(n16435), .B2(n16433), .A(n16434), .ZN(n16583) );
  AOI22_X1 U19863 ( .A1(n16583), .A2(n16497), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n16503), .ZN(n16436) );
  OAI21_X1 U19864 ( .B1(n16437), .B2(n16503), .A(n16436), .ZN(P2_U2866) );
  INV_X1 U19865 ( .A(n16438), .ZN(n16445) );
  NOR2_X1 U19866 ( .A1(n16439), .A2(n16440), .ZN(n16458) );
  NAND2_X1 U19867 ( .A1(n16451), .A2(n16447), .ZN(n16446) );
  INV_X1 U19868 ( .A(n16441), .ZN(n16443) );
  INV_X1 U19869 ( .A(n16433), .ZN(n16442) );
  AOI21_X1 U19870 ( .B1(n16446), .B2(n16443), .A(n16442), .ZN(n16589) );
  AOI22_X1 U19871 ( .A1(n16589), .A2(n16497), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n16503), .ZN(n16444) );
  OAI21_X1 U19872 ( .B1(n16445), .B2(n16503), .A(n16444), .ZN(P2_U2867) );
  OAI21_X1 U19873 ( .B1(n16451), .B2(n16447), .A(n16446), .ZN(n16599) );
  INV_X1 U19874 ( .A(n16599), .ZN(n16448) );
  AOI22_X1 U19875 ( .A1(n16448), .A2(n16497), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n16503), .ZN(n16449) );
  OAI21_X1 U19876 ( .B1(n17065), .B2(n16503), .A(n16449), .ZN(P2_U2868) );
  INV_X1 U19877 ( .A(n16450), .ZN(n16453) );
  INV_X1 U19878 ( .A(n16458), .ZN(n16452) );
  AOI21_X1 U19879 ( .B1(n16453), .B2(n16452), .A(n16451), .ZN(n16606) );
  AOI22_X1 U19880 ( .A1(n16606), .A2(n16497), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n16503), .ZN(n16454) );
  OAI21_X1 U19881 ( .B1(n16455), .B2(n16503), .A(n16454), .ZN(P2_U2869) );
  INV_X1 U19882 ( .A(n16439), .ZN(n16473) );
  NAND2_X1 U19883 ( .A1(n16473), .A2(n16472), .ZN(n16471) );
  INV_X1 U19884 ( .A(n16456), .ZN(n16467) );
  NOR2_X1 U19885 ( .A1(n16471), .A2(n16467), .ZN(n16466) );
  NAND2_X1 U19886 ( .A1(n16466), .A2(n16462), .ZN(n16461) );
  INV_X1 U19887 ( .A(n16457), .ZN(n16459) );
  AOI21_X1 U19888 ( .B1(n16461), .B2(n16459), .A(n16458), .ZN(n16612) );
  AOI22_X1 U19889 ( .A1(n16612), .A2(n16497), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n16503), .ZN(n16460) );
  OAI21_X1 U19890 ( .B1(n17089), .B2(n16503), .A(n16460), .ZN(P2_U2870) );
  OAI21_X1 U19891 ( .B1(n16466), .B2(n16462), .A(n16461), .ZN(n16624) );
  INV_X1 U19892 ( .A(n16624), .ZN(n16463) );
  AOI22_X1 U19893 ( .A1(n16463), .A2(n16497), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n16503), .ZN(n16464) );
  OAI21_X1 U19894 ( .B1(n17101), .B2(n16503), .A(n16464), .ZN(P2_U2871) );
  AOI21_X1 U19895 ( .B1(n16465), .B2(n15824), .A(n15798), .ZN(n20042) );
  INV_X1 U19896 ( .A(n20042), .ZN(n16470) );
  AOI211_X1 U19897 ( .C1(n16467), .C2(n16471), .A(n20076), .B(n16466), .ZN(
        n16468) );
  AOI21_X1 U19898 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(n16503), .A(n16468), .ZN(
        n16469) );
  OAI21_X1 U19899 ( .B1(n16470), .B2(n16503), .A(n16469), .ZN(P2_U2872) );
  NAND2_X1 U19900 ( .A1(n17119), .A2(n20082), .ZN(n16475) );
  OAI211_X1 U19901 ( .C1(n16473), .C2(n16472), .A(n16471), .B(n16497), .ZN(
        n16474) );
  OAI211_X1 U19902 ( .C1(n20082), .C2(n16476), .A(n16475), .B(n16474), .ZN(
        P2_U2873) );
  INV_X1 U19903 ( .A(n16477), .ZN(n20078) );
  NAND2_X1 U19904 ( .A1(n20075), .A2(n16489), .ZN(n16483) );
  INV_X1 U19905 ( .A(n16484), .ZN(n16478) );
  NOR2_X1 U19906 ( .A1(n16483), .A2(n16478), .ZN(n16480) );
  OAI211_X1 U19907 ( .C1(n16480), .C2(n16479), .A(n16497), .B(n16439), .ZN(
        n16482) );
  NAND2_X1 U19908 ( .A1(n16503), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n16481) );
  OAI211_X1 U19909 ( .C1(n17132), .C2(n16503), .A(n16482), .B(n16481), .ZN(
        P2_U2874) );
  XOR2_X1 U19910 ( .A(n16484), .B(n16483), .Z(n16488) );
  MUX2_X1 U19911 ( .A(n16486), .B(n16485), .S(n16503), .Z(n16487) );
  OAI21_X1 U19912 ( .B1(n16488), .B2(n20076), .A(n16487), .ZN(P2_U2875) );
  XNOR2_X1 U19913 ( .A(n20075), .B(n16489), .ZN(n16492) );
  NOR2_X1 U19914 ( .A1(n17150), .A2(n16503), .ZN(n16490) );
  AOI21_X1 U19915 ( .B1(P2_EBX_REG_11__SCAN_IN), .B2(n16503), .A(n16490), .ZN(
        n16491) );
  OAI21_X1 U19916 ( .B1(n16492), .B2(n20076), .A(n16491), .ZN(P2_U2876) );
  NAND2_X1 U19917 ( .A1(n16493), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n16502) );
  NOR2_X1 U19918 ( .A1(n16502), .A2(n16494), .ZN(n16499) );
  INV_X1 U19919 ( .A(n16495), .ZN(n16496) );
  OAI211_X1 U19920 ( .C1(n16499), .C2(n16498), .A(n16497), .B(n16496), .ZN(
        n16501) );
  NAND2_X1 U19921 ( .A1(n16503), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n16500) );
  OAI211_X1 U19922 ( .C1(n17187), .C2(n16503), .A(n16501), .B(n16500), .ZN(
        P2_U2879) );
  XOR2_X1 U19923 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n16502), .Z(n16506)
         );
  INV_X1 U19924 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n16504) );
  MUX2_X1 U19925 ( .A(n17208), .B(n16504), .S(n16503), .Z(n16505) );
  OAI21_X1 U19926 ( .B1(n16506), .B2(n20076), .A(n16505), .ZN(P2_U2880) );
  INV_X1 U19927 ( .A(n16615), .ZN(n16604) );
  INV_X1 U19928 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16509) );
  AOI22_X1 U19929 ( .A1(n16618), .A2(n16507), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n20093), .ZN(n16508) );
  OAI21_X1 U19930 ( .B1(n16604), .B2(n16509), .A(n16508), .ZN(n16510) );
  INV_X1 U19931 ( .A(n16616), .ZN(n16512) );
  INV_X1 U19932 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n16511) );
  NOR2_X1 U19933 ( .A1(n16512), .A2(n16511), .ZN(n16513) );
  INV_X1 U19934 ( .A(n16516), .ZN(n16517) );
  OAI21_X1 U19935 ( .B1(n16518), .B2(n16625), .A(n16517), .ZN(P2_U2889) );
  NAND3_X1 U19936 ( .A1(n16520), .A2(n22058), .A3(n16519), .ZN(n16526) );
  NAND2_X1 U19937 ( .A1(n16616), .A2(BUF2_REG_29__SCAN_IN), .ZN(n16524) );
  NAND2_X1 U19938 ( .A1(n16615), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16523) );
  AOI22_X1 U19939 ( .A1(n16618), .A2(n16521), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n20093), .ZN(n16522) );
  AND3_X1 U19940 ( .A1(n16524), .A2(n16523), .A3(n16522), .ZN(n16525) );
  OAI211_X1 U19941 ( .C1(n20085), .C2(n16950), .A(n16526), .B(n16525), .ZN(
        P2_U2890) );
  NAND2_X1 U19942 ( .A1(n16615), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16529) );
  AOI22_X1 U19943 ( .A1(n16618), .A2(n16527), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n20093), .ZN(n16528) );
  NAND2_X1 U19944 ( .A1(n16529), .A2(n16528), .ZN(n16531) );
  NOR2_X1 U19945 ( .A1(n16963), .A2(n20085), .ZN(n16530) );
  AOI211_X1 U19946 ( .C1(n16616), .C2(BUF2_REG_28__SCAN_IN), .A(n16531), .B(
        n16530), .ZN(n16532) );
  OAI21_X1 U19947 ( .B1(n16533), .B2(n16625), .A(n16532), .ZN(P2_U2891) );
  INV_X1 U19948 ( .A(n16534), .ZN(n16541) );
  NAND2_X1 U19949 ( .A1(n16615), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16537) );
  AOI22_X1 U19950 ( .A1(n16618), .A2(n16535), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n20093), .ZN(n16536) );
  NAND2_X1 U19951 ( .A1(n16537), .A2(n16536), .ZN(n16539) );
  NOR2_X1 U19952 ( .A1(n16970), .A2(n20085), .ZN(n16538) );
  AOI211_X1 U19953 ( .C1(n16616), .C2(BUF2_REG_27__SCAN_IN), .A(n16539), .B(
        n16538), .ZN(n16540) );
  OAI21_X1 U19954 ( .B1(n16541), .B2(n16625), .A(n16540), .ZN(P2_U2892) );
  INV_X1 U19955 ( .A(n16542), .ZN(n16549) );
  NAND2_X1 U19956 ( .A1(n16615), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16545) );
  AOI22_X1 U19957 ( .A1(n16618), .A2(n16543), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n20093), .ZN(n16544) );
  NAND2_X1 U19958 ( .A1(n16545), .A2(n16544), .ZN(n16547) );
  NOR2_X1 U19959 ( .A1(n16991), .A2(n20085), .ZN(n16546) );
  AOI211_X1 U19960 ( .C1(n16616), .C2(BUF2_REG_26__SCAN_IN), .A(n16547), .B(
        n16546), .ZN(n16548) );
  OAI21_X1 U19961 ( .B1(n16549), .B2(n16625), .A(n16548), .ZN(P2_U2893) );
  NAND2_X1 U19962 ( .A1(n16615), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16552) );
  AOI22_X1 U19963 ( .A1(n16618), .A2(n16550), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n20093), .ZN(n16551) );
  NAND2_X1 U19964 ( .A1(n16552), .A2(n16551), .ZN(n16554) );
  NOR2_X1 U19965 ( .A1(n17003), .A2(n20085), .ZN(n16553) );
  AOI211_X1 U19966 ( .C1(n16616), .C2(BUF2_REG_25__SCAN_IN), .A(n16554), .B(
        n16553), .ZN(n16555) );
  OAI21_X1 U19967 ( .B1(n16625), .B2(n16556), .A(n16555), .ZN(P2_U2894) );
  NAND2_X1 U19968 ( .A1(n16615), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16559) );
  AOI22_X1 U19969 ( .A1(n16618), .A2(n16557), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n20093), .ZN(n16558) );
  NAND2_X1 U19970 ( .A1(n16559), .A2(n16558), .ZN(n16561) );
  NOR2_X1 U19971 ( .A1(n17014), .A2(n20085), .ZN(n16560) );
  AOI211_X1 U19972 ( .C1(n16616), .C2(BUF2_REG_24__SCAN_IN), .A(n16561), .B(
        n16560), .ZN(n16564) );
  NAND3_X1 U19973 ( .A1(n16416), .A2(n16562), .A3(n22058), .ZN(n16563) );
  NAND2_X1 U19974 ( .A1(n16564), .A2(n16563), .ZN(P2_U2895) );
  NAND2_X1 U19975 ( .A1(n16616), .A2(BUF2_REG_23__SCAN_IN), .ZN(n16567) );
  AOI22_X1 U19976 ( .A1(n16618), .A2(n16565), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n20093), .ZN(n16566) );
  NAND2_X1 U19977 ( .A1(n16567), .A2(n16566), .ZN(n16569) );
  NOR2_X1 U19978 ( .A1(n17023), .A2(n20085), .ZN(n16568) );
  AOI211_X1 U19979 ( .C1(BUF1_REG_23__SCAN_IN), .C2(n16615), .A(n16569), .B(
        n16568), .ZN(n16570) );
  OAI21_X1 U19980 ( .B1(n16625), .B2(n16571), .A(n16570), .ZN(P2_U2896) );
  INV_X1 U19981 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16575) );
  INV_X1 U19982 ( .A(n17309), .ZN(n16572) );
  AOI22_X1 U19983 ( .A1(n16618), .A2(n16572), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n20093), .ZN(n16574) );
  NAND2_X1 U19984 ( .A1(n16615), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16573) );
  OAI211_X1 U19985 ( .C1(n16512), .C2(n16575), .A(n16574), .B(n16573), .ZN(
        n16576) );
  AOI21_X1 U19986 ( .B1(n16577), .B2(n22058), .A(n16576), .ZN(n16578) );
  OAI21_X1 U19987 ( .B1(n17036), .B2(n20085), .A(n16578), .ZN(P2_U2897) );
  INV_X1 U19988 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16581) );
  AOI22_X1 U19989 ( .A1(n16618), .A2(n20168), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n20093), .ZN(n16580) );
  NAND2_X1 U19990 ( .A1(n16615), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16579) );
  OAI211_X1 U19991 ( .C1(n16512), .C2(n16581), .A(n16580), .B(n16579), .ZN(
        n16582) );
  AOI21_X1 U19992 ( .B1(n16583), .B2(n22058), .A(n16582), .ZN(n16584) );
  OAI21_X1 U19993 ( .B1(n17052), .B2(n20085), .A(n16584), .ZN(P2_U2898) );
  INV_X1 U19994 ( .A(n20163), .ZN(n16585) );
  AOI22_X1 U19995 ( .A1(n16618), .A2(n16585), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n20093), .ZN(n16587) );
  NAND2_X1 U19996 ( .A1(n16616), .A2(BUF2_REG_20__SCAN_IN), .ZN(n16586) );
  OAI211_X1 U19997 ( .C1(n16604), .C2(n21081), .A(n16587), .B(n16586), .ZN(
        n16588) );
  AOI21_X1 U19998 ( .B1(n16589), .B2(n22058), .A(n16588), .ZN(n16590) );
  OAI21_X1 U19999 ( .B1(n16591), .B2(n20085), .A(n16590), .ZN(P2_U2899) );
  NAND2_X1 U20000 ( .A1(n17063), .A2(n22053), .ZN(n16598) );
  INV_X1 U20001 ( .A(n16618), .ZN(n16593) );
  OAI22_X1 U20002 ( .A1(n16593), .A2(n22063), .B1(n20084), .B2(n16592), .ZN(
        n16596) );
  NOR2_X1 U20003 ( .A1(n16604), .A2(n16594), .ZN(n16595) );
  AOI211_X1 U20004 ( .C1(n16616), .C2(BUF2_REG_19__SCAN_IN), .A(n16596), .B(
        n16595), .ZN(n16597) );
  OAI211_X1 U20005 ( .C1(n16599), .C2(n16625), .A(n16598), .B(n16597), .ZN(
        P2_U2900) );
  INV_X1 U20006 ( .A(n16600), .ZN(n17074) );
  AOI22_X1 U20007 ( .A1(n16618), .A2(n16601), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n20093), .ZN(n16603) );
  NAND2_X1 U20008 ( .A1(n16616), .A2(BUF2_REG_18__SCAN_IN), .ZN(n16602) );
  OAI211_X1 U20009 ( .C1(n16604), .C2(n21067), .A(n16603), .B(n16602), .ZN(
        n16605) );
  AOI21_X1 U20010 ( .B1(n16606), .B2(n22058), .A(n16605), .ZN(n16607) );
  OAI21_X1 U20011 ( .B1(n17074), .B2(n20085), .A(n16607), .ZN(P2_U2901) );
  NAND2_X1 U20012 ( .A1(n16615), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16611) );
  NAND2_X1 U20013 ( .A1(n16616), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16610) );
  AOI22_X1 U20014 ( .A1(n16618), .A2(n16608), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n20093), .ZN(n16609) );
  AND3_X1 U20015 ( .A1(n16611), .A2(n16610), .A3(n16609), .ZN(n16614) );
  NAND2_X1 U20016 ( .A1(n16612), .A2(n22058), .ZN(n16613) );
  OAI211_X1 U20017 ( .C1(n17085), .C2(n20085), .A(n16614), .B(n16613), .ZN(
        P2_U2902) );
  NAND2_X1 U20018 ( .A1(n16615), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16621) );
  NAND2_X1 U20019 ( .A1(n16616), .A2(BUF2_REG_16__SCAN_IN), .ZN(n16620) );
  AOI22_X1 U20020 ( .A1(n16618), .A2(n16617), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n20093), .ZN(n16619) );
  NAND3_X1 U20021 ( .A1(n16621), .A2(n16620), .A3(n16619), .ZN(n16622) );
  AOI21_X1 U20022 ( .B1(n17099), .B2(n22053), .A(n16622), .ZN(n16623) );
  OAI21_X1 U20023 ( .B1(n16625), .B2(n16624), .A(n16623), .ZN(P2_U2903) );
  XOR2_X1 U20024 ( .A(n14366), .B(n16626), .Z(n20039) );
  INV_X1 U20025 ( .A(n20039), .ZN(n16628) );
  OAI222_X1 U20026 ( .A1(n20084), .A2(n13856), .B1(n16628), .B2(n16637), .C1(
        n22062), .C2(n16627), .ZN(P2_U2904) );
  INV_X1 U20027 ( .A(n17257), .ZN(n22054) );
  INV_X1 U20028 ( .A(n20199), .ZN(n20805) );
  XOR2_X1 U20029 ( .A(n17257), .B(n20199), .Z(n22057) );
  INV_X1 U20030 ( .A(n20817), .ZN(n16631) );
  OAI21_X1 U20031 ( .B1(n16631), .B2(n16630), .A(n16629), .ZN(n22056) );
  NAND2_X1 U20032 ( .A1(n22057), .A2(n22056), .ZN(n22055) );
  OAI21_X1 U20033 ( .B1(n22054), .B2(n20805), .A(n22055), .ZN(n16632) );
  NAND2_X1 U20034 ( .A1(n16632), .A2(n20086), .ZN(n20089) );
  INV_X1 U20035 ( .A(n20088), .ZN(n16633) );
  NAND3_X1 U20036 ( .A1(n20089), .A2(n16633), .A3(n22058), .ZN(n16636) );
  AOI22_X1 U20037 ( .A1(n16634), .A2(n20168), .B1(n20093), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n16635) );
  OAI211_X1 U20038 ( .C1(n17233), .C2(n16637), .A(n16636), .B(n16635), .ZN(
        P2_U2914) );
  NAND2_X1 U20039 ( .A1(n16639), .A2(n16638), .ZN(n16640) );
  NOR2_X1 U20040 ( .A1(n16877), .A2(n20776), .ZN(n16945) );
  AOI21_X1 U20041 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16945), .ZN(n16642) );
  OAI21_X1 U20042 ( .B1(n16643), .B2(n16933), .A(n16642), .ZN(n16644) );
  OAI21_X1 U20043 ( .B1(n9855), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16647), .ZN(n16969) );
  INV_X1 U20044 ( .A(n16662), .ZN(n16648) );
  NOR2_X1 U20045 ( .A1(n16650), .A2(n16649), .ZN(n16653) );
  XNOR2_X1 U20046 ( .A(n16651), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16652) );
  XNOR2_X1 U20047 ( .A(n16653), .B(n16652), .ZN(n16967) );
  INV_X1 U20048 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n16654) );
  NOR2_X1 U20049 ( .A1(n16877), .A2(n16654), .ZN(n16957) );
  AOI21_X1 U20050 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16957), .ZN(n16657) );
  NAND2_X1 U20051 ( .A1(n16655), .A2(n16924), .ZN(n16656) );
  OAI211_X1 U20052 ( .C1(n16964), .C2(n17306), .A(n16657), .B(n16656), .ZN(
        n16658) );
  AOI21_X1 U20053 ( .B1(n16899), .B2(n16967), .A(n16658), .ZN(n16659) );
  OAI21_X1 U20054 ( .B1(n16911), .B2(n16969), .A(n16659), .ZN(P2_U2986) );
  NOR2_X1 U20055 ( .A1(n16661), .A2(n16660), .ZN(n16664) );
  XNOR2_X1 U20056 ( .A(n16662), .B(n16974), .ZN(n16663) );
  XNOR2_X1 U20057 ( .A(n16664), .B(n16663), .ZN(n16983) );
  INV_X1 U20058 ( .A(n16665), .ZN(n16978) );
  NOR2_X1 U20059 ( .A1(n16877), .A2(n20774), .ZN(n16971) );
  AOI21_X1 U20060 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16971), .ZN(n16666) );
  OAI21_X1 U20061 ( .B1(n16667), .B2(n16933), .A(n16666), .ZN(n16668) );
  AOI21_X1 U20062 ( .B1(n16978), .B2(n16935), .A(n16668), .ZN(n16671) );
  INV_X1 U20063 ( .A(n9855), .ZN(n16980) );
  NAND2_X1 U20064 ( .A1(n16669), .A2(n16974), .ZN(n16979) );
  NAND3_X1 U20065 ( .A1(n16980), .A2(n16939), .A3(n16979), .ZN(n16670) );
  OAI211_X1 U20066 ( .C1(n16983), .C2(n16942), .A(n16671), .B(n16670), .ZN(
        P2_U2987) );
  INV_X1 U20067 ( .A(n16686), .ZN(n16675) );
  NOR2_X1 U20068 ( .A1(n16877), .A2(n16677), .ZN(n16985) );
  NOR2_X1 U20069 ( .A1(n16678), .A2(n16933), .ZN(n16679) );
  AOI211_X1 U20070 ( .C1(n16930), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16985), .B(n16679), .ZN(n16680) );
  OAI21_X1 U20071 ( .B1(n16681), .B2(n17306), .A(n16680), .ZN(n16682) );
  AOI21_X1 U20072 ( .B1(n16899), .B2(n16993), .A(n16682), .ZN(n16683) );
  OAI21_X1 U20073 ( .B1(n16911), .B2(n16994), .A(n16683), .ZN(P2_U2988) );
  XNOR2_X1 U20074 ( .A(n16684), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17007) );
  NOR2_X1 U20075 ( .A1(n16686), .A2(n16685), .ZN(n16687) );
  XNOR2_X1 U20076 ( .A(n16674), .B(n16687), .ZN(n17005) );
  NAND2_X1 U20077 ( .A1(n16995), .A2(n16935), .ZN(n16689) );
  NOR2_X1 U20078 ( .A1(n16877), .A2(n21909), .ZN(n16996) );
  AOI21_X1 U20079 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16996), .ZN(n16688) );
  OAI211_X1 U20080 ( .C1(n16933), .C2(n16690), .A(n16689), .B(n16688), .ZN(
        n16691) );
  AOI21_X1 U20081 ( .B1(n16899), .B2(n17005), .A(n16691), .ZN(n16692) );
  OAI21_X1 U20082 ( .B1(n16911), .B2(n17007), .A(n16692), .ZN(P2_U2989) );
  OAI21_X1 U20083 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16706), .A(
        n16694), .ZN(n17018) );
  INV_X1 U20084 ( .A(n16696), .ZN(n16697) );
  XNOR2_X1 U20085 ( .A(n16696), .B(n21939), .ZN(n16710) );
  INV_X1 U20086 ( .A(n16698), .ZN(n16699) );
  NAND2_X1 U20087 ( .A1(n17008), .A2(n16935), .ZN(n16702) );
  NOR2_X1 U20088 ( .A1(n16877), .A2(n20769), .ZN(n17010) );
  AOI21_X1 U20089 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n17010), .ZN(n16701) );
  OAI211_X1 U20090 ( .C1(n16933), .C2(n16703), .A(n16702), .B(n16701), .ZN(
        n16704) );
  AOI21_X1 U20091 ( .B1(n16899), .B2(n17016), .A(n16704), .ZN(n16705) );
  OAI21_X1 U20092 ( .B1(n16911), .B2(n17018), .A(n16705), .ZN(P2_U2990) );
  OAI21_X1 U20093 ( .B1(n16714), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16693), .ZN(n17030) );
  NOR2_X1 U20094 ( .A1(n16877), .A2(n20767), .ZN(n17019) );
  AOI21_X1 U20095 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17019), .ZN(n16707) );
  OAI21_X1 U20096 ( .B1(n16708), .B2(n16933), .A(n16707), .ZN(n16712) );
  NOR3_X1 U20097 ( .A1(n17025), .A2(n17024), .A3(n16942), .ZN(n16711) );
  AOI211_X1 U20098 ( .C1(n16935), .C2(n17028), .A(n16712), .B(n16711), .ZN(
        n16713) );
  OAI21_X1 U20099 ( .B1(n17030), .B2(n16911), .A(n16713), .ZN(P2_U2991) );
  OAI21_X1 U20100 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16734), .A(
        n16715), .ZN(n17042) );
  INV_X1 U20101 ( .A(n16716), .ZN(n17038) );
  INV_X1 U20102 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16717) );
  NOR2_X1 U20103 ( .A1(n16877), .A2(n16717), .ZN(n17031) );
  AOI21_X1 U20104 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17031), .ZN(n16718) );
  OAI21_X1 U20105 ( .B1(n16719), .B2(n16933), .A(n16718), .ZN(n16720) );
  AOI21_X1 U20106 ( .B1(n17038), .B2(n16935), .A(n16720), .ZN(n16726) );
  NAND2_X1 U20107 ( .A1(n16722), .A2(n16721), .ZN(n16723) );
  XNOR2_X1 U20108 ( .A(n16724), .B(n16723), .ZN(n17039) );
  NAND2_X1 U20109 ( .A1(n17039), .A2(n16899), .ZN(n16725) );
  OAI211_X1 U20110 ( .C1(n17042), .C2(n16911), .A(n16726), .B(n16725), .ZN(
        P2_U2992) );
  INV_X1 U20111 ( .A(n16727), .ZN(n16728) );
  NAND2_X1 U20112 ( .A1(n16732), .A2(n16731), .ZN(n16733) );
  NAND2_X1 U20113 ( .A1(n17043), .A2(n16935), .ZN(n16737) );
  NOR2_X1 U20114 ( .A1(n16877), .A2(n20764), .ZN(n17047) );
  AOI21_X1 U20115 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n17047), .ZN(n16736) );
  OAI211_X1 U20116 ( .C1(n16933), .C2(n16738), .A(n16737), .B(n16736), .ZN(
        n16739) );
  OAI21_X1 U20117 ( .B1(n17056), .B2(n16942), .A(n16740), .ZN(P2_U2993) );
  NAND2_X1 U20118 ( .A1(n16742), .A2(n16741), .ZN(n16746) );
  INV_X1 U20119 ( .A(n16743), .ZN(n16752) );
  XOR2_X1 U20120 ( .A(n16746), .B(n16745), .Z(n17069) );
  XNOR2_X1 U20121 ( .A(n16756), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17067) );
  NOR2_X1 U20122 ( .A1(n16877), .A2(n20760), .ZN(n17058) );
  NOR2_X1 U20123 ( .A1(n16747), .A2(n16933), .ZN(n16748) );
  AOI211_X1 U20124 ( .C1(n16930), .C2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n17058), .B(n16748), .ZN(n16749) );
  OAI21_X1 U20125 ( .B1(n17065), .B2(n17306), .A(n16749), .ZN(n16750) );
  AOI21_X1 U20126 ( .B1(n17067), .B2(n16939), .A(n16750), .ZN(n16751) );
  OAI21_X1 U20127 ( .B1(n17069), .B2(n16942), .A(n16751), .ZN(P2_U2995) );
  NOR2_X1 U20128 ( .A1(n16753), .A2(n16752), .ZN(n16754) );
  XNOR2_X1 U20129 ( .A(n16755), .B(n16754), .ZN(n17079) );
  INV_X1 U20130 ( .A(n16756), .ZN(n16758) );
  AOI21_X1 U20131 ( .B1(n16765), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16757) );
  NAND2_X1 U20132 ( .A1(n16759), .A2(n16924), .ZN(n16760) );
  NAND2_X1 U20133 ( .A1(n20033), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n17073) );
  OAI211_X1 U20134 ( .C1(n16921), .C2(n16761), .A(n16760), .B(n17073), .ZN(
        n16762) );
  AOI21_X1 U20135 ( .B1(n17076), .B2(n16935), .A(n16762), .ZN(n16763) );
  OAI211_X1 U20136 ( .C1(n17079), .C2(n16942), .A(n16764), .B(n16763), .ZN(
        P2_U2996) );
  XNOR2_X1 U20137 ( .A(n16765), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16771) );
  NAND2_X1 U20138 ( .A1(n20033), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17084) );
  NAND2_X1 U20139 ( .A1(n16930), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16766) );
  OAI211_X1 U20140 ( .C1(n16767), .C2(n16933), .A(n17084), .B(n16766), .ZN(
        n16770) );
  XNOR2_X1 U20141 ( .A(n17092), .B(n17103), .ZN(n16781) );
  INV_X1 U20142 ( .A(n17101), .ZN(n16775) );
  NOR2_X1 U20143 ( .A1(n16877), .A2(n20755), .ZN(n17098) );
  AOI21_X1 U20144 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17098), .ZN(n16772) );
  OAI21_X1 U20145 ( .B1(n16933), .B2(n16773), .A(n16772), .ZN(n16774) );
  AOI21_X1 U20146 ( .B1(n16775), .B2(n16935), .A(n16774), .ZN(n16780) );
  OR2_X1 U20147 ( .A1(n16777), .A2(n16776), .ZN(n17097) );
  NAND3_X1 U20148 ( .A1(n17097), .A2(n16778), .A3(n16899), .ZN(n16779) );
  OAI211_X1 U20149 ( .C1(n16781), .C2(n16911), .A(n16780), .B(n16779), .ZN(
        P2_U2998) );
  INV_X1 U20150 ( .A(n16806), .ZN(n16784) );
  NAND2_X1 U20151 ( .A1(n16792), .A2(n16796), .ZN(n16788) );
  NAND2_X1 U20152 ( .A1(n16786), .A2(n16785), .ZN(n16787) );
  XNOR2_X1 U20153 ( .A(n16788), .B(n16787), .ZN(n17110) );
  NOR2_X1 U20154 ( .A1(n16877), .A2(n16789), .ZN(n17104) );
  AOI21_X1 U20155 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n17104), .ZN(n16790) );
  OAI21_X1 U20156 ( .B1(n16933), .B2(n20045), .A(n16790), .ZN(n16791) );
  INV_X1 U20157 ( .A(n16792), .ZN(n16797) );
  AOI21_X1 U20158 ( .B1(n16794), .B2(n16796), .A(n16793), .ZN(n16795) );
  AOI21_X1 U20159 ( .B1(n16797), .B2(n16796), .A(n16795), .ZN(n17123) );
  NAND2_X1 U20160 ( .A1(n16924), .A2(n16798), .ZN(n16799) );
  NAND2_X1 U20161 ( .A1(n20033), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n17114) );
  OAI211_X1 U20162 ( .C1(n16921), .C2(n16800), .A(n16799), .B(n17114), .ZN(
        n16801) );
  AOI21_X1 U20163 ( .B1(n17119), .B2(n16935), .A(n16801), .ZN(n16803) );
  OAI211_X1 U20164 ( .C1(n17123), .C2(n16942), .A(n16803), .B(n16802), .ZN(
        P2_U3000) );
  NAND2_X1 U20165 ( .A1(n16806), .A2(n16805), .ZN(n16807) );
  XNOR2_X1 U20166 ( .A(n16808), .B(n16807), .ZN(n17134) );
  NOR2_X1 U20167 ( .A1(n16877), .A2(n16809), .ZN(n17127) );
  NOR2_X1 U20168 ( .A1(n16933), .A2(n16810), .ZN(n16811) );
  AOI211_X1 U20169 ( .C1(n16930), .C2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n17127), .B(n16811), .ZN(n16812) );
  OAI21_X1 U20170 ( .B1(n17132), .B2(n17306), .A(n16812), .ZN(n16813) );
  AOI21_X1 U20171 ( .B1(n17134), .B2(n16899), .A(n16813), .ZN(n16814) );
  OAI21_X1 U20172 ( .B1(n17136), .B2(n16911), .A(n16814), .ZN(P2_U3001) );
  OR2_X1 U20173 ( .A1(n10356), .A2(n16816), .ZN(n16817) );
  XNOR2_X1 U20174 ( .A(n9894), .B(n16817), .ZN(n17149) );
  NAND2_X1 U20175 ( .A1(n16823), .A2(n17142), .ZN(n17137) );
  NAND2_X1 U20176 ( .A1(n20033), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n17140) );
  NAND2_X1 U20177 ( .A1(n16930), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16818) );
  OAI211_X1 U20178 ( .C1(n16933), .C2(n16819), .A(n17140), .B(n16818), .ZN(
        n16820) );
  AOI21_X1 U20179 ( .B1(n17146), .B2(n16935), .A(n16820), .ZN(n16821) );
  OAI211_X1 U20180 ( .C1(n17149), .C2(n16942), .A(n16822), .B(n16821), .ZN(
        P2_U3002) );
  INV_X1 U20181 ( .A(n16838), .ZN(n16827) );
  OAI21_X1 U20182 ( .B1(n16854), .B2(n16827), .A(n16826), .ZN(n16831) );
  NAND2_X1 U20183 ( .A1(n16829), .A2(n16828), .ZN(n16830) );
  XNOR2_X1 U20184 ( .A(n16831), .B(n16830), .ZN(n17159) );
  NAND2_X1 U20185 ( .A1(n20033), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n17154) );
  OAI21_X1 U20186 ( .B1(n16921), .B2(n10659), .A(n17154), .ZN(n16832) );
  AOI21_X1 U20187 ( .B1(n16924), .B2(n16833), .A(n16832), .ZN(n16834) );
  OAI21_X1 U20188 ( .B1(n17150), .B2(n17306), .A(n16834), .ZN(n16835) );
  AOI21_X1 U20189 ( .B1(n17159), .B2(n16899), .A(n16835), .ZN(n16836) );
  OAI21_X1 U20190 ( .B1(n17162), .B2(n16911), .A(n16836), .ZN(P2_U3003) );
  NAND2_X1 U20191 ( .A1(n16838), .A2(n16837), .ZN(n16840) );
  NAND2_X1 U20192 ( .A1(n16854), .A2(n16849), .ZN(n16839) );
  XOR2_X1 U20193 ( .A(n16840), .B(n16839), .Z(n17174) );
  NAND2_X1 U20194 ( .A1(n17163), .A2(n16939), .ZN(n16847) );
  OR2_X1 U20195 ( .A1(n16877), .A2(n16841), .ZN(n17166) );
  OAI21_X1 U20196 ( .B1(n16921), .B2(n16842), .A(n17166), .ZN(n16844) );
  NOR2_X1 U20197 ( .A1(n20074), .A2(n17306), .ZN(n16843) );
  AOI211_X1 U20198 ( .C1(n16924), .C2(n16845), .A(n16844), .B(n16843), .ZN(
        n16846) );
  INV_X1 U20199 ( .A(n16849), .ZN(n16853) );
  NAND2_X1 U20200 ( .A1(n16849), .A2(n16848), .ZN(n16850) );
  NAND2_X1 U20201 ( .A1(n16851), .A2(n16850), .ZN(n16852) );
  OAI21_X1 U20202 ( .B1(n16854), .B2(n16853), .A(n16852), .ZN(n17186) );
  INV_X1 U20203 ( .A(n16855), .ZN(n16858) );
  NAND2_X1 U20204 ( .A1(n17175), .A2(n16939), .ZN(n16864) );
  NOR2_X1 U20205 ( .A1(n16877), .A2(n20745), .ZN(n17177) );
  INV_X1 U20206 ( .A(n17177), .ZN(n16860) );
  NAND2_X1 U20207 ( .A1(n16930), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16859) );
  OAI211_X1 U20208 ( .C1(n16933), .C2(n16861), .A(n16860), .B(n16859), .ZN(
        n16862) );
  AOI21_X1 U20209 ( .B1(n17183), .B2(n16935), .A(n16862), .ZN(n16863) );
  OAI211_X1 U20210 ( .C1(n16942), .C2(n17186), .A(n16864), .B(n16863), .ZN(
        P2_U3005) );
  XNOR2_X1 U20211 ( .A(n16866), .B(n16867), .ZN(n16883) );
  AOI22_X1 U20212 ( .A1(n16883), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16866), .B2(n16868), .ZN(n16869) );
  XOR2_X1 U20213 ( .A(n16870), .B(n16869), .Z(n17200) );
  NAND2_X1 U20214 ( .A1(n16872), .A2(n16871), .ZN(n16876) );
  INV_X1 U20215 ( .A(n16885), .ZN(n16874) );
  AOI21_X1 U20216 ( .B1(n16873), .B2(n16884), .A(n16874), .ZN(n16875) );
  XOR2_X1 U20217 ( .A(n16876), .B(n16875), .Z(n17198) );
  NOR2_X1 U20218 ( .A1(n16877), .A2(n20743), .ZN(n17193) );
  NOR2_X1 U20219 ( .A1(n16933), .A2(n16878), .ZN(n16879) );
  AOI211_X1 U20220 ( .C1(n16930), .C2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17193), .B(n16879), .ZN(n16880) );
  OAI21_X1 U20221 ( .B1(n17187), .B2(n17306), .A(n16880), .ZN(n16881) );
  AOI21_X1 U20222 ( .B1(n17198), .B2(n16899), .A(n16881), .ZN(n16882) );
  OAI21_X1 U20223 ( .B1(n17200), .B2(n16911), .A(n16882), .ZN(P2_U3006) );
  XNOR2_X1 U20224 ( .A(n16883), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17212) );
  NAND2_X1 U20225 ( .A1(n16885), .A2(n16884), .ZN(n16886) );
  XNOR2_X1 U20226 ( .A(n16873), .B(n16886), .ZN(n17210) );
  NAND2_X1 U20227 ( .A1(n20033), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n17202) );
  OAI21_X1 U20228 ( .B1(n16921), .B2(n16887), .A(n17202), .ZN(n16888) );
  AOI21_X1 U20229 ( .B1(n16924), .B2(n16889), .A(n16888), .ZN(n16890) );
  OAI21_X1 U20230 ( .B1(n17208), .B2(n17306), .A(n16890), .ZN(n16891) );
  AOI21_X1 U20231 ( .B1(n17210), .B2(n16899), .A(n16891), .ZN(n16892) );
  OAI21_X1 U20232 ( .B1(n17212), .B2(n16911), .A(n16892), .ZN(P2_U3007) );
  XNOR2_X1 U20233 ( .A(n16893), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17224) );
  XNOR2_X1 U20234 ( .A(n16895), .B(n16894), .ZN(n17222) );
  NAND2_X1 U20235 ( .A1(n20033), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n17214) );
  OAI21_X1 U20236 ( .B1(n16921), .B2(n10665), .A(n17214), .ZN(n16896) );
  AOI21_X1 U20237 ( .B1(n16924), .B2(n20061), .A(n16896), .ZN(n16897) );
  OAI21_X1 U20238 ( .B1(n20067), .B2(n17306), .A(n16897), .ZN(n16898) );
  AOI21_X1 U20239 ( .B1(n17222), .B2(n16899), .A(n16898), .ZN(n16900) );
  OAI21_X1 U20240 ( .B1(n17224), .B2(n16911), .A(n16900), .ZN(P2_U3008) );
  XNOR2_X1 U20241 ( .A(n16901), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16902) );
  XNOR2_X1 U20242 ( .A(n16903), .B(n16902), .ZN(n17240) );
  NOR2_X1 U20243 ( .A1(n20051), .A2(n16904), .ZN(n17231) );
  AOI21_X1 U20244 ( .B1(n16930), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n17231), .ZN(n16905) );
  OAI21_X1 U20245 ( .B1(n16933), .B2(n16906), .A(n16905), .ZN(n16913) );
  OAI21_X1 U20246 ( .B1(n16910), .B2(n16908), .A(n16907), .ZN(n16909) );
  NOR2_X1 U20247 ( .A1(n17235), .A2(n16911), .ZN(n16912) );
  AOI211_X1 U20248 ( .C1(n16935), .C2(n17238), .A(n16913), .B(n16912), .ZN(
        n16914) );
  OAI21_X1 U20249 ( .B1(n16942), .B2(n17240), .A(n16914), .ZN(P2_U3009) );
  XNOR2_X1 U20250 ( .A(n16915), .B(n17253), .ZN(n16929) );
  AOI22_X1 U20251 ( .A1(n16929), .A2(n16928), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16915), .ZN(n16918) );
  XNOR2_X1 U20252 ( .A(n16916), .B(n17228), .ZN(n16917) );
  XNOR2_X1 U20253 ( .A(n16918), .B(n16917), .ZN(n17252) );
  XNOR2_X1 U20254 ( .A(n16919), .B(n17228), .ZN(n17250) );
  NAND2_X1 U20255 ( .A1(n20033), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n17246) );
  OAI21_X1 U20256 ( .B1(n16921), .B2(n16920), .A(n17246), .ZN(n16922) );
  AOI21_X1 U20257 ( .B1(n16924), .B2(n16923), .A(n16922), .ZN(n16925) );
  OAI21_X1 U20258 ( .B1(n17242), .B2(n17306), .A(n16925), .ZN(n16926) );
  AOI21_X1 U20259 ( .B1(n17250), .B2(n16939), .A(n16926), .ZN(n16927) );
  OAI21_X1 U20260 ( .B1(n17252), .B2(n16942), .A(n16927), .ZN(P2_U3010) );
  XNOR2_X1 U20261 ( .A(n16929), .B(n16928), .ZN(n17267) );
  AOI22_X1 U20262 ( .A1(n16930), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n20033), .ZN(n16931) );
  OAI21_X1 U20263 ( .B1(n16933), .B2(n16932), .A(n16931), .ZN(n16934) );
  AOI21_X1 U20264 ( .B1(n15957), .B2(n16935), .A(n16934), .ZN(n16941) );
  OR2_X1 U20265 ( .A1(n16937), .A2(n16936), .ZN(n17263) );
  NAND3_X1 U20266 ( .A1(n17263), .A2(n16939), .A3(n17261), .ZN(n16940) );
  OAI211_X1 U20267 ( .C1(n17267), .C2(n16942), .A(n16941), .B(n16940), .ZN(
        P2_U3011) );
  NAND2_X1 U20268 ( .A1(n16943), .A2(n16974), .ZN(n16944) );
  OR2_X1 U20269 ( .A1(n16998), .A2(n16944), .ZN(n16973) );
  NAND2_X1 U20270 ( .A1(n16975), .A2(n16973), .ZN(n16961) );
  XNOR2_X1 U20271 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16947) );
  INV_X1 U20272 ( .A(n16945), .ZN(n16946) );
  OAI21_X1 U20273 ( .B1(n16959), .B2(n16947), .A(n16946), .ZN(n16948) );
  AOI21_X1 U20274 ( .B1(n16961), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16948), .ZN(n16949) );
  OAI21_X1 U20275 ( .B1(n16950), .B2(n17256), .A(n16949), .ZN(n16951) );
  AOI21_X1 U20276 ( .B1(n16952), .B2(n17260), .A(n16951), .ZN(n16955) );
  NAND2_X1 U20277 ( .A1(n16953), .A2(n17262), .ZN(n16954) );
  OAI211_X1 U20278 ( .C1(n16956), .C2(n17266), .A(n16955), .B(n16954), .ZN(
        P2_U3017) );
  INV_X1 U20279 ( .A(n16957), .ZN(n16958) );
  OAI21_X1 U20280 ( .B1(n16959), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16958), .ZN(n16960) );
  AOI21_X1 U20281 ( .B1(n16961), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16960), .ZN(n16962) );
  OAI21_X1 U20282 ( .B1(n16963), .B2(n17256), .A(n16962), .ZN(n16966) );
  NOR2_X1 U20283 ( .A1(n16964), .A2(n17241), .ZN(n16965) );
  NOR2_X1 U20284 ( .A1(n16970), .A2(n17256), .ZN(n16977) );
  INV_X1 U20285 ( .A(n16971), .ZN(n16972) );
  OAI211_X1 U20286 ( .C1(n16975), .C2(n16974), .A(n16973), .B(n16972), .ZN(
        n16976) );
  NAND3_X1 U20287 ( .A1(n16980), .A2(n17262), .A3(n16979), .ZN(n16981) );
  OAI211_X1 U20288 ( .C1(n16983), .C2(n17266), .A(n16982), .B(n16981), .ZN(
        P2_U3019) );
  NAND2_X1 U20289 ( .A1(n16984), .A2(n17260), .ZN(n16990) );
  XNOR2_X1 U20290 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16987) );
  INV_X1 U20291 ( .A(n16985), .ZN(n16986) );
  OAI21_X1 U20292 ( .B1(n16998), .B2(n16987), .A(n16986), .ZN(n16988) );
  AOI21_X1 U20293 ( .B1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17000), .A(
        n16988), .ZN(n16989) );
  OAI211_X1 U20294 ( .C1(n17256), .C2(n16991), .A(n16990), .B(n16989), .ZN(
        n16992) );
  NAND2_X1 U20295 ( .A1(n16995), .A2(n17260), .ZN(n17002) );
  INV_X1 U20296 ( .A(n16996), .ZN(n16997) );
  OAI21_X1 U20297 ( .B1(n16998), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16997), .ZN(n16999) );
  AOI21_X1 U20298 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17000), .A(
        n16999), .ZN(n17001) );
  OAI211_X1 U20299 ( .C1(n17256), .C2(n17003), .A(n17002), .B(n17001), .ZN(
        n17004) );
  AOI21_X1 U20300 ( .B1(n17221), .B2(n17005), .A(n17004), .ZN(n17006) );
  OAI21_X1 U20301 ( .B1(n17234), .B2(n17007), .A(n17006), .ZN(P2_U3021) );
  NAND2_X1 U20302 ( .A1(n17008), .A2(n17260), .ZN(n17013) );
  AOI211_X1 U20303 ( .C1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n17011), .A(
        n17010), .B(n17009), .ZN(n17012) );
  OAI211_X1 U20304 ( .C1(n17256), .C2(n17014), .A(n17013), .B(n17012), .ZN(
        n17015) );
  AOI21_X1 U20305 ( .B1(n17221), .B2(n17016), .A(n17015), .ZN(n17017) );
  OAI21_X1 U20306 ( .B1(n17234), .B2(n17018), .A(n17017), .ZN(P2_U3022) );
  AOI21_X1 U20307 ( .B1(n17049), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17019), .ZN(n17022) );
  OAI211_X1 U20308 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17033), .B(n17020), .ZN(
        n17021) );
  OAI211_X1 U20309 ( .C1(n17023), .C2(n17256), .A(n17022), .B(n17021), .ZN(
        n17027) );
  NOR3_X1 U20310 ( .A1(n17025), .A2(n17024), .A3(n17266), .ZN(n17026) );
  AOI211_X1 U20311 ( .C1(n17028), .C2(n17260), .A(n17027), .B(n17026), .ZN(
        n17029) );
  OAI21_X1 U20312 ( .B1(n17030), .B2(n17234), .A(n17029), .ZN(P2_U3023) );
  AOI21_X1 U20313 ( .B1(n17049), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n17031), .ZN(n17035) );
  NAND2_X1 U20314 ( .A1(n17033), .A2(n17032), .ZN(n17034) );
  OAI211_X1 U20315 ( .C1(n17036), .C2(n17256), .A(n17035), .B(n17034), .ZN(
        n17037) );
  AOI21_X1 U20316 ( .B1(n17038), .B2(n17260), .A(n17037), .ZN(n17041) );
  NAND2_X1 U20317 ( .A1(n17039), .A2(n17221), .ZN(n17040) );
  OAI211_X1 U20318 ( .C1(n17042), .C2(n17234), .A(n17041), .B(n17040), .ZN(
        P2_U3024) );
  NAND2_X1 U20319 ( .A1(n17043), .A2(n17260), .ZN(n17051) );
  OAI21_X1 U20320 ( .B1(n17046), .B2(n17045), .A(n17044), .ZN(n17048) );
  AOI21_X1 U20321 ( .B1(n17049), .B2(n17048), .A(n17047), .ZN(n17050) );
  OAI211_X1 U20322 ( .C1(n17256), .C2(n17052), .A(n17051), .B(n17050), .ZN(
        n17053) );
  AOI21_X1 U20323 ( .B1(n17054), .B2(n17262), .A(n17053), .ZN(n17055) );
  NAND2_X1 U20324 ( .A1(n17057), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17060) );
  INV_X1 U20325 ( .A(n17058), .ZN(n17059) );
  OAI211_X1 U20326 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17061), .A(
        n17060), .B(n17059), .ZN(n17062) );
  AOI21_X1 U20327 ( .B1(n17063), .B2(n12994), .A(n17062), .ZN(n17064) );
  OAI21_X1 U20328 ( .B1(n17065), .B2(n17241), .A(n17064), .ZN(n17066) );
  AOI21_X1 U20329 ( .B1(n17067), .B2(n17262), .A(n17066), .ZN(n17068) );
  OAI21_X1 U20330 ( .B1(n17069), .B2(n17266), .A(n17068), .ZN(P2_U3027) );
  OAI21_X1 U20331 ( .B1(n17071), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17070), .ZN(n17072) );
  OAI211_X1 U20332 ( .C1(n17074), .C2(n17256), .A(n17073), .B(n17072), .ZN(
        n17075) );
  AOI21_X1 U20333 ( .B1(n17076), .B2(n17260), .A(n17075), .ZN(n17077) );
  OAI211_X1 U20334 ( .C1(n17079), .C2(n17266), .A(n17078), .B(n17077), .ZN(
        P2_U3028) );
  INV_X1 U20335 ( .A(n17105), .ZN(n17081) );
  AOI21_X1 U20336 ( .B1(n17103), .B2(n17225), .A(n17096), .ZN(n17095) );
  INV_X1 U20337 ( .A(n17083), .ZN(n17089) );
  OAI21_X1 U20338 ( .B1(n17085), .B2(n17256), .A(n17084), .ZN(n17086) );
  INV_X1 U20339 ( .A(n17086), .ZN(n17088) );
  INV_X1 U20340 ( .A(n17090), .ZN(n17093) );
  AOI21_X1 U20341 ( .B1(n17099), .B2(n12994), .A(n17098), .ZN(n17100) );
  NAND2_X1 U20342 ( .A1(n20039), .A2(n12994), .ZN(n17107) );
  AOI21_X1 U20343 ( .B1(n17105), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17104), .ZN(n17106) );
  OAI211_X1 U20344 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n17108), .A(
        n17107), .B(n17106), .ZN(n17109) );
  NOR2_X1 U20345 ( .A1(n17111), .A2(n17256), .ZN(n17118) );
  NAND2_X1 U20346 ( .A1(n17124), .A2(n17142), .ZN(n17141) );
  NAND2_X1 U20347 ( .A1(n17143), .A2(n17141), .ZN(n17128) );
  AOI21_X1 U20348 ( .B1(n17124), .B2(n10058), .A(n17128), .ZN(n17116) );
  NAND2_X1 U20349 ( .A1(n17112), .A2(n17115), .ZN(n17113) );
  OAI211_X1 U20350 ( .C1(n17116), .C2(n17115), .A(n17114), .B(n17113), .ZN(
        n17117) );
  AOI211_X1 U20351 ( .C1(n17119), .C2(n17260), .A(n17118), .B(n17117), .ZN(
        n17122) );
  NAND2_X1 U20352 ( .A1(n17120), .A2(n17262), .ZN(n17121) );
  OAI211_X1 U20353 ( .C1(n17123), .C2(n17266), .A(n17122), .B(n17121), .ZN(
        P2_U3032) );
  INV_X1 U20354 ( .A(n17124), .ZN(n17125) );
  NOR3_X1 U20355 ( .A1(n17125), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n17142), .ZN(n17126) );
  AOI211_X1 U20356 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n17128), .A(
        n17127), .B(n17126), .ZN(n17131) );
  NAND2_X1 U20357 ( .A1(n17129), .A2(n12994), .ZN(n17130) );
  OAI211_X1 U20358 ( .C1(n17132), .C2(n17241), .A(n17131), .B(n17130), .ZN(
        n17133) );
  AOI21_X1 U20359 ( .B1(n17134), .B2(n17221), .A(n17133), .ZN(n17135) );
  NAND3_X1 U20360 ( .A1(n17138), .A2(n17262), .A3(n17137), .ZN(n17148) );
  NOR2_X1 U20361 ( .A1(n17139), .A2(n17256), .ZN(n17145) );
  OAI211_X1 U20362 ( .C1(n17143), .C2(n17142), .A(n17141), .B(n17140), .ZN(
        n17144) );
  AOI211_X1 U20363 ( .C1(n17146), .C2(n17260), .A(n17145), .B(n17144), .ZN(
        n17147) );
  OAI211_X1 U20364 ( .C1(n17149), .C2(n17266), .A(n17148), .B(n17147), .ZN(
        P2_U3034) );
  INV_X1 U20365 ( .A(n17150), .ZN(n17158) );
  NOR2_X1 U20366 ( .A1(n17151), .A2(n17256), .ZN(n17157) );
  OAI211_X1 U20367 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17164), .B(n17152), .ZN(
        n17153) );
  OAI211_X1 U20368 ( .C1(n17168), .C2(n17155), .A(n17154), .B(n17153), .ZN(
        n17156) );
  AOI211_X1 U20369 ( .C1(n17158), .C2(n17260), .A(n17157), .B(n17156), .ZN(
        n17161) );
  NAND2_X1 U20370 ( .A1(n17159), .A2(n17221), .ZN(n17160) );
  OAI211_X1 U20371 ( .C1(n17162), .C2(n17234), .A(n17161), .B(n17160), .ZN(
        P2_U3035) );
  NAND2_X1 U20372 ( .A1(n17163), .A2(n17262), .ZN(n17173) );
  NAND2_X1 U20373 ( .A1(n17164), .A2(n17167), .ZN(n17165) );
  OAI211_X1 U20374 ( .C1(n17168), .C2(n17167), .A(n17166), .B(n17165), .ZN(
        n17170) );
  NOR2_X1 U20375 ( .A1(n20074), .A2(n17241), .ZN(n17169) );
  AOI211_X1 U20376 ( .C1(n12994), .C2(n17171), .A(n17170), .B(n17169), .ZN(
        n17172) );
  OAI211_X1 U20377 ( .C1(n17174), .C2(n17266), .A(n17173), .B(n17172), .ZN(
        P2_U3036) );
  NAND2_X1 U20378 ( .A1(n17175), .A2(n17262), .ZN(n17185) );
  INV_X1 U20379 ( .A(n17176), .ZN(n17178) );
  AOI21_X1 U20380 ( .B1(n17178), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17177), .ZN(n17180) );
  OAI211_X1 U20381 ( .C1(n17181), .C2(n17256), .A(n17180), .B(n17179), .ZN(
        n17182) );
  AOI21_X1 U20382 ( .B1(n17183), .B2(n17260), .A(n17182), .ZN(n17184) );
  OAI211_X1 U20383 ( .C1(n17186), .C2(n17266), .A(n17185), .B(n17184), .ZN(
        P2_U3037) );
  NOR2_X1 U20384 ( .A1(n17187), .A2(n17241), .ZN(n17197) );
  INV_X1 U20385 ( .A(n17216), .ZN(n17201) );
  INV_X1 U20386 ( .A(n17188), .ZN(n17189) );
  AOI211_X1 U20387 ( .C1(n17191), .C2(n17190), .A(n17189), .B(n17204), .ZN(
        n17192) );
  AOI211_X1 U20388 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n17201), .A(
        n17193), .B(n17192), .ZN(n17194) );
  OAI21_X1 U20389 ( .B1(n17256), .B2(n17195), .A(n17194), .ZN(n17196) );
  AOI211_X1 U20390 ( .C1(n17198), .C2(n17221), .A(n17197), .B(n17196), .ZN(
        n17199) );
  OAI21_X1 U20391 ( .B1(n17200), .B2(n17234), .A(n17199), .ZN(P2_U3038) );
  NAND2_X1 U20392 ( .A1(n17201), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17203) );
  OAI211_X1 U20393 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17204), .A(
        n17203), .B(n17202), .ZN(n17205) );
  AOI21_X1 U20394 ( .B1(n12994), .B2(n17206), .A(n17205), .ZN(n17207) );
  OAI21_X1 U20395 ( .B1(n17208), .B2(n17241), .A(n17207), .ZN(n17209) );
  AOI21_X1 U20396 ( .B1(n17210), .B2(n17221), .A(n17209), .ZN(n17211) );
  OAI21_X1 U20397 ( .B1(n17212), .B2(n17234), .A(n17211), .ZN(P2_U3039) );
  AOI21_X1 U20398 ( .B1(n17254), .B2(n17213), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17215) );
  OAI21_X1 U20399 ( .B1(n17216), .B2(n17215), .A(n17214), .ZN(n17217) );
  AOI21_X1 U20400 ( .B1(n12994), .B2(n17218), .A(n17217), .ZN(n17219) );
  OAI21_X1 U20401 ( .B1(n20067), .B2(n17241), .A(n17219), .ZN(n17220) );
  AOI21_X1 U20402 ( .B1(n17222), .B2(n17221), .A(n17220), .ZN(n17223) );
  OAI21_X1 U20403 ( .B1(n17224), .B2(n17234), .A(n17223), .ZN(P2_U3040) );
  INV_X1 U20404 ( .A(n17255), .ZN(n17227) );
  NAND2_X1 U20405 ( .A1(n17225), .A2(n17253), .ZN(n17226) );
  NAND2_X1 U20406 ( .A1(n17227), .A2(n17226), .ZN(n17243) );
  NAND2_X1 U20407 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17254), .ZN(
        n17245) );
  AOI221_X1 U20408 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n17229), .C2(n17228), .A(
        n17245), .ZN(n17230) );
  AOI211_X1 U20409 ( .C1(n17243), .C2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n17231), .B(n17230), .ZN(n17232) );
  OAI21_X1 U20410 ( .B1(n17233), .B2(n17256), .A(n17232), .ZN(n17237) );
  NOR2_X1 U20411 ( .A1(n17235), .A2(n17234), .ZN(n17236) );
  AOI211_X1 U20412 ( .C1(n17238), .C2(n17260), .A(n17237), .B(n17236), .ZN(
        n17239) );
  OAI21_X1 U20413 ( .B1(n17266), .B2(n17240), .A(n17239), .ZN(P2_U3041) );
  NOR2_X1 U20414 ( .A1(n17242), .A2(n17241), .ZN(n17249) );
  INV_X1 U20415 ( .A(n17243), .ZN(n17244) );
  MUX2_X1 U20416 ( .A(n17245), .B(n17244), .S(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n17247) );
  OAI211_X1 U20417 ( .C1(n17256), .C2(n20086), .A(n17247), .B(n17246), .ZN(
        n17248) );
  AOI211_X1 U20418 ( .C1(n17250), .C2(n17262), .A(n17249), .B(n17248), .ZN(
        n17251) );
  OAI21_X1 U20419 ( .B1(n17252), .B2(n17266), .A(n17251), .ZN(P2_U3042) );
  MUX2_X1 U20420 ( .A(n17255), .B(n17254), .S(n17253), .Z(n17259) );
  OAI22_X1 U20421 ( .A1(n17257), .A2(n17256), .B1(n20736), .B2(n20051), .ZN(
        n17258) );
  AOI211_X1 U20422 ( .C1(n15957), .C2(n17260), .A(n17259), .B(n17258), .ZN(
        n17265) );
  NAND3_X1 U20423 ( .A1(n17263), .A2(n17262), .A3(n17261), .ZN(n17264) );
  OAI211_X1 U20424 ( .C1(n17267), .C2(n17266), .A(n17265), .B(n17264), .ZN(
        P2_U3043) );
  INV_X1 U20425 ( .A(n17268), .ZN(n20823) );
  AOI22_X1 U20426 ( .A1(n17271), .A2(n17270), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n17269), .ZN(n17272) );
  OAI21_X1 U20427 ( .B1(n20133), .B2(n20823), .A(n17272), .ZN(n17276) );
  NAND2_X1 U20428 ( .A1(n20835), .A2(n17273), .ZN(n17274) );
  NAND2_X1 U20429 ( .A1(n17274), .A2(n17610), .ZN(n17275) );
  AND2_X1 U20430 ( .A1(n17275), .A2(n20555), .ZN(n20832) );
  MUX2_X1 U20431 ( .A(n17276), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(
        n20832), .Z(P2_U3605) );
  INV_X1 U20432 ( .A(n17277), .ZN(n17278) );
  MUX2_X1 U20433 ( .A(n17278), .B(n17327), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n17279) );
  AOI21_X1 U20434 ( .B1(n17281), .B2(n17280), .A(n17279), .ZN(n17314) );
  OAI222_X1 U20435 ( .A1(n20797), .A2(n17283), .B1(n20803), .B2(n17314), .C1(
        n17365), .C2(n17282), .ZN(n17284) );
  MUX2_X1 U20436 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n17284), .S(
        n17298), .Z(P2_U3601) );
  OR2_X1 U20437 ( .A1(n14213), .A2(n17319), .ZN(n17296) );
  NAND2_X1 U20438 ( .A1(n9919), .A2(n17285), .ZN(n17332) );
  OAI21_X1 U20439 ( .B1(n16378), .B2(n11015), .A(n11252), .ZN(n17294) );
  NAND2_X1 U20440 ( .A1(n17347), .A2(n17346), .ZN(n17323) );
  NAND2_X1 U20441 ( .A1(n17286), .A2(n17335), .ZN(n17321) );
  XNOR2_X1 U20442 ( .A(n17321), .B(n11015), .ZN(n17287) );
  NAND2_X1 U20443 ( .A1(n17323), .A2(n17287), .ZN(n17292) );
  AOI21_X1 U20444 ( .B1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17288) );
  NOR2_X1 U20445 ( .A1(n17289), .A2(n17288), .ZN(n17290) );
  NAND2_X1 U20446 ( .A1(n17327), .A2(n17290), .ZN(n17291) );
  NAND2_X1 U20447 ( .A1(n17292), .A2(n17291), .ZN(n17293) );
  AOI21_X1 U20448 ( .B1(n17332), .B2(n17294), .A(n17293), .ZN(n17295) );
  NAND2_X1 U20449 ( .A1(n17296), .A2(n17295), .ZN(n17313) );
  INV_X1 U20450 ( .A(n17313), .ZN(n17297) );
  OAI22_X1 U20451 ( .A1(n20199), .A2(n20797), .B1(n17297), .B2(n20803), .ZN(
        n17299) );
  MUX2_X1 U20452 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17299), .S(
        n17298), .Z(P2_U3596) );
  OR2_X1 U20453 ( .A1(n20199), .A2(n20481), .ZN(n20656) );
  NAND3_X1 U20454 ( .A1(n20831), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20550) );
  OAI21_X1 U20455 ( .B1(n20656), .B2(n20327), .A(n20550), .ZN(n17304) );
  INV_X1 U20456 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n17300) );
  INV_X1 U20457 ( .A(n20550), .ZN(n17301) );
  NAND2_X1 U20458 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n17301), .ZN(
        n20612) );
  AOI21_X1 U20459 ( .B1(n17302), .B2(n20612), .A(n20555), .ZN(n17303) );
  INV_X1 U20460 ( .A(n20605), .ZN(n20585) );
  INV_X1 U20461 ( .A(n20175), .ZN(n20177) );
  OAI22_X1 U20462 ( .A1(n16511), .A2(n20177), .B1(n16509), .B2(n20179), .ZN(
        n20698) );
  INV_X1 U20463 ( .A(n20644), .ZN(n20581) );
  AOI22_X1 U20464 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20175), .ZN(n20703) );
  INV_X1 U20465 ( .A(n20703), .ZN(n20572) );
  AOI22_X1 U20466 ( .A1(n20604), .A2(n20698), .B1(n20581), .B2(n20572), .ZN(
        n17311) );
  INV_X1 U20467 ( .A(n20612), .ZN(n20615) );
  NOR2_X2 U20468 ( .A1(n17309), .A2(n20555), .ZN(n20697) );
  NAND2_X1 U20469 ( .A1(n20660), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20151) );
  NOR2_X2 U20470 ( .A1(n13989), .A2(n20151), .ZN(n20696) );
  AOI22_X1 U20471 ( .A1(n20602), .A2(n20697), .B1(n20615), .B2(n20696), .ZN(
        n17310) );
  OAI211_X1 U20472 ( .C1(n20585), .C2(n17312), .A(n17311), .B(n17310), .ZN(
        P2_U3158) );
  MUX2_X1 U20473 ( .A(n17313), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17336), .Z(n17344) );
  INV_X1 U20474 ( .A(n17344), .ZN(n17341) );
  INV_X1 U20475 ( .A(n20253), .ZN(n20515) );
  OAI22_X1 U20476 ( .A1(n17315), .A2(n20515), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17317) );
  AOI21_X1 U20477 ( .B1(n17315), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17314), .ZN(n17316) );
  OAI21_X1 U20478 ( .B1(n17317), .B2(n17316), .A(n17361), .ZN(n17318) );
  INV_X1 U20479 ( .A(n17318), .ZN(n17338) );
  OR2_X1 U20480 ( .A1(n17320), .A2(n17319), .ZN(n17334) );
  INV_X1 U20481 ( .A(n17322), .ZN(n17331) );
  NAND2_X1 U20482 ( .A1(n17323), .A2(n17322), .ZN(n17329) );
  INV_X1 U20483 ( .A(n17324), .ZN(n17325) );
  OAI21_X1 U20484 ( .B1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n21769), .A(
        n17325), .ZN(n17326) );
  NAND2_X1 U20485 ( .A1(n17327), .A2(n17326), .ZN(n17328) );
  NAND2_X1 U20486 ( .A1(n17329), .A2(n17328), .ZN(n17330) );
  AOI21_X1 U20487 ( .B1(n17332), .B2(n17331), .A(n17330), .ZN(n17333) );
  AND2_X1 U20488 ( .A1(n17334), .A2(n17333), .ZN(n20796) );
  AND2_X1 U20489 ( .A1(n17336), .A2(n17335), .ZN(n17337) );
  AOI21_X1 U20490 ( .B1(n20796), .B2(n17361), .A(n17337), .ZN(n17343) );
  OAI21_X1 U20491 ( .B1(n17338), .B2(n20821), .A(n17343), .ZN(n17339) );
  NAND2_X1 U20492 ( .A1(n17338), .A2(n20821), .ZN(n17340) );
  AND3_X1 U20493 ( .A1(n17341), .A2(n17339), .A3(n17340), .ZN(n17342) );
  OAI22_X1 U20494 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17342), .B1(
        n17341), .B2(n17340), .ZN(n17364) );
  NAND2_X1 U20495 ( .A1(n17344), .A2(n17343), .ZN(n17360) );
  MUX2_X1 U20496 ( .A(n17347), .B(n17346), .S(n17345), .Z(n17351) );
  NAND2_X1 U20497 ( .A1(n17349), .A2(n17348), .ZN(n17350) );
  NAND2_X1 U20498 ( .A1(n17351), .A2(n17350), .ZN(n20834) );
  NOR2_X1 U20499 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n17356) );
  INV_X1 U20500 ( .A(n17352), .ZN(n17353) );
  NAND2_X1 U20501 ( .A1(n17353), .A2(n20851), .ZN(n17354) );
  OAI211_X1 U20502 ( .C1(n17357), .C2(n17356), .A(n17355), .B(n17354), .ZN(
        n17358) );
  NOR2_X1 U20503 ( .A1(n20834), .A2(n17358), .ZN(n17359) );
  OAI211_X1 U20504 ( .C1(n17362), .C2(n17361), .A(n17360), .B(n17359), .ZN(
        n17363) );
  AOI21_X1 U20505 ( .B1(n17364), .B2(n17534), .A(n17363), .ZN(n17618) );
  NAND2_X1 U20506 ( .A1(n17618), .A2(n17365), .ZN(n17370) );
  NOR2_X1 U20507 ( .A1(n17366), .A2(n17300), .ZN(n20848) );
  OAI21_X1 U20508 ( .B1(n17368), .B2(n17367), .A(n20848), .ZN(n17369) );
  NOR3_X1 U20509 ( .A1(n10286), .A2(n20844), .A3(n20803), .ZN(n17371) );
  NOR2_X1 U20510 ( .A1(n17372), .A2(n17371), .ZN(n17374) );
  NOR2_X1 U20511 ( .A1(n10286), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17606) );
  OAI211_X1 U20512 ( .C1(n17612), .C2(n17606), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n20844), .ZN(n17373) );
  OAI211_X1 U20513 ( .C1(n17612), .C2(n17374), .A(n17373), .B(n20062), .ZN(
        P2_U3177) );
  INV_X1 U20514 ( .A(n17612), .ZN(n17378) );
  INV_X1 U20515 ( .A(n17375), .ZN(n17377) );
  OAI211_X1 U20516 ( .C1(n17378), .C2(n20814), .A(n17377), .B(n17376), .ZN(
        P2_U3593) );
  INV_X1 U20517 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n18096) );
  AOI22_X1 U20518 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U20519 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U20520 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U20521 ( .A1(n18315), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17379) );
  NAND4_X1 U20522 ( .A1(n17382), .A2(n17381), .A3(n17380), .A4(n17379), .ZN(
        n17388) );
  AOI22_X1 U20523 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U20524 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U20525 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U20526 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17383) );
  NAND4_X1 U20527 ( .A1(n17386), .A2(n17385), .A3(n17384), .A4(n17383), .ZN(
        n17387) );
  NOR2_X1 U20528 ( .A1(n17388), .A2(n17387), .ZN(n18131) );
  AOI22_X1 U20529 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20530 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20531 ( .A1(n12808), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20532 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17389) );
  NAND4_X1 U20533 ( .A1(n17392), .A2(n17391), .A3(n17390), .A4(n17389), .ZN(
        n17398) );
  AOI22_X1 U20534 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U20535 ( .A1(n18314), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20536 ( .A1(n18333), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U20537 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17393) );
  NAND4_X1 U20538 ( .A1(n17396), .A2(n17395), .A3(n17394), .A4(n17393), .ZN(
        n17397) );
  NOR2_X1 U20539 ( .A1(n17398), .A2(n17397), .ZN(n18141) );
  AOI22_X1 U20540 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18334), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n18322), .ZN(n17402) );
  AOI22_X1 U20541 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18341), .ZN(n17401) );
  AOI22_X1 U20542 ( .A1(n18314), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17456), .ZN(n17400) );
  AOI22_X1 U20543 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18315), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18333), .ZN(n17399) );
  NAND4_X1 U20544 ( .A1(n17402), .A2(n17401), .A3(n17400), .A4(n17399), .ZN(
        n17408) );
  AOI22_X1 U20545 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17439), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n18312), .ZN(n17406) );
  AOI22_X1 U20546 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U20547 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18340), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17404) );
  AOI22_X1 U20548 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18297), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17403) );
  NAND4_X1 U20549 ( .A1(n17406), .A2(n17405), .A3(n17404), .A4(n17403), .ZN(
        n17407) );
  NOR2_X1 U20550 ( .A1(n17408), .A2(n17407), .ZN(n18149) );
  AOI22_X1 U20551 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20552 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17417) );
  INV_X1 U20553 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n21848) );
  AOI22_X1 U20554 ( .A1(n18314), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20555 ( .B1(n9732), .B2(n21848), .A(n17409), .ZN(n17415) );
  AOI22_X1 U20556 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U20557 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U20558 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U20559 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17410) );
  NAND4_X1 U20560 ( .A1(n17413), .A2(n17412), .A3(n17411), .A4(n17410), .ZN(
        n17414) );
  AOI211_X1 U20561 ( .C1(n18320), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17415), .B(n17414), .ZN(n17416) );
  NAND3_X1 U20562 ( .A1(n17418), .A2(n17417), .A3(n17416), .ZN(n18154) );
  AOI22_X1 U20563 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20564 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17427) );
  INV_X1 U20565 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18357) );
  AOI22_X1 U20566 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17419) );
  OAI21_X1 U20567 ( .B1(n9747), .B2(n18357), .A(n17419), .ZN(n17425) );
  AOI22_X1 U20568 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17423) );
  AOI22_X1 U20569 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20570 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17421) );
  AOI22_X1 U20571 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17420) );
  NAND4_X1 U20572 ( .A1(n17423), .A2(n17422), .A3(n17421), .A4(n17420), .ZN(
        n17424) );
  AOI211_X1 U20573 ( .C1(n18320), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n17425), .B(n17424), .ZN(n17426) );
  NAND3_X1 U20574 ( .A1(n17428), .A2(n17427), .A3(n17426), .ZN(n18155) );
  NAND2_X1 U20575 ( .A1(n18154), .A2(n18155), .ZN(n18153) );
  NOR2_X1 U20576 ( .A1(n18149), .A2(n18153), .ZN(n18146) );
  AOI22_X1 U20577 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U20578 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U20579 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17429) );
  OAI21_X1 U20580 ( .B1(n18106), .B2(n18381), .A(n17429), .ZN(n17435) );
  AOI22_X1 U20581 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17433) );
  AOI22_X1 U20582 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20583 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20584 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17430) );
  NAND4_X1 U20585 ( .A1(n17433), .A2(n17432), .A3(n17431), .A4(n17430), .ZN(
        n17434) );
  AOI211_X1 U20586 ( .C1(n18345), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n17435), .B(n17434), .ZN(n17436) );
  NAND3_X1 U20587 ( .A1(n17438), .A2(n17437), .A3(n17436), .ZN(n18145) );
  NAND2_X1 U20588 ( .A1(n18146), .A2(n18145), .ZN(n18144) );
  NOR2_X1 U20589 ( .A1(n18141), .A2(n18144), .ZN(n18138) );
  AOI22_X1 U20590 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17439), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U20591 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U20592 ( .A1(n18333), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17440) );
  OAI21_X1 U20593 ( .B1(n18106), .B2(n18370), .A(n17440), .ZN(n17446) );
  AOI22_X1 U20594 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20595 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20596 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U20597 ( .A1(n12808), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17441) );
  NAND4_X1 U20598 ( .A1(n17444), .A2(n17443), .A3(n17442), .A4(n17441), .ZN(
        n17445) );
  AOI211_X1 U20599 ( .C1(n18344), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n17446), .B(n17445), .ZN(n17447) );
  NAND3_X1 U20600 ( .A1(n17449), .A2(n17448), .A3(n17447), .ZN(n18137) );
  NAND2_X1 U20601 ( .A1(n18138), .A2(n18137), .ZN(n18136) );
  XNOR2_X1 U20602 ( .A(n18131), .B(n18136), .ZN(n18412) );
  NAND3_X1 U20603 ( .A1(n18130), .A2(P3_EBX_REG_28__SCAN_IN), .A3(n18379), 
        .ZN(n17450) );
  OAI221_X1 U20604 ( .B1(n18130), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n18379), 
        .C2(n18412), .A(n17450), .ZN(P3_U2675) );
  AOI22_X1 U20605 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20606 ( .A1(n12808), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U20607 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20608 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17451) );
  NAND4_X1 U20609 ( .A1(n17454), .A2(n17453), .A3(n17452), .A4(n17451), .ZN(
        n17462) );
  AOI22_X1 U20610 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20611 ( .A1(n18333), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17459) );
  AOI22_X1 U20612 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U20613 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17439), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17457) );
  NAND4_X1 U20614 ( .A1(n17460), .A2(n17459), .A3(n17458), .A4(n17457), .ZN(
        n17461) );
  NOR2_X1 U20615 ( .A1(n17462), .A2(n17461), .ZN(n18485) );
  NAND2_X1 U20616 ( .A1(n18379), .A2(n17463), .ZN(n18282) );
  INV_X1 U20617 ( .A(n18282), .ZN(n18295) );
  NAND2_X1 U20618 ( .A1(n19375), .A2(n18390), .ZN(n18385) );
  INV_X1 U20619 ( .A(n18385), .ZN(n18386) );
  NAND2_X1 U20620 ( .A1(n18386), .A2(n17925), .ZN(n18281) );
  NAND2_X1 U20621 ( .A1(n17465), .A2(n17464), .ZN(n18308) );
  NOR3_X1 U20622 ( .A1(n17466), .A2(n18281), .A3(n18308), .ZN(n17467) );
  AOI22_X1 U20623 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18295), .B1(
        P3_EBX_REG_12__SCAN_IN), .B2(n17467), .ZN(n17468) );
  OAI21_X1 U20624 ( .B1(n18485), .B2(n18379), .A(n17468), .ZN(P3_U2690) );
  INV_X1 U20625 ( .A(n19685), .ZN(n19629) );
  NAND3_X1 U20626 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19935)
         );
  INV_X1 U20627 ( .A(n19935), .ZN(n17469) );
  NAND3_X1 U20628 ( .A1(n17484), .A2(n9747), .A3(n19824), .ZN(n19337) );
  INV_X1 U20629 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19338) );
  NOR2_X1 U20630 ( .A1(n19338), .A2(n19935), .ZN(n17482) );
  AOI211_X1 U20631 ( .C1(n17469), .C2(n19337), .A(n19632), .B(n17482), .ZN(
        n17475) );
  INV_X1 U20632 ( .A(n17475), .ZN(n19344) );
  NAND2_X1 U20633 ( .A1(n19629), .A2(n19344), .ZN(n17471) );
  NAND2_X1 U20634 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19797), .ZN(n19339) );
  NAND2_X1 U20635 ( .A1(n19339), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19422) );
  NAND2_X1 U20636 ( .A1(n18981), .A2(n17470), .ZN(n17473) );
  NAND2_X1 U20637 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19346) );
  AOI21_X1 U20638 ( .B1(n17473), .B2(n19346), .A(n17475), .ZN(n17476) );
  OAI22_X1 U20639 ( .A1(n17471), .A2(n19422), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17476), .ZN(n17472) );
  INV_X1 U20640 ( .A(n17472), .ZN(P3_U2864) );
  NOR2_X1 U20641 ( .A1(n19799), .A2(n19803), .ZN(n19513) );
  AOI22_X1 U20642 ( .A1(n19513), .A2(n19339), .B1(n19937), .B2(n17473), .ZN(
        n17474) );
  NOR2_X1 U20643 ( .A1(n17475), .A2(n17474), .ZN(n19343) );
  AOI22_X1 U20644 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17476), .B1(
        n19685), .B2(n19344), .ZN(n19342) );
  AOI22_X1 U20645 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19343), .B1(
        n19342), .B2(n19803), .ZN(P3_U2865) );
  NOR4_X1 U20646 ( .A1(n19990), .A2(n17478), .A3(n18545), .A4(n19986), .ZN(
        n17480) );
  INV_X1 U20647 ( .A(n19802), .ZN(n19823) );
  NOR2_X1 U20648 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19937), .ZN(n19348) );
  INV_X1 U20649 ( .A(n19968), .ZN(n19965) );
  AOI21_X1 U20650 ( .B1(n17484), .B2(n19824), .A(n17483), .ZN(n19819) );
  NAND3_X1 U20651 ( .A1(n19965), .A2(n20002), .A3(n19819), .ZN(n17485) );
  OAI21_X1 U20652 ( .B1(n19965), .B2(n19824), .A(n17485), .ZN(P3_U3284) );
  INV_X1 U20653 ( .A(n19214), .ZN(n17487) );
  INV_X1 U20654 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n19022) );
  AOI211_X1 U20655 ( .C1(n17487), .C2(n19022), .A(n19325), .B(n17486), .ZN(
        n17638) );
  OAI21_X1 U20656 ( .B1(n19317), .B2(n17638), .A(n17488), .ZN(n17489) );
  AOI21_X1 U20657 ( .B1(n19321), .B2(n18655), .A(n17489), .ZN(n17493) );
  NOR2_X1 U20658 ( .A1(n9755), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17647) );
  AOI21_X1 U20659 ( .B1(n17636), .B2(n17490), .A(n17647), .ZN(n17491) );
  XNOR2_X1 U20660 ( .A(n17491), .B(n17631), .ZN(n17628) );
  AOI22_X1 U20661 ( .A1(n19317), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n19239), 
        .B2(n17628), .ZN(n17492) );
  OAI221_X1 U20662 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17494), 
        .C1(n17631), .C2(n17493), .A(n17492), .ZN(P3_U2833) );
  INV_X1 U20663 ( .A(n17495), .ZN(n17496) );
  OAI211_X1 U20664 ( .C1(n17498), .C2(n17497), .A(n17496), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17503) );
  INV_X1 U20665 ( .A(n17503), .ZN(n17501) );
  OAI22_X1 U20666 ( .A1(n17501), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n17500), .B2(n17499), .ZN(n17502) );
  OAI21_X1 U20667 ( .B1(n17503), .B2(n21468), .A(n17502), .ZN(n17506) );
  INV_X1 U20668 ( .A(n17504), .ZN(n17505) );
  AOI222_X1 U20669 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17506), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17505), .C1(n17506), 
        .C2(n17505), .ZN(n17508) );
  OR2_X1 U20670 ( .A1(n17508), .A2(n17507), .ZN(n17509) );
  AOI22_X1 U20671 ( .A1(n21385), .A2(n17509), .B1(n17508), .B2(n17507), .ZN(
        n17516) );
  OR2_X1 U20672 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n17513) );
  INV_X1 U20673 ( .A(n17510), .ZN(n17512) );
  AOI211_X1 U20674 ( .C1(n17514), .C2(n17513), .A(n17512), .B(n17511), .ZN(
        n17515) );
  OAI21_X1 U20675 ( .B1(n17516), .B2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n17515), .ZN(n17517) );
  NOR3_X1 U20676 ( .A1(n17519), .A2(n17518), .A3(n17517), .ZN(n17533) );
  NOR3_X1 U20677 ( .A1(n17522), .A2(n17521), .A3(n17520), .ZN(n17523) );
  AOI221_X1 U20678 ( .B1(n17525), .B2(n17524), .C1(n21653), .C2(n17524), .A(
        n17523), .ZN(n17599) );
  AOI21_X1 U20679 ( .B1(n17533), .B2(n17599), .A(n21645), .ZN(n17605) );
  OAI21_X1 U20680 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21653), .A(n17605), 
        .ZN(n17603) );
  INV_X1 U20681 ( .A(n17599), .ZN(n17526) );
  OAI222_X1 U20682 ( .A1(n17530), .A2(n17529), .B1(n17603), .B2(n17528), .C1(
        n17527), .C2(n17526), .ZN(n17531) );
  OAI211_X1 U20683 ( .C1(n17533), .C2(n20866), .A(n17532), .B(n17531), .ZN(
        P1_U3161) );
  INV_X1 U20684 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17723) );
  NOR2_X1 U20685 ( .A1(n20985), .A2(n17723), .ZN(P1_U2905) );
  INV_X1 U20686 ( .A(n20832), .ZN(n20829) );
  NOR2_X1 U20687 ( .A1(n17534), .A2(n20829), .ZN(P2_U3047) );
  NAND2_X1 U20688 ( .A1(n19375), .A2(n18392), .ZN(n18539) );
  AOI22_X1 U20689 ( .A1(n18538), .A2(BUF2_REG_0__SCAN_IN), .B1(n18537), .B2(
        n9733), .ZN(n17538) );
  OAI221_X1 U20690 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n18539), .C1(n18594), 
        .C2(n18392), .A(n17538), .ZN(P3_U2735) );
  AOI22_X1 U20691 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n21051), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17545) );
  NAND2_X1 U20692 ( .A1(n17540), .A2(n17539), .ZN(n17541) );
  XNOR2_X1 U20693 ( .A(n17542), .B(n17541), .ZN(n17572) );
  INV_X1 U20694 ( .A(n20908), .ZN(n17543) );
  AOI22_X1 U20695 ( .A1(n21001), .A2(n17572), .B1(n17543), .B2(n21000), .ZN(
        n17544) );
  OAI211_X1 U20696 ( .C1(n21006), .C2(n20906), .A(n17545), .B(n17544), .ZN(
        P1_U2992) );
  AOI22_X1 U20697 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n21051), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17550) );
  XNOR2_X1 U20698 ( .A(n17546), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17547) );
  XNOR2_X1 U20699 ( .A(n17548), .B(n17547), .ZN(n17578) );
  AOI22_X1 U20700 ( .A1(n20971), .A2(n21000), .B1(n17578), .B2(n21001), .ZN(
        n17549) );
  OAI211_X1 U20701 ( .C1(n21006), .C2(n20915), .A(n17550), .B(n17549), .ZN(
        P1_U2993) );
  AOI22_X1 U20702 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n21051), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n17555) );
  XNOR2_X1 U20703 ( .A(n17551), .B(n21018), .ZN(n20993) );
  NAND2_X1 U20704 ( .A1(n20993), .A2(n20994), .ZN(n20998) );
  OAI21_X1 U20705 ( .B1(n21018), .B2(n10364), .A(n20998), .ZN(n17553) );
  XNOR2_X1 U20706 ( .A(n12420), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17552) );
  XNOR2_X1 U20707 ( .A(n17553), .B(n17552), .ZN(n17588) );
  AOI22_X1 U20708 ( .A1(n17588), .A2(n21001), .B1(n21000), .B2(n20931), .ZN(
        n17554) );
  OAI211_X1 U20709 ( .C1(n21006), .C2(n20934), .A(n17555), .B(n17554), .ZN(
        P1_U2994) );
  NAND2_X1 U20710 ( .A1(n21011), .A2(n17585), .ZN(n17584) );
  OAI21_X1 U20711 ( .B1(n17556), .B2(n21008), .A(n21030), .ZN(n17557) );
  AOI21_X1 U20712 ( .B1(n17559), .B2(n17558), .A(n17557), .ZN(n17586) );
  OAI21_X1 U20713 ( .B1(n17560), .B2(n17584), .A(n17586), .ZN(n17579) );
  AOI21_X1 U20714 ( .B1(n21843), .B2(n17561), .A(n17579), .ZN(n17574) );
  AOI22_X1 U20715 ( .A1(n21051), .A2(P1_REIP_REG_8__SCAN_IN), .B1(n21027), 
        .B2(n17562), .ZN(n17568) );
  NAND2_X1 U20716 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17563), .ZN(
        n17576) );
  AOI221_X1 U20717 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n17569), .C2(n17575), .A(
        n17576), .ZN(n17566) );
  AND2_X1 U20718 ( .A1(n17564), .A2(n21042), .ZN(n17565) );
  NOR2_X1 U20719 ( .A1(n17566), .A2(n17565), .ZN(n17567) );
  OAI211_X1 U20720 ( .C1(n17574), .C2(n17569), .A(n17568), .B(n17567), .ZN(
        P1_U3023) );
  OAI22_X1 U20721 ( .A1(n21054), .A2(n20912), .B1(n21674), .B2(n17570), .ZN(
        n17571) );
  AOI21_X1 U20722 ( .B1(n17572), .B2(n21042), .A(n17571), .ZN(n17573) );
  OAI221_X1 U20723 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17576), .C1(
        n17575), .C2(n17574), .A(n17573), .ZN(P1_U3024) );
  AOI21_X1 U20724 ( .B1(n17577), .B2(n14955), .A(n9926), .ZN(n20970) );
  AOI22_X1 U20725 ( .A1(n21051), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n21027), 
        .B2(n20970), .ZN(n17581) );
  AOI22_X1 U20726 ( .A1(n17579), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n21042), .B2(n17578), .ZN(n17580) );
  OAI211_X1 U20727 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n17582), .A(
        n17581), .B(n17580), .ZN(P1_U3025) );
  NAND2_X1 U20728 ( .A1(n21007), .A2(n17583), .ZN(n21024) );
  OAI22_X1 U20729 ( .A1(n17586), .A2(n17585), .B1(n17584), .B2(n21024), .ZN(
        n17587) );
  AOI21_X1 U20730 ( .B1(n21042), .B2(n17588), .A(n17587), .ZN(n17590) );
  NAND2_X1 U20731 ( .A1(n21051), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n17589) );
  OAI211_X1 U20732 ( .C1(n21054), .C2(n20926), .A(n17590), .B(n17589), .ZN(
        P1_U3026) );
  INV_X1 U20733 ( .A(n17591), .ZN(n17594) );
  NAND4_X1 U20734 ( .A1(n17594), .A2(n17593), .A3(n17592), .A4(n20942), .ZN(
        n17595) );
  OAI21_X1 U20735 ( .B1(n17597), .B2(n17596), .A(n17595), .ZN(P1_U3468) );
  NOR2_X1 U20736 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21739), .ZN(n17598) );
  OAI221_X1 U20737 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n21645), .C2(n17598), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21646) );
  AOI21_X1 U20738 ( .B1(n21646), .B2(n17600), .A(n17599), .ZN(n17602) );
  AOI211_X1 U20739 ( .C1(n21644), .C2(n17603), .A(n17602), .B(n17601), .ZN(
        P1_U3162) );
  OAI21_X1 U20740 ( .B1(n17605), .B2(n21474), .A(n17604), .ZN(P1_U3466) );
  INV_X1 U20741 ( .A(n17606), .ZN(n17608) );
  OAI21_X1 U20742 ( .B1(n17608), .B2(n20850), .A(n17607), .ZN(n17609) );
  AOI21_X1 U20743 ( .B1(n20835), .B2(n17610), .A(n17609), .ZN(n17616) );
  MUX2_X1 U20744 ( .A(n20797), .B(n17612), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n17614) );
  INV_X1 U20745 ( .A(n17611), .ZN(n20849) );
  NAND3_X1 U20746 ( .A1(n17612), .A2(n20844), .A3(n10286), .ZN(n17613) );
  OAI21_X1 U20747 ( .B1(n17614), .B2(n20849), .A(n17613), .ZN(n17615) );
  OAI211_X1 U20748 ( .C1(n17618), .C2(n17617), .A(n17616), .B(n17615), .ZN(
        P2_U3176) );
  INV_X1 U20749 ( .A(n17637), .ZN(n17630) );
  AOI21_X1 U20750 ( .B1(n17631), .B2(n17641), .A(n17619), .ZN(n17627) );
  AOI22_X1 U20751 ( .A1(n19317), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17620), .ZN(n17623) );
  OAI21_X1 U20752 ( .B1(n18865), .B2(n17621), .A(n17749), .ZN(n17622) );
  OAI211_X1 U20753 ( .C1(n17625), .C2(n17624), .A(n17623), .B(n17622), .ZN(
        n17626) );
  AOI211_X1 U20754 ( .C1(n17628), .C2(n18921), .A(n17627), .B(n17626), .ZN(
        n17629) );
  OAI221_X1 U20755 ( .B1(n17632), .B2(n17631), .C1(n17632), .C2(n17630), .A(
        n17629), .ZN(P3_U2801) );
  OAI21_X1 U20756 ( .B1(n17633), .B2(n9755), .A(n18670), .ZN(n18660) );
  AOI22_X1 U20757 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18920), .B1(
        n9755), .B2(n18655), .ZN(n18661) );
  NAND4_X1 U20758 ( .A1(n19810), .A2(n17636), .A3(n17635), .A4(n18659), .ZN(
        n17643) );
  NAND2_X1 U20759 ( .A1(n19810), .A2(n18510), .ZN(n19182) );
  OR2_X1 U20760 ( .A1(n17637), .A2(n19182), .ZN(n17639) );
  NAND2_X1 U20761 ( .A1(n17639), .A2(n17638), .ZN(n17640) );
  NAND2_X1 U20762 ( .A1(n17644), .A2(n19328), .ZN(n17651) );
  INV_X1 U20763 ( .A(n19182), .ZN(n19073) );
  AOI22_X1 U20764 ( .A1(n19811), .A2(n18877), .B1(n19177), .B2(n19073), .ZN(
        n19119) );
  OAI21_X1 U20765 ( .B1(n19775), .B2(n19964), .A(n19794), .ZN(n19304) );
  AOI21_X1 U20766 ( .B1(n19068), .B2(n19304), .A(n17645), .ZN(n19038) );
  OAI21_X1 U20767 ( .B1(n19119), .B2(n19120), .A(n19038), .ZN(n19078) );
  NAND2_X1 U20768 ( .A1(n19327), .A2(n19078), .ZN(n19086) );
  NOR2_X1 U20769 ( .A1(n19015), .A2(n19086), .ZN(n19058) );
  NOR2_X1 U20770 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17646), .ZN(
        n18658) );
  INV_X1 U20771 ( .A(n19297), .ZN(n19331) );
  AND3_X1 U20772 ( .A1(n17633), .A2(n19331), .A3(n17647), .ZN(n17648) );
  INV_X1 U20773 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19916) );
  NOR2_X1 U20774 ( .A1(n19328), .A2(n19916), .ZN(n18652) );
  AOI211_X1 U20775 ( .C1(n19058), .C2(n18658), .A(n17648), .B(n18652), .ZN(
        n17650) );
  INV_X1 U20776 ( .A(n19239), .ZN(n19171) );
  NOR3_X1 U20777 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_0__SCAN_IN), .ZN(n17653) );
  NOR4_X1 U20778 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17652) );
  NAND4_X1 U20779 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17653), .A3(n17652), .A4(
        U215), .ZN(U213) );
  INV_X1 U20780 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20100) );
  NAND2_X2 U20781 ( .A1(U214), .A2(n17654), .ZN(n17692) );
  OAI222_X1 U20782 ( .A1(U212), .A2(n20100), .B1(n17692), .B2(n21103), .C1(
        U214), .C2(n17723), .ZN(U216) );
  OAI222_X1 U20783 ( .A1(U212), .A2(n17720), .B1(n17692), .B2(n16509), .C1(
        U214), .C2(n14116), .ZN(U217) );
  INV_X1 U20784 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n21089) );
  AOI22_X1 U20785 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17687), .ZN(n17655) );
  OAI21_X1 U20786 ( .B1(n21089), .B2(n17692), .A(n17655), .ZN(U218) );
  AOI22_X1 U20787 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17687), .ZN(n17656) );
  OAI21_X1 U20788 ( .B1(n21082), .B2(n17692), .A(n17656), .ZN(U219) );
  INV_X1 U20789 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n21077) );
  AOI22_X1 U20790 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17687), .ZN(n17657) );
  OAI21_X1 U20791 ( .B1(n21077), .B2(n17692), .A(n17657), .ZN(U220) );
  AOI22_X1 U20792 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17687), .ZN(n17658) );
  OAI21_X1 U20793 ( .B1(n21068), .B2(n17692), .A(n17658), .ZN(U221) );
  INV_X1 U20794 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n17717) );
  INV_X1 U20795 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n21059) );
  OAI222_X1 U20796 ( .A1(U212), .A2(n17717), .B1(n17692), .B2(n21059), .C1(
        U214), .C2(n14112), .ZN(U222) );
  AOI22_X1 U20797 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17687), .ZN(n17659) );
  OAI21_X1 U20798 ( .B1(n17660), .B2(n17692), .A(n17659), .ZN(U223) );
  INV_X1 U20799 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n21101) );
  AOI22_X1 U20800 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17687), .ZN(n17661) );
  OAI21_X1 U20801 ( .B1(n21101), .B2(n17692), .A(n17661), .ZN(U224) );
  INV_X1 U20802 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n21096) );
  AOI22_X1 U20803 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17687), .ZN(n17662) );
  OAI21_X1 U20804 ( .B1(n21096), .B2(n17692), .A(n17662), .ZN(U225) );
  INV_X1 U20805 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n21088) );
  OAI222_X1 U20806 ( .A1(U212), .A2(n17713), .B1(n17692), .B2(n21088), .C1(
        U214), .C2(n14101), .ZN(U226) );
  AOI22_X1 U20807 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17687), .ZN(n17663) );
  OAI21_X1 U20808 ( .B1(n21081), .B2(n17692), .A(n17663), .ZN(U227) );
  AOI22_X1 U20809 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17687), .ZN(n17664) );
  OAI21_X1 U20810 ( .B1(n16594), .B2(n17692), .A(n17664), .ZN(U228) );
  AOI22_X1 U20811 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17687), .ZN(n17665) );
  OAI21_X1 U20812 ( .B1(n21067), .B2(n17692), .A(n17665), .ZN(U229) );
  INV_X1 U20813 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n21064) );
  AOI22_X1 U20814 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17687), .ZN(n17666) );
  OAI21_X1 U20815 ( .B1(n21064), .B2(n17692), .A(n17666), .ZN(U230) );
  AOI22_X1 U20816 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17687), .ZN(n17667) );
  OAI21_X1 U20817 ( .B1(n22004), .B2(n17692), .A(n17667), .ZN(U231) );
  AOI22_X1 U20818 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17687), .ZN(n17668) );
  OAI21_X1 U20819 ( .B1(n14162), .B2(n17692), .A(n17668), .ZN(U232) );
  AOI22_X1 U20820 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17687), .ZN(n17669) );
  OAI21_X1 U20821 ( .B1(n14220), .B2(n17692), .A(n17669), .ZN(U233) );
  INV_X1 U20822 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n17705) );
  INV_X1 U20823 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n21907) );
  OAI222_X1 U20824 ( .A1(U212), .A2(n17705), .B1(n17692), .B2(n14089), .C1(
        U214), .C2(n21907), .ZN(U234) );
  AOI22_X1 U20825 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17687), .ZN(n17670) );
  OAI21_X1 U20826 ( .B1(n17671), .B2(n17692), .A(n17670), .ZN(U235) );
  AOI22_X1 U20827 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17687), .ZN(n17672) );
  OAI21_X1 U20828 ( .B1(n17673), .B2(n17692), .A(n17672), .ZN(U236) );
  AOI22_X1 U20829 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17687), .ZN(n17674) );
  OAI21_X1 U20830 ( .B1(n17675), .B2(n17692), .A(n17674), .ZN(U237) );
  AOI22_X1 U20831 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17687), .ZN(n17676) );
  OAI21_X1 U20832 ( .B1(n14074), .B2(n17692), .A(n17676), .ZN(U238) );
  AOI22_X1 U20833 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17687), .ZN(n17677) );
  OAI21_X1 U20834 ( .B1(n14240), .B2(n17692), .A(n17677), .ZN(U239) );
  INV_X1 U20835 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n17679) );
  AOI22_X1 U20836 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n17687), .ZN(n17678) );
  OAI21_X1 U20837 ( .B1(n17679), .B2(n17692), .A(n17678), .ZN(U240) );
  AOI22_X1 U20838 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17687), .ZN(n17680) );
  OAI21_X1 U20839 ( .B1(n13838), .B2(n17692), .A(n17680), .ZN(U241) );
  INV_X1 U20840 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n17682) );
  AOI22_X1 U20841 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17687), .ZN(n17681) );
  OAI21_X1 U20842 ( .B1(n17682), .B2(n17692), .A(n17681), .ZN(U242) );
  INV_X1 U20843 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17683) );
  OAI222_X1 U20844 ( .A1(U212), .A2(n13892), .B1(n17692), .B2(n17683), .C1(
        U214), .C2(n21879), .ZN(U243) );
  INV_X1 U20845 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n17685) );
  AOI22_X1 U20846 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n17687), .ZN(n17684) );
  OAI21_X1 U20847 ( .B1(n17685), .B2(n17692), .A(n17684), .ZN(U244) );
  INV_X1 U20848 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17695) );
  INV_X1 U20849 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17686) );
  OAI222_X1 U20850 ( .A1(U212), .A2(n17695), .B1(n17692), .B2(n17686), .C1(
        U214), .C2(n22038), .ZN(U245) );
  INV_X1 U20851 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n17690) );
  AOI22_X1 U20852 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17688), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17687), .ZN(n17689) );
  OAI21_X1 U20853 ( .B1(n17690), .B2(n17692), .A(n17689), .ZN(U246) );
  INV_X1 U20854 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17693) );
  INV_X1 U20855 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n17691) );
  OAI222_X1 U20856 ( .A1(U212), .A2(n17693), .B1(n17692), .B2(n17691), .C1(
        U214), .C2(n21830), .ZN(U247) );
  AOI22_X1 U20857 ( .A1(n17721), .A2(n17693), .B1(n19345), .B2(U215), .ZN(U251) );
  OAI22_X1 U20858 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17721), .ZN(n17694) );
  INV_X1 U20859 ( .A(n17694), .ZN(U252) );
  AOI22_X1 U20860 ( .A1(n17721), .A2(n17695), .B1(n19354), .B2(U215), .ZN(U253) );
  INV_X1 U20861 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17696) );
  INV_X1 U20862 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19358) );
  AOI22_X1 U20863 ( .A1(n17721), .A2(n17696), .B1(n19358), .B2(U215), .ZN(U254) );
  INV_X1 U20864 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19362) );
  AOI22_X1 U20865 ( .A1(n17721), .A2(n13892), .B1(n19362), .B2(U215), .ZN(U255) );
  INV_X1 U20866 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17697) );
  AOI22_X1 U20867 ( .A1(n17721), .A2(n17697), .B1(n13829), .B2(U215), .ZN(U256) );
  INV_X1 U20868 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17698) );
  AOI22_X1 U20869 ( .A1(n17722), .A2(n17698), .B1(n13839), .B2(U215), .ZN(U257) );
  INV_X1 U20870 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17699) );
  AOI22_X1 U20871 ( .A1(n17722), .A2(n17699), .B1(n13920), .B2(U215), .ZN(U258) );
  OAI22_X1 U20872 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17721), .ZN(n17700) );
  INV_X1 U20873 ( .A(n17700), .ZN(U259) );
  INV_X1 U20874 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17701) );
  AOI22_X1 U20875 ( .A1(n17722), .A2(n17701), .B1(n13821), .B2(U215), .ZN(U260) );
  INV_X1 U20876 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17702) );
  AOI22_X1 U20877 ( .A1(n17721), .A2(n17702), .B1(n18639), .B2(U215), .ZN(U261) );
  INV_X1 U20878 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17703) );
  AOI22_X1 U20879 ( .A1(n17722), .A2(n17703), .B1(n13817), .B2(U215), .ZN(U262) );
  INV_X1 U20880 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U20881 ( .A1(n17721), .A2(n17704), .B1(n18642), .B2(U215), .ZN(U263) );
  AOI22_X1 U20882 ( .A1(n17722), .A2(n17705), .B1(n13833), .B2(U215), .ZN(U264) );
  OAI22_X1 U20883 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17721), .ZN(n17706) );
  INV_X1 U20884 ( .A(n17706), .ZN(U265) );
  INV_X1 U20885 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n17707) );
  AOI22_X1 U20886 ( .A1(n17722), .A2(n17707), .B1(n13855), .B2(U215), .ZN(U266) );
  OAI22_X1 U20887 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17721), .ZN(n17708) );
  INV_X1 U20888 ( .A(n17708), .ZN(U267) );
  OAI22_X1 U20889 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17721), .ZN(n17709) );
  INV_X1 U20890 ( .A(n17709), .ZN(U268) );
  OAI22_X1 U20891 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17722), .ZN(n17710) );
  INV_X1 U20892 ( .A(n17710), .ZN(U269) );
  OAI22_X1 U20893 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17722), .ZN(n17711) );
  INV_X1 U20894 ( .A(n17711), .ZN(U270) );
  OAI22_X1 U20895 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17722), .ZN(n17712) );
  INV_X1 U20896 ( .A(n17712), .ZN(U271) );
  AOI22_X1 U20897 ( .A1(n17721), .A2(n17713), .B1(n16581), .B2(U215), .ZN(U272) );
  OAI22_X1 U20898 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17721), .ZN(n17714) );
  INV_X1 U20899 ( .A(n17714), .ZN(U273) );
  OAI22_X1 U20900 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17721), .ZN(n17715) );
  INV_X1 U20901 ( .A(n17715), .ZN(U274) );
  OAI22_X1 U20902 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17721), .ZN(n17716) );
  INV_X1 U20903 ( .A(n17716), .ZN(U275) );
  INV_X1 U20904 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n22030) );
  AOI22_X1 U20905 ( .A1(n17721), .A2(n17717), .B1(n22030), .B2(U215), .ZN(U276) );
  AOI22_X1 U20906 ( .A1(n17721), .A2(n13899), .B1(n21883), .B2(U215), .ZN(U277) );
  OAI22_X1 U20907 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17721), .ZN(n17718) );
  INV_X1 U20908 ( .A(n17718), .ZN(U278) );
  INV_X1 U20909 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n20160) );
  AOI22_X1 U20910 ( .A1(n17721), .A2(n13897), .B1(n20160), .B2(U215), .ZN(U279) );
  OAI22_X1 U20911 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17721), .ZN(n17719) );
  INV_X1 U20912 ( .A(n17719), .ZN(U280) );
  AOI22_X1 U20913 ( .A1(n17721), .A2(n17720), .B1(n16511), .B2(U215), .ZN(U281) );
  INV_X1 U20914 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n20178) );
  AOI22_X1 U20915 ( .A1(n17722), .A2(n20100), .B1(n20178), .B2(U215), .ZN(U282) );
  INV_X1 U20916 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n22005) );
  AOI222_X1 U20917 ( .A1(n20100), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17723), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n22005), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17724) );
  INV_X2 U20918 ( .A(n17724), .ZN(n17726) );
  INV_X2 U20919 ( .A(n17726), .ZN(n17725) );
  INV_X1 U20920 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19881) );
  INV_X1 U20921 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20747) );
  AOI22_X1 U20922 ( .A1(n17725), .A2(n19881), .B1(n20747), .B2(n17726), .ZN(
        U347) );
  INV_X1 U20923 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19879) );
  INV_X1 U20924 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20746) );
  AOI22_X1 U20925 ( .A1(n17725), .A2(n19879), .B1(n20746), .B2(n17726), .ZN(
        U348) );
  INV_X1 U20926 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n21953) );
  INV_X1 U20927 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20744) );
  AOI22_X1 U20928 ( .A1(n17725), .A2(n21953), .B1(n20744), .B2(n17726), .ZN(
        U349) );
  INV_X1 U20929 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19876) );
  INV_X1 U20930 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20742) );
  AOI22_X1 U20931 ( .A1(n17725), .A2(n19876), .B1(n20742), .B2(n17726), .ZN(
        U350) );
  INV_X1 U20932 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19874) );
  INV_X1 U20933 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20740) );
  AOI22_X1 U20934 ( .A1(n17725), .A2(n19874), .B1(n20740), .B2(n17726), .ZN(
        U351) );
  INV_X1 U20935 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19871) );
  INV_X1 U20936 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20739) );
  AOI22_X1 U20937 ( .A1(n17725), .A2(n19871), .B1(n20739), .B2(n17726), .ZN(
        U352) );
  INV_X1 U20938 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19870) );
  INV_X1 U20939 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n21832) );
  AOI22_X1 U20940 ( .A1(n17725), .A2(n19870), .B1(n21832), .B2(n17726), .ZN(
        U353) );
  INV_X1 U20941 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19868) );
  INV_X1 U20942 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20737) );
  AOI22_X1 U20943 ( .A1(n17725), .A2(n19868), .B1(n20737), .B2(n17726), .ZN(
        U354) );
  INV_X1 U20944 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19920) );
  INV_X1 U20945 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20780) );
  AOI22_X1 U20946 ( .A1(n17725), .A2(n19920), .B1(n20780), .B2(n17726), .ZN(
        U355) );
  INV_X1 U20947 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19918) );
  INV_X1 U20948 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n21809) );
  AOI22_X1 U20949 ( .A1(n17725), .A2(n19918), .B1(n21809), .B2(n17726), .ZN(
        U356) );
  INV_X1 U20950 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19915) );
  AOI22_X1 U20951 ( .A1(n17725), .A2(n19915), .B1(n20775), .B2(n17726), .ZN(
        U357) );
  INV_X1 U20952 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19914) );
  INV_X1 U20953 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20773) );
  AOI22_X1 U20954 ( .A1(n17725), .A2(n19914), .B1(n20773), .B2(n17726), .ZN(
        U358) );
  INV_X1 U20955 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19912) );
  INV_X1 U20956 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20772) );
  AOI22_X1 U20957 ( .A1(n17725), .A2(n19912), .B1(n20772), .B2(n17726), .ZN(
        U359) );
  INV_X1 U20958 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19910) );
  INV_X1 U20959 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20771) );
  AOI22_X1 U20960 ( .A1(n17725), .A2(n19910), .B1(n20771), .B2(n17726), .ZN(
        U360) );
  INV_X1 U20961 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19907) );
  INV_X1 U20962 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20770) );
  AOI22_X1 U20963 ( .A1(n17725), .A2(n19907), .B1(n20770), .B2(n17726), .ZN(
        U361) );
  INV_X1 U20964 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19905) );
  INV_X1 U20965 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20768) );
  AOI22_X1 U20966 ( .A1(n17725), .A2(n19905), .B1(n20768), .B2(n17726), .ZN(
        U362) );
  INV_X1 U20967 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19903) );
  INV_X1 U20968 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20766) );
  AOI22_X1 U20969 ( .A1(n17725), .A2(n19903), .B1(n20766), .B2(n17726), .ZN(
        U363) );
  INV_X1 U20970 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19901) );
  INV_X1 U20971 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20765) );
  AOI22_X1 U20972 ( .A1(n17725), .A2(n19901), .B1(n20765), .B2(n17726), .ZN(
        U364) );
  INV_X1 U20973 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19866) );
  INV_X1 U20974 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20735) );
  AOI22_X1 U20975 ( .A1(n17725), .A2(n19866), .B1(n20735), .B2(n17726), .ZN(
        U365) );
  INV_X1 U20976 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19899) );
  INV_X1 U20977 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20763) );
  AOI22_X1 U20978 ( .A1(n17725), .A2(n19899), .B1(n20763), .B2(n17726), .ZN(
        U366) );
  INV_X1 U20979 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19897) );
  INV_X1 U20980 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20761) );
  AOI22_X1 U20981 ( .A1(n17725), .A2(n19897), .B1(n20761), .B2(n17726), .ZN(
        U367) );
  INV_X1 U20982 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19895) );
  INV_X1 U20983 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20759) );
  AOI22_X1 U20984 ( .A1(n17725), .A2(n19895), .B1(n20759), .B2(n17726), .ZN(
        U368) );
  INV_X1 U20985 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19893) );
  INV_X1 U20986 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20758) );
  AOI22_X1 U20987 ( .A1(n17725), .A2(n19893), .B1(n20758), .B2(n17726), .ZN(
        U369) );
  INV_X1 U20988 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19891) );
  INV_X1 U20989 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20756) );
  AOI22_X1 U20990 ( .A1(n17725), .A2(n19891), .B1(n20756), .B2(n17726), .ZN(
        U370) );
  INV_X1 U20991 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19890) );
  INV_X1 U20992 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20754) );
  AOI22_X1 U20993 ( .A1(n17725), .A2(n19890), .B1(n20754), .B2(n17726), .ZN(
        U371) );
  INV_X1 U20994 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19888) );
  INV_X1 U20995 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20753) );
  AOI22_X1 U20996 ( .A1(n17724), .A2(n19888), .B1(n20753), .B2(n17726), .ZN(
        U372) );
  INV_X1 U20997 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19886) );
  INV_X1 U20998 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20752) );
  AOI22_X1 U20999 ( .A1(n17725), .A2(n19886), .B1(n20752), .B2(n17726), .ZN(
        U373) );
  INV_X1 U21000 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19884) );
  INV_X1 U21001 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20751) );
  AOI22_X1 U21002 ( .A1(n17724), .A2(n19884), .B1(n20751), .B2(n17726), .ZN(
        U374) );
  INV_X1 U21003 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19883) );
  INV_X1 U21004 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20749) );
  AOI22_X1 U21005 ( .A1(n17725), .A2(n19883), .B1(n20749), .B2(n17726), .ZN(
        U375) );
  INV_X1 U21006 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19864) );
  INV_X1 U21007 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20733) );
  AOI22_X1 U21008 ( .A1(n17725), .A2(n19864), .B1(n20733), .B2(n17726), .ZN(
        U376) );
  INV_X1 U21009 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17727) );
  INV_X1 U21010 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19863) );
  NAND2_X1 U21011 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19863), .ZN(n19852) );
  AOI22_X1 U21012 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19852), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19861), .ZN(n19934) );
  OAI21_X1 U21013 ( .B1(n19861), .B2(n17727), .A(n19931), .ZN(P3_U2633) );
  INV_X1 U21014 ( .A(n17733), .ZN(n17728) );
  OAI21_X1 U21015 ( .B1(n17728), .B2(n18598), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17729) );
  OAI21_X1 U21016 ( .B1(n17730), .B2(n19841), .A(n17729), .ZN(P3_U2634) );
  AOI21_X1 U21017 ( .B1(n19861), .B2(n19863), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17731) );
  AOI22_X1 U21018 ( .A1(n19928), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17731), 
        .B2(n19999), .ZN(P3_U2635) );
  NOR2_X1 U21019 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19849) );
  OAI21_X1 U21020 ( .B1(n19849), .B2(BS16), .A(n19934), .ZN(n19932) );
  OAI21_X1 U21021 ( .B1(n19934), .B2(n19988), .A(n19932), .ZN(P3_U2636) );
  AND3_X1 U21022 ( .A1(n17733), .A2(n19814), .A3(n17732), .ZN(n19820) );
  NOR2_X1 U21023 ( .A1(n19820), .A2(n19836), .ZN(n19979) );
  OAI21_X1 U21024 ( .B1(n19979), .B2(n19338), .A(n17734), .ZN(P3_U2637) );
  NOR4_X1 U21025 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17738) );
  NOR4_X1 U21026 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n17737) );
  NOR4_X1 U21027 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17736) );
  NOR4_X1 U21028 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17735) );
  NAND4_X1 U21029 ( .A1(n17738), .A2(n17737), .A3(n17736), .A4(n17735), .ZN(
        n17744) );
  NOR4_X1 U21030 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n17742) );
  AOI211_X1 U21031 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_4__SCAN_IN), .B(
        P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n17741) );
  NOR4_X1 U21032 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n17740) );
  NOR4_X1 U21033 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17739) );
  NAND4_X1 U21034 ( .A1(n17742), .A2(n17741), .A3(n17740), .A4(n17739), .ZN(
        n17743) );
  NOR2_X1 U21035 ( .A1(n17744), .A2(n17743), .ZN(n19973) );
  INV_X1 U21036 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19926) );
  NOR3_X1 U21037 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17746) );
  OAI21_X1 U21038 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17746), .A(n19973), .ZN(
        n17745) );
  OAI21_X1 U21039 ( .B1(n19973), .B2(n19926), .A(n17745), .ZN(P3_U2638) );
  INV_X1 U21040 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19969) );
  INV_X1 U21041 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19933) );
  AOI21_X1 U21042 ( .B1(n19969), .B2(n19933), .A(n17746), .ZN(n17747) );
  INV_X1 U21043 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19924) );
  INV_X1 U21044 ( .A(n19973), .ZN(n19976) );
  AOI22_X1 U21045 ( .A1(n19973), .A2(n17747), .B1(n19924), .B2(n19976), .ZN(
        P3_U2639) );
  INV_X1 U21046 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19917) );
  NAND2_X1 U21047 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n17761), .ZN(n17750) );
  OAI22_X1 U21048 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17750), .B1(n21895), 
        .B2(n18076), .ZN(n17751) );
  INV_X1 U21049 ( .A(n17752), .ZN(n17753) );
  OAI21_X1 U21050 ( .B1(n17758), .B2(n18098), .A(n17753), .ZN(n17754) );
  AOI22_X1 U21051 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n17771), .B1(n18074), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17763) );
  AOI211_X1 U21052 ( .C1(n18654), .C2(n17757), .A(n17756), .B(n10977), .ZN(
        n17760) );
  AOI211_X1 U21053 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17772), .A(n17758), .B(
        n18080), .ZN(n17759) );
  AOI211_X1 U21054 ( .C1(n17761), .C2(n19916), .A(n17760), .B(n17759), .ZN(
        n17762) );
  OAI211_X1 U21055 ( .C1(n17764), .C2(n18076), .A(n17763), .B(n17762), .ZN(
        P3_U2643) );
  AOI22_X1 U21056 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18005), .B1(
        n18074), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n17776) );
  NAND2_X1 U21057 ( .A1(n17765), .A2(n19913), .ZN(n17770) );
  AOI211_X1 U21058 ( .C1(n17768), .C2(n17767), .A(n17766), .B(n10977), .ZN(
        n17769) );
  AOI21_X1 U21059 ( .B1(n17771), .B2(n17770), .A(n17769), .ZN(n17775) );
  OAI211_X1 U21060 ( .C1(n17781), .C2(n17773), .A(n18090), .B(n17772), .ZN(
        n17774) );
  NAND3_X1 U21061 ( .A1(n17776), .A2(n17775), .A3(n17774), .ZN(P3_U2644) );
  AOI22_X1 U21062 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18005), .B1(
        n18074), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17786) );
  AOI221_X1 U21063 ( .B1(n18081), .B2(n19911), .C1(n17778), .C2(n19911), .A(
        n17777), .ZN(n17784) );
  AOI211_X1 U21064 ( .C1(n18684), .C2(n17780), .A(n17779), .B(n10977), .ZN(
        n17783) );
  AOI211_X1 U21065 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17791), .A(n17781), .B(
        n18080), .ZN(n17782) );
  AOI211_X1 U21066 ( .C1(n17784), .C2(n18089), .A(n17783), .B(n17782), .ZN(
        n17785) );
  NAND2_X1 U21067 ( .A1(n17786), .A2(n17785), .ZN(P3_U2645) );
  AOI22_X1 U21068 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18005), .B1(
        n18074), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n17797) );
  NOR2_X1 U21069 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18081), .ZN(n17798) );
  NAND2_X1 U21070 ( .A1(n18055), .A2(n17787), .ZN(n17810) );
  NAND2_X1 U21071 ( .A1(n18091), .A2(n17810), .ZN(n17807) );
  AOI211_X1 U21072 ( .C1(n18698), .C2(n17789), .A(n17788), .B(n10977), .ZN(
        n17790) );
  AOI221_X1 U21073 ( .B1(n17798), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n17807), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n17790), .ZN(n17796) );
  OAI211_X1 U21074 ( .C1(n17800), .C2(n17792), .A(n18090), .B(n17791), .ZN(
        n17795) );
  INV_X1 U21075 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19909) );
  NAND3_X1 U21076 ( .A1(n18055), .A2(n17793), .A3(n19909), .ZN(n17794) );
  NAND4_X1 U21077 ( .A1(n17797), .A2(n17796), .A3(n17795), .A4(n17794), .ZN(
        P3_U2646) );
  AOI22_X1 U21078 ( .A1(n18074), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17799), 
        .B2(n17798), .ZN(n17806) );
  AOI211_X1 U21079 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17814), .A(n17800), .B(
        n18080), .ZN(n17804) );
  AOI211_X1 U21080 ( .C1(n18713), .C2(n17802), .A(n17801), .B(n10977), .ZN(
        n17803) );
  AOI211_X1 U21081 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n17807), .A(n17804), 
        .B(n17803), .ZN(n17805) );
  OAI211_X1 U21082 ( .C1(n18710), .C2(n18076), .A(n17806), .B(n17805), .ZN(
        P3_U2647) );
  INV_X1 U21083 ( .A(n17807), .ZN(n17817) );
  AOI211_X1 U21084 ( .C1(n18722), .C2(n17809), .A(n17808), .B(n10977), .ZN(
        n17813) );
  OAI22_X1 U21085 ( .A1(n18694), .A2(n18076), .B1(n17811), .B2(n17810), .ZN(
        n17812) );
  AOI211_X1 U21086 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n18074), .A(n17813), .B(
        n17812), .ZN(n17816) );
  OAI211_X1 U21087 ( .C1(n17820), .C2(n18097), .A(n18090), .B(n17814), .ZN(
        n17815) );
  OAI211_X1 U21088 ( .C1(n17817), .C2(n19904), .A(n17816), .B(n17815), .ZN(
        P3_U2648) );
  NOR3_X1 U21089 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n18081), .A3(n17818), 
        .ZN(n17819) );
  AOI21_X1 U21090 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18074), .A(n17819), .ZN(
        n17829) );
  OAI221_X1 U21091 ( .B1(n18081), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n18081), 
        .C2(n17836), .A(n18091), .ZN(n17827) );
  AOI211_X1 U21092 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17832), .A(n17820), .B(
        n18080), .ZN(n17826) );
  INV_X1 U21093 ( .A(n17821), .ZN(n17824) );
  INV_X1 U21094 ( .A(n17822), .ZN(n17823) );
  AOI211_X1 U21095 ( .C1(n18738), .C2(n17824), .A(n17823), .B(n10977), .ZN(
        n17825) );
  AOI211_X1 U21096 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17827), .A(n17826), 
        .B(n17825), .ZN(n17828) );
  OAI211_X1 U21097 ( .C1(n18735), .C2(n18076), .A(n17829), .B(n17828), .ZN(
        P3_U2649) );
  OAI21_X1 U21098 ( .B1(n17836), .B2(n18081), .A(n18091), .ZN(n17844) );
  AOI211_X1 U21099 ( .C1(n18750), .C2(n17831), .A(n17830), .B(n10977), .ZN(
        n17835) );
  OAI211_X1 U21100 ( .C1(n17841), .C2(n18182), .A(n18090), .B(n17832), .ZN(
        n17833) );
  OAI21_X1 U21101 ( .B1(n18182), .B2(n18059), .A(n17833), .ZN(n17834) );
  AOI211_X1 U21102 ( .C1(n17844), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17835), 
        .B(n17834), .ZN(n17838) );
  INV_X1 U21103 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19900) );
  NAND3_X1 U21104 ( .A1(n18055), .A2(n17836), .A3(n19900), .ZN(n17837) );
  OAI211_X1 U21105 ( .C1(n18076), .C2(n18747), .A(n17838), .B(n17837), .ZN(
        P3_U2650) );
  AOI211_X1 U21106 ( .C1(n17840), .C2(n17839), .A(n9934), .B(n10977), .ZN(
        n17843) );
  AOI211_X1 U21107 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17857), .A(n17841), .B(
        n18080), .ZN(n17842) );
  AOI211_X1 U21108 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n18074), .A(n17843), .B(
        n17842), .ZN(n17846) );
  NAND4_X1 U21109 ( .A1(n18055), .A2(P3_REIP_REG_16__SCAN_IN), .A3(
        P3_REIP_REG_17__SCAN_IN), .A4(n17871), .ZN(n17848) );
  NOR2_X1 U21110 ( .A1(n19894), .A2(n17848), .ZN(n17856) );
  OAI221_X1 U21111 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(P3_REIP_REG_19__SCAN_IN), .C1(P3_REIP_REG_20__SCAN_IN), .C2(n17856), .A(n17844), .ZN(n17845) );
  OAI211_X1 U21112 ( .C1(n18076), .C2(n18759), .A(n17846), .B(n17845), .ZN(
        P3_U2651) );
  AOI22_X1 U21113 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18005), .B1(
        n18074), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n17860) );
  AOI21_X1 U21114 ( .B1(n18055), .B2(n17847), .A(n18073), .ZN(n17875) );
  OR2_X1 U21115 ( .A1(n17848), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17867) );
  NAND2_X1 U21116 ( .A1(n17875), .A2(n17867), .ZN(n17855) );
  INV_X1 U21117 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17862) );
  NOR2_X1 U21118 ( .A1(n17862), .A2(n17863), .ZN(n17850) );
  INV_X1 U21119 ( .A(n17849), .ZN(n18731) );
  OAI21_X1 U21120 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17850), .A(
        n18731), .ZN(n18775) );
  AOI22_X1 U21121 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17863), .B1(
        n18771), .B2(n17862), .ZN(n18785) );
  OAI211_X1 U21122 ( .C1(n18771), .C2(n18043), .A(n17851), .B(n18785), .ZN(
        n17864) );
  NAND2_X1 U21123 ( .A1(n18017), .A2(n17864), .ZN(n17853) );
  OAI21_X1 U21124 ( .B1(n18775), .B2(n17853), .A(n18067), .ZN(n17852) );
  AOI21_X1 U21125 ( .B1(n18775), .B2(n17853), .A(n17852), .ZN(n17854) );
  AOI221_X1 U21126 ( .B1(n17856), .B2(n19896), .C1(n17855), .C2(
        P3_REIP_REG_19__SCAN_IN), .A(n17854), .ZN(n17859) );
  OAI211_X1 U21127 ( .C1(n17861), .C2(n18195), .A(n18090), .B(n17857), .ZN(
        n17858) );
  NAND4_X1 U21128 ( .A1(n17860), .A2(n17859), .A3(n19328), .A4(n17858), .ZN(
        P3_U2652) );
  AOI211_X1 U21129 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17878), .A(n17861), .B(
        n18080), .ZN(n17870) );
  OAI22_X1 U21130 ( .A1(n17862), .A2(n18076), .B1(n18059), .B2(n18224), .ZN(
        n17869) );
  INV_X1 U21131 ( .A(n17851), .ZN(n17885) );
  AOI21_X1 U21132 ( .B1(n18017), .B2(n17863), .A(n17885), .ZN(n17865) );
  OAI211_X1 U21133 ( .C1(n17865), .C2(n18785), .A(n18067), .B(n17864), .ZN(
        n17866) );
  OAI211_X1 U21134 ( .C1(n17875), .C2(n19894), .A(n17867), .B(n17866), .ZN(
        n17868) );
  OR4_X1 U21135 ( .A1(n19317), .A2(n17870), .A3(n17869), .A4(n17868), .ZN(
        P3_U2653) );
  AND2_X1 U21136 ( .A1(n18055), .A2(n17871), .ZN(n17881) );
  AOI21_X1 U21137 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n17881), .A(
        P3_REIP_REG_17__SCAN_IN), .ZN(n17876) );
  INV_X1 U21138 ( .A(n17895), .ZN(n17883) );
  NAND2_X1 U21139 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17883), .ZN(
        n17882) );
  AOI21_X1 U21140 ( .B1(n18796), .B2(n17882), .A(n18771), .ZN(n18800) );
  INV_X1 U21141 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18078) );
  NAND2_X1 U21142 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18078), .ZN(
        n18065) );
  OAI21_X1 U21143 ( .B1(n17872), .B2(n18065), .A(n18017), .ZN(n17873) );
  XOR2_X1 U21144 ( .A(n18800), .B(n17873), .Z(n17874) );
  OAI22_X1 U21145 ( .A1(n17876), .A2(n17875), .B1(n10977), .B2(n17874), .ZN(
        n17877) );
  AOI211_X1 U21146 ( .C1(n18074), .C2(P3_EBX_REG_17__SCAN_IN), .A(n19317), .B(
        n17877), .ZN(n17880) );
  OAI211_X1 U21147 ( .C1(n17886), .C2(n18235), .A(n18090), .B(n17878), .ZN(
        n17879) );
  OAI211_X1 U21148 ( .C1(n18076), .C2(n18796), .A(n17880), .B(n17879), .ZN(
        P3_U2654) );
  INV_X1 U21149 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n22035) );
  AOI22_X1 U21150 ( .A1(n18074), .A2(P3_EBX_REG_16__SCAN_IN), .B1(n17881), 
        .B2(n22035), .ZN(n17893) );
  OAI21_X1 U21151 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17883), .A(
        n17882), .ZN(n18815) );
  INV_X1 U21152 ( .A(n18815), .ZN(n17884) );
  AOI221_X1 U21153 ( .B1(n17851), .B2(n18815), .C1(n17885), .C2(n17884), .A(
        n10977), .ZN(n17888) );
  AOI211_X1 U21154 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17898), .A(n17886), .B(
        n18080), .ZN(n17887) );
  AOI211_X1 U21155 ( .C1(n18005), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17888), .B(n17887), .ZN(n17892) );
  NOR2_X1 U21156 ( .A1(n18073), .A2(n17890), .ZN(n17908) );
  NOR2_X1 U21157 ( .A1(n17889), .A2(n17908), .ZN(n17913) );
  NOR3_X1 U21158 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n18081), .A3(n17890), 
        .ZN(n17894) );
  OAI21_X1 U21159 ( .B1(n17913), .B2(n17894), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n17891) );
  NAND4_X1 U21160 ( .A1(n17893), .A2(n17892), .A3(n19328), .A4(n17891), .ZN(
        P3_U2655) );
  INV_X1 U21161 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18823) );
  AOI21_X1 U21162 ( .B1(n17913), .B2(P3_REIP_REG_15__SCAN_IN), .A(n17894), 
        .ZN(n17905) );
  NOR2_X1 U21163 ( .A1(n17851), .A2(n10977), .ZN(n17903) );
  OAI21_X1 U21164 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18810), .A(
        n17895), .ZN(n18820) );
  INV_X1 U21165 ( .A(n18810), .ZN(n17897) );
  NAND2_X1 U21166 ( .A1(n18017), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17896) );
  NAND2_X1 U21167 ( .A1(n18067), .A2(n17896), .ZN(n18075) );
  AOI211_X1 U21168 ( .C1(n18017), .C2(n17897), .A(n18820), .B(n18075), .ZN(
        n17902) );
  OAI211_X1 U21169 ( .C1(n17906), .C2(n17900), .A(n18090), .B(n17898), .ZN(
        n17899) );
  OAI211_X1 U21170 ( .C1(n18059), .C2(n17900), .A(n19328), .B(n17899), .ZN(
        n17901) );
  AOI211_X1 U21171 ( .C1(n17903), .C2(n18820), .A(n17902), .B(n17901), .ZN(
        n17904) );
  OAI211_X1 U21172 ( .C1(n18823), .C2(n18076), .A(n17905), .B(n17904), .ZN(
        P3_U2656) );
  AOI211_X1 U21173 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17924), .A(n17906), .B(
        n18080), .ZN(n17907) );
  AOI21_X1 U21174 ( .B1(n18005), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17907), .ZN(n17917) );
  NOR2_X1 U21175 ( .A1(n17908), .A2(n18081), .ZN(n17909) );
  AOI22_X1 U21176 ( .A1(n18074), .A2(P3_EBX_REG_14__SCAN_IN), .B1(n17910), 
        .B2(n17909), .ZN(n17916) );
  INV_X1 U21177 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17911) );
  INV_X1 U21178 ( .A(n17944), .ZN(n18848) );
  NAND2_X1 U21179 ( .A1(n18847), .A2(n18848), .ZN(n17921) );
  AOI21_X1 U21180 ( .B1(n17911), .B2(n17921), .A(n18810), .ZN(n18835) );
  OAI21_X1 U21181 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17921), .A(
        n18017), .ZN(n17912) );
  XNOR2_X1 U21182 ( .A(n18835), .B(n17912), .ZN(n17914) );
  AOI22_X1 U21183 ( .A1(n18067), .A2(n17914), .B1(P3_REIP_REG_14__SCAN_IN), 
        .B2(n17913), .ZN(n17915) );
  NAND4_X1 U21184 ( .A1(n17917), .A2(n17916), .A3(n17915), .A4(n19328), .ZN(
        P3_U2657) );
  NOR3_X1 U21185 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n18081), .A3(n17918), 
        .ZN(n17919) );
  AOI211_X1 U21186 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18005), .A(
        n19317), .B(n17919), .ZN(n17929) );
  NOR2_X1 U21187 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17921), .ZN(
        n17920) );
  NOR2_X1 U21188 ( .A1(n17920), .A2(n18077), .ZN(n17922) );
  NOR2_X1 U21189 ( .A1(n18861), .A2(n17944), .ZN(n17934) );
  OAI21_X1 U21190 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17934), .A(
        n17921), .ZN(n18850) );
  AOI22_X1 U21191 ( .A1(n18074), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n17922), 
        .B2(n18850), .ZN(n17928) );
  OAI21_X1 U21192 ( .B1(n17933), .B2(n18081), .A(n18091), .ZN(n17953) );
  NOR2_X1 U21193 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18081), .ZN(n17932) );
  AOI211_X1 U21194 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18017), .A(
        n18850), .B(n18075), .ZN(n17923) );
  AOI221_X1 U21195 ( .B1(n17953), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n17932), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n17923), .ZN(n17927) );
  OAI211_X1 U21196 ( .C1(n17930), .C2(n17925), .A(n18090), .B(n17924), .ZN(
        n17926) );
  NAND4_X1 U21197 ( .A1(n17929), .A2(n17928), .A3(n17927), .A4(n17926), .ZN(
        P3_U2658) );
  AOI211_X1 U21198 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17947), .A(n17930), .B(
        n18080), .ZN(n17931) );
  AOI21_X1 U21199 ( .B1(n18005), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17931), .ZN(n17940) );
  AOI22_X1 U21200 ( .A1(n18074), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n17933), 
        .B2(n17932), .ZN(n17939) );
  AOI21_X1 U21201 ( .B1(n18861), .B2(n17944), .A(n17934), .ZN(n18864) );
  OAI21_X1 U21202 ( .B1(n17935), .B2(n18065), .A(n18017), .ZN(n17936) );
  XNOR2_X1 U21203 ( .A(n18864), .B(n17936), .ZN(n17937) );
  AOI22_X1 U21204 ( .A1(n18067), .A2(n17937), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n17953), .ZN(n17938) );
  NAND4_X1 U21205 ( .A1(n17940), .A2(n17939), .A3(n17938), .A4(n19328), .ZN(
        P3_U2659) );
  OR2_X1 U21206 ( .A1(n18081), .A2(n17959), .ZN(n17957) );
  OAI21_X1 U21207 ( .B1(n17941), .B2(n17957), .A(n19882), .ZN(n17952) );
  NOR2_X1 U21208 ( .A1(n17942), .A2(n18065), .ZN(n17994) );
  NAND2_X1 U21209 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17994), .ZN(
        n17983) );
  OAI21_X1 U21210 ( .B1(n17943), .B2(n17983), .A(n18017), .ZN(n17946) );
  INV_X1 U21211 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21923) );
  NAND3_X1 U21212 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(n17993), .ZN(n17967) );
  NOR2_X1 U21213 ( .A1(n21923), .A2(n17967), .ZN(n17956) );
  OAI21_X1 U21214 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17956), .A(
        n17944), .ZN(n18872) );
  AOI21_X1 U21215 ( .B1(n17946), .B2(n18872), .A(n10977), .ZN(n17945) );
  OAI21_X1 U21216 ( .B1(n17946), .B2(n18872), .A(n17945), .ZN(n17949) );
  OAI211_X1 U21217 ( .C1(n17961), .C2(n17955), .A(n18090), .B(n17947), .ZN(
        n17948) );
  OAI211_X1 U21218 ( .C1(n18076), .C2(n17950), .A(n17949), .B(n17948), .ZN(
        n17951) );
  AOI21_X1 U21219 ( .B1(n17953), .B2(n17952), .A(n17951), .ZN(n17954) );
  OAI211_X1 U21220 ( .C1(n18059), .C2(n17955), .A(n17954), .B(n19328), .ZN(
        P3_U2660) );
  AOI21_X1 U21221 ( .B1(n21923), .B2(n17967), .A(n17956), .ZN(n18885) );
  OAI21_X1 U21222 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17967), .A(
        n18017), .ZN(n17970) );
  XOR2_X1 U21223 ( .A(n18885), .B(n17970), .Z(n17966) );
  INV_X1 U21224 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19878) );
  NOR3_X1 U21225 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n19878), .A3(n17957), 
        .ZN(n17958) );
  AOI211_X1 U21226 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18005), .A(
        n19317), .B(n17958), .ZN(n17965) );
  AOI21_X1 U21227 ( .B1(n18055), .B2(n17959), .A(n18073), .ZN(n17991) );
  NOR3_X1 U21228 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17959), .A3(n18081), .ZN(
        n17971) );
  INV_X1 U21229 ( .A(n17971), .ZN(n17960) );
  INV_X1 U21230 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19880) );
  AOI21_X1 U21231 ( .B1(n17991), .B2(n17960), .A(n19880), .ZN(n17963) );
  AOI211_X1 U21232 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17972), .A(n17961), .B(
        n18080), .ZN(n17962) );
  AOI211_X1 U21233 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n18074), .A(n17963), .B(
        n17962), .ZN(n17964) );
  OAI211_X1 U21234 ( .C1(n10977), .C2(n17966), .A(n17965), .B(n17964), .ZN(
        P3_U2661) );
  INV_X1 U21235 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18913) );
  INV_X1 U21236 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17975) );
  OAI21_X1 U21237 ( .B1(n18913), .B2(n17982), .A(n17975), .ZN(n17968) );
  NAND2_X1 U21238 ( .A1(n17967), .A2(n17968), .ZN(n18902) );
  AND2_X1 U21239 ( .A1(n17967), .A2(n18017), .ZN(n17969) );
  AOI22_X1 U21240 ( .A1(n17970), .A2(n18902), .B1(n17969), .B2(n17968), .ZN(
        n17978) );
  NOR3_X1 U21241 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18913), .A3(
        n17983), .ZN(n17977) );
  AOI211_X1 U21242 ( .C1(n18074), .C2(P3_EBX_REG_9__SCAN_IN), .A(n19317), .B(
        n17971), .ZN(n17974) );
  OAI211_X1 U21243 ( .C1(n17986), .C2(n18309), .A(n18090), .B(n17972), .ZN(
        n17973) );
  OAI211_X1 U21244 ( .C1(n18076), .C2(n17975), .A(n17974), .B(n17973), .ZN(
        n17976) );
  AOI221_X1 U21245 ( .B1(n17978), .B2(n18067), .C1(n17977), .C2(n18067), .A(
        n17976), .ZN(n17979) );
  OAI21_X1 U21246 ( .B1(n19878), .B2(n17991), .A(n17979), .ZN(P3_U2662) );
  INV_X1 U21247 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19877) );
  NAND2_X1 U21248 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n17980) );
  NAND2_X1 U21249 ( .A1(n18055), .A2(n17992), .ZN(n17995) );
  NOR3_X1 U21250 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17980), .A3(n17995), .ZN(
        n17981) );
  AOI211_X1 U21251 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18005), .A(
        n19317), .B(n17981), .ZN(n17990) );
  AOI22_X1 U21252 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17982), .B1(
        n17993), .B2(n18913), .ZN(n18915) );
  NAND2_X1 U21253 ( .A1(n18017), .A2(n17983), .ZN(n17985) );
  OAI21_X1 U21254 ( .B1(n18915), .B2(n17985), .A(n18067), .ZN(n17984) );
  AOI21_X1 U21255 ( .B1(n18915), .B2(n17985), .A(n17984), .ZN(n17988) );
  AOI211_X1 U21256 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n18000), .A(n17986), .B(
        n18080), .ZN(n17987) );
  AOI211_X1 U21257 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n18074), .A(n17988), .B(
        n17987), .ZN(n17989) );
  OAI211_X1 U21258 ( .C1(n19877), .C2(n17991), .A(n17990), .B(n17989), .ZN(
        P3_U2663) );
  OAI21_X1 U21259 ( .B1(n17992), .B2(n18081), .A(n18091), .ZN(n18015) );
  NOR2_X1 U21260 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17995), .ZN(n18004) );
  NAND3_X1 U21261 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18941), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18008) );
  AOI21_X1 U21262 ( .B1(n18930), .B2(n18008), .A(n17993), .ZN(n18935) );
  NOR2_X1 U21263 ( .A1(n17994), .A2(n18043), .ZN(n18010) );
  XNOR2_X1 U21264 ( .A(n18935), .B(n18010), .ZN(n17998) );
  NOR2_X1 U21265 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17995), .ZN(n17996) );
  AOI22_X1 U21266 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18005), .B1(
        P3_REIP_REG_6__SCAN_IN), .B2(n17996), .ZN(n17997) );
  OAI211_X1 U21267 ( .C1(n10977), .C2(n17998), .A(n17997), .B(n19328), .ZN(
        n17999) );
  AOI221_X1 U21268 ( .B1(n18015), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n18004), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n17999), .ZN(n18002) );
  OAI211_X1 U21269 ( .C1(n18006), .C2(n18003), .A(n18090), .B(n18000), .ZN(
        n18001) );
  OAI211_X1 U21270 ( .C1(n18003), .C2(n18059), .A(n18002), .B(n18001), .ZN(
        P3_U2664) );
  AOI211_X1 U21271 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18005), .A(
        n19317), .B(n18004), .ZN(n18014) );
  AOI211_X1 U21272 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18022), .A(n18006), .B(
        n18080), .ZN(n18007) );
  AOI21_X1 U21273 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18074), .A(n18007), .ZN(
        n18013) );
  AND2_X1 U21274 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18941), .ZN(
        n18016) );
  OAI21_X1 U21275 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18016), .A(
        n18008), .ZN(n18944) );
  AOI211_X1 U21276 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18017), .A(
        n18944), .B(n18075), .ZN(n18009) );
  AOI21_X1 U21277 ( .B1(n18015), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18009), .ZN(
        n18012) );
  NAND3_X1 U21278 ( .A1(n18067), .A2(n18010), .A3(n18944), .ZN(n18011) );
  NAND4_X1 U21279 ( .A1(n18014), .A2(n18013), .A3(n18012), .A4(n18011), .ZN(
        P3_U2665) );
  NOR2_X1 U21280 ( .A1(n18081), .A2(n18040), .ZN(n18027) );
  AOI21_X1 U21281 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n18027), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18020) );
  INV_X1 U21282 ( .A(n18015), .ZN(n18019) );
  OR2_X1 U21283 ( .A1(n19006), .A2(n18957), .ZN(n18029) );
  AOI21_X1 U21284 ( .B1(n18956), .B2(n18029), .A(n18016), .ZN(n18958) );
  OAI21_X1 U21285 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18029), .A(
        n18017), .ZN(n18030) );
  XOR2_X1 U21286 ( .A(n18958), .B(n18030), .Z(n18018) );
  OAI22_X1 U21287 ( .A1(n18020), .A2(n18019), .B1(n10977), .B2(n18018), .ZN(
        n18021) );
  AOI211_X1 U21288 ( .C1(n18074), .C2(P3_EBX_REG_5__SCAN_IN), .A(n19317), .B(
        n18021), .ZN(n18024) );
  OAI211_X1 U21289 ( .C1(n18032), .C2(n18356), .A(n18090), .B(n18022), .ZN(
        n18023) );
  OAI211_X1 U21290 ( .C1(n18076), .C2(n18956), .A(n18024), .B(n18023), .ZN(
        P3_U2666) );
  AOI21_X1 U21291 ( .B1(n18055), .B2(n18040), .A(n18073), .ZN(n18052) );
  INV_X1 U21292 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21945) );
  INV_X1 U21293 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n18025) );
  OAI22_X1 U21294 ( .A1(n21945), .A2(n18076), .B1(n18059), .B2(n18025), .ZN(
        n18026) );
  AOI21_X1 U21295 ( .B1(n18027), .B2(n19869), .A(n18026), .ZN(n18038) );
  AND2_X1 U21296 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18028), .ZN(
        n18045) );
  OAI21_X1 U21297 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18045), .A(
        n18029), .ZN(n18973) );
  INV_X1 U21298 ( .A(n18973), .ZN(n18031) );
  NAND2_X1 U21299 ( .A1(n18028), .A2(n21945), .ZN(n18966) );
  OAI22_X1 U21300 ( .A1(n18031), .A2(n18030), .B1(n18065), .B2(n18966), .ZN(
        n18036) );
  AOI211_X1 U21301 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18046), .A(n18032), .B(
        n18080), .ZN(n18035) );
  NAND2_X1 U21302 ( .A1(n18067), .A2(n18043), .ZN(n18071) );
  NAND2_X1 U21303 ( .A1(n19349), .A2(n20004), .ZN(n18087) );
  INV_X1 U21304 ( .A(n18087), .ZN(n20005) );
  OAI21_X1 U21305 ( .B1(n18039), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20005), .ZN(n18033) );
  OAI211_X1 U21306 ( .C1(n18973), .C2(n18071), .A(n19328), .B(n18033), .ZN(
        n18034) );
  AOI211_X1 U21307 ( .C1(n18067), .C2(n18036), .A(n18035), .B(n18034), .ZN(
        n18037) );
  OAI211_X1 U21308 ( .C1(n18052), .C2(n19869), .A(n18038), .B(n18037), .ZN(
        P3_U2667) );
  INV_X1 U21309 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19867) );
  NOR2_X1 U21310 ( .A1(n19961), .A2(n19953), .ZN(n19786) );
  NAND2_X1 U21311 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19786), .ZN(
        n19777) );
  AOI21_X1 U21312 ( .B1(n10623), .B2(n19777), .A(n18039), .ZN(n19939) );
  NAND2_X1 U21313 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n18056) );
  NAND2_X1 U21314 ( .A1(n18055), .A2(n18040), .ZN(n18041) );
  OAI22_X1 U21315 ( .A1(n21906), .A2(n18076), .B1(n18056), .B2(n18041), .ZN(
        n18042) );
  AOI21_X1 U21316 ( .B1(n20005), .B2(n19939), .A(n18042), .ZN(n18051) );
  NAND2_X1 U21317 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18053) );
  INV_X1 U21318 ( .A(n18053), .ZN(n18044) );
  AOI21_X1 U21319 ( .B1(n18044), .B2(n18078), .A(n18043), .ZN(n18066) );
  AOI21_X1 U21320 ( .B1(n21906), .B2(n18053), .A(n18045), .ZN(n18982) );
  XOR2_X1 U21321 ( .A(n18066), .B(n18982), .Z(n18049) );
  OAI211_X1 U21322 ( .C1(n18054), .C2(n18371), .A(n18090), .B(n18046), .ZN(
        n18047) );
  OAI21_X1 U21323 ( .B1(n18371), .B2(n18059), .A(n18047), .ZN(n18048) );
  AOI21_X1 U21324 ( .B1(n18049), .B2(n18067), .A(n18048), .ZN(n18050) );
  OAI211_X1 U21325 ( .C1(n18052), .C2(n19867), .A(n18051), .B(n18050), .ZN(
        P3_U2668) );
  OAI21_X1 U21326 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18053), .ZN(n18993) );
  INV_X1 U21327 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18389) );
  INV_X1 U21328 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18383) );
  NAND2_X1 U21329 ( .A1(n18389), .A2(n18383), .ZN(n18079) );
  AOI211_X1 U21330 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18079), .A(n18054), .B(
        n18080), .ZN(n18064) );
  OAI211_X1 U21331 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n18056), .B(n18055), .ZN(n18057) );
  INV_X1 U21332 ( .A(n18057), .ZN(n18063) );
  INV_X1 U21333 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19865) );
  OAI22_X1 U21334 ( .A1(n18059), .A2(n18058), .B1(n18091), .B2(n19865), .ZN(
        n18062) );
  NAND2_X1 U21335 ( .A1(n19787), .A2(n19953), .ZN(n19776) );
  NAND2_X1 U21336 ( .A1(n19777), .A2(n19776), .ZN(n19947) );
  OAI22_X1 U21337 ( .A1(n18060), .A2(n18076), .B1(n19947), .B2(n18087), .ZN(
        n18061) );
  NOR4_X1 U21338 ( .A1(n18064), .A2(n18063), .A3(n18062), .A4(n18061), .ZN(
        n18070) );
  INV_X1 U21339 ( .A(n18065), .ZN(n18068) );
  OAI211_X1 U21340 ( .C1(n18068), .C2(n18993), .A(n18067), .B(n18066), .ZN(
        n18069) );
  OAI211_X1 U21341 ( .C1(n18071), .C2(n18993), .A(n18070), .B(n18069), .ZN(
        P3_U2669) );
  NAND2_X1 U21342 ( .A1(n19787), .A2(n18072), .ZN(n19954) );
  AOI22_X1 U21343 ( .A1(n18074), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n18073), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18086) );
  INV_X1 U21344 ( .A(n18075), .ZN(n18084) );
  OAI21_X1 U21345 ( .B1(n18078), .B2(n18077), .A(n18076), .ZN(n18083) );
  NAND2_X1 U21346 ( .A1(n18079), .A2(n18376), .ZN(n18384) );
  OAI22_X1 U21347 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18081), .B1(n18080), 
        .B2(n18384), .ZN(n18082) );
  AOI221_X1 U21348 ( .B1(n18084), .B2(n19006), .C1(n18083), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n18082), .ZN(n18085) );
  OAI211_X1 U21349 ( .C1(n19954), .C2(n18087), .A(n18086), .B(n18085), .ZN(
        P3_U2670) );
  AOI22_X1 U21350 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n18089), .B1(n20005), 
        .B2(n19967), .ZN(n18094) );
  OAI21_X1 U21351 ( .B1(n18074), .B2(n18090), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n18093) );
  NAND3_X1 U21352 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19949), .A3(
        n18091), .ZN(n18092) );
  NAND3_X1 U21353 ( .A1(n18094), .A2(n18093), .A3(n18092), .ZN(P3_U2671) );
  NAND4_X1 U21354 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n18095)
         );
  NOR4_X1 U21355 ( .A1(n18098), .A2(n18097), .A3(n18096), .A4(n18095), .ZN(
        n18099) );
  NAND4_X1 U21356 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n18181), .A4(n18099), .ZN(n18102) );
  NAND2_X1 U21357 ( .A1(n18379), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18101) );
  NAND2_X1 U21358 ( .A1(n18129), .A2(n19375), .ZN(n18100) );
  OAI22_X1 U21359 ( .A1(n18129), .A2(n18101), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18100), .ZN(P3_U2672) );
  NAND2_X1 U21360 ( .A1(n18103), .A2(n18102), .ZN(n18104) );
  NAND2_X1 U21361 ( .A1(n18104), .A2(n18379), .ZN(n18128) );
  AOI22_X1 U21362 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18115) );
  AOI22_X1 U21363 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18114) );
  AOI22_X1 U21364 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18105) );
  OAI21_X1 U21365 ( .B1(n18106), .B2(n18357), .A(n18105), .ZN(n18112) );
  AOI22_X1 U21366 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18110) );
  AOI22_X1 U21367 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18109) );
  AOI22_X1 U21368 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18108) );
  AOI22_X1 U21369 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18107) );
  NAND4_X1 U21370 ( .A1(n18110), .A2(n18109), .A3(n18108), .A4(n18107), .ZN(
        n18111) );
  AOI211_X1 U21371 ( .C1(n18320), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n18112), .B(n18111), .ZN(n18113) );
  NAND3_X1 U21372 ( .A1(n18115), .A2(n18114), .A3(n18113), .ZN(n18127) );
  AOI22_X1 U21373 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18125) );
  AOI22_X1 U21374 ( .A1(n18312), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18343), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18124) );
  AOI22_X1 U21375 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18116) );
  OAI21_X1 U21376 ( .B1(n9732), .B2(n21817), .A(n18116), .ZN(n18122) );
  AOI22_X1 U21377 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18120) );
  AOI22_X1 U21378 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18119) );
  AOI22_X1 U21379 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18118) );
  AOI22_X1 U21380 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18117) );
  NAND4_X1 U21381 ( .A1(n18120), .A2(n18119), .A3(n18118), .A4(n18117), .ZN(
        n18121) );
  AOI211_X1 U21382 ( .C1(n18313), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n18122), .B(n18121), .ZN(n18123) );
  AND3_X1 U21383 ( .A1(n18125), .A2(n18124), .A3(n18123), .ZN(n18132) );
  NOR3_X1 U21384 ( .A1(n18132), .A2(n18131), .A3(n18136), .ZN(n18126) );
  XNOR2_X1 U21385 ( .A(n18127), .B(n18126), .ZN(n18400) );
  OAI22_X1 U21386 ( .A1(n18129), .A2(n18128), .B1(n18400), .B2(n18379), .ZN(
        P3_U2673) );
  NAND2_X1 U21387 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18140), .ZN(n18135) );
  NOR2_X1 U21388 ( .A1(n18136), .A2(n18131), .ZN(n18133) );
  XOR2_X1 U21389 ( .A(n18133), .B(n18132), .Z(n18408) );
  NAND3_X1 U21390 ( .A1(n18135), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n18379), 
        .ZN(n18134) );
  OAI221_X1 U21391 ( .B1(n18135), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n18379), 
        .C2(n18408), .A(n18134), .ZN(P3_U2674) );
  AOI21_X1 U21392 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18379), .A(n18143), .ZN(
        n18139) );
  OAI21_X1 U21393 ( .B1(n18138), .B2(n18137), .A(n18136), .ZN(n18416) );
  OAI22_X1 U21394 ( .A1(n18140), .A2(n18139), .B1(n18379), .B2(n18416), .ZN(
        P3_U2676) );
  AOI21_X1 U21395 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18379), .A(n18148), .ZN(
        n18142) );
  XNOR2_X1 U21396 ( .A(n18141), .B(n18144), .ZN(n18420) );
  OAI22_X1 U21397 ( .A1(n18143), .A2(n18142), .B1(n18379), .B2(n18420), .ZN(
        P3_U2677) );
  AOI21_X1 U21398 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18379), .A(n18151), .ZN(
        n18147) );
  OAI21_X1 U21399 ( .B1(n18146), .B2(n18145), .A(n18144), .ZN(n18425) );
  OAI22_X1 U21400 ( .A1(n18148), .A2(n18147), .B1(n18379), .B2(n18425), .ZN(
        P3_U2678) );
  AOI21_X1 U21401 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18379), .A(n18157), .ZN(
        n18150) );
  XNOR2_X1 U21402 ( .A(n18149), .B(n18153), .ZN(n18431) );
  OAI22_X1 U21403 ( .A1(n18151), .A2(n18150), .B1(n18379), .B2(n18431), .ZN(
        P3_U2679) );
  INV_X1 U21404 ( .A(n18170), .ZN(n18152) );
  AOI22_X1 U21405 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n18379), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n18152), .ZN(n18156) );
  OAI21_X1 U21406 ( .B1(n18155), .B2(n18154), .A(n18153), .ZN(n18437) );
  OAI22_X1 U21407 ( .A1(n18157), .A2(n18156), .B1(n18379), .B2(n18437), .ZN(
        P3_U2680) );
  AOI22_X1 U21408 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18167) );
  AOI22_X1 U21409 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18343), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18166) );
  AOI22_X1 U21410 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18158) );
  OAI21_X1 U21411 ( .B1(n18239), .B2(n21817), .A(n18158), .ZN(n18164) );
  AOI22_X1 U21412 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18162) );
  AOI22_X1 U21413 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U21414 ( .A1(n18315), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18160) );
  AOI22_X1 U21415 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18159) );
  NAND4_X1 U21416 ( .A1(n18162), .A2(n18161), .A3(n18160), .A4(n18159), .ZN(
        n18163) );
  AOI211_X1 U21417 ( .C1(n18334), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n18164), .B(n18163), .ZN(n18165) );
  NAND3_X1 U21418 ( .A1(n18167), .A2(n18166), .A3(n18165), .ZN(n18438) );
  INV_X1 U21419 ( .A(n18438), .ZN(n18169) );
  NAND3_X1 U21420 ( .A1(n18170), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n18379), 
        .ZN(n18168) );
  OAI221_X1 U21421 ( .B1(n18170), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n18379), 
        .C2(n18169), .A(n18168), .ZN(P3_U2681) );
  AOI22_X1 U21422 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18174) );
  AOI22_X1 U21423 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18345), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18173) );
  AOI22_X1 U21424 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18172) );
  AOI22_X1 U21425 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18171) );
  NAND4_X1 U21426 ( .A1(n18174), .A2(n18173), .A3(n18172), .A4(n18171), .ZN(
        n18180) );
  AOI22_X1 U21427 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18178) );
  AOI22_X1 U21428 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18177) );
  AOI22_X1 U21429 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18313), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18176) );
  AOI22_X1 U21430 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18175) );
  NAND4_X1 U21431 ( .A1(n18178), .A2(n18177), .A3(n18176), .A4(n18175), .ZN(
        n18179) );
  NOR2_X1 U21432 ( .A1(n18180), .A2(n18179), .ZN(n18445) );
  NOR2_X1 U21433 ( .A1(n18387), .A2(n18181), .ZN(n18196) );
  AOI22_X1 U21434 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18196), .B1(n18183), 
        .B2(n18182), .ZN(n18184) );
  OAI21_X1 U21435 ( .B1(n18445), .B2(n18379), .A(n18184), .ZN(P3_U2682) );
  AOI22_X1 U21436 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18188) );
  AOI22_X1 U21437 ( .A1(n12808), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17439), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18187) );
  AOI22_X1 U21438 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18186) );
  AOI22_X1 U21439 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9743), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18185) );
  NAND4_X1 U21440 ( .A1(n18188), .A2(n18187), .A3(n18186), .A4(n18185), .ZN(
        n18194) );
  AOI22_X1 U21441 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18192) );
  AOI22_X1 U21442 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U21443 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18312), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18190) );
  AOI22_X1 U21444 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18189) );
  NAND4_X1 U21445 ( .A1(n18192), .A2(n18191), .A3(n18190), .A4(n18189), .ZN(
        n18193) );
  NOR2_X1 U21446 ( .A1(n18194), .A2(n18193), .ZN(n18452) );
  NOR2_X1 U21447 ( .A1(n18195), .A2(n18224), .ZN(n18197) );
  NOR2_X1 U21448 ( .A1(n18501), .A2(n9832), .ZN(n18222) );
  OAI221_X1 U21449 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18197), .C1(
        P3_EBX_REG_20__SCAN_IN), .C2(n18222), .A(n18196), .ZN(n18198) );
  OAI21_X1 U21450 ( .B1(n18452), .B2(n18379), .A(n18198), .ZN(P3_U2683) );
  AOI22_X1 U21451 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18379), .B1(
        P3_EBX_REG_18__SCAN_IN), .B2(n18222), .ZN(n18209) );
  AOI22_X1 U21452 ( .A1(n18312), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U21453 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18201) );
  AOI22_X1 U21454 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12810), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18200) );
  AOI22_X1 U21455 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18199) );
  NAND4_X1 U21456 ( .A1(n18202), .A2(n18201), .A3(n18200), .A4(n18199), .ZN(
        n18208) );
  AOI22_X1 U21457 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18206) );
  AOI22_X1 U21458 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18343), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18205) );
  AOI22_X1 U21459 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18204) );
  AOI22_X1 U21460 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18203) );
  NAND4_X1 U21461 ( .A1(n18206), .A2(n18205), .A3(n18204), .A4(n18203), .ZN(
        n18207) );
  NOR2_X1 U21462 ( .A1(n18208), .A2(n18207), .ZN(n18457) );
  OAI22_X1 U21463 ( .A1(n18210), .A2(n18209), .B1(n18457), .B2(n18379), .ZN(
        P3_U2684) );
  NAND2_X1 U21464 ( .A1(n18379), .A2(n9832), .ZN(n18236) );
  AOI22_X1 U21465 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18221) );
  AOI22_X1 U21466 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18220) );
  AOI22_X1 U21467 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18211) );
  OAI21_X1 U21468 ( .B1(n9747), .B2(n18381), .A(n18211), .ZN(n18218) );
  AOI22_X1 U21469 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U21470 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18215) );
  AOI22_X1 U21471 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18214) );
  AOI22_X1 U21472 ( .A1(n18212), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18213) );
  NAND4_X1 U21473 ( .A1(n18216), .A2(n18215), .A3(n18214), .A4(n18213), .ZN(
        n18217) );
  AOI211_X1 U21474 ( .C1(n18334), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n18218), .B(n18217), .ZN(n18219) );
  NAND3_X1 U21475 ( .A1(n18221), .A2(n18220), .A3(n18219), .ZN(n18458) );
  AOI22_X1 U21476 ( .A1(n18387), .A2(n18458), .B1(n18222), .B2(n18224), .ZN(
        n18223) );
  OAI21_X1 U21477 ( .B1(n18224), .B2(n18236), .A(n18223), .ZN(P3_U2685) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18333), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18228) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18320), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18227) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18312), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18297), .ZN(n18226) );
  AOI22_X1 U21481 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18315), .ZN(n18225) );
  NAND4_X1 U21482 ( .A1(n18228), .A2(n18227), .A3(n18226), .A4(n18225), .ZN(
        n18234) );
  AOI22_X1 U21483 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U21484 ( .A1(n12808), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n18268), .ZN(n18231) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18322), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18230) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17456), .B1(
        n17439), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18229) );
  NAND4_X1 U21487 ( .A1(n18232), .A2(n18231), .A3(n18230), .A4(n18229), .ZN(
        n18233) );
  NOR2_X1 U21488 ( .A1(n18234), .A2(n18233), .ZN(n18469) );
  AND2_X1 U21489 ( .A1(n18235), .A2(n18249), .ZN(n18237) );
  OAI22_X1 U21490 ( .A1(n18469), .A2(n18379), .B1(n18237), .B2(n18236), .ZN(
        P3_U2686) );
  AOI22_X1 U21491 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18248) );
  AOI22_X1 U21492 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18247) );
  AOI22_X1 U21493 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18238) );
  OAI21_X1 U21494 ( .B1(n18239), .B2(n21848), .A(n18238), .ZN(n18245) );
  AOI22_X1 U21495 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18243) );
  AOI22_X1 U21496 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18242) );
  AOI22_X1 U21497 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18241) );
  AOI22_X1 U21498 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18240) );
  NAND4_X1 U21499 ( .A1(n18243), .A2(n18242), .A3(n18241), .A4(n18240), .ZN(
        n18244) );
  AOI211_X1 U21500 ( .C1(n18340), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n18245), .B(n18244), .ZN(n18246) );
  NAND3_X1 U21501 ( .A1(n18248), .A2(n18247), .A3(n18246), .ZN(n18470) );
  INV_X1 U21502 ( .A(n18470), .ZN(n18251) );
  OAI21_X1 U21503 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18265), .A(n18249), .ZN(
        n18250) );
  AOI22_X1 U21504 ( .A1(n18387), .A2(n18251), .B1(n18250), .B2(n18379), .ZN(
        P3_U2687) );
  INV_X1 U21505 ( .A(n18252), .ZN(n18253) );
  OAI21_X1 U21506 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n18253), .A(n18379), .ZN(
        n18264) );
  AOI22_X1 U21507 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U21508 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18256) );
  AOI22_X1 U21509 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18255) );
  AOI22_X1 U21510 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12810), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18254) );
  NAND4_X1 U21511 ( .A1(n18257), .A2(n18256), .A3(n18255), .A4(n18254), .ZN(
        n18263) );
  AOI22_X1 U21512 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18261) );
  AOI22_X1 U21513 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18260) );
  AOI22_X1 U21514 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18259) );
  AOI22_X1 U21515 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18258) );
  NAND4_X1 U21516 ( .A1(n18261), .A2(n18260), .A3(n18259), .A4(n18258), .ZN(
        n18262) );
  NOR2_X1 U21517 ( .A1(n18263), .A2(n18262), .ZN(n18479) );
  OAI22_X1 U21518 ( .A1(n18265), .A2(n18264), .B1(n18479), .B2(n18379), .ZN(
        P3_U2688) );
  INV_X1 U21519 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18283) );
  AOI22_X1 U21520 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18340), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18277) );
  AOI22_X1 U21521 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18276) );
  AOI22_X1 U21522 ( .A1(n18314), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18266) );
  OAI21_X1 U21523 ( .B1(n18267), .B2(n21817), .A(n18266), .ZN(n18274) );
  AOI22_X1 U21524 ( .A1(n18268), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18272) );
  AOI22_X1 U21525 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18271) );
  AOI22_X1 U21526 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U21527 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18269) );
  NAND4_X1 U21528 ( .A1(n18272), .A2(n18271), .A3(n18270), .A4(n18269), .ZN(
        n18273) );
  AOI211_X1 U21529 ( .C1(n18313), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n18274), .B(n18273), .ZN(n18275) );
  NAND3_X1 U21530 ( .A1(n18277), .A2(n18276), .A3(n18275), .ZN(n18480) );
  NOR2_X1 U21531 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18501), .ZN(n18278) );
  AOI22_X1 U21532 ( .A1(n18387), .A2(n18480), .B1(n18279), .B2(n18278), .ZN(
        n18280) );
  OAI221_X1 U21533 ( .B1(n18283), .B2(n18282), .C1(n18283), .C2(n18281), .A(
        n18280), .ZN(P3_U2689) );
  AOI22_X1 U21534 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18288) );
  AOI22_X1 U21535 ( .A1(n18284), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18287) );
  AOI22_X1 U21536 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18312), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18286) );
  AOI22_X1 U21537 ( .A1(n18341), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12810), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18285) );
  NAND4_X1 U21538 ( .A1(n18288), .A2(n18287), .A3(n18286), .A4(n18285), .ZN(
        n18294) );
  AOI22_X1 U21539 ( .A1(n12808), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18292) );
  AOI22_X1 U21540 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18291) );
  AOI22_X1 U21541 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18290) );
  AOI22_X1 U21542 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18314), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18289) );
  NAND4_X1 U21543 ( .A1(n18292), .A2(n18291), .A3(n18290), .A4(n18289), .ZN(
        n18293) );
  NOR2_X1 U21544 ( .A1(n18294), .A2(n18293), .ZN(n18489) );
  OAI21_X1 U21545 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n9936), .A(n18295), .ZN(
        n18296) );
  OAI21_X1 U21546 ( .B1(n18489), .B2(n18379), .A(n18296), .ZN(P3_U2691) );
  AOI22_X1 U21547 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18301) );
  AOI22_X1 U21548 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18300) );
  AOI22_X1 U21549 ( .A1(n18297), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18333), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18299) );
  AOI22_X1 U21550 ( .A1(n18320), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18315), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18298) );
  NAND4_X1 U21551 ( .A1(n18301), .A2(n18300), .A3(n18299), .A4(n18298), .ZN(
        n18307) );
  AOI22_X1 U21552 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18305) );
  AOI22_X1 U21553 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18304) );
  AOI22_X1 U21554 ( .A1(n12808), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18344), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18303) );
  AOI22_X1 U21555 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18302) );
  NAND4_X1 U21556 ( .A1(n18305), .A2(n18304), .A3(n18303), .A4(n18302), .ZN(
        n18306) );
  NOR2_X1 U21557 ( .A1(n18307), .A2(n18306), .ZN(n18498) );
  AOI21_X1 U21558 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18330), .A(n18387), .ZN(
        n18329) );
  NOR3_X1 U21559 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18309), .A3(n18308), .ZN(
        n18310) );
  AOI22_X1 U21560 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18329), .B1(n18386), 
        .B2(n18310), .ZN(n18311) );
  OAI21_X1 U21561 ( .B1(n18498), .B2(n18379), .A(n18311), .ZN(P3_U2693) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18313), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18312), .ZN(n18319) );
  AOI22_X1 U21563 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18341), .ZN(n18318) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18314), .B1(
        n18343), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18317) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9744), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17456), .ZN(n18316) );
  NAND4_X1 U21566 ( .A1(n18319), .A2(n18318), .A3(n18317), .A4(n18316), .ZN(
        n18328) );
  AOI22_X1 U21567 ( .A1(n18039), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18326) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18340), .B1(
        n18320), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18325) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18333), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18324) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18322), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18323) );
  NAND4_X1 U21571 ( .A1(n18326), .A2(n18325), .A3(n18324), .A4(n18323), .ZN(
        n18327) );
  NOR2_X1 U21572 ( .A1(n18328), .A2(n18327), .ZN(n18502) );
  OAI21_X1 U21573 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18330), .A(n18329), .ZN(
        n18331) );
  OAI21_X1 U21574 ( .B1(n18502), .B2(n18379), .A(n18331), .ZN(P3_U2694) );
  AOI22_X1 U21575 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18322), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U21576 ( .A1(n18333), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18332), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18338) );
  AOI22_X1 U21577 ( .A1(n18335), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18337) );
  AOI22_X1 U21578 ( .A1(n18313), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9744), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18336) );
  NAND4_X1 U21579 ( .A1(n18339), .A2(n18338), .A3(n18337), .A4(n18336), .ZN(
        n18351) );
  AOI22_X1 U21580 ( .A1(n18340), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18321), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18349) );
  AOI22_X1 U21581 ( .A1(n18342), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18341), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18348) );
  AOI22_X1 U21582 ( .A1(n18344), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18343), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18347) );
  AOI22_X1 U21583 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18268), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18346) );
  NAND4_X1 U21584 ( .A1(n18349), .A2(n18348), .A3(n18347), .A4(n18346), .ZN(
        n18350) );
  NOR2_X1 U21585 ( .A1(n18351), .A2(n18350), .ZN(n18508) );
  NOR2_X1 U21586 ( .A1(n18353), .A2(n18352), .ZN(n18359) );
  OAI21_X1 U21587 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n18359), .A(n18354), .ZN(
        n18355) );
  AOI22_X1 U21588 ( .A1(n18387), .A2(n18508), .B1(n18355), .B2(n18379), .ZN(
        P3_U2695) );
  NAND2_X1 U21589 ( .A1(n19375), .A2(n18364), .ZN(n18368) );
  NOR2_X1 U21590 ( .A1(n18356), .A2(n18368), .ZN(n18360) );
  AOI22_X1 U21591 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n18379), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n18360), .ZN(n18358) );
  OAI22_X1 U21592 ( .A1(n18359), .A2(n18358), .B1(n18357), .B2(n18379), .ZN(
        P3_U2696) );
  INV_X1 U21593 ( .A(n18360), .ZN(n18363) );
  INV_X1 U21594 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18362) );
  NAND3_X1 U21595 ( .A1(n18363), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n18379), .ZN(
        n18361) );
  OAI221_X1 U21596 ( .B1(n18363), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n18379), 
        .C2(n18362), .A(n18361), .ZN(P3_U2697) );
  INV_X1 U21597 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18366) );
  OAI211_X1 U21598 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n18364), .A(n18363), .B(
        n18379), .ZN(n18365) );
  OAI21_X1 U21599 ( .B1(n18379), .B2(n18366), .A(n18365), .ZN(P3_U2698) );
  NAND2_X1 U21600 ( .A1(n18367), .A2(n18386), .ZN(n18377) );
  NOR2_X1 U21601 ( .A1(n18371), .A2(n18377), .ZN(n18375) );
  OAI211_X1 U21602 ( .C1(n18375), .C2(P3_EBX_REG_4__SCAN_IN), .A(n18379), .B(
        n18368), .ZN(n18369) );
  OAI21_X1 U21603 ( .B1(n18379), .B2(n18370), .A(n18369), .ZN(P3_U2699) );
  OAI21_X1 U21604 ( .B1(n18371), .B2(n18387), .A(n18377), .ZN(n18372) );
  INV_X1 U21605 ( .A(n18372), .ZN(n18374) );
  INV_X1 U21606 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18373) );
  OAI22_X1 U21607 ( .A1(n18375), .A2(n18374), .B1(n18373), .B2(n18379), .ZN(
        P3_U2700) );
  INV_X1 U21608 ( .A(n18376), .ZN(n18378) );
  OAI221_X1 U21609 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n18390), .C1(
        P3_EBX_REG_2__SCAN_IN), .C2(n18378), .A(n18377), .ZN(n18380) );
  AOI22_X1 U21610 ( .A1(n18387), .A2(n18381), .B1(n18380), .B2(n18379), .ZN(
        P3_U2701) );
  INV_X1 U21611 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18382) );
  OAI222_X1 U21612 ( .A1(n18385), .A2(n18384), .B1(n18383), .B2(n18390), .C1(
        n18382), .C2(n18379), .ZN(P3_U2702) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18387), .B1(
        n18386), .B2(n18389), .ZN(n18388) );
  OAI21_X1 U21614 ( .B1(n18390), .B2(n18389), .A(n18388), .ZN(P3_U2703) );
  NAND2_X1 U21615 ( .A1(n18531), .A2(n18391), .ZN(n18444) );
  INV_X1 U21616 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18619) );
  INV_X1 U21617 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18616) );
  INV_X1 U21618 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18614) );
  INV_X1 U21619 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18565) );
  NAND2_X1 U21620 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n18509) );
  NAND4_X1 U21621 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n18394)
         );
  NAND3_X1 U21622 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_13__SCAN_IN), .ZN(n18393) );
  AND4_X1 U21623 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n18440)
         );
  INV_X1 U21624 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18612) );
  NAND2_X1 U21625 ( .A1(n19375), .A2(n18432), .ZN(n18426) );
  NAND2_X1 U21626 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18405), .ZN(n18404) );
  NOR2_X1 U21627 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n18404), .ZN(n18397) );
  NAND2_X1 U21628 ( .A1(n18523), .A2(n18404), .ZN(n18403) );
  OAI21_X1 U21629 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18539), .A(n18403), .ZN(
        n18396) );
  AOI22_X1 U21630 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18397), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18396), .ZN(n18398) );
  OAI21_X1 U21631 ( .B1(n20178), .B2(n18444), .A(n18398), .ZN(P3_U2704) );
  INV_X1 U21632 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18624) );
  OAI22_X1 U21633 ( .A1(n18400), .A2(n18525), .B1(n16511), .B2(n18444), .ZN(
        n18401) );
  AOI21_X1 U21634 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18463), .A(n18401), .ZN(
        n18402) );
  OAI221_X1 U21635 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18404), .C1(n18624), 
        .C2(n18403), .A(n18402), .ZN(P3_U2705) );
  AOI22_X1 U21636 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18463), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18471), .ZN(n18407) );
  OAI211_X1 U21637 ( .C1(n18405), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18523), .B(
        n18404), .ZN(n18406) );
  OAI211_X1 U21638 ( .C1(n18525), .C2(n18408), .A(n18407), .B(n18406), .ZN(
        P3_U2706) );
  AOI22_X1 U21639 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18463), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18471), .ZN(n18411) );
  OAI211_X1 U21640 ( .C1(n9837), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18523), .B(
        n18409), .ZN(n18410) );
  OAI211_X1 U21641 ( .C1(n18525), .C2(n18412), .A(n18411), .B(n18410), .ZN(
        P3_U2707) );
  AOI22_X1 U21642 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18463), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18471), .ZN(n18415) );
  AOI211_X1 U21643 ( .C1(n18619), .C2(n18417), .A(n9837), .B(n18531), .ZN(
        n18413) );
  INV_X1 U21644 ( .A(n18413), .ZN(n18414) );
  OAI211_X1 U21645 ( .C1(n18416), .C2(n18525), .A(n18415), .B(n18414), .ZN(
        P3_U2708) );
  AOI22_X1 U21646 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18463), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18471), .ZN(n18419) );
  OAI211_X1 U21647 ( .C1(n18421), .C2(P3_EAX_REG_26__SCAN_IN), .A(n18523), .B(
        n18417), .ZN(n18418) );
  OAI211_X1 U21648 ( .C1(n18420), .C2(n18525), .A(n18419), .B(n18418), .ZN(
        P3_U2709) );
  AOI22_X1 U21649 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18463), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18471), .ZN(n18424) );
  AOI211_X1 U21650 ( .C1(n18616), .C2(n18427), .A(n18421), .B(n18531), .ZN(
        n18422) );
  INV_X1 U21651 ( .A(n18422), .ZN(n18423) );
  OAI211_X1 U21652 ( .C1(n18425), .C2(n18525), .A(n18424), .B(n18423), .ZN(
        P3_U2710) );
  AOI22_X1 U21653 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18463), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18471), .ZN(n18430) );
  OAI21_X1 U21654 ( .B1(n18614), .B2(n18531), .A(n18426), .ZN(n18428) );
  NAND2_X1 U21655 ( .A1(n18428), .A2(n18427), .ZN(n18429) );
  OAI211_X1 U21656 ( .C1(n18431), .C2(n18525), .A(n18430), .B(n18429), .ZN(
        P3_U2711) );
  AOI211_X1 U21657 ( .C1(n18612), .C2(n18433), .A(n18531), .B(n18432), .ZN(
        n18434) );
  AOI21_X1 U21658 ( .B1(n18471), .B2(BUF2_REG_23__SCAN_IN), .A(n18434), .ZN(
        n18436) );
  NAND2_X1 U21659 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18463), .ZN(n18435) );
  OAI211_X1 U21660 ( .C1(n18437), .C2(n18525), .A(n18436), .B(n18435), .ZN(
        P3_U2712) );
  INV_X1 U21661 ( .A(n18463), .ZN(n18475) );
  AOI22_X1 U21662 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18471), .B1(n18537), .B2(
        n18438), .ZN(n18443) );
  INV_X1 U21663 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18605) );
  INV_X1 U21664 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18601) );
  NAND2_X1 U21665 ( .A1(n19375), .A2(n9833), .ZN(n18464) );
  NAND2_X1 U21666 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18460), .ZN(n18459) );
  NAND2_X1 U21667 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18453), .ZN(n18449) );
  NAND2_X1 U21668 ( .A1(n18523), .A2(n18449), .ZN(n18448) );
  OAI21_X1 U21669 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18539), .A(n18448), .ZN(
        n18441) );
  INV_X1 U21670 ( .A(n18460), .ZN(n18465) );
  NOR2_X1 U21671 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18465), .ZN(n18439) );
  AOI22_X1 U21672 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18441), .B1(n18440), 
        .B2(n18439), .ZN(n18442) );
  OAI211_X1 U21673 ( .C1(n13839), .C2(n18475), .A(n18443), .B(n18442), .ZN(
        P3_U2713) );
  INV_X1 U21674 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18608) );
  OAI22_X1 U21675 ( .A1(n18445), .A2(n18525), .B1(n16581), .B2(n18444), .ZN(
        n18446) );
  AOI21_X1 U21676 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n18463), .A(n18446), .ZN(
        n18447) );
  OAI221_X1 U21677 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18449), .C1(n18608), 
        .C2(n18448), .A(n18447), .ZN(P3_U2714) );
  AOI22_X1 U21678 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18463), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18471), .ZN(n18451) );
  OAI211_X1 U21679 ( .C1(n18453), .C2(P3_EAX_REG_20__SCAN_IN), .A(n18523), .B(
        n18449), .ZN(n18450) );
  OAI211_X1 U21680 ( .C1(n18452), .C2(n18525), .A(n18451), .B(n18450), .ZN(
        P3_U2715) );
  AOI22_X1 U21681 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18463), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18471), .ZN(n18456) );
  AOI211_X1 U21682 ( .C1(n18605), .C2(n18459), .A(n18453), .B(n18531), .ZN(
        n18454) );
  INV_X1 U21683 ( .A(n18454), .ZN(n18455) );
  OAI211_X1 U21684 ( .C1(n18457), .C2(n18525), .A(n18456), .B(n18455), .ZN(
        P3_U2716) );
  AOI22_X1 U21685 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n18471), .B1(n18537), .B2(
        n18458), .ZN(n18462) );
  OAI211_X1 U21686 ( .C1(n18460), .C2(P3_EAX_REG_18__SCAN_IN), .A(n18523), .B(
        n18459), .ZN(n18461) );
  OAI211_X1 U21687 ( .C1(n18475), .C2(n19354), .A(n18462), .B(n18461), .ZN(
        P3_U2717) );
  AOI22_X1 U21688 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18463), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18471), .ZN(n18468) );
  OAI21_X1 U21689 ( .B1(n18601), .B2(n18531), .A(n18464), .ZN(n18466) );
  NAND2_X1 U21690 ( .A1(n18466), .A2(n18465), .ZN(n18467) );
  OAI211_X1 U21691 ( .C1(n18469), .C2(n18525), .A(n18468), .B(n18467), .ZN(
        P3_U2718) );
  AOI22_X1 U21692 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n18471), .B1(n18537), .B2(
        n18470), .ZN(n18474) );
  AOI211_X1 U21693 ( .C1(n18565), .C2(n18476), .A(n18531), .B(n9833), .ZN(
        n18472) );
  INV_X1 U21694 ( .A(n18472), .ZN(n18473) );
  OAI211_X1 U21695 ( .C1(n18475), .C2(n19345), .A(n18474), .B(n18473), .ZN(
        P3_U2719) );
  OAI211_X1 U21696 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n18481), .A(n18523), .B(
        n18476), .ZN(n18478) );
  NAND2_X1 U21697 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18538), .ZN(n18477) );
  OAI211_X1 U21698 ( .C1(n18479), .C2(n18525), .A(n18478), .B(n18477), .ZN(
        P3_U2720) );
  INV_X1 U21699 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18573) );
  INV_X1 U21700 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18577) );
  NAND4_X1 U21701 ( .A1(n19375), .A2(n18500), .A3(P3_EAX_REG_9__SCAN_IN), .A4(
        P3_EAX_REG_8__SCAN_IN), .ZN(n18499) );
  NAND2_X1 U21702 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18495), .ZN(n18488) );
  NOR2_X1 U21703 ( .A1(n18573), .A2(n18488), .ZN(n18491) );
  NAND2_X1 U21704 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18491), .ZN(n18484) );
  AOI22_X1 U21705 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18538), .B1(n18537), .B2(
        n18480), .ZN(n18483) );
  INV_X1 U21706 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18647) );
  OR3_X1 U21707 ( .A1(n18647), .A2(n18531), .A3(n18481), .ZN(n18482) );
  OAI211_X1 U21708 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n18484), .A(n18483), .B(
        n18482), .ZN(P3_U2721) );
  INV_X1 U21709 ( .A(n18484), .ZN(n18487) );
  AOI21_X1 U21710 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18523), .A(n18491), .ZN(
        n18486) );
  OAI222_X1 U21711 ( .A1(n18528), .A2(n13833), .B1(n18487), .B2(n18486), .C1(
        n18525), .C2(n18485), .ZN(P3_U2722) );
  INV_X1 U21712 ( .A(n18488), .ZN(n18494) );
  AOI21_X1 U21713 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18523), .A(n18494), .ZN(
        n18490) );
  OAI222_X1 U21714 ( .A1(n18528), .A2(n18642), .B1(n18491), .B2(n18490), .C1(
        n18525), .C2(n18489), .ZN(P3_U2723) );
  AOI21_X1 U21715 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18523), .A(n18495), .ZN(
        n18493) );
  OAI222_X1 U21716 ( .A1(n18528), .A2(n13817), .B1(n18494), .B2(n18493), .C1(
        n18525), .C2(n18492), .ZN(P3_U2724) );
  AOI211_X1 U21717 ( .C1(n18577), .C2(n18499), .A(n18531), .B(n18495), .ZN(
        n18496) );
  AOI21_X1 U21718 ( .B1(n18538), .B2(BUF2_REG_10__SCAN_IN), .A(n18496), .ZN(
        n18497) );
  OAI21_X1 U21719 ( .B1(n18498), .B2(n18525), .A(n18497), .ZN(P3_U2725) );
  INV_X1 U21720 ( .A(n18499), .ZN(n18504) );
  INV_X1 U21721 ( .A(n18500), .ZN(n18505) );
  NOR2_X1 U21722 ( .A1(n18501), .A2(n18505), .ZN(n18512) );
  AOI22_X1 U21723 ( .A1(n18512), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n18523), .ZN(n18503) );
  OAI222_X1 U21724 ( .A1(n18528), .A2(n13821), .B1(n18504), .B2(n18503), .C1(
        n18525), .C2(n18502), .ZN(P3_U2726) );
  INV_X1 U21725 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18635) );
  AOI22_X1 U21726 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18538), .B1(n18512), .B2(
        n18635), .ZN(n18507) );
  NAND3_X1 U21727 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18523), .A3(n18505), .ZN(
        n18506) );
  OAI211_X1 U21728 ( .C1(n18508), .C2(n18525), .A(n18507), .B(n18506), .ZN(
        P3_U2727) );
  INV_X1 U21729 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18590) );
  NOR2_X1 U21730 ( .A1(n18594), .A2(n18539), .ZN(n18542) );
  NAND2_X1 U21731 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n18542), .ZN(n18530) );
  NAND2_X1 U21732 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18529), .ZN(n18519) );
  NOR2_X1 U21733 ( .A1(n18509), .A2(n18519), .ZN(n18518) );
  AOI22_X1 U21734 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18523), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n18518), .ZN(n18511) );
  OAI222_X1 U21735 ( .A1(n18528), .A2(n13920), .B1(n18512), .B2(n18511), .C1(
        n18525), .C2(n18510), .ZN(P3_U2728) );
  AOI21_X1 U21736 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18523), .A(n18518), .ZN(
        n18515) );
  AND2_X1 U21737 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18518), .ZN(n18514) );
  OAI222_X1 U21738 ( .A1(n18528), .A2(n13839), .B1(n18515), .B2(n18514), .C1(
        n18525), .C2(n18513), .ZN(P3_U2729) );
  INV_X1 U21739 ( .A(n18519), .ZN(n18527) );
  AOI22_X1 U21740 ( .A1(n18527), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n18523), .ZN(n18517) );
  OAI222_X1 U21741 ( .A1(n13829), .A2(n18528), .B1(n18518), .B2(n18517), .C1(
        n18525), .C2(n18516), .ZN(P3_U2730) );
  INV_X1 U21742 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18587) );
  NOR2_X1 U21743 ( .A1(n18587), .A2(n18519), .ZN(n18522) );
  AOI21_X1 U21744 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18523), .A(n18527), .ZN(
        n18521) );
  OAI222_X1 U21745 ( .A1(n19362), .A2(n18528), .B1(n18522), .B2(n18521), .C1(
        n18525), .C2(n18520), .ZN(P3_U2731) );
  AOI21_X1 U21746 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18523), .A(n18529), .ZN(
        n18526) );
  OAI222_X1 U21747 ( .A1(n19358), .A2(n18528), .B1(n18527), .B2(n18526), .C1(
        n18525), .C2(n18524), .ZN(P3_U2732) );
  INV_X1 U21748 ( .A(n18529), .ZN(n18534) );
  OAI21_X1 U21749 ( .B1(n18590), .B2(n18531), .A(n18530), .ZN(n18533) );
  AOI222_X1 U21750 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18538), .B1(n18534), .B2(
        n18533), .C1(n18537), .C2(n18532), .ZN(n18535) );
  INV_X1 U21751 ( .A(n18535), .ZN(P3_U2733) );
  AOI22_X1 U21752 ( .A1(n18538), .A2(BUF2_REG_1__SCAN_IN), .B1(n18537), .B2(
        n18536), .ZN(n18544) );
  NOR2_X1 U21753 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18539), .ZN(n18541) );
  OAI22_X1 U21754 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n18542), .B1(n18541), .B2(
        n18540), .ZN(n18543) );
  NAND2_X1 U21755 ( .A1(n18544), .A2(n18543), .ZN(P3_U2734) );
  INV_X2 U21756 ( .A(n18559), .ZN(n19982) );
  NOR2_X1 U21757 ( .A1(n22005), .A2(n18567), .ZN(P3_U2736) );
  NAND2_X1 U21758 ( .A1(n18568), .A2(n18546), .ZN(n18564) );
  AOI22_X1 U21759 ( .A1(n19982), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18547) );
  OAI21_X1 U21760 ( .B1(n18624), .B2(n18564), .A(n18547), .ZN(P3_U2737) );
  INV_X1 U21761 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n21889) );
  INV_X1 U21762 ( .A(n18564), .ZN(n18557) );
  AOI22_X1 U21763 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18557), .B1(n19982), 
        .B2(P3_UWORD_REG_13__SCAN_IN), .ZN(n18548) );
  OAI21_X1 U21764 ( .B1(n21889), .B2(n18567), .A(n18548), .ZN(P3_U2738) );
  INV_X1 U21765 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18621) );
  AOI22_X1 U21766 ( .A1(n19982), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18549) );
  OAI21_X1 U21767 ( .B1(n18621), .B2(n18564), .A(n18549), .ZN(P3_U2739) );
  AOI22_X1 U21768 ( .A1(n19982), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18550) );
  OAI21_X1 U21769 ( .B1(n18619), .B2(n18564), .A(n18550), .ZN(P3_U2740) );
  AOI22_X1 U21770 ( .A1(P3_DATAO_REG_26__SCAN_IN), .A2(n9750), .B1(n19982), 
        .B2(P3_UWORD_REG_10__SCAN_IN), .ZN(n18551) );
  OAI21_X1 U21771 ( .B1(n10331), .B2(n18564), .A(n18551), .ZN(P3_U2741) );
  AOI22_X1 U21772 ( .A1(n19982), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18552) );
  OAI21_X1 U21773 ( .B1(n18616), .B2(n18564), .A(n18552), .ZN(P3_U2742) );
  AOI22_X1 U21774 ( .A1(n19982), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18553) );
  OAI21_X1 U21775 ( .B1(n18614), .B2(n18564), .A(n18553), .ZN(P3_U2743) );
  AOI22_X1 U21776 ( .A1(n19982), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18554) );
  OAI21_X1 U21777 ( .B1(n18612), .B2(n18564), .A(n18554), .ZN(P3_U2744) );
  INV_X1 U21778 ( .A(P3_UWORD_REG_6__SCAN_IN), .ZN(n21845) );
  AOI22_X1 U21779 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18557), .B1(n9750), .B2(
        P3_DATAO_REG_22__SCAN_IN), .ZN(n18555) );
  OAI21_X1 U21780 ( .B1(n21845), .B2(n18559), .A(n18555), .ZN(P3_U2745) );
  AOI22_X1 U21781 ( .A1(n19982), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18556) );
  OAI21_X1 U21782 ( .B1(n18608), .B2(n18564), .A(n18556), .ZN(P3_U2746) );
  INV_X1 U21783 ( .A(P3_UWORD_REG_4__SCAN_IN), .ZN(n21952) );
  AOI22_X1 U21784 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18557), .B1(n9750), .B2(
        P3_DATAO_REG_20__SCAN_IN), .ZN(n18558) );
  OAI21_X1 U21785 ( .B1(n21952), .B2(n18559), .A(n18558), .ZN(P3_U2747) );
  AOI22_X1 U21786 ( .A1(n19982), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18560) );
  OAI21_X1 U21787 ( .B1(n18605), .B2(n18564), .A(n18560), .ZN(P3_U2748) );
  INV_X1 U21788 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18603) );
  AOI22_X1 U21789 ( .A1(n19982), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18561) );
  OAI21_X1 U21790 ( .B1(n18603), .B2(n18564), .A(n18561), .ZN(P3_U2749) );
  AOI22_X1 U21791 ( .A1(n19982), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18562) );
  OAI21_X1 U21792 ( .B1(n18601), .B2(n18564), .A(n18562), .ZN(P3_U2750) );
  AOI22_X1 U21793 ( .A1(P3_UWORD_REG_0__SCAN_IN), .A2(n19982), .B1(n9750), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18563) );
  OAI21_X1 U21794 ( .B1(n18565), .B2(n18564), .A(n18563), .ZN(P3_U2751) );
  INV_X1 U21795 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n21801) );
  AOI22_X1 U21796 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n18568), .B1(n19982), 
        .B2(P3_LWORD_REG_15__SCAN_IN), .ZN(n18566) );
  OAI21_X1 U21797 ( .B1(n21801), .B2(n18567), .A(n18566), .ZN(P3_U2752) );
  AOI22_X1 U21798 ( .A1(n19982), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18569) );
  OAI21_X1 U21799 ( .B1(n18647), .B2(n18593), .A(n18569), .ZN(P3_U2753) );
  INV_X1 U21800 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18571) );
  AOI22_X1 U21801 ( .A1(n19982), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18570) );
  OAI21_X1 U21802 ( .B1(n18571), .B2(n18593), .A(n18570), .ZN(P3_U2754) );
  AOI22_X1 U21803 ( .A1(n19982), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18572) );
  OAI21_X1 U21804 ( .B1(n18573), .B2(n18593), .A(n18572), .ZN(P3_U2755) );
  INV_X1 U21805 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18575) );
  AOI22_X1 U21806 ( .A1(n19982), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18574) );
  OAI21_X1 U21807 ( .B1(n18575), .B2(n18593), .A(n18574), .ZN(P3_U2756) );
  AOI22_X1 U21808 ( .A1(n19982), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18576) );
  OAI21_X1 U21809 ( .B1(n18577), .B2(n18593), .A(n18576), .ZN(P3_U2757) );
  INV_X1 U21810 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18579) );
  AOI22_X1 U21811 ( .A1(n19982), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18578) );
  OAI21_X1 U21812 ( .B1(n18579), .B2(n18593), .A(n18578), .ZN(P3_U2758) );
  AOI22_X1 U21813 ( .A1(n19982), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18580) );
  OAI21_X1 U21814 ( .B1(n18635), .B2(n18593), .A(n18580), .ZN(P3_U2759) );
  INV_X1 U21815 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n21827) );
  AOI22_X1 U21816 ( .A1(n19982), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18581) );
  OAI21_X1 U21817 ( .B1(n21827), .B2(n18593), .A(n18581), .ZN(P3_U2760) );
  INV_X1 U21818 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18583) );
  AOI22_X1 U21819 ( .A1(n19982), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18582) );
  OAI21_X1 U21820 ( .B1(n18583), .B2(n18593), .A(n18582), .ZN(P3_U2761) );
  INV_X1 U21821 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18585) );
  AOI22_X1 U21822 ( .A1(n19982), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18584) );
  OAI21_X1 U21823 ( .B1(n18585), .B2(n18593), .A(n18584), .ZN(P3_U2762) );
  AOI22_X1 U21824 ( .A1(n19982), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18586) );
  OAI21_X1 U21825 ( .B1(n18587), .B2(n18593), .A(n18586), .ZN(P3_U2763) );
  INV_X1 U21826 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n21833) );
  AOI22_X1 U21827 ( .A1(n19982), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18588) );
  OAI21_X1 U21828 ( .B1(n21833), .B2(n18593), .A(n18588), .ZN(P3_U2764) );
  AOI22_X1 U21829 ( .A1(n19982), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18589) );
  OAI21_X1 U21830 ( .B1(n18590), .B2(n18593), .A(n18589), .ZN(P3_U2765) );
  INV_X1 U21831 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18627) );
  AOI22_X1 U21832 ( .A1(n19982), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18591) );
  OAI21_X1 U21833 ( .B1(n18627), .B2(n18593), .A(n18591), .ZN(P3_U2766) );
  AOI22_X1 U21834 ( .A1(n19982), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n9750), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18592) );
  OAI21_X1 U21835 ( .B1(n18594), .B2(n18593), .A(n18592), .ZN(P3_U2767) );
  INV_X1 U21836 ( .A(P3_UWORD_REG_0__SCAN_IN), .ZN(n21922) );
  NOR2_X2 U21837 ( .A1(n19987), .A2(n18637), .ZN(n18644) );
  NAND2_X1 U21838 ( .A1(n19987), .A2(n18597), .ZN(n19828) );
  AOI22_X1 U21839 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18644), .B1(
        P3_EAX_REG_16__SCAN_IN), .B2(n18649), .ZN(n18599) );
  OAI21_X1 U21840 ( .B1(n18610), .B2(n21922), .A(n18599), .ZN(P3_U2768) );
  AOI22_X1 U21841 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18637), .ZN(n18600) );
  OAI21_X1 U21842 ( .B1(n18601), .B2(n18646), .A(n18600), .ZN(P3_U2769) );
  AOI22_X1 U21843 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18637), .ZN(n18602) );
  OAI21_X1 U21844 ( .B1(n18603), .B2(n18646), .A(n18602), .ZN(P3_U2770) );
  AOI22_X1 U21845 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18637), .ZN(n18604) );
  OAI21_X1 U21846 ( .B1(n18605), .B2(n18646), .A(n18604), .ZN(P3_U2771) );
  AOI22_X1 U21847 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18644), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n18649), .ZN(n18606) );
  OAI21_X1 U21848 ( .B1(n18610), .B2(n21952), .A(n18606), .ZN(P3_U2772) );
  AOI22_X1 U21849 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18637), .ZN(n18607) );
  OAI21_X1 U21850 ( .B1(n18608), .B2(n18646), .A(n18607), .ZN(P3_U2773) );
  AOI22_X1 U21851 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18644), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n18649), .ZN(n18609) );
  OAI21_X1 U21852 ( .B1(n18610), .B2(n21845), .A(n18609), .ZN(P3_U2774) );
  AOI22_X1 U21853 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18637), .ZN(n18611) );
  OAI21_X1 U21854 ( .B1(n18612), .B2(n18646), .A(n18611), .ZN(P3_U2775) );
  AOI22_X1 U21855 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18637), .ZN(n18613) );
  OAI21_X1 U21856 ( .B1(n18614), .B2(n18646), .A(n18613), .ZN(P3_U2776) );
  AOI22_X1 U21857 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18637), .ZN(n18615) );
  OAI21_X1 U21858 ( .B1(n18616), .B2(n18646), .A(n18615), .ZN(P3_U2777) );
  AOI22_X1 U21859 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18637), .ZN(n18617) );
  OAI21_X1 U21860 ( .B1(n10331), .B2(n18646), .A(n18617), .ZN(P3_U2778) );
  AOI22_X1 U21861 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18637), .ZN(n18618) );
  OAI21_X1 U21862 ( .B1(n18619), .B2(n18646), .A(n18618), .ZN(P3_U2779) );
  AOI22_X1 U21863 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18637), .ZN(n18620) );
  OAI21_X1 U21864 ( .B1(n18621), .B2(n18646), .A(n18620), .ZN(P3_U2780) );
  AOI22_X1 U21865 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18649), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18637), .ZN(n18622) );
  OAI21_X1 U21866 ( .B1(n13833), .B2(n18651), .A(n18622), .ZN(P3_U2781) );
  AOI22_X1 U21867 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18644), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18648), .ZN(n18623) );
  OAI21_X1 U21868 ( .B1(n18624), .B2(n18646), .A(n18623), .ZN(P3_U2782) );
  AOI22_X1 U21869 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18648), .ZN(n18625) );
  OAI21_X1 U21870 ( .B1(n19345), .B2(n18651), .A(n18625), .ZN(P3_U2783) );
  AOI22_X1 U21871 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18644), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18648), .ZN(n18626) );
  OAI21_X1 U21872 ( .B1(n18627), .B2(n18646), .A(n18626), .ZN(P3_U2784) );
  AOI22_X1 U21873 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18648), .ZN(n18628) );
  OAI21_X1 U21874 ( .B1(n19354), .B2(n18651), .A(n18628), .ZN(P3_U2785) );
  AOI22_X1 U21875 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18648), .ZN(n18629) );
  OAI21_X1 U21876 ( .B1(n19358), .B2(n18651), .A(n18629), .ZN(P3_U2786) );
  AOI22_X1 U21877 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18648), .ZN(n18630) );
  OAI21_X1 U21878 ( .B1(n19362), .B2(n18651), .A(n18630), .ZN(P3_U2787) );
  AOI22_X1 U21879 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18637), .ZN(n18631) );
  OAI21_X1 U21880 ( .B1(n13829), .B2(n18651), .A(n18631), .ZN(P3_U2788) );
  AOI22_X1 U21881 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18637), .ZN(n18632) );
  OAI21_X1 U21882 ( .B1(n13839), .B2(n18651), .A(n18632), .ZN(P3_U2789) );
  AOI22_X1 U21883 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18637), .ZN(n18633) );
  OAI21_X1 U21884 ( .B1(n13920), .B2(n18651), .A(n18633), .ZN(P3_U2790) );
  AOI22_X1 U21885 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18644), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18637), .ZN(n18634) );
  OAI21_X1 U21886 ( .B1(n18635), .B2(n18646), .A(n18634), .ZN(P3_U2791) );
  AOI22_X1 U21887 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18637), .ZN(n18636) );
  OAI21_X1 U21888 ( .B1(n13821), .B2(n18651), .A(n18636), .ZN(P3_U2792) );
  AOI22_X1 U21889 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18637), .ZN(n18638) );
  OAI21_X1 U21890 ( .B1(n18639), .B2(n18651), .A(n18638), .ZN(P3_U2793) );
  AOI22_X1 U21891 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18648), .ZN(n18640) );
  OAI21_X1 U21892 ( .B1(n13817), .B2(n18651), .A(n18640), .ZN(P3_U2794) );
  AOI22_X1 U21893 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18648), .ZN(n18641) );
  OAI21_X1 U21894 ( .B1(n18642), .B2(n18651), .A(n18641), .ZN(P3_U2795) );
  AOI22_X1 U21895 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18648), .ZN(n18643) );
  OAI21_X1 U21896 ( .B1(n13833), .B2(n18651), .A(n18643), .ZN(P3_U2796) );
  AOI22_X1 U21897 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18644), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18648), .ZN(n18645) );
  OAI21_X1 U21898 ( .B1(n18647), .B2(n18646), .A(n18645), .ZN(P3_U2797) );
  AOI22_X1 U21899 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n18649), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18648), .ZN(n18650) );
  OAI21_X1 U21900 ( .B1(n13855), .B2(n18651), .A(n18650), .ZN(P3_U2798) );
  NOR3_X1 U21901 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18846), .A3(
        n10842), .ZN(n18653) );
  AOI211_X1 U21902 ( .C1(n18865), .C2(n18654), .A(n18653), .B(n18652), .ZN(
        n18669) );
  NOR2_X1 U21903 ( .A1(n19015), .A2(n18819), .ZN(n18729) );
  NOR2_X1 U21904 ( .A1(n18999), .A2(n18922), .ZN(n18765) );
  NOR2_X1 U21905 ( .A1(n18765), .A2(n18655), .ZN(n18657) );
  AOI22_X1 U21906 ( .A1(n18999), .A2(n19020), .B1(n18922), .B2(n19019), .ZN(
        n18689) );
  NAND2_X1 U21907 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18689), .ZN(
        n18677) );
  AOI22_X1 U21908 ( .A1(n18658), .A2(n18729), .B1(n18657), .B2(n18677), .ZN(
        n18668) );
  OAI211_X1 U21909 ( .C1(n18661), .C2(n18660), .A(n18921), .B(n18659), .ZN(
        n18667) );
  NOR3_X1 U21910 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18846), .A3(
        n18662), .ZN(n18675) );
  OAI21_X1 U21911 ( .B1(n18663), .B2(n18981), .A(n19009), .ZN(n18664) );
  AOI21_X1 U21912 ( .B1(n18732), .B2(n18665), .A(n18664), .ZN(n18681) );
  OAI21_X1 U21913 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18692), .A(
        n18681), .ZN(n18676) );
  OAI21_X1 U21914 ( .B1(n18675), .B2(n18676), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18666) );
  NAND4_X1 U21915 ( .A1(n18669), .A2(n18668), .A3(n18667), .A4(n18666), .ZN(
        P3_U2802) );
  NAND2_X1 U21916 ( .A1(n18671), .A2(n18670), .ZN(n18672) );
  XNOR2_X1 U21917 ( .A(n18672), .B(n18920), .ZN(n19028) );
  INV_X1 U21918 ( .A(n18921), .ZN(n18840) );
  OAI22_X1 U21919 ( .A1(n19328), .A2(n19913), .B1(n18851), .B2(n18673), .ZN(
        n18674) );
  AOI211_X1 U21920 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n18676), .A(
        n18675), .B(n18674), .ZN(n18680) );
  NOR2_X1 U21921 ( .A1(n19024), .A2(n18819), .ZN(n18678) );
  OAI21_X1 U21922 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18678), .A(
        n18677), .ZN(n18679) );
  OAI211_X1 U21923 ( .C1(n19028), .C2(n18840), .A(n18680), .B(n18679), .ZN(
        P3_U2803) );
  NAND2_X2 U21924 ( .A1(n18851), .A2(n18692), .ZN(n19002) );
  AOI221_X1 U21925 ( .B1(n18682), .B2(n22029), .C1(n19369), .C2(n22029), .A(
        n18681), .ZN(n18683) );
  NOR2_X1 U21926 ( .A1(n19328), .A2(n19911), .ZN(n19033) );
  AOI211_X1 U21927 ( .C1(n18684), .C2(n19002), .A(n18683), .B(n19033), .ZN(
        n18688) );
  XNOR2_X1 U21928 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n18685), .ZN(
        n19032) );
  NOR2_X1 U21929 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18686), .ZN(
        n19030) );
  AOI22_X1 U21930 ( .A1(n18921), .A2(n19032), .B1(n18729), .B2(n19030), .ZN(
        n18687) );
  OAI211_X1 U21931 ( .C1(n18689), .C2(n12851), .A(n18688), .B(n18687), .ZN(
        P3_U2804) );
  INV_X1 U21932 ( .A(n18922), .ZN(n18878) );
  NAND3_X1 U21933 ( .A1(n19141), .A2(n18714), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18690) );
  XNOR2_X1 U21934 ( .A(n18690), .B(n19042), .ZN(n19039) );
  NAND2_X1 U21935 ( .A1(n18691), .A2(n18772), .ZN(n18711) );
  AOI221_X1 U21936 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C1(n18710), .C2(n18695), .A(
        n18711), .ZN(n18697) );
  INV_X1 U21937 ( .A(n18692), .ZN(n18760) );
  OR2_X1 U21938 ( .A1(n19369), .A2(n18691), .ZN(n18726) );
  OAI211_X1 U21939 ( .C1(n18693), .C2(n19848), .A(n19009), .B(n18726), .ZN(
        n18723) );
  AOI21_X1 U21940 ( .B1(n18760), .B2(n18694), .A(n18723), .ZN(n18709) );
  OAI22_X1 U21941 ( .A1(n18709), .A2(n18695), .B1(n19328), .B2(n19909), .ZN(
        n18696) );
  AOI211_X1 U21942 ( .C1(n18698), .C2(n18865), .A(n18697), .B(n18696), .ZN(
        n18706) );
  NAND2_X1 U21943 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18714), .ZN(
        n19037) );
  NOR2_X1 U21944 ( .A1(n19149), .A2(n19037), .ZN(n18699) );
  XNOR2_X1 U21945 ( .A(n18699), .B(n19042), .ZN(n19045) );
  INV_X1 U21946 ( .A(n18707), .ZN(n18703) );
  INV_X1 U21947 ( .A(n18701), .ZN(n18702) );
  AOI21_X1 U21948 ( .B1(n18703), .B2(n9755), .A(n18702), .ZN(n18704) );
  XNOR2_X1 U21949 ( .A(n18704), .B(n19042), .ZN(n19044) );
  AOI22_X1 U21950 ( .A1(n18999), .A2(n19045), .B1(n18921), .B2(n19044), .ZN(
        n18705) );
  OAI211_X1 U21951 ( .C1(n18878), .C2(n19039), .A(n18706), .B(n18705), .ZN(
        P3_U2805) );
  AOI21_X1 U21952 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18708), .A(
        n18707), .ZN(n19061) );
  NAND2_X1 U21953 ( .A1(n19317), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n19059) );
  OAI221_X1 U21954 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18711), .C1(
        n18710), .C2(n18709), .A(n19059), .ZN(n18712) );
  AOI21_X1 U21955 ( .B1(n18865), .B2(n18713), .A(n18712), .ZN(n18717) );
  INV_X1 U21956 ( .A(n19141), .ZN(n19072) );
  INV_X1 U21957 ( .A(n18714), .ZN(n18715) );
  NOR2_X1 U21958 ( .A1(n19072), .A2(n18715), .ZN(n19050) );
  NOR2_X1 U21959 ( .A1(n19149), .A2(n18715), .ZN(n19049) );
  OAI22_X1 U21960 ( .A1(n19050), .A2(n18878), .B1(n19049), .B2(n19013), .ZN(
        n18728) );
  NOR2_X1 U21961 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n19014), .ZN(
        n19057) );
  AOI22_X1 U21962 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18728), .B1(
        n18729), .B2(n19057), .ZN(n18716) );
  OAI211_X1 U21963 ( .C1(n19061), .C2(n18840), .A(n18717), .B(n18716), .ZN(
        P3_U2806) );
  AOI22_X1 U21964 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n9755), .B1(
        n18719), .B2(n18740), .ZN(n18720) );
  NAND2_X1 U21965 ( .A1(n18766), .A2(n18720), .ZN(n18721) );
  XNOR2_X1 U21966 ( .A(n18721), .B(n19014), .ZN(n19066) );
  AOI22_X1 U21967 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18723), .B1(
        n18722), .B2(n19002), .ZN(n18724) );
  NAND2_X1 U21968 ( .A1(n19317), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n19065) );
  OAI211_X1 U21969 ( .C1(n18726), .C2(n18725), .A(n18724), .B(n19065), .ZN(
        n18727) );
  AOI221_X1 U21970 ( .B1(n18729), .B2(n19014), .C1(n18728), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n18727), .ZN(n18730) );
  OAI21_X1 U21971 ( .B1(n18840), .B2(n19066), .A(n18730), .ZN(P3_U2807) );
  NAND2_X1 U21972 ( .A1(n18734), .A2(n18772), .ZN(n18748) );
  AOI221_X1 U21973 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n18747), .C2(n18735), .A(
        n18748), .ZN(n18737) );
  NAND2_X1 U21974 ( .A1(n18732), .A2(n18731), .ZN(n18733) );
  OAI211_X1 U21975 ( .C1(n18734), .C2(n18981), .A(n19009), .B(n18733), .ZN(
        n18764) );
  AOI21_X1 U21976 ( .B1(n18760), .B2(n18759), .A(n18764), .ZN(n18746) );
  OAI22_X1 U21977 ( .A1(n18746), .A2(n18735), .B1(n19328), .B2(n19902), .ZN(
        n18736) );
  AOI211_X1 U21978 ( .C1(n18738), .C2(n18865), .A(n18737), .B(n18736), .ZN(
        n18745) );
  AOI22_X1 U21979 ( .A1(n18999), .A2(n19149), .B1(n18922), .B2(n19072), .ZN(
        n18818) );
  OAI21_X1 U21980 ( .B1(n19077), .B2(n18765), .A(n18818), .ZN(n18756) );
  INV_X1 U21981 ( .A(n18766), .ZN(n18739) );
  AOI221_X1 U21982 ( .B1(n18741), .B2(n18740), .C1(n18751), .C2(n18740), .A(
        n18739), .ZN(n18742) );
  XNOR2_X1 U21983 ( .A(n18742), .B(n19084), .ZN(n19067) );
  AOI22_X1 U21984 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18756), .B1(
        n18921), .B2(n19067), .ZN(n18744) );
  NAND3_X1 U21985 ( .A1(n19077), .A2(n18794), .A3(n19084), .ZN(n18743) );
  NAND3_X1 U21986 ( .A1(n18745), .A2(n18744), .A3(n18743), .ZN(P3_U2808) );
  NAND2_X1 U21987 ( .A1(n18754), .A2(n21959), .ZN(n19097) );
  INV_X1 U21988 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21874) );
  NOR2_X1 U21989 ( .A1(n19113), .A2(n21874), .ZN(n19087) );
  NAND2_X1 U21990 ( .A1(n18794), .A2(n19087), .ZN(n18783) );
  NAND2_X1 U21991 ( .A1(n19317), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n19095) );
  OAI221_X1 U21992 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18748), .C1(
        n18747), .C2(n18746), .A(n19095), .ZN(n18749) );
  AOI21_X1 U21993 ( .B1(n18865), .B2(n18750), .A(n18749), .ZN(n18758) );
  NOR3_X1 U21994 ( .A1(n21874), .A2(n9755), .A3(n18751), .ZN(n18778) );
  AOI22_X1 U21995 ( .A1(n18754), .A2(n18778), .B1(n18752), .B2(n18753), .ZN(
        n18755) );
  XNOR2_X1 U21996 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18755), .ZN(
        n19094) );
  AOI22_X1 U21997 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18756), .B1(
        n18921), .B2(n19094), .ZN(n18757) );
  OAI211_X1 U21998 ( .C1(n19097), .C2(n18783), .A(n18758), .B(n18757), .ZN(
        P3_U2809) );
  NAND2_X1 U21999 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19070), .ZN(
        n19105) );
  OAI21_X1 U22000 ( .B1(n9949), .B2(n19369), .A(n18759), .ZN(n18763) );
  NAND2_X1 U22001 ( .A1(n19317), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n19103) );
  OAI221_X1 U22002 ( .B1(n18761), .B2(n18851), .C1(n18761), .C2(n18692), .A(
        n19103), .ZN(n18762) );
  AOI21_X1 U22003 ( .B1(n18764), .B2(n18763), .A(n18762), .ZN(n18769) );
  INV_X1 U22004 ( .A(n19087), .ZN(n19085) );
  NOR2_X1 U22005 ( .A1(n21877), .A2(n19085), .ZN(n19100) );
  OAI21_X1 U22006 ( .B1(n18765), .B2(n19100), .A(n18818), .ZN(n18780) );
  OAI221_X1 U22007 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18790), 
        .C1(n21877), .C2(n18778), .A(n18766), .ZN(n18767) );
  XNOR2_X1 U22008 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18767), .ZN(
        n19102) );
  AOI22_X1 U22009 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18780), .B1(
        n18921), .B2(n19102), .ZN(n18768) );
  OAI211_X1 U22010 ( .C1(n18783), .C2(n19105), .A(n18769), .B(n18768), .ZN(
        P3_U2810) );
  OAI21_X1 U22011 ( .B1(n18980), .B2(n18770), .A(n18901), .ZN(n18795) );
  OAI21_X1 U22012 ( .B1(n18771), .B2(n19848), .A(n18795), .ZN(n18789) );
  NOR2_X1 U22013 ( .A1(n19328), .A2(n19896), .ZN(n18777) );
  NAND2_X1 U22014 ( .A1(n10844), .A2(n18772), .ZN(n18786) );
  OAI21_X1 U22015 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18773), .ZN(n18774) );
  OAI22_X1 U22016 ( .A1(n18851), .A2(n18775), .B1(n18786), .B2(n18774), .ZN(
        n18776) );
  AOI211_X1 U22017 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n18789), .A(
        n18777), .B(n18776), .ZN(n18782) );
  AOI21_X1 U22018 ( .B1(n18790), .B2(n18752), .A(n18778), .ZN(n18779) );
  XNOR2_X1 U22019 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n18779), .ZN(
        n19106) );
  AOI22_X1 U22020 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18780), .B1(
        n18921), .B2(n19106), .ZN(n18781) );
  OAI211_X1 U22021 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18783), .A(
        n18782), .B(n18781), .ZN(P3_U2811) );
  INV_X1 U22022 ( .A(n18818), .ZN(n18784) );
  AOI21_X1 U22023 ( .B1(n18794), .B2(n19113), .A(n18784), .ZN(n18804) );
  NOR2_X1 U22024 ( .A1(n19328), .A2(n19894), .ZN(n18788) );
  OAI22_X1 U22025 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18786), .B1(
        n18851), .B2(n18785), .ZN(n18787) );
  AOI211_X1 U22026 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18789), .A(
        n18788), .B(n18787), .ZN(n18793) );
  AOI21_X1 U22027 ( .B1(n18920), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n18790), .ZN(n18791) );
  XOR2_X1 U22028 ( .A(n18791), .B(n18752), .Z(n19122) );
  NOR2_X1 U22029 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n19113), .ZN(
        n19121) );
  AOI22_X1 U22030 ( .A1(n18921), .A2(n19122), .B1(n18794), .B2(n19121), .ZN(
        n18792) );
  OAI211_X1 U22031 ( .C1(n18804), .C2(n21874), .A(n18793), .B(n18792), .ZN(
        P3_U2812) );
  AOI21_X1 U22032 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18794), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18803) );
  AOI221_X1 U22033 ( .B1(n17872), .B2(n18796), .C1(n19369), .C2(n18796), .A(
        n18795), .ZN(n18797) );
  AOI21_X1 U22034 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n19317), .A(n18797), 
        .ZN(n18802) );
  OAI21_X1 U22035 ( .B1(n18799), .B2(n19127), .A(n18798), .ZN(n19125) );
  AOI22_X1 U22036 ( .A1(n18921), .A2(n19125), .B1(n18800), .B2(n19002), .ZN(
        n18801) );
  OAI211_X1 U22037 ( .C1(n18804), .C2(n18803), .A(n18802), .B(n18801), .ZN(
        P3_U2813) );
  AOI21_X1 U22038 ( .B1(n18920), .B2(n18806), .A(n18805), .ZN(n18807) );
  XNOR2_X1 U22039 ( .A(n18807), .B(n19136), .ZN(n19138) );
  INV_X1 U22040 ( .A(n18981), .ZN(n18912) );
  INV_X1 U22041 ( .A(n18808), .ZN(n18809) );
  AOI21_X1 U22042 ( .B1(n18912), .B2(n18809), .A(n18980), .ZN(n18845) );
  OAI21_X1 U22043 ( .B1(n18810), .B2(n19848), .A(n18845), .ZN(n18822) );
  AOI22_X1 U22044 ( .A1(n19317), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18822), .ZN(n18814) );
  NOR3_X1 U22045 ( .A1(n18846), .A2(n18811), .A3(n17935), .ZN(n18824) );
  OAI211_X1 U22046 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18824), .B(n18812), .ZN(n18813) );
  OAI211_X1 U22047 ( .C1(n18851), .C2(n18815), .A(n18814), .B(n18813), .ZN(
        n18816) );
  AOI21_X1 U22048 ( .B1(n18921), .B2(n19138), .A(n18816), .ZN(n18817) );
  OAI221_X1 U22049 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18819), 
        .C1(n19136), .C2(n18818), .A(n18817), .ZN(P3_U2814) );
  NOR2_X1 U22050 ( .A1(n22014), .A2(n19163), .ZN(n18827) );
  NAND2_X1 U22051 ( .A1(n19183), .A2(n18877), .ZN(n19185) );
  INV_X1 U22052 ( .A(n19185), .ZN(n18855) );
  NOR2_X1 U22053 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18836), .ZN(
        n19148) );
  NAND2_X1 U22054 ( .A1(n18999), .A2(n19149), .ZN(n18833) );
  OAI22_X1 U22055 ( .A1(n19328), .A2(n19889), .B1(n18851), .B2(n18820), .ZN(
        n18821) );
  AOI221_X1 U22056 ( .B1(n18824), .B2(n18823), .C1(n18822), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18821), .ZN(n18832) );
  NOR2_X1 U22057 ( .A1(n19181), .A2(n18825), .ZN(n18857) );
  NAND2_X1 U22058 ( .A1(n18826), .A2(n9755), .ZN(n18896) );
  NOR3_X1 U22059 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18891), .A3(
        n18896), .ZN(n18866) );
  AOI22_X1 U22060 ( .A1(n18857), .A2(n18827), .B1(n18866), .B2(n22014), .ZN(
        n18828) );
  AOI221_X1 U22061 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n19174), 
        .C1(n9755), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n18828), .ZN(
        n18829) );
  XNOR2_X1 U22062 ( .A(n18829), .B(n19143), .ZN(n19151) );
  NOR2_X1 U22063 ( .A1(n19141), .A2(n18878), .ZN(n18830) );
  NAND2_X1 U22064 ( .A1(n19143), .A2(n18839), .ZN(n19146) );
  AOI22_X1 U22065 ( .A1(n18921), .A2(n19151), .B1(n18830), .B2(n19146), .ZN(
        n18831) );
  OAI211_X1 U22066 ( .C1(n19148), .C2(n18833), .A(n18832), .B(n18831), .ZN(
        P3_U2815) );
  NAND2_X1 U22067 ( .A1(n10852), .A2(n19659), .ZN(n18914) );
  NOR2_X1 U22068 ( .A1(n10577), .A2(n18914), .ZN(n18874) );
  AOI21_X1 U22069 ( .B1(n18847), .B2(n18874), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18844) );
  AOI22_X1 U22070 ( .A1(n19317), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n18835), 
        .B2(n19002), .ZN(n18843) );
  AOI221_X1 U22071 ( .B1(n22014), .B2(n19163), .C1(n19185), .C2(n19163), .A(
        n18836), .ZN(n19167) );
  NAND2_X1 U22072 ( .A1(n18866), .A2(n22014), .ZN(n18837) );
  NAND2_X1 U22073 ( .A1(n19183), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n19161) );
  NAND2_X1 U22074 ( .A1(n18920), .A2(n19177), .ZN(n18897) );
  OAI22_X1 U22075 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18837), .B1(
        n19161), .B2(n18897), .ZN(n18838) );
  XNOR2_X1 U22076 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18838), .ZN(
        n19172) );
  AND2_X1 U22077 ( .A1(n19183), .A2(n19177), .ZN(n18854) );
  OAI221_X1 U22078 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18854), .A(n18839), .ZN(
        n19166) );
  OAI22_X1 U22079 ( .A1(n19172), .A2(n18840), .B1(n18878), .B2(n19166), .ZN(
        n18841) );
  AOI21_X1 U22080 ( .B1(n18999), .B2(n19167), .A(n18841), .ZN(n18842) );
  OAI211_X1 U22081 ( .C1(n18845), .C2(n18844), .A(n18843), .B(n18842), .ZN(
        P3_U2816) );
  NAND2_X1 U22082 ( .A1(n19183), .A2(n22014), .ZN(n19190) );
  OAI21_X1 U22083 ( .B1(n18848), .B2(n19848), .A(n19009), .ZN(n18849) );
  AOI21_X1 U22084 ( .B1(n18912), .B2(n17935), .A(n18849), .ZN(n18860) );
  OAI22_X1 U22085 ( .A1(n18860), .A2(n18852), .B1(n18851), .B2(n18850), .ZN(
        n18853) );
  OAI22_X1 U22086 ( .A1(n18855), .A2(n19013), .B1(n18854), .B2(n18878), .ZN(
        n18868) );
  NOR2_X1 U22087 ( .A1(n19174), .A2(n9755), .ZN(n18856) );
  OAI22_X1 U22088 ( .A1(n18857), .A2(n19174), .B1(n18866), .B2(n18856), .ZN(
        n18858) );
  XNOR2_X1 U22089 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18858), .ZN(
        n19173) );
  AOI22_X1 U22090 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18868), .B1(
        n18921), .B2(n19173), .ZN(n18859) );
  NOR3_X1 U22091 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18909), .A3(
        n19181), .ZN(n18863) );
  NAND2_X1 U22092 ( .A1(n19317), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n19198) );
  OAI221_X1 U22093 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9790), .C1(
        n18861), .C2(n18860), .A(n19198), .ZN(n18862) );
  AOI211_X1 U22094 ( .C1(n18865), .C2(n18864), .A(n18863), .B(n18862), .ZN(
        n18870) );
  INV_X1 U22095 ( .A(n19181), .ZN(n19196) );
  INV_X1 U22096 ( .A(n18897), .ZN(n18888) );
  AOI21_X1 U22097 ( .B1(n19196), .B2(n18888), .A(n18866), .ZN(n18867) );
  XNOR2_X1 U22098 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18867), .ZN(
        n19197) );
  AOI22_X1 U22099 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18868), .B1(
        n18921), .B2(n19197), .ZN(n18869) );
  NAND2_X1 U22100 ( .A1(n18870), .A2(n18869), .ZN(P3_U2818) );
  INV_X1 U22101 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n19175) );
  NAND2_X1 U22102 ( .A1(n19207), .A2(n19175), .ZN(n19212) );
  NAND2_X1 U22103 ( .A1(n19207), .A2(n18888), .ZN(n18886) );
  OAI21_X1 U22104 ( .B1(n18891), .B2(n18896), .A(n18886), .ZN(n18871) );
  XNOR2_X1 U22105 ( .A(n18871), .B(n19175), .ZN(n19201) );
  NOR2_X1 U22106 ( .A1(n19328), .A2(n19882), .ZN(n18876) );
  NOR2_X1 U22107 ( .A1(n18913), .A2(n18914), .ZN(n18900) );
  NAND2_X1 U22108 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18900), .ZN(
        n18899) );
  NOR2_X1 U22109 ( .A1(n21923), .A2(n18899), .ZN(n18882) );
  AOI21_X1 U22110 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18901), .A(
        n18882), .ZN(n18873) );
  OAI22_X1 U22111 ( .A1(n18874), .A2(n18873), .B1(n18994), .B2(n18872), .ZN(
        n18875) );
  AOI211_X1 U22112 ( .C1(n18921), .C2(n19201), .A(n18876), .B(n18875), .ZN(
        n18880) );
  NOR2_X1 U22113 ( .A1(n19207), .A2(n18909), .ZN(n18892) );
  OAI22_X1 U22114 ( .A1(n19177), .A2(n18878), .B1(n19013), .B2(n18877), .ZN(
        n18881) );
  OAI21_X1 U22115 ( .B1(n18892), .B2(n18881), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18879) );
  OAI211_X1 U22116 ( .C1(n18909), .C2(n19212), .A(n18880), .B(n18879), .ZN(
        P3_U2819) );
  INV_X1 U22117 ( .A(n18881), .ZN(n18908) );
  INV_X1 U22118 ( .A(n18901), .ZN(n19007) );
  AOI211_X1 U22119 ( .C1(n18899), .C2(n21923), .A(n19007), .B(n18882), .ZN(
        n18884) );
  NOR2_X1 U22120 ( .A1(n19328), .A2(n19880), .ZN(n18883) );
  AOI211_X1 U22121 ( .C1(n18885), .C2(n19002), .A(n18884), .B(n18883), .ZN(
        n18894) );
  INV_X1 U22122 ( .A(n18891), .ZN(n18890) );
  NAND2_X1 U22123 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18895), .ZN(
        n19219) );
  NAND4_X1 U22124 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18826), .A3(
        n19227), .A4(n9755), .ZN(n18887) );
  OAI211_X1 U22125 ( .C1(n18888), .C2(n19219), .A(n18887), .B(n18886), .ZN(
        n18889) );
  AOI21_X1 U22126 ( .B1(n18890), .B2(n18896), .A(n18889), .ZN(n19213) );
  AOI22_X1 U22127 ( .A1(n18921), .A2(n19213), .B1(n18892), .B2(n18891), .ZN(
        n18893) );
  OAI211_X1 U22128 ( .C1(n18908), .C2(n18895), .A(n18894), .B(n18893), .ZN(
        P3_U2820) );
  NAND2_X1 U22129 ( .A1(n18897), .A2(n18896), .ZN(n18898) );
  XNOR2_X1 U22130 ( .A(n18898), .B(n19227), .ZN(n19224) );
  NOR2_X1 U22131 ( .A1(n19328), .A2(n19878), .ZN(n18906) );
  INV_X1 U22132 ( .A(n18899), .ZN(n18904) );
  AOI21_X1 U22133 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18901), .A(
        n18900), .ZN(n18903) );
  OAI22_X1 U22134 ( .A1(n18904), .A2(n18903), .B1(n18994), .B2(n18902), .ZN(
        n18905) );
  AOI211_X1 U22135 ( .C1(n18921), .C2(n19224), .A(n18906), .B(n18905), .ZN(
        n18907) );
  OAI221_X1 U22136 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18909), .C1(
        n19227), .C2(n18908), .A(n18907), .ZN(P3_U2821) );
  OAI21_X1 U22137 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18911), .A(
        n18910), .ZN(n19243) );
  AOI21_X1 U22138 ( .B1(n18912), .B2(n17942), .A(n18980), .ZN(n18931) );
  NAND2_X1 U22139 ( .A1(n19659), .A2(n18930), .ZN(n18929) );
  AOI21_X1 U22140 ( .B1(n18931), .B2(n18929), .A(n18913), .ZN(n18917) );
  OAI22_X1 U22141 ( .A1(n18994), .A2(n18915), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18914), .ZN(n18916) );
  AOI211_X1 U22142 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n19317), .A(n18917), .B(
        n18916), .ZN(n18924) );
  OAI21_X1 U22143 ( .B1(n18920), .B2(n18918), .A(n18919), .ZN(n19238) );
  AOI22_X1 U22144 ( .A1(n18922), .A2(n18918), .B1(n18921), .B2(n19238), .ZN(
        n18923) );
  OAI211_X1 U22145 ( .C1(n19013), .C2(n19243), .A(n18924), .B(n18923), .ZN(
        P3_U2822) );
  OAI21_X1 U22146 ( .B1(n18927), .B2(n18926), .A(n18925), .ZN(n18928) );
  XNOR2_X1 U22147 ( .A(n18928), .B(n19251), .ZN(n19246) );
  OAI22_X1 U22148 ( .A1(n18931), .A2(n18930), .B1(n17942), .B2(n18929), .ZN(
        n18932) );
  AOI21_X1 U22149 ( .B1(n19317), .B2(P3_REIP_REG_7__SCAN_IN), .A(n18932), .ZN(
        n18937) );
  AOI21_X1 U22150 ( .B1(n19251), .B2(n18934), .A(n18933), .ZN(n19245) );
  AOI22_X1 U22151 ( .A1(n19003), .A2(n19245), .B1(n18935), .B2(n19002), .ZN(
        n18936) );
  OAI211_X1 U22152 ( .C1(n19013), .C2(n19246), .A(n18937), .B(n18936), .ZN(
        P3_U2823) );
  NAND2_X1 U22153 ( .A1(n18941), .A2(n19659), .ZN(n18948) );
  AOI21_X1 U22154 ( .B1(n18940), .B2(n18939), .A(n18938), .ZN(n19258) );
  AOI22_X1 U22155 ( .A1(n19003), .A2(n19258), .B1(n19317), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n18947) );
  AOI21_X1 U22156 ( .B1(n18941), .B2(n19659), .A(n19007), .ZN(n18960) );
  OAI21_X1 U22157 ( .B1(n18943), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n18942), .ZN(n19260) );
  OAI22_X1 U22158 ( .A1(n18994), .A2(n18944), .B1(n19013), .B2(n19260), .ZN(
        n18945) );
  AOI21_X1 U22159 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18960), .A(
        n18945), .ZN(n18946) );
  OAI211_X1 U22160 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18948), .A(
        n18947), .B(n18946), .ZN(P3_U2824) );
  OAI21_X1 U22161 ( .B1(n18951), .B2(n18950), .A(n18949), .ZN(n19268) );
  OAI21_X1 U22162 ( .B1(n18954), .B2(n18953), .A(n18952), .ZN(n18955) );
  XNOR2_X1 U22163 ( .A(n18955), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19266) );
  AOI22_X1 U22164 ( .A1(n19003), .A2(n19266), .B1(n19317), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18962) );
  OAI21_X1 U22165 ( .B1(n18980), .B2(n18957), .A(n18956), .ZN(n18959) );
  AOI22_X1 U22166 ( .A1(n18960), .A2(n18959), .B1(n18958), .B2(n19002), .ZN(
        n18961) );
  OAI211_X1 U22167 ( .C1(n19013), .C2(n19268), .A(n18962), .B(n18961), .ZN(
        P3_U2825) );
  OAI21_X1 U22168 ( .B1(n18965), .B2(n18964), .A(n18963), .ZN(n19283) );
  OAI22_X1 U22169 ( .A1(n19013), .A2(n19283), .B1(n19369), .B2(n18966), .ZN(
        n18967) );
  AOI21_X1 U22170 ( .B1(n19317), .B2(P3_REIP_REG_4__SCAN_IN), .A(n18967), .ZN(
        n18972) );
  AOI21_X1 U22171 ( .B1(n18970), .B2(n18969), .A(n18968), .ZN(n19281) );
  OAI21_X1 U22172 ( .B1(n18028), .B2(n18981), .A(n19009), .ZN(n18978) );
  AOI22_X1 U22173 ( .A1(n19003), .A2(n19281), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18978), .ZN(n18971) );
  OAI211_X1 U22174 ( .C1(n18994), .C2(n18973), .A(n18972), .B(n18971), .ZN(
        P3_U2826) );
  OAI21_X1 U22175 ( .B1(n18976), .B2(n18975), .A(n18974), .ZN(n18977) );
  XOR2_X1 U22176 ( .A(n18977), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n19296) );
  INV_X1 U22177 ( .A(n19296), .ZN(n18979) );
  AOI22_X1 U22178 ( .A1(n19003), .A2(n18979), .B1(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18978), .ZN(n18986) );
  NOR2_X1 U22179 ( .A1(n18980), .A2(n18060), .ZN(n18997) );
  NOR2_X1 U22180 ( .A1(n18028), .A2(n18981), .ZN(n18983) );
  AOI22_X1 U22181 ( .A1(n18997), .A2(n18983), .B1(n18982), .B2(n19002), .ZN(
        n18985) );
  NAND2_X1 U22182 ( .A1(n19317), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19294) );
  OAI211_X1 U22183 ( .C1(n19286), .C2(n19285), .A(n18999), .B(n19284), .ZN(
        n18984) );
  NAND4_X1 U22184 ( .A1(n18986), .A2(n18985), .A3(n19294), .A4(n18984), .ZN(
        P3_U2827) );
  AOI21_X1 U22185 ( .B1(n18989), .B2(n18988), .A(n18987), .ZN(n19311) );
  NOR2_X1 U22186 ( .A1(n19328), .A2(n19865), .ZN(n19312) );
  OAI21_X1 U22187 ( .B1(n18992), .B2(n18991), .A(n18990), .ZN(n19308) );
  OAI22_X1 U22188 ( .A1(n18994), .A2(n18993), .B1(n19013), .B2(n19308), .ZN(
        n18995) );
  AOI211_X1 U22189 ( .C1(n19003), .C2(n19311), .A(n19312), .B(n18995), .ZN(
        n18996) );
  OAI221_X1 U22190 ( .B1(n18997), .B2(n18060), .C1(n18997), .C2(n19369), .A(
        n18996), .ZN(P3_U2828) );
  NOR2_X1 U22191 ( .A1(n9733), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18998) );
  XNOR2_X1 U22192 ( .A(n18998), .B(n19001), .ZN(n19319) );
  AOI22_X1 U22193 ( .A1(n18999), .A2(n19319), .B1(n19317), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n19005) );
  AOI21_X1 U22194 ( .B1(n19001), .B2(n19008), .A(n19000), .ZN(n19316) );
  AOI22_X1 U22195 ( .A1(n19003), .A2(n19316), .B1(n19006), .B2(n19002), .ZN(
        n19004) );
  OAI211_X1 U22196 ( .C1(n19007), .C2(n19006), .A(n19005), .B(n19004), .ZN(
        P3_U2829) );
  OAI21_X1 U22197 ( .B1(n9733), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19008), .ZN(n19332) );
  INV_X1 U22198 ( .A(n19332), .ZN(n19330) );
  NAND3_X1 U22199 ( .A1(n19946), .A2(n19009), .A3(n19848), .ZN(n19010) );
  AOI22_X1 U22200 ( .A1(n19317), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19010), .ZN(n19011) );
  OAI221_X1 U22201 ( .B1(n19330), .B2(n19013), .C1(n19332), .C2(n19012), .A(
        n19011), .ZN(P3_U2830) );
  INV_X1 U22202 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n19054) );
  AOI221_X1 U22203 ( .B1(n19812), .B2(n19015), .C1(n19812), .C2(n19112), .A(
        n19014), .ZN(n19053) );
  INV_X1 U22204 ( .A(n19053), .ZN(n19017) );
  NOR2_X1 U22205 ( .A1(n19775), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19302) );
  NOR2_X1 U22206 ( .A1(n19302), .A2(n19016), .ZN(n19110) );
  NOR2_X1 U22207 ( .A1(n19326), .A2(n19792), .ZN(n19300) );
  AOI21_X1 U22208 ( .B1(n19029), .B2(n19110), .A(n19300), .ZN(n19052) );
  AOI221_X1 U22209 ( .B1(n19054), .B2(n19270), .C1(n19017), .C2(n19270), .A(
        n19052), .ZN(n19040) );
  NAND2_X1 U22210 ( .A1(n19775), .A2(n19299), .ZN(n19156) );
  AOI22_X1 U22211 ( .A1(n19326), .A2(n19042), .B1(n19018), .B2(n19156), .ZN(
        n19021) );
  NOR2_X1 U22212 ( .A1(n19023), .A2(n19022), .ZN(n19026) );
  NOR3_X1 U22213 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n19024), .A3(
        n19086), .ZN(n19025) );
  AOI221_X1 U22214 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n19317), .C1(n19026), 
        .C2(n19328), .A(n19025), .ZN(n19027) );
  OAI21_X1 U22215 ( .B1(n19028), .B2(n19171), .A(n19027), .ZN(P3_U2835) );
  AND2_X1 U22216 ( .A1(n19078), .A2(n19029), .ZN(n19063) );
  AOI22_X1 U22217 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n19031), .B1(
        n19030), .B2(n19063), .ZN(n19036) );
  AOI22_X1 U22218 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n19325), .B1(
        n19239), .B2(n19032), .ZN(n19035) );
  INV_X1 U22219 ( .A(n19033), .ZN(n19034) );
  OAI211_X1 U22220 ( .C1(n19036), .C2(n19314), .A(n19035), .B(n19034), .ZN(
        P3_U2836) );
  NOR2_X1 U22221 ( .A1(n19038), .A2(n19037), .ZN(n19043) );
  OAI22_X1 U22222 ( .A1(n19040), .A2(n19042), .B1(n19182), .B2(n19039), .ZN(
        n19041) );
  AOI21_X1 U22223 ( .B1(n19043), .B2(n19042), .A(n19041), .ZN(n19048) );
  AOI22_X1 U22224 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19325), .B1(
        n19317), .B2(P3_REIP_REG_25__SCAN_IN), .ZN(n19047) );
  AOI22_X1 U22225 ( .A1(n19333), .A2(n19045), .B1(n19239), .B2(n19044), .ZN(
        n19046) );
  OAI211_X1 U22226 ( .C1(n19048), .C2(n19314), .A(n19047), .B(n19046), .ZN(
        P3_U2837) );
  INV_X1 U22227 ( .A(n19811), .ZN(n19307) );
  OAI22_X1 U22228 ( .A1(n19050), .A2(n19182), .B1(n19049), .B2(n19307), .ZN(
        n19051) );
  NOR3_X1 U22229 ( .A1(n19325), .A2(n19052), .A3(n19051), .ZN(n19055) );
  AOI21_X1 U22230 ( .B1(n19053), .B2(n19055), .A(n19317), .ZN(n19062) );
  AOI21_X1 U22231 ( .B1(n19234), .B2(n19055), .A(n19054), .ZN(n19056) );
  AOI22_X1 U22232 ( .A1(n19058), .A2(n19057), .B1(n19062), .B2(n19056), .ZN(
        n19060) );
  OAI211_X1 U22233 ( .C1(n19061), .C2(n19171), .A(n19060), .B(n19059), .ZN(
        P3_U2838) );
  INV_X1 U22234 ( .A(n19325), .ZN(n19318) );
  OAI221_X1 U22235 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n19063), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n19318), .A(n19062), .ZN(
        n19064) );
  OAI211_X1 U22236 ( .C1(n19066), .C2(n19171), .A(n19065), .B(n19064), .ZN(
        P3_U2839) );
  AOI22_X1 U22237 ( .A1(n19317), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n19239), 
        .B2(n19067), .ZN(n19083) );
  NOR2_X1 U22238 ( .A1(n19811), .A2(n19073), .ZN(n19206) );
  AOI21_X1 U22239 ( .B1(n19068), .B2(n19100), .A(n19794), .ZN(n19069) );
  AOI221_X1 U22240 ( .B1(n19112), .B2(n19812), .C1(n19085), .C2(n19812), .A(
        n19069), .ZN(n19099) );
  NAND2_X1 U22241 ( .A1(n19326), .A2(n19070), .ZN(n19071) );
  OAI211_X1 U22242 ( .C1(n19077), .C2(n19206), .A(n19099), .B(n19071), .ZN(
        n19090) );
  OAI21_X1 U22243 ( .B1(n19084), .B2(n19792), .A(n19074), .ZN(n19075) );
  OAI211_X1 U22244 ( .C1(n19214), .C2(n19076), .A(n19088), .B(n19075), .ZN(
        n19081) );
  AOI21_X1 U22245 ( .B1(n19078), .B2(n19077), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19079) );
  INV_X1 U22246 ( .A(n19079), .ZN(n19080) );
  OAI211_X1 U22247 ( .C1(n19090), .C2(n19081), .A(n19327), .B(n19080), .ZN(
        n19082) );
  OAI211_X1 U22248 ( .C1(n19318), .C2(n19084), .A(n19083), .B(n19082), .ZN(
        P3_U2840) );
  AOI21_X1 U22249 ( .B1(n19131), .B2(n19087), .A(n19775), .ZN(n19089) );
  NOR2_X1 U22250 ( .A1(n19089), .A2(n19135), .ZN(n19098) );
  AOI21_X1 U22251 ( .B1(n19091), .B2(n19156), .A(n19090), .ZN(n19092) );
  AOI211_X1 U22252 ( .C1(n19098), .C2(n19092), .A(n19317), .B(n21959), .ZN(
        n19093) );
  AOI21_X1 U22253 ( .B1(n19239), .B2(n19094), .A(n19093), .ZN(n19096) );
  OAI211_X1 U22254 ( .C1(n19097), .C2(n19109), .A(n19096), .B(n19095), .ZN(
        P3_U2841) );
  NAND3_X1 U22255 ( .A1(n21877), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n19156), 
        .ZN(n19101) );
  OAI211_X1 U22256 ( .C1(n19109), .C2(n19105), .A(n19104), .B(n19103), .ZN(
        P3_U2842) );
  AOI22_X1 U22257 ( .A1(n19317), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n19239), 
        .B2(n19106), .ZN(n19107) );
  OAI221_X1 U22258 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n19109), 
        .C1(n21877), .C2(n19108), .A(n19107), .ZN(P3_U2843) );
  INV_X1 U22259 ( .A(n19135), .ZN(n19115) );
  AOI21_X1 U22260 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19110), .A(
        n19300), .ZN(n19111) );
  AOI221_X1 U22261 ( .B1(n19113), .B2(n19812), .C1(n19112), .C2(n19812), .A(
        n19111), .ZN(n19114) );
  OAI211_X1 U22262 ( .C1(n19116), .C2(n19206), .A(n19115), .B(n19114), .ZN(
        n19126) );
  INV_X1 U22263 ( .A(n19300), .ZN(n19273) );
  OAI221_X1 U22264 ( .B1(n19126), .B2(n19127), .C1(n19126), .C2(n19273), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19124) );
  AOI22_X1 U22265 ( .A1(n19272), .A2(n19812), .B1(n19271), .B2(n19304), .ZN(
        n19117) );
  NAND2_X1 U22266 ( .A1(n19118), .A2(n19292), .ZN(n19142) );
  NAND2_X1 U22267 ( .A1(n19119), .A2(n19142), .ZN(n19195) );
  NAND2_X1 U22268 ( .A1(n19327), .A2(n19195), .ZN(n19228) );
  NOR2_X1 U22269 ( .A1(n19120), .A2(n19228), .ZN(n19137) );
  AOI22_X1 U22270 ( .A1(n19239), .A2(n19122), .B1(n19137), .B2(n19121), .ZN(
        n19123) );
  OAI221_X1 U22271 ( .B1(n19317), .B2(n19124), .C1(n19328), .C2(n19894), .A(
        n19123), .ZN(P3_U2844) );
  AOI22_X1 U22272 ( .A1(n19317), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n19239), 
        .B2(n19125), .ZN(n19130) );
  NAND3_X1 U22273 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n19328), .A3(
        n19126), .ZN(n19129) );
  NAND3_X1 U22274 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19137), .A3(
        n19127), .ZN(n19128) );
  NAND3_X1 U22275 ( .A1(n19130), .A2(n19129), .A3(n19128), .ZN(P3_U2845) );
  NAND2_X1 U22276 ( .A1(n19326), .A2(n19178), .ZN(n19220) );
  OAI211_X1 U22277 ( .C1(n19775), .C2(n19131), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n19220), .ZN(n19132) );
  INV_X1 U22278 ( .A(n19132), .ZN(n19133) );
  NAND2_X1 U22279 ( .A1(n19812), .A2(n19157), .ZN(n19176) );
  OAI211_X1 U22280 ( .C1(n19214), .C2(n19134), .A(n19133), .B(n19176), .ZN(
        n19145) );
  OAI221_X1 U22281 ( .B1(n19135), .B2(n19270), .C1(n19135), .C2(n19145), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n19140) );
  AOI22_X1 U22282 ( .A1(n19138), .A2(n19239), .B1(n19137), .B2(n19136), .ZN(
        n19139) );
  OAI221_X1 U22283 ( .B1(n19317), .B2(n19140), .C1(n19328), .C2(n22035), .A(
        n19139), .ZN(P3_U2846) );
  NOR2_X1 U22284 ( .A1(n19141), .A2(n19182), .ZN(n19147) );
  OR2_X1 U22285 ( .A1(n19142), .A2(n19161), .ZN(n19155) );
  OAI21_X1 U22286 ( .B1(n19163), .B2(n19155), .A(n19143), .ZN(n19144) );
  AOI22_X1 U22287 ( .A1(n19147), .A2(n19146), .B1(n19145), .B2(n19144), .ZN(
        n19154) );
  AOI22_X1 U22288 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19325), .B1(
        n19317), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n19153) );
  NOR2_X1 U22289 ( .A1(n19148), .A2(n19288), .ZN(n19150) );
  AOI22_X1 U22290 ( .A1(n19151), .A2(n19239), .B1(n19150), .B2(n19149), .ZN(
        n19152) );
  OAI211_X1 U22291 ( .C1(n19154), .C2(n19314), .A(n19153), .B(n19152), .ZN(
        P3_U2847) );
  NAND2_X1 U22292 ( .A1(n19163), .A2(n19155), .ZN(n19165) );
  NAND2_X1 U22293 ( .A1(n19327), .A2(n19156), .ZN(n19336) );
  NOR2_X1 U22294 ( .A1(n19964), .A2(n19178), .ZN(n19222) );
  INV_X1 U22295 ( .A(n19222), .ZN(n19204) );
  NOR2_X1 U22296 ( .A1(n19158), .A2(n19204), .ZN(n19193) );
  OR2_X1 U22297 ( .A1(n19775), .A2(n19193), .ZN(n19186) );
  OAI21_X1 U22298 ( .B1(n19158), .B2(n19157), .A(n19812), .ZN(n19159) );
  NAND4_X1 U22299 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19186), .A3(
        n19220), .A4(n19159), .ZN(n19160) );
  AOI21_X1 U22300 ( .B1(n19326), .B2(n19161), .A(n19160), .ZN(n19162) );
  OAI222_X1 U22301 ( .A1(n19163), .A2(n19318), .B1(n19336), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(n19314), .C2(n19162), .ZN(
        n19164) );
  AOI22_X1 U22302 ( .A1(n19317), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n19165), 
        .B2(n19164), .ZN(n19170) );
  INV_X1 U22303 ( .A(n19166), .ZN(n19168) );
  AOI22_X1 U22304 ( .A1(n19240), .A2(n19168), .B1(n19333), .B2(n19167), .ZN(
        n19169) );
  OAI211_X1 U22305 ( .C1(n19172), .C2(n19171), .A(n19170), .B(n19169), .ZN(
        P3_U2848) );
  AOI22_X1 U22306 ( .A1(n19317), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n19239), 
        .B2(n19173), .ZN(n19189) );
  AOI21_X1 U22307 ( .B1(n19326), .B2(n19175), .A(n19174), .ZN(n19192) );
  OAI21_X1 U22308 ( .B1(n19177), .B2(n19182), .A(n19176), .ZN(n19202) );
  INV_X1 U22309 ( .A(n19178), .ZN(n19179) );
  AOI21_X1 U22310 ( .B1(n19207), .B2(n19179), .A(n19794), .ZN(n19180) );
  AOI21_X1 U22311 ( .B1(n19812), .B2(n19181), .A(n19180), .ZN(n19208) );
  OAI21_X1 U22312 ( .B1(n19183), .B2(n19182), .A(n19208), .ZN(n19184) );
  AOI211_X1 U22313 ( .C1(n19811), .C2(n19185), .A(n19202), .B(n19184), .ZN(
        n19191) );
  OAI211_X1 U22314 ( .C1(n19214), .C2(n19192), .A(n19191), .B(n19186), .ZN(
        n19187) );
  OAI211_X1 U22315 ( .C1(n19314), .C2(n19187), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19328), .ZN(n19188) );
  OAI211_X1 U22316 ( .C1(n19228), .C2(n19190), .A(n19189), .B(n19188), .ZN(
        P3_U2849) );
  OAI211_X1 U22317 ( .C1(n19193), .C2(n19775), .A(n19192), .B(n19191), .ZN(
        n19194) );
  OAI221_X1 U22318 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n19196), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n19195), .A(n19194), .ZN(
        n19200) );
  AOI22_X1 U22319 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19325), .B1(
        n19239), .B2(n19197), .ZN(n19199) );
  OAI211_X1 U22320 ( .C1(n19314), .C2(n19200), .A(n19199), .B(n19198), .ZN(
        P3_U2850) );
  AOI22_X1 U22321 ( .A1(n19317), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n19239), 
        .B2(n19201), .ZN(n19211) );
  AOI211_X1 U22322 ( .C1(n19811), .C2(n19203), .A(n19314), .B(n19202), .ZN(
        n19221) );
  OAI21_X1 U22323 ( .B1(n19227), .B2(n19204), .A(n19792), .ZN(n19205) );
  OAI211_X1 U22324 ( .C1(n19207), .C2(n19206), .A(n19221), .B(n19205), .ZN(
        n19215) );
  OAI21_X1 U22325 ( .B1(n19775), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n19208), .ZN(n19209) );
  OAI211_X1 U22326 ( .C1(n19215), .C2(n19209), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19328), .ZN(n19210) );
  OAI211_X1 U22327 ( .C1(n19212), .C2(n19228), .A(n19211), .B(n19210), .ZN(
        P3_U2851) );
  AOI22_X1 U22328 ( .A1(n19317), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n19239), 
        .B2(n19213), .ZN(n19218) );
  AOI21_X1 U22329 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19220), .A(
        n19214), .ZN(n19216) );
  OAI211_X1 U22330 ( .C1(n19216), .C2(n19215), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n19328), .ZN(n19217) );
  OAI211_X1 U22331 ( .C1(n19219), .C2(n19228), .A(n19218), .B(n19217), .ZN(
        P3_U2852) );
  OAI211_X1 U22332 ( .C1(n19775), .C2(n19222), .A(n19221), .B(n19220), .ZN(
        n19223) );
  NAND2_X1 U22333 ( .A1(n19328), .A2(n19223), .ZN(n19226) );
  AOI22_X1 U22334 ( .A1(n19317), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n19239), 
        .B2(n19224), .ZN(n19225) );
  OAI221_X1 U22335 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19228), .C1(
        n19227), .C2(n19226), .A(n19225), .ZN(P3_U2853) );
  INV_X1 U22336 ( .A(n19229), .ZN(n19235) );
  INV_X1 U22337 ( .A(n19272), .ZN(n19230) );
  AOI221_X1 U22338 ( .B1(n19230), .B2(n19812), .C1(n19229), .C2(n19812), .A(
        n19302), .ZN(n19231) );
  OAI221_X1 U22339 ( .B1(n19300), .B2(n19271), .C1(n19300), .C2(n19235), .A(
        n19231), .ZN(n19253) );
  NOR2_X1 U22340 ( .A1(n19251), .A2(n19253), .ZN(n19244) );
  OAI21_X1 U22341 ( .B1(n19244), .B2(n19314), .A(n19318), .ZN(n19232) );
  AOI21_X1 U22342 ( .B1(n19321), .B2(n19255), .A(n19232), .ZN(n19252) );
  AOI211_X1 U22343 ( .C1(n19234), .C2(n19318), .A(n19252), .B(n19233), .ZN(
        n19237) );
  NAND3_X1 U22344 ( .A1(n19235), .A2(n19327), .A3(n19292), .ZN(n19256) );
  NOR4_X1 U22345 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19255), .A3(
        n19251), .A4(n19256), .ZN(n19236) );
  AOI211_X1 U22346 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n19317), .A(n19237), .B(
        n19236), .ZN(n19242) );
  AOI22_X1 U22347 ( .A1(n18918), .A2(n19240), .B1(n19239), .B2(n19238), .ZN(
        n19241) );
  OAI211_X1 U22348 ( .C1(n19288), .C2(n19243), .A(n19242), .B(n19241), .ZN(
        P3_U2854) );
  NOR3_X1 U22349 ( .A1(n19244), .A2(n19255), .A3(n19256), .ZN(n19249) );
  INV_X1 U22350 ( .A(n19245), .ZN(n19247) );
  OAI22_X1 U22351 ( .A1(n19297), .A2(n19247), .B1(n19288), .B2(n19246), .ZN(
        n19248) );
  AOI211_X1 U22352 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n19317), .A(n19249), .B(
        n19248), .ZN(n19250) );
  OAI21_X1 U22353 ( .B1(n19252), .B2(n19251), .A(n19250), .ZN(P3_U2855) );
  OAI21_X1 U22354 ( .B1(n19314), .B2(n19253), .A(n19328), .ZN(n19261) );
  NAND2_X1 U22355 ( .A1(n19317), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n19254) );
  OAI221_X1 U22356 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19256), .C1(
        n19255), .C2(n19261), .A(n19254), .ZN(n19257) );
  AOI21_X1 U22357 ( .B1(n19331), .B2(n19258), .A(n19257), .ZN(n19259) );
  OAI21_X1 U22358 ( .B1(n19288), .B2(n19260), .A(n19259), .ZN(P3_U2856) );
  NOR2_X1 U22359 ( .A1(n19328), .A2(n19872), .ZN(n19265) );
  NAND3_X1 U22360 ( .A1(n19327), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n19292), .ZN(n19269) );
  NOR2_X1 U22361 ( .A1(n10406), .A2(n19269), .ZN(n19263) );
  INV_X1 U22362 ( .A(n19261), .ZN(n19262) );
  MUX2_X1 U22363 ( .A(n19263), .B(n19262), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n19264) );
  AOI211_X1 U22364 ( .C1(n19331), .C2(n19266), .A(n19265), .B(n19264), .ZN(
        n19267) );
  OAI21_X1 U22365 ( .B1(n19288), .B2(n19268), .A(n19267), .ZN(P3_U2857) );
  NOR2_X1 U22366 ( .A1(n19328), .A2(n19869), .ZN(n19280) );
  INV_X1 U22367 ( .A(n19269), .ZN(n19278) );
  NOR2_X1 U22368 ( .A1(n19325), .A2(n19270), .ZN(n19276) );
  INV_X1 U22369 ( .A(n19271), .ZN(n19274) );
  NOR2_X1 U22370 ( .A1(n19299), .A2(n19272), .ZN(n19310) );
  AOI211_X1 U22371 ( .C1(n19274), .C2(n19273), .A(n19310), .B(n19302), .ZN(
        n19275) );
  AOI21_X1 U22372 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19275), .A(
        n19314), .ZN(n19293) );
  NOR2_X1 U22373 ( .A1(n19325), .A2(n19293), .ZN(n19290) );
  NOR2_X1 U22374 ( .A1(n19276), .A2(n19290), .ZN(n19277) );
  MUX2_X1 U22375 ( .A(n19278), .B(n19277), .S(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n19279) );
  AOI211_X1 U22376 ( .C1(n19281), .C2(n19331), .A(n19280), .B(n19279), .ZN(
        n19282) );
  OAI21_X1 U22377 ( .B1(n19288), .B2(n19283), .A(n19282), .ZN(P3_U2858) );
  OAI21_X1 U22378 ( .B1(n19286), .B2(n19285), .A(n19284), .ZN(n19287) );
  OAI22_X1 U22379 ( .A1(n19290), .A2(n19289), .B1(n19288), .B2(n19287), .ZN(
        n19291) );
  AOI21_X1 U22380 ( .B1(n19293), .B2(n19292), .A(n19291), .ZN(n19295) );
  OAI211_X1 U22381 ( .C1(n19297), .C2(n19296), .A(n19295), .B(n19294), .ZN(
        P3_U2859) );
  NAND2_X1 U22382 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19298) );
  OAI22_X1 U22383 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19300), .B1(
        n19299), .B2(n19298), .ZN(n19301) );
  OAI21_X1 U22384 ( .B1(n19302), .B2(n19301), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19306) );
  NAND3_X1 U22385 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19304), .A3(
        n19303), .ZN(n19305) );
  OAI211_X1 U22386 ( .C1(n19308), .C2(n19307), .A(n19306), .B(n19305), .ZN(
        n19309) );
  AOI211_X1 U22387 ( .C1(n19311), .C2(n19810), .A(n19310), .B(n19309), .ZN(
        n19315) );
  AOI21_X1 U22388 ( .B1(n19325), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n19312), .ZN(n19313) );
  OAI21_X1 U22389 ( .B1(n19315), .B2(n19314), .A(n19313), .ZN(P3_U2860) );
  AOI22_X1 U22390 ( .A1(n19317), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n19331), 
        .B2(n19316), .ZN(n19324) );
  OAI21_X1 U22391 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19336), .A(
        n19318), .ZN(n19320) );
  AOI22_X1 U22392 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19320), .B1(
        n19333), .B2(n19319), .ZN(n19323) );
  OAI211_X1 U22393 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19326), .A(
        n19321), .B(n10622), .ZN(n19322) );
  NAND3_X1 U22394 ( .A1(n19324), .A2(n19323), .A3(n19322), .ZN(P3_U2861) );
  AOI21_X1 U22395 ( .B1(n19327), .B2(n19326), .A(n19325), .ZN(n19335) );
  INV_X1 U22396 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19975) );
  NOR2_X1 U22397 ( .A1(n19328), .A2(n19975), .ZN(n19329) );
  AOI221_X1 U22398 ( .B1(n19333), .B2(n19332), .C1(n19331), .C2(n19330), .A(
        n19329), .ZN(n19334) );
  OAI221_X1 U22399 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19336), .C1(
        n19964), .C2(n19335), .A(n19334), .ZN(P3_U2862) );
  AOI211_X1 U22400 ( .C1(n19338), .C2(n19337), .A(n20001), .B(n19946), .ZN(
        n19830) );
  INV_X1 U22401 ( .A(n19339), .ZN(n19379) );
  OAI21_X1 U22402 ( .B1(n19830), .B2(n19379), .A(n19344), .ZN(n19340) );
  OAI221_X1 U22403 ( .B1(n19797), .B2(n19984), .C1(n19797), .C2(n19344), .A(
        n19340), .ZN(P3_U2863) );
  NOR2_X1 U22404 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19803), .ZN(
        n19514) );
  NOR2_X1 U22405 ( .A1(n19604), .A2(n19514), .ZN(n19341) );
  OAI22_X1 U22406 ( .A1(n19343), .A2(n19805), .B1(n19342), .B2(n19341), .ZN(
        P3_U2866) );
  NOR2_X1 U22407 ( .A1(n19806), .A2(n19344), .ZN(P3_U2867) );
  NAND2_X1 U22408 ( .A1(n19659), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19725) );
  NOR2_X1 U22409 ( .A1(n19803), .A2(n19805), .ZN(n19721) );
  INV_X1 U22410 ( .A(n19721), .ZN(n19656) );
  NAND2_X1 U22411 ( .A1(n19797), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19580) );
  NOR2_X2 U22412 ( .A1(n19656), .A2(n19580), .ZN(n19713) );
  NAND2_X1 U22413 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19799), .ZN(
        n19559) );
  NOR2_X2 U22414 ( .A1(n19656), .A2(n19559), .ZN(n19758) );
  NAND2_X1 U22415 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19659), .ZN(n19689) );
  INV_X1 U22416 ( .A(n19689), .ZN(n19719) );
  NOR2_X2 U22417 ( .A1(n19421), .A2(n19345), .ZN(n19718) );
  NAND2_X1 U22418 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19513), .ZN(
        n19717) );
  NOR2_X2 U22419 ( .A1(n19797), .A2(n19717), .ZN(n19769) );
  NAND2_X1 U22420 ( .A1(n19799), .A2(n19797), .ZN(n19800) );
  NAND2_X1 U22421 ( .A1(n19803), .A2(n19805), .ZN(n19424) );
  NOR2_X2 U22422 ( .A1(n19800), .A2(n19424), .ZN(n19438) );
  NAND2_X1 U22423 ( .A1(n19416), .A2(n19445), .ZN(n19400) );
  AOI22_X1 U22424 ( .A1(n19758), .A2(n19719), .B1(n19718), .B2(n19373), .ZN(
        n19351) );
  INV_X1 U22425 ( .A(n19758), .ZN(n19774) );
  NAND2_X1 U22426 ( .A1(n19399), .A2(n19774), .ZN(n19686) );
  NAND2_X1 U22427 ( .A1(n19632), .A2(n19346), .ZN(n19534) );
  INV_X1 U22428 ( .A(n19534), .ZN(n19683) );
  AOI22_X1 U22429 ( .A1(n19659), .A2(n19686), .B1(n19683), .B2(n19400), .ZN(
        n19376) );
  NAND2_X1 U22430 ( .A1(n19348), .A2(n19347), .ZN(n19374) );
  NOR2_X2 U22431 ( .A1(n19349), .A2(n19374), .ZN(n19722) );
  AOI22_X1 U22432 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19376), .B1(
        n19438), .B2(n19722), .ZN(n19350) );
  OAI211_X1 U22433 ( .C1(n19725), .C2(n19399), .A(n19351), .B(n19350), .ZN(
        P3_U2868) );
  NAND2_X1 U22434 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19659), .ZN(n19693) );
  NAND2_X1 U22435 ( .A1(n19659), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19731) );
  INV_X1 U22436 ( .A(n19731), .ZN(n19690) );
  AND2_X1 U22437 ( .A1(n19632), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19726) );
  AOI22_X1 U22438 ( .A1(n19713), .A2(n19690), .B1(n19373), .B2(n19726), .ZN(
        n19353) );
  NOR2_X2 U22439 ( .A1(n19987), .A2(n19374), .ZN(n19728) );
  AOI22_X1 U22440 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19376), .B1(
        n19438), .B2(n19728), .ZN(n19352) );
  OAI211_X1 U22441 ( .C1(n19774), .C2(n19693), .A(n19353), .B(n19352), .ZN(
        P3_U2869) );
  NAND2_X1 U22442 ( .A1(n19659), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19737) );
  NOR2_X1 U22443 ( .A1(n21883), .A2(n19369), .ZN(n19732) );
  NOR2_X2 U22444 ( .A1(n19421), .A2(n19354), .ZN(n19733) );
  AOI22_X1 U22445 ( .A1(n19758), .A2(n19732), .B1(n19373), .B2(n19733), .ZN(
        n19357) );
  NOR2_X2 U22446 ( .A1(n19355), .A2(n19374), .ZN(n19734) );
  AOI22_X1 U22447 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19376), .B1(
        n19438), .B2(n19734), .ZN(n19356) );
  OAI211_X1 U22448 ( .C1(n19399), .C2(n19737), .A(n19357), .B(n19356), .ZN(
        P3_U2870) );
  NAND2_X1 U22449 ( .A1(n19659), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19743) );
  NAND2_X1 U22450 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19659), .ZN(n19701) );
  INV_X1 U22451 ( .A(n19701), .ZN(n19738) );
  NOR2_X2 U22452 ( .A1(n19421), .A2(n19358), .ZN(n19739) );
  AOI22_X1 U22453 ( .A1(n19758), .A2(n19738), .B1(n19373), .B2(n19739), .ZN(
        n19361) );
  NOR2_X2 U22454 ( .A1(n19359), .A2(n19374), .ZN(n19740) );
  AOI22_X1 U22455 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19376), .B1(
        n19438), .B2(n19740), .ZN(n19360) );
  OAI211_X1 U22456 ( .C1(n19399), .C2(n19743), .A(n19361), .B(n19360), .ZN(
        P3_U2871) );
  NAND2_X1 U22457 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19659), .ZN(n19617) );
  NAND2_X1 U22458 ( .A1(n19659), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19749) );
  INV_X1 U22459 ( .A(n19749), .ZN(n19613) );
  NOR2_X2 U22460 ( .A1(n19421), .A2(n19362), .ZN(n19744) );
  AOI22_X1 U22461 ( .A1(n19713), .A2(n19613), .B1(n19373), .B2(n19744), .ZN(
        n19365) );
  NOR2_X2 U22462 ( .A1(n19363), .A2(n19374), .ZN(n19746) );
  AOI22_X1 U22463 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19376), .B1(
        n19438), .B2(n19746), .ZN(n19364) );
  OAI211_X1 U22464 ( .C1(n19774), .C2(n19617), .A(n19365), .B(n19364), .ZN(
        P3_U2872) );
  NAND2_X1 U22465 ( .A1(n19659), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19755) );
  NAND2_X1 U22466 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19659), .ZN(n19707) );
  INV_X1 U22467 ( .A(n19707), .ZN(n19750) );
  NOR2_X2 U22468 ( .A1(n19421), .A2(n13829), .ZN(n19751) );
  AOI22_X1 U22469 ( .A1(n19758), .A2(n19750), .B1(n19373), .B2(n19751), .ZN(
        n19368) );
  NOR2_X2 U22470 ( .A1(n19366), .A2(n19374), .ZN(n19752) );
  AOI22_X1 U22471 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19376), .B1(
        n19438), .B2(n19752), .ZN(n19367) );
  OAI211_X1 U22472 ( .C1(n19399), .C2(n19755), .A(n19368), .B(n19367), .ZN(
        P3_U2873) );
  NAND2_X1 U22473 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19659), .ZN(n19623) );
  NOR2_X1 U22474 ( .A1(n16511), .A2(n19369), .ZN(n19620) );
  NOR2_X2 U22475 ( .A1(n13839), .A2(n19421), .ZN(n19756) );
  AOI22_X1 U22476 ( .A1(n19758), .A2(n19620), .B1(n19373), .B2(n19756), .ZN(
        n19372) );
  NOR2_X2 U22477 ( .A1(n19370), .A2(n19374), .ZN(n19759) );
  AOI22_X1 U22478 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19376), .B1(
        n19438), .B2(n19759), .ZN(n19371) );
  OAI211_X1 U22479 ( .C1(n19399), .C2(n19623), .A(n19372), .B(n19371), .ZN(
        P3_U2874) );
  NAND2_X1 U22480 ( .A1(n19659), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19654) );
  NAND2_X1 U22481 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19659), .ZN(n19773) );
  INV_X1 U22482 ( .A(n19773), .ZN(n19648) );
  NOR2_X2 U22483 ( .A1(n13920), .A2(n19421), .ZN(n19765) );
  AOI22_X1 U22484 ( .A1(n19713), .A2(n19648), .B1(n19373), .B2(n19765), .ZN(
        n19378) );
  NOR2_X2 U22485 ( .A1(n19375), .A2(n19374), .ZN(n19768) );
  AOI22_X1 U22486 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19376), .B1(
        n19438), .B2(n19768), .ZN(n19377) );
  OAI211_X1 U22487 ( .C1(n19774), .C2(n19654), .A(n19378), .B(n19377), .ZN(
        P3_U2875) );
  NAND2_X1 U22488 ( .A1(n19799), .A2(n19680), .ZN(n19655) );
  NOR2_X1 U22489 ( .A1(n19424), .A2(n19655), .ZN(n19395) );
  AOI22_X1 U22490 ( .A1(n19713), .A2(n19719), .B1(n19718), .B2(n19395), .ZN(
        n19382) );
  INV_X1 U22491 ( .A(n19717), .ZN(n19380) );
  INV_X1 U22492 ( .A(n19424), .ZN(n19423) );
  NOR3_X1 U22493 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19379), .A3(
        n19421), .ZN(n19657) );
  AOI22_X1 U22494 ( .A1(n19659), .A2(n19380), .B1(n19423), .B2(n19657), .ZN(
        n19396) );
  NOR2_X2 U22495 ( .A1(n19424), .A2(n19559), .ZN(n19464) );
  AOI22_X1 U22496 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19396), .B1(
        n19722), .B2(n19464), .ZN(n19381) );
  OAI211_X1 U22497 ( .C1(n19725), .C2(n19416), .A(n19382), .B(n19381), .ZN(
        P3_U2876) );
  INV_X1 U22498 ( .A(n19693), .ZN(n19727) );
  AOI22_X1 U22499 ( .A1(n19713), .A2(n19727), .B1(n19726), .B2(n19395), .ZN(
        n19384) );
  AOI22_X1 U22500 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19396), .B1(
        n19728), .B2(n19464), .ZN(n19383) );
  OAI211_X1 U22501 ( .C1(n19416), .C2(n19731), .A(n19384), .B(n19383), .ZN(
        P3_U2877) );
  AOI22_X1 U22502 ( .A1(n19713), .A2(n19732), .B1(n19733), .B2(n19395), .ZN(
        n19386) );
  AOI22_X1 U22503 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19396), .B1(
        n19734), .B2(n19464), .ZN(n19385) );
  OAI211_X1 U22504 ( .C1(n19416), .C2(n19737), .A(n19386), .B(n19385), .ZN(
        P3_U2878) );
  AOI22_X1 U22505 ( .A1(n19713), .A2(n19738), .B1(n19739), .B2(n19395), .ZN(
        n19388) );
  AOI22_X1 U22506 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19396), .B1(
        n19740), .B2(n19464), .ZN(n19387) );
  OAI211_X1 U22507 ( .C1(n19416), .C2(n19743), .A(n19388), .B(n19387), .ZN(
        P3_U2879) );
  AOI22_X1 U22508 ( .A1(n19769), .A2(n19613), .B1(n19744), .B2(n19395), .ZN(
        n19390) );
  AOI22_X1 U22509 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19396), .B1(
        n19746), .B2(n19464), .ZN(n19389) );
  OAI211_X1 U22510 ( .C1(n19399), .C2(n19617), .A(n19390), .B(n19389), .ZN(
        P3_U2880) );
  INV_X1 U22511 ( .A(n19755), .ZN(n19704) );
  AOI22_X1 U22512 ( .A1(n19769), .A2(n19704), .B1(n19751), .B2(n19395), .ZN(
        n19392) );
  AOI22_X1 U22513 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19396), .B1(
        n19752), .B2(n19464), .ZN(n19391) );
  OAI211_X1 U22514 ( .C1(n19399), .C2(n19707), .A(n19392), .B(n19391), .ZN(
        P3_U2881) );
  AOI22_X1 U22515 ( .A1(n19713), .A2(n19620), .B1(n19756), .B2(n19395), .ZN(
        n19394) );
  AOI22_X1 U22516 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19396), .B1(
        n19759), .B2(n19464), .ZN(n19393) );
  OAI211_X1 U22517 ( .C1(n19416), .C2(n19623), .A(n19394), .B(n19393), .ZN(
        P3_U2882) );
  AOI22_X1 U22518 ( .A1(n19769), .A2(n19648), .B1(n19765), .B2(n19395), .ZN(
        n19398) );
  AOI22_X1 U22519 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19396), .B1(
        n19768), .B2(n19464), .ZN(n19397) );
  OAI211_X1 U22520 ( .C1(n19399), .C2(n19654), .A(n19398), .B(n19397), .ZN(
        P3_U2883) );
  NOR2_X2 U22521 ( .A1(n19580), .A2(n19424), .ZN(n19481) );
  NOR2_X1 U22522 ( .A1(n19464), .A2(n19481), .ZN(n19446) );
  NOR2_X1 U22523 ( .A1(n19839), .A2(n19446), .ZN(n19417) );
  AOI22_X1 U22524 ( .A1(n19769), .A2(n19719), .B1(n19718), .B2(n19417), .ZN(
        n19403) );
  INV_X1 U22525 ( .A(n19446), .ZN(n19401) );
  OAI221_X1 U22526 ( .B1(n19401), .B2(n19685), .C1(n19401), .C2(n19400), .A(
        n19683), .ZN(n19418) );
  AOI22_X1 U22527 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19418), .B1(
        n19722), .B2(n19481), .ZN(n19402) );
  OAI211_X1 U22528 ( .C1(n19725), .C2(n19445), .A(n19403), .B(n19402), .ZN(
        P3_U2884) );
  AOI22_X1 U22529 ( .A1(n19769), .A2(n19727), .B1(n19726), .B2(n19417), .ZN(
        n19405) );
  AOI22_X1 U22530 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19418), .B1(
        n19728), .B2(n19481), .ZN(n19404) );
  OAI211_X1 U22531 ( .C1(n19445), .C2(n19731), .A(n19405), .B(n19404), .ZN(
        P3_U2885) );
  AOI22_X1 U22532 ( .A1(n19769), .A2(n19732), .B1(n19733), .B2(n19417), .ZN(
        n19407) );
  AOI22_X1 U22533 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19418), .B1(
        n19734), .B2(n19481), .ZN(n19406) );
  OAI211_X1 U22534 ( .C1(n19445), .C2(n19737), .A(n19407), .B(n19406), .ZN(
        P3_U2886) );
  AOI22_X1 U22535 ( .A1(n19769), .A2(n19738), .B1(n19739), .B2(n19417), .ZN(
        n19409) );
  AOI22_X1 U22536 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19418), .B1(
        n19740), .B2(n19481), .ZN(n19408) );
  OAI211_X1 U22537 ( .C1(n19445), .C2(n19743), .A(n19409), .B(n19408), .ZN(
        P3_U2887) );
  INV_X1 U22538 ( .A(n19617), .ZN(n19745) );
  AOI22_X1 U22539 ( .A1(n19769), .A2(n19745), .B1(n19744), .B2(n19417), .ZN(
        n19411) );
  AOI22_X1 U22540 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19418), .B1(
        n19746), .B2(n19481), .ZN(n19410) );
  OAI211_X1 U22541 ( .C1(n19445), .C2(n19749), .A(n19411), .B(n19410), .ZN(
        P3_U2888) );
  AOI22_X1 U22542 ( .A1(n19769), .A2(n19750), .B1(n19751), .B2(n19417), .ZN(
        n19413) );
  AOI22_X1 U22543 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19418), .B1(
        n19752), .B2(n19481), .ZN(n19412) );
  OAI211_X1 U22544 ( .C1(n19445), .C2(n19755), .A(n19413), .B(n19412), .ZN(
        P3_U2889) );
  INV_X1 U22545 ( .A(n19620), .ZN(n19763) );
  AOI22_X1 U22546 ( .A1(n19438), .A2(n19757), .B1(n19756), .B2(n19417), .ZN(
        n19415) );
  AOI22_X1 U22547 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19418), .B1(
        n19759), .B2(n19481), .ZN(n19414) );
  OAI211_X1 U22548 ( .C1(n19416), .C2(n19763), .A(n19415), .B(n19414), .ZN(
        P3_U2890) );
  INV_X1 U22549 ( .A(n19654), .ZN(n19767) );
  AOI22_X1 U22550 ( .A1(n19769), .A2(n19767), .B1(n19765), .B2(n19417), .ZN(
        n19420) );
  AOI22_X1 U22551 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19418), .B1(
        n19768), .B2(n19481), .ZN(n19419) );
  OAI211_X1 U22552 ( .C1(n19445), .C2(n19773), .A(n19420), .B(n19419), .ZN(
        P3_U2891) );
  AOI21_X1 U22553 ( .B1(n19629), .B2(n19422), .A(n19421), .ZN(n19720) );
  NAND2_X1 U22554 ( .A1(n19720), .A2(n19423), .ZN(n19442) );
  INV_X1 U22555 ( .A(n19442), .ZN(n19433) );
  NOR2_X1 U22556 ( .A1(n19799), .A2(n19424), .ZN(n19468) );
  AND2_X1 U22557 ( .A1(n19680), .A2(n19468), .ZN(n19441) );
  AOI22_X1 U22558 ( .A1(n19681), .A2(n19464), .B1(n19718), .B2(n19441), .ZN(
        n19426) );
  NAND2_X1 U22559 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19468), .ZN(
        n19504) );
  AOI22_X1 U22560 ( .A1(n19438), .A2(n19719), .B1(n19722), .B2(n19508), .ZN(
        n19425) );
  OAI211_X1 U22561 ( .C1(n19433), .C2(n21848), .A(n19426), .B(n19425), .ZN(
        P3_U2892) );
  INV_X1 U22562 ( .A(n19464), .ZN(n19462) );
  AOI22_X1 U22563 ( .A1(n19438), .A2(n19727), .B1(n19726), .B2(n19441), .ZN(
        n19428) );
  AOI22_X1 U22564 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19442), .B1(
        n19728), .B2(n19508), .ZN(n19427) );
  OAI211_X1 U22565 ( .C1(n19731), .C2(n19462), .A(n19428), .B(n19427), .ZN(
        P3_U2893) );
  INV_X1 U22566 ( .A(n19737), .ZN(n19694) );
  AOI22_X1 U22567 ( .A1(n19694), .A2(n19464), .B1(n19733), .B2(n19441), .ZN(
        n19430) );
  AOI22_X1 U22568 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19442), .B1(
        n19734), .B2(n19508), .ZN(n19429) );
  OAI211_X1 U22569 ( .C1(n19445), .C2(n19697), .A(n19430), .B(n19429), .ZN(
        P3_U2894) );
  INV_X1 U22570 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n22016) );
  INV_X1 U22571 ( .A(n19743), .ZN(n19698) );
  AOI22_X1 U22572 ( .A1(n19698), .A2(n19464), .B1(n19739), .B2(n19441), .ZN(
        n19432) );
  AOI22_X1 U22573 ( .A1(n19438), .A2(n19738), .B1(n19740), .B2(n19508), .ZN(
        n19431) );
  OAI211_X1 U22574 ( .C1(n19433), .C2(n22016), .A(n19432), .B(n19431), .ZN(
        P3_U2895) );
  AOI22_X1 U22575 ( .A1(n19438), .A2(n19745), .B1(n19744), .B2(n19441), .ZN(
        n19435) );
  AOI22_X1 U22576 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19442), .B1(
        n19746), .B2(n19508), .ZN(n19434) );
  OAI211_X1 U22577 ( .C1(n19749), .C2(n19462), .A(n19435), .B(n19434), .ZN(
        P3_U2896) );
  AOI22_X1 U22578 ( .A1(n19704), .A2(n19464), .B1(n19751), .B2(n19441), .ZN(
        n19437) );
  AOI22_X1 U22579 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19442), .B1(
        n19752), .B2(n19508), .ZN(n19436) );
  OAI211_X1 U22580 ( .C1(n19445), .C2(n19707), .A(n19437), .B(n19436), .ZN(
        P3_U2897) );
  AOI22_X1 U22581 ( .A1(n19438), .A2(n19620), .B1(n19756), .B2(n19441), .ZN(
        n19440) );
  AOI22_X1 U22582 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19442), .B1(
        n19759), .B2(n19508), .ZN(n19439) );
  OAI211_X1 U22583 ( .C1(n19623), .C2(n19462), .A(n19440), .B(n19439), .ZN(
        P3_U2898) );
  AOI22_X1 U22584 ( .A1(n19765), .A2(n19441), .B1(n19648), .B2(n19464), .ZN(
        n19444) );
  AOI22_X1 U22585 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19442), .B1(
        n19768), .B2(n19508), .ZN(n19443) );
  OAI211_X1 U22586 ( .C1(n19445), .C2(n19654), .A(n19444), .B(n19443), .ZN(
        P3_U2899) );
  NOR2_X1 U22587 ( .A1(n19508), .A2(n9731), .ZN(n19490) );
  NOR2_X1 U22588 ( .A1(n19839), .A2(n19490), .ZN(n19463) );
  AOI22_X1 U22589 ( .A1(n19681), .A2(n19481), .B1(n19718), .B2(n19463), .ZN(
        n19449) );
  OAI21_X1 U22590 ( .B1(n19446), .B2(n19629), .A(n19490), .ZN(n19447) );
  OAI211_X1 U22591 ( .C1(n9731), .C2(n19937), .A(n19632), .B(n19447), .ZN(
        n19465) );
  AOI22_X1 U22592 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19465), .B1(
        n19722), .B2(n9731), .ZN(n19448) );
  OAI211_X1 U22593 ( .C1(n19689), .C2(n19462), .A(n19449), .B(n19448), .ZN(
        P3_U2900) );
  AOI22_X1 U22594 ( .A1(n19727), .A2(n19464), .B1(n19726), .B2(n19463), .ZN(
        n19451) );
  AOI22_X1 U22595 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19465), .B1(
        n19728), .B2(n9731), .ZN(n19450) );
  OAI211_X1 U22596 ( .C1(n19731), .C2(n19488), .A(n19451), .B(n19450), .ZN(
        P3_U2901) );
  AOI22_X1 U22597 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19465), .B1(
        n19733), .B2(n19463), .ZN(n19453) );
  AOI22_X1 U22598 ( .A1(n19734), .A2(n9731), .B1(n19732), .B2(n19464), .ZN(
        n19452) );
  OAI211_X1 U22599 ( .C1(n19737), .C2(n19488), .A(n19453), .B(n19452), .ZN(
        P3_U2902) );
  AOI22_X1 U22600 ( .A1(n19698), .A2(n19481), .B1(n19739), .B2(n19463), .ZN(
        n19455) );
  AOI22_X1 U22601 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19465), .B1(
        n19740), .B2(n9731), .ZN(n19454) );
  OAI211_X1 U22602 ( .C1(n19701), .C2(n19462), .A(n19455), .B(n19454), .ZN(
        P3_U2903) );
  AOI22_X1 U22603 ( .A1(n19745), .A2(n19464), .B1(n19744), .B2(n19463), .ZN(
        n19457) );
  AOI22_X1 U22604 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19465), .B1(
        n19746), .B2(n9731), .ZN(n19456) );
  OAI211_X1 U22605 ( .C1(n19749), .C2(n19488), .A(n19457), .B(n19456), .ZN(
        P3_U2904) );
  AOI22_X1 U22606 ( .A1(n19751), .A2(n19463), .B1(n19750), .B2(n19464), .ZN(
        n19459) );
  AOI22_X1 U22607 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19465), .B1(
        n19752), .B2(n9731), .ZN(n19458) );
  OAI211_X1 U22608 ( .C1(n19755), .C2(n19488), .A(n19459), .B(n19458), .ZN(
        P3_U2905) );
  AOI22_X1 U22609 ( .A1(n19757), .A2(n19481), .B1(n19756), .B2(n19463), .ZN(
        n19461) );
  AOI22_X1 U22610 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19465), .B1(
        n19759), .B2(n9731), .ZN(n19460) );
  OAI211_X1 U22611 ( .C1(n19763), .C2(n19462), .A(n19461), .B(n19460), .ZN(
        P3_U2906) );
  AOI22_X1 U22612 ( .A1(n19767), .A2(n19464), .B1(n19765), .B2(n19463), .ZN(
        n19467) );
  AOI22_X1 U22613 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19465), .B1(
        n19768), .B2(n9731), .ZN(n19466) );
  OAI211_X1 U22614 ( .C1(n19773), .C2(n19488), .A(n19467), .B(n19466), .ZN(
        P3_U2907) );
  NOR2_X1 U22615 ( .A1(n19489), .A2(n19655), .ZN(n19484) );
  AOI22_X1 U22616 ( .A1(n19681), .A2(n19508), .B1(n19718), .B2(n19484), .ZN(
        n19470) );
  AOI22_X1 U22617 ( .A1(n19659), .A2(n19468), .B1(n19514), .B2(n19657), .ZN(
        n19485) );
  NOR2_X2 U22618 ( .A1(n19489), .A2(n19559), .ZN(n19549) );
  AOI22_X1 U22619 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19485), .B1(
        n19722), .B2(n19549), .ZN(n19469) );
  OAI211_X1 U22620 ( .C1(n19689), .C2(n19488), .A(n19470), .B(n19469), .ZN(
        P3_U2908) );
  AOI22_X1 U22621 ( .A1(n19727), .A2(n19481), .B1(n19726), .B2(n19484), .ZN(
        n19472) );
  AOI22_X1 U22622 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19485), .B1(
        n19728), .B2(n19549), .ZN(n19471) );
  OAI211_X1 U22623 ( .C1(n19731), .C2(n19504), .A(n19472), .B(n19471), .ZN(
        P3_U2909) );
  AOI22_X1 U22624 ( .A1(n19694), .A2(n19508), .B1(n19733), .B2(n19484), .ZN(
        n19474) );
  AOI22_X1 U22625 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19485), .B1(
        n19734), .B2(n19549), .ZN(n19473) );
  OAI211_X1 U22626 ( .C1(n19697), .C2(n19488), .A(n19474), .B(n19473), .ZN(
        P3_U2910) );
  AOI22_X1 U22627 ( .A1(n19739), .A2(n19484), .B1(n19738), .B2(n19481), .ZN(
        n19476) );
  AOI22_X1 U22628 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19485), .B1(
        n19740), .B2(n19549), .ZN(n19475) );
  OAI211_X1 U22629 ( .C1(n19743), .C2(n19504), .A(n19476), .B(n19475), .ZN(
        P3_U2911) );
  AOI22_X1 U22630 ( .A1(n19613), .A2(n19508), .B1(n19744), .B2(n19484), .ZN(
        n19478) );
  AOI22_X1 U22631 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19485), .B1(
        n19746), .B2(n19549), .ZN(n19477) );
  OAI211_X1 U22632 ( .C1(n19617), .C2(n19488), .A(n19478), .B(n19477), .ZN(
        P3_U2912) );
  AOI22_X1 U22633 ( .A1(n19704), .A2(n19508), .B1(n19751), .B2(n19484), .ZN(
        n19480) );
  AOI22_X1 U22634 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19485), .B1(
        n19752), .B2(n19549), .ZN(n19479) );
  OAI211_X1 U22635 ( .C1(n19707), .C2(n19488), .A(n19480), .B(n19479), .ZN(
        P3_U2913) );
  AOI22_X1 U22636 ( .A1(n19756), .A2(n19484), .B1(n19620), .B2(n19481), .ZN(
        n19483) );
  AOI22_X1 U22637 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19485), .B1(
        n19759), .B2(n19549), .ZN(n19482) );
  OAI211_X1 U22638 ( .C1(n19623), .C2(n19504), .A(n19483), .B(n19482), .ZN(
        P3_U2914) );
  AOI22_X1 U22639 ( .A1(n19765), .A2(n19484), .B1(n19648), .B2(n19508), .ZN(
        n19487) );
  AOI22_X1 U22640 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19485), .B1(
        n19768), .B2(n19549), .ZN(n19486) );
  OAI211_X1 U22641 ( .C1(n19654), .C2(n19488), .A(n19487), .B(n19486), .ZN(
        P3_U2915) );
  NOR2_X2 U22642 ( .A1(n19489), .A2(n19580), .ZN(n19576) );
  NOR2_X1 U22643 ( .A1(n19549), .A2(n19576), .ZN(n19535) );
  NOR2_X1 U22644 ( .A1(n19839), .A2(n19535), .ZN(n19507) );
  AOI22_X1 U22645 ( .A1(n19681), .A2(n9731), .B1(n19718), .B2(n19507), .ZN(
        n19493) );
  OAI21_X1 U22646 ( .B1(n19490), .B2(n19629), .A(n19535), .ZN(n19491) );
  OAI211_X1 U22647 ( .C1(n19576), .C2(n19937), .A(n19632), .B(n19491), .ZN(
        n19509) );
  AOI22_X1 U22648 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19509), .B1(
        n19722), .B2(n19576), .ZN(n19492) );
  OAI211_X1 U22649 ( .C1(n19689), .C2(n19504), .A(n19493), .B(n19492), .ZN(
        P3_U2916) );
  INV_X1 U22650 ( .A(n9731), .ZN(n19512) );
  AOI22_X1 U22651 ( .A1(n19727), .A2(n19508), .B1(n19726), .B2(n19507), .ZN(
        n19495) );
  AOI22_X1 U22652 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19509), .B1(
        n19728), .B2(n19576), .ZN(n19494) );
  OAI211_X1 U22653 ( .C1(n19731), .C2(n19512), .A(n19495), .B(n19494), .ZN(
        P3_U2917) );
  AOI22_X1 U22654 ( .A1(n19733), .A2(n19507), .B1(n19732), .B2(n19508), .ZN(
        n19497) );
  AOI22_X1 U22655 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19509), .B1(
        n19734), .B2(n19576), .ZN(n19496) );
  OAI211_X1 U22656 ( .C1(n19737), .C2(n19512), .A(n19497), .B(n19496), .ZN(
        P3_U2918) );
  AOI22_X1 U22657 ( .A1(n19739), .A2(n19507), .B1(n19738), .B2(n19508), .ZN(
        n19499) );
  AOI22_X1 U22658 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19509), .B1(
        n19740), .B2(n19576), .ZN(n19498) );
  OAI211_X1 U22659 ( .C1(n19743), .C2(n19512), .A(n19499), .B(n19498), .ZN(
        P3_U2919) );
  AOI22_X1 U22660 ( .A1(n19613), .A2(n9731), .B1(n19744), .B2(n19507), .ZN(
        n19501) );
  AOI22_X1 U22661 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19509), .B1(
        n19746), .B2(n19576), .ZN(n19500) );
  OAI211_X1 U22662 ( .C1(n19617), .C2(n19504), .A(n19501), .B(n19500), .ZN(
        P3_U2920) );
  AOI22_X1 U22663 ( .A1(n19704), .A2(n9731), .B1(n19751), .B2(n19507), .ZN(
        n19503) );
  AOI22_X1 U22664 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19509), .B1(
        n19752), .B2(n19576), .ZN(n19502) );
  OAI211_X1 U22665 ( .C1(n19707), .C2(n19504), .A(n19503), .B(n19502), .ZN(
        P3_U2921) );
  AOI22_X1 U22666 ( .A1(n19756), .A2(n19507), .B1(n19620), .B2(n19508), .ZN(
        n19506) );
  AOI22_X1 U22667 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19509), .B1(
        n19759), .B2(n19576), .ZN(n19505) );
  OAI211_X1 U22668 ( .C1(n19623), .C2(n19512), .A(n19506), .B(n19505), .ZN(
        P3_U2922) );
  AOI22_X1 U22669 ( .A1(n19767), .A2(n19508), .B1(n19765), .B2(n19507), .ZN(
        n19511) );
  AOI22_X1 U22670 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19509), .B1(
        n19768), .B2(n19576), .ZN(n19510) );
  OAI211_X1 U22671 ( .C1(n19773), .C2(n19512), .A(n19511), .B(n19510), .ZN(
        P3_U2923) );
  NAND2_X1 U22672 ( .A1(n19513), .A2(n19805), .ZN(n19557) );
  NOR2_X1 U22673 ( .A1(n19839), .A2(n19557), .ZN(n19530) );
  AOI22_X1 U22674 ( .A1(n19719), .A2(n9731), .B1(n19718), .B2(n19530), .ZN(
        n19516) );
  NAND2_X1 U22675 ( .A1(n19514), .A2(n19720), .ZN(n19531) );
  NOR2_X2 U22676 ( .A1(n19797), .A2(n19557), .ZN(n19599) );
  AOI22_X1 U22677 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19531), .B1(
        n19722), .B2(n19599), .ZN(n19515) );
  OAI211_X1 U22678 ( .C1(n19725), .C2(n19556), .A(n19516), .B(n19515), .ZN(
        P3_U2924) );
  AOI22_X1 U22679 ( .A1(n19727), .A2(n9731), .B1(n19726), .B2(n19530), .ZN(
        n19518) );
  AOI22_X1 U22680 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19531), .B1(
        n19728), .B2(n19599), .ZN(n19517) );
  OAI211_X1 U22681 ( .C1(n19731), .C2(n19556), .A(n19518), .B(n19517), .ZN(
        P3_U2925) );
  AOI22_X1 U22682 ( .A1(n19733), .A2(n19530), .B1(n19732), .B2(n9731), .ZN(
        n19520) );
  AOI22_X1 U22683 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19531), .B1(
        n19734), .B2(n19599), .ZN(n19519) );
  OAI211_X1 U22684 ( .C1(n19737), .C2(n19556), .A(n19520), .B(n19519), .ZN(
        P3_U2926) );
  AOI22_X1 U22685 ( .A1(n19739), .A2(n19530), .B1(n19738), .B2(n9731), .ZN(
        n19523) );
  AOI22_X1 U22686 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19531), .B1(
        n19740), .B2(n19599), .ZN(n19522) );
  OAI211_X1 U22687 ( .C1(n19743), .C2(n19556), .A(n19523), .B(n19522), .ZN(
        P3_U2927) );
  AOI22_X1 U22688 ( .A1(n19745), .A2(n9731), .B1(n19744), .B2(n19530), .ZN(
        n19525) );
  AOI22_X1 U22689 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19531), .B1(
        n19746), .B2(n19599), .ZN(n19524) );
  OAI211_X1 U22690 ( .C1(n19749), .C2(n19556), .A(n19525), .B(n19524), .ZN(
        P3_U2928) );
  AOI22_X1 U22691 ( .A1(n19751), .A2(n19530), .B1(n19750), .B2(n9731), .ZN(
        n19527) );
  AOI22_X1 U22692 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19531), .B1(
        n19752), .B2(n19599), .ZN(n19526) );
  OAI211_X1 U22693 ( .C1(n19755), .C2(n19556), .A(n19527), .B(n19526), .ZN(
        P3_U2929) );
  AOI22_X1 U22694 ( .A1(n19756), .A2(n19530), .B1(n19620), .B2(n9731), .ZN(
        n19529) );
  AOI22_X1 U22695 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19531), .B1(
        n19759), .B2(n19599), .ZN(n19528) );
  OAI211_X1 U22696 ( .C1(n19623), .C2(n19556), .A(n19529), .B(n19528), .ZN(
        P3_U2930) );
  AOI22_X1 U22697 ( .A1(n19767), .A2(n9731), .B1(n19765), .B2(n19530), .ZN(
        n19533) );
  AOI22_X1 U22698 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19531), .B1(
        n19768), .B2(n19599), .ZN(n19532) );
  OAI211_X1 U22699 ( .C1(n19773), .C2(n19556), .A(n19533), .B(n19532), .ZN(
        P3_U2931) );
  INV_X1 U22700 ( .A(n19576), .ZN(n19574) );
  INV_X1 U22701 ( .A(n19604), .ZN(n19603) );
  NOR2_X2 U22702 ( .A1(n19800), .A2(n19603), .ZN(n19625) );
  NOR2_X1 U22703 ( .A1(n19599), .A2(n19625), .ZN(n19581) );
  NOR2_X1 U22704 ( .A1(n19839), .A2(n19581), .ZN(n19552) );
  AOI22_X1 U22705 ( .A1(n19719), .A2(n19549), .B1(n19718), .B2(n19552), .ZN(
        n19538) );
  AOI221_X1 U22706 ( .B1(n19581), .B2(n19629), .C1(n19581), .C2(n19535), .A(
        n19534), .ZN(n19536) );
  INV_X1 U22707 ( .A(n19536), .ZN(n19553) );
  AOI22_X1 U22708 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19553), .B1(
        n19722), .B2(n19625), .ZN(n19537) );
  OAI211_X1 U22709 ( .C1(n19725), .C2(n19574), .A(n19538), .B(n19537), .ZN(
        P3_U2932) );
  AOI22_X1 U22710 ( .A1(n19727), .A2(n19549), .B1(n19726), .B2(n19552), .ZN(
        n19540) );
  AOI22_X1 U22711 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19553), .B1(
        n19728), .B2(n19625), .ZN(n19539) );
  OAI211_X1 U22712 ( .C1(n19731), .C2(n19574), .A(n19540), .B(n19539), .ZN(
        P3_U2933) );
  AOI22_X1 U22713 ( .A1(n19694), .A2(n19576), .B1(n19733), .B2(n19552), .ZN(
        n19542) );
  AOI22_X1 U22714 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19553), .B1(
        n19734), .B2(n19625), .ZN(n19541) );
  OAI211_X1 U22715 ( .C1(n19697), .C2(n19556), .A(n19542), .B(n19541), .ZN(
        P3_U2934) );
  AOI22_X1 U22716 ( .A1(n19698), .A2(n19576), .B1(n19739), .B2(n19552), .ZN(
        n19544) );
  AOI22_X1 U22717 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19553), .B1(
        n19740), .B2(n19625), .ZN(n19543) );
  OAI211_X1 U22718 ( .C1(n19701), .C2(n19556), .A(n19544), .B(n19543), .ZN(
        P3_U2935) );
  AOI22_X1 U22719 ( .A1(n19745), .A2(n19549), .B1(n19744), .B2(n19552), .ZN(
        n19546) );
  AOI22_X1 U22720 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19553), .B1(
        n19746), .B2(n19625), .ZN(n19545) );
  OAI211_X1 U22721 ( .C1(n19749), .C2(n19574), .A(n19546), .B(n19545), .ZN(
        P3_U2936) );
  AOI22_X1 U22722 ( .A1(n19751), .A2(n19552), .B1(n19750), .B2(n19549), .ZN(
        n19548) );
  AOI22_X1 U22723 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19553), .B1(
        n19752), .B2(n19625), .ZN(n19547) );
  OAI211_X1 U22724 ( .C1(n19755), .C2(n19574), .A(n19548), .B(n19547), .ZN(
        P3_U2937) );
  AOI22_X1 U22725 ( .A1(n19756), .A2(n19552), .B1(n19620), .B2(n19549), .ZN(
        n19551) );
  AOI22_X1 U22726 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19553), .B1(
        n19759), .B2(n19625), .ZN(n19550) );
  OAI211_X1 U22727 ( .C1(n19623), .C2(n19574), .A(n19551), .B(n19550), .ZN(
        P3_U2938) );
  AOI22_X1 U22728 ( .A1(n19765), .A2(n19552), .B1(n19648), .B2(n19576), .ZN(
        n19555) );
  AOI22_X1 U22729 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19553), .B1(
        n19768), .B2(n19625), .ZN(n19554) );
  OAI211_X1 U22730 ( .C1(n19654), .C2(n19556), .A(n19555), .B(n19554), .ZN(
        P3_U2939) );
  NOR2_X1 U22731 ( .A1(n19603), .A2(n19655), .ZN(n19575) );
  AOI22_X1 U22732 ( .A1(n19719), .A2(n19576), .B1(n19718), .B2(n19575), .ZN(
        n19561) );
  INV_X1 U22733 ( .A(n19557), .ZN(n19558) );
  AOI22_X1 U22734 ( .A1(n19659), .A2(n19558), .B1(n19604), .B2(n19657), .ZN(
        n19577) );
  NOR2_X2 U22735 ( .A1(n19603), .A2(n19559), .ZN(n19643) );
  AOI22_X1 U22736 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19577), .B1(
        n19722), .B2(n19643), .ZN(n19560) );
  OAI211_X1 U22737 ( .C1(n19725), .C2(n19597), .A(n19561), .B(n19560), .ZN(
        P3_U2940) );
  AOI22_X1 U22738 ( .A1(n19690), .A2(n19599), .B1(n19726), .B2(n19575), .ZN(
        n19563) );
  AOI22_X1 U22739 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19577), .B1(
        n19728), .B2(n19643), .ZN(n19562) );
  OAI211_X1 U22740 ( .C1(n19693), .C2(n19574), .A(n19563), .B(n19562), .ZN(
        P3_U2941) );
  AOI22_X1 U22741 ( .A1(n19733), .A2(n19575), .B1(n19732), .B2(n19576), .ZN(
        n19565) );
  AOI22_X1 U22742 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19577), .B1(
        n19734), .B2(n19643), .ZN(n19564) );
  OAI211_X1 U22743 ( .C1(n19737), .C2(n19597), .A(n19565), .B(n19564), .ZN(
        P3_U2942) );
  AOI22_X1 U22744 ( .A1(n19698), .A2(n19599), .B1(n19739), .B2(n19575), .ZN(
        n19567) );
  AOI22_X1 U22745 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19577), .B1(
        n19740), .B2(n19643), .ZN(n19566) );
  OAI211_X1 U22746 ( .C1(n19701), .C2(n19574), .A(n19567), .B(n19566), .ZN(
        P3_U2943) );
  AOI22_X1 U22747 ( .A1(n19745), .A2(n19576), .B1(n19744), .B2(n19575), .ZN(
        n19569) );
  AOI22_X1 U22748 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19577), .B1(
        n19746), .B2(n19643), .ZN(n19568) );
  OAI211_X1 U22749 ( .C1(n19749), .C2(n19597), .A(n19569), .B(n19568), .ZN(
        P3_U2944) );
  AOI22_X1 U22750 ( .A1(n19751), .A2(n19575), .B1(n19750), .B2(n19576), .ZN(
        n19571) );
  AOI22_X1 U22751 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19577), .B1(
        n19752), .B2(n19643), .ZN(n19570) );
  OAI211_X1 U22752 ( .C1(n19755), .C2(n19597), .A(n19571), .B(n19570), .ZN(
        P3_U2945) );
  AOI22_X1 U22753 ( .A1(n19757), .A2(n19599), .B1(n19756), .B2(n19575), .ZN(
        n19573) );
  AOI22_X1 U22754 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19577), .B1(
        n19759), .B2(n19643), .ZN(n19572) );
  OAI211_X1 U22755 ( .C1(n19763), .C2(n19574), .A(n19573), .B(n19572), .ZN(
        P3_U2946) );
  AOI22_X1 U22756 ( .A1(n19767), .A2(n19576), .B1(n19765), .B2(n19575), .ZN(
        n19579) );
  AOI22_X1 U22757 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19577), .B1(
        n19768), .B2(n19643), .ZN(n19578) );
  OAI211_X1 U22758 ( .C1(n19773), .C2(n19597), .A(n19579), .B(n19578), .ZN(
        P3_U2947) );
  NOR2_X2 U22759 ( .A1(n19603), .A2(n19580), .ZN(n19676) );
  NOR2_X1 U22760 ( .A1(n19643), .A2(n19676), .ZN(n19630) );
  NOR2_X1 U22761 ( .A1(n19839), .A2(n19630), .ZN(n19598) );
  AOI22_X1 U22762 ( .A1(n19681), .A2(n19625), .B1(n19718), .B2(n19598), .ZN(
        n19584) );
  OAI21_X1 U22763 ( .B1(n19581), .B2(n19629), .A(n19630), .ZN(n19582) );
  OAI211_X1 U22764 ( .C1(n19676), .C2(n19937), .A(n19632), .B(n19582), .ZN(
        n19600) );
  AOI22_X1 U22765 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19600), .B1(
        n19722), .B2(n19676), .ZN(n19583) );
  OAI211_X1 U22766 ( .C1(n19689), .C2(n19597), .A(n19584), .B(n19583), .ZN(
        P3_U2948) );
  INV_X1 U22767 ( .A(n19625), .ZN(n19616) );
  AOI22_X1 U22768 ( .A1(n19727), .A2(n19599), .B1(n19726), .B2(n19598), .ZN(
        n19586) );
  AOI22_X1 U22769 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19600), .B1(
        n19728), .B2(n19676), .ZN(n19585) );
  OAI211_X1 U22770 ( .C1(n19731), .C2(n19616), .A(n19586), .B(n19585), .ZN(
        P3_U2949) );
  AOI22_X1 U22771 ( .A1(n19694), .A2(n19625), .B1(n19733), .B2(n19598), .ZN(
        n19588) );
  AOI22_X1 U22772 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19600), .B1(
        n19734), .B2(n19676), .ZN(n19587) );
  OAI211_X1 U22773 ( .C1(n19697), .C2(n19597), .A(n19588), .B(n19587), .ZN(
        P3_U2950) );
  AOI22_X1 U22774 ( .A1(n19739), .A2(n19598), .B1(n19738), .B2(n19599), .ZN(
        n19590) );
  AOI22_X1 U22775 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19600), .B1(
        n19740), .B2(n19676), .ZN(n19589) );
  OAI211_X1 U22776 ( .C1(n19743), .C2(n19616), .A(n19590), .B(n19589), .ZN(
        P3_U2951) );
  AOI22_X1 U22777 ( .A1(n19745), .A2(n19599), .B1(n19744), .B2(n19598), .ZN(
        n19592) );
  AOI22_X1 U22778 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19600), .B1(
        n19746), .B2(n19676), .ZN(n19591) );
  OAI211_X1 U22779 ( .C1(n19749), .C2(n19616), .A(n19592), .B(n19591), .ZN(
        P3_U2952) );
  AOI22_X1 U22780 ( .A1(n19751), .A2(n19598), .B1(n19750), .B2(n19599), .ZN(
        n19594) );
  AOI22_X1 U22781 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19600), .B1(
        n19752), .B2(n19676), .ZN(n19593) );
  OAI211_X1 U22782 ( .C1(n19755), .C2(n19616), .A(n19594), .B(n19593), .ZN(
        P3_U2953) );
  AOI22_X1 U22783 ( .A1(n19757), .A2(n19625), .B1(n19756), .B2(n19598), .ZN(
        n19596) );
  AOI22_X1 U22784 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19600), .B1(
        n19759), .B2(n19676), .ZN(n19595) );
  OAI211_X1 U22785 ( .C1(n19763), .C2(n19597), .A(n19596), .B(n19595), .ZN(
        P3_U2954) );
  AOI22_X1 U22786 ( .A1(n19767), .A2(n19599), .B1(n19765), .B2(n19598), .ZN(
        n19602) );
  AOI22_X1 U22787 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19600), .B1(
        n19768), .B2(n19676), .ZN(n19601) );
  OAI211_X1 U22788 ( .C1(n19773), .C2(n19616), .A(n19602), .B(n19601), .ZN(
        P3_U2955) );
  NOR2_X1 U22789 ( .A1(n19799), .A2(n19603), .ZN(n19658) );
  AND2_X1 U22790 ( .A1(n19680), .A2(n19658), .ZN(n19624) );
  AOI22_X1 U22791 ( .A1(n19681), .A2(n19643), .B1(n19718), .B2(n19624), .ZN(
        n19606) );
  NAND2_X1 U22792 ( .A1(n19604), .A2(n19720), .ZN(n19626) );
  NAND2_X1 U22793 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19658), .ZN(
        n19710) );
  INV_X1 U22794 ( .A(n19710), .ZN(n19712) );
  AOI22_X1 U22795 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19626), .B1(
        n19722), .B2(n19712), .ZN(n19605) );
  OAI211_X1 U22796 ( .C1(n19689), .C2(n19616), .A(n19606), .B(n19605), .ZN(
        P3_U2956) );
  AOI22_X1 U22797 ( .A1(n19727), .A2(n19625), .B1(n19726), .B2(n19624), .ZN(
        n19608) );
  AOI22_X1 U22798 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19626), .B1(
        n19728), .B2(n19712), .ZN(n19607) );
  OAI211_X1 U22799 ( .C1(n19731), .C2(n19653), .A(n19608), .B(n19607), .ZN(
        P3_U2957) );
  AOI22_X1 U22800 ( .A1(n19694), .A2(n19643), .B1(n19733), .B2(n19624), .ZN(
        n19610) );
  AOI22_X1 U22801 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19626), .B1(
        n19734), .B2(n19712), .ZN(n19609) );
  OAI211_X1 U22802 ( .C1(n19697), .C2(n19616), .A(n19610), .B(n19609), .ZN(
        P3_U2958) );
  AOI22_X1 U22803 ( .A1(n19739), .A2(n19624), .B1(n19738), .B2(n19625), .ZN(
        n19612) );
  AOI22_X1 U22804 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19626), .B1(
        n19740), .B2(n19712), .ZN(n19611) );
  OAI211_X1 U22805 ( .C1(n19743), .C2(n19653), .A(n19612), .B(n19611), .ZN(
        P3_U2959) );
  AOI22_X1 U22806 ( .A1(n19613), .A2(n19643), .B1(n19744), .B2(n19624), .ZN(
        n19615) );
  AOI22_X1 U22807 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19626), .B1(
        n19746), .B2(n19712), .ZN(n19614) );
  OAI211_X1 U22808 ( .C1(n19617), .C2(n19616), .A(n19615), .B(n19614), .ZN(
        P3_U2960) );
  AOI22_X1 U22809 ( .A1(n19751), .A2(n19624), .B1(n19750), .B2(n19625), .ZN(
        n19619) );
  AOI22_X1 U22810 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19626), .B1(
        n19752), .B2(n19712), .ZN(n19618) );
  OAI211_X1 U22811 ( .C1(n19755), .C2(n19653), .A(n19619), .B(n19618), .ZN(
        P3_U2961) );
  AOI22_X1 U22812 ( .A1(n19756), .A2(n19624), .B1(n19620), .B2(n19625), .ZN(
        n19622) );
  AOI22_X1 U22813 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19626), .B1(
        n19759), .B2(n19712), .ZN(n19621) );
  OAI211_X1 U22814 ( .C1(n19623), .C2(n19653), .A(n19622), .B(n19621), .ZN(
        P3_U2962) );
  AOI22_X1 U22815 ( .A1(n19767), .A2(n19625), .B1(n19765), .B2(n19624), .ZN(
        n19628) );
  AOI22_X1 U22816 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19626), .B1(
        n19768), .B2(n19712), .ZN(n19627) );
  OAI211_X1 U22817 ( .C1(n19773), .C2(n19653), .A(n19628), .B(n19627), .ZN(
        P3_U2963) );
  INV_X1 U22818 ( .A(n19762), .ZN(n19766) );
  NOR2_X1 U22819 ( .A1(n19712), .A2(n19766), .ZN(n19682) );
  OAI21_X1 U22820 ( .B1(n19630), .B2(n19629), .A(n19682), .ZN(n19631) );
  OAI211_X1 U22821 ( .C1(n19766), .C2(n19937), .A(n19632), .B(n19631), .ZN(
        n19650) );
  NOR2_X1 U22822 ( .A1(n19839), .A2(n19682), .ZN(n19649) );
  AOI22_X1 U22823 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19650), .B1(
        n19718), .B2(n19649), .ZN(n19634) );
  AOI22_X1 U22824 ( .A1(n19681), .A2(n19676), .B1(n19722), .B2(n19766), .ZN(
        n19633) );
  OAI211_X1 U22825 ( .C1(n19689), .C2(n19653), .A(n19634), .B(n19633), .ZN(
        P3_U2964) );
  AOI22_X1 U22826 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19650), .B1(
        n19726), .B2(n19649), .ZN(n19636) );
  AOI22_X1 U22827 ( .A1(n19728), .A2(n19766), .B1(n19690), .B2(n19676), .ZN(
        n19635) );
  OAI211_X1 U22828 ( .C1(n19693), .C2(n19653), .A(n19636), .B(n19635), .ZN(
        P3_U2965) );
  INV_X1 U22829 ( .A(n19676), .ZN(n19674) );
  AOI22_X1 U22830 ( .A1(n19733), .A2(n19649), .B1(n19732), .B2(n19643), .ZN(
        n19638) );
  AOI22_X1 U22831 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19650), .B1(
        n19734), .B2(n19766), .ZN(n19637) );
  OAI211_X1 U22832 ( .C1(n19737), .C2(n19674), .A(n19638), .B(n19637), .ZN(
        P3_U2966) );
  AOI22_X1 U22833 ( .A1(n19739), .A2(n19649), .B1(n19738), .B2(n19643), .ZN(
        n19640) );
  AOI22_X1 U22834 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19650), .B1(
        n19740), .B2(n19766), .ZN(n19639) );
  OAI211_X1 U22835 ( .C1(n19743), .C2(n19674), .A(n19640), .B(n19639), .ZN(
        P3_U2967) );
  AOI22_X1 U22836 ( .A1(n19745), .A2(n19643), .B1(n19744), .B2(n19649), .ZN(
        n19642) );
  AOI22_X1 U22837 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19650), .B1(
        n19746), .B2(n19766), .ZN(n19641) );
  OAI211_X1 U22838 ( .C1(n19749), .C2(n19674), .A(n19642), .B(n19641), .ZN(
        P3_U2968) );
  AOI22_X1 U22839 ( .A1(n19751), .A2(n19649), .B1(n19750), .B2(n19643), .ZN(
        n19645) );
  AOI22_X1 U22840 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19650), .B1(
        n19752), .B2(n19766), .ZN(n19644) );
  OAI211_X1 U22841 ( .C1(n19755), .C2(n19674), .A(n19645), .B(n19644), .ZN(
        P3_U2969) );
  AOI22_X1 U22842 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19650), .B1(
        n19756), .B2(n19649), .ZN(n19647) );
  AOI22_X1 U22843 ( .A1(n19757), .A2(n19676), .B1(n19759), .B2(n19766), .ZN(
        n19646) );
  OAI211_X1 U22844 ( .C1(n19763), .C2(n19653), .A(n19647), .B(n19646), .ZN(
        P3_U2970) );
  AOI22_X1 U22845 ( .A1(n19765), .A2(n19649), .B1(n19648), .B2(n19676), .ZN(
        n19652) );
  AOI22_X1 U22846 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19650), .B1(
        n19768), .B2(n19766), .ZN(n19651) );
  OAI211_X1 U22847 ( .C1(n19654), .C2(n19653), .A(n19652), .B(n19651), .ZN(
        P3_U2971) );
  NOR2_X1 U22848 ( .A1(n19656), .A2(n19655), .ZN(n19675) );
  AOI22_X1 U22849 ( .A1(n19681), .A2(n19712), .B1(n19718), .B2(n19675), .ZN(
        n19661) );
  AOI22_X1 U22850 ( .A1(n19659), .A2(n19658), .B1(n19721), .B2(n19657), .ZN(
        n19677) );
  AOI22_X1 U22851 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19677), .B1(
        n19758), .B2(n19722), .ZN(n19660) );
  OAI211_X1 U22852 ( .C1(n19689), .C2(n19674), .A(n19661), .B(n19660), .ZN(
        P3_U2972) );
  AOI22_X1 U22853 ( .A1(n19727), .A2(n19676), .B1(n19726), .B2(n19675), .ZN(
        n19663) );
  AOI22_X1 U22854 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19677), .B1(
        n19758), .B2(n19728), .ZN(n19662) );
  OAI211_X1 U22855 ( .C1(n19731), .C2(n19710), .A(n19663), .B(n19662), .ZN(
        P3_U2973) );
  AOI22_X1 U22856 ( .A1(n19733), .A2(n19675), .B1(n19732), .B2(n19676), .ZN(
        n19665) );
  AOI22_X1 U22857 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19677), .B1(
        n19758), .B2(n19734), .ZN(n19664) );
  OAI211_X1 U22858 ( .C1(n19737), .C2(n19710), .A(n19665), .B(n19664), .ZN(
        P3_U2974) );
  AOI22_X1 U22859 ( .A1(n19739), .A2(n19675), .B1(n19738), .B2(n19676), .ZN(
        n19667) );
  AOI22_X1 U22860 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19677), .B1(
        n19758), .B2(n19740), .ZN(n19666) );
  OAI211_X1 U22861 ( .C1(n19743), .C2(n19710), .A(n19667), .B(n19666), .ZN(
        P3_U2975) );
  AOI22_X1 U22862 ( .A1(n19745), .A2(n19676), .B1(n19744), .B2(n19675), .ZN(
        n19669) );
  AOI22_X1 U22863 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19677), .B1(
        n19758), .B2(n19746), .ZN(n19668) );
  OAI211_X1 U22864 ( .C1(n19749), .C2(n19710), .A(n19669), .B(n19668), .ZN(
        P3_U2976) );
  AOI22_X1 U22865 ( .A1(n19704), .A2(n19712), .B1(n19751), .B2(n19675), .ZN(
        n19671) );
  AOI22_X1 U22866 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19677), .B1(
        n19758), .B2(n19752), .ZN(n19670) );
  OAI211_X1 U22867 ( .C1(n19707), .C2(n19674), .A(n19671), .B(n19670), .ZN(
        P3_U2977) );
  AOI22_X1 U22868 ( .A1(n19757), .A2(n19712), .B1(n19756), .B2(n19675), .ZN(
        n19673) );
  AOI22_X1 U22869 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19677), .B1(
        n19758), .B2(n19759), .ZN(n19672) );
  OAI211_X1 U22870 ( .C1(n19763), .C2(n19674), .A(n19673), .B(n19672), .ZN(
        P3_U2978) );
  AOI22_X1 U22871 ( .A1(n19767), .A2(n19676), .B1(n19765), .B2(n19675), .ZN(
        n19679) );
  AOI22_X1 U22872 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19677), .B1(
        n19758), .B2(n19768), .ZN(n19678) );
  OAI211_X1 U22873 ( .C1(n19773), .C2(n19710), .A(n19679), .B(n19678), .ZN(
        P3_U2979) );
  AOI22_X1 U22874 ( .A1(n19681), .A2(n19766), .B1(n19718), .B2(n19711), .ZN(
        n19688) );
  INV_X1 U22875 ( .A(n19682), .ZN(n19684) );
  OAI221_X1 U22876 ( .B1(n19686), .B2(n19685), .C1(n19686), .C2(n19684), .A(
        n19683), .ZN(n19714) );
  AOI22_X1 U22877 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19722), .ZN(n19687) );
  OAI211_X1 U22878 ( .C1(n19689), .C2(n19710), .A(n19688), .B(n19687), .ZN(
        P3_U2980) );
  AOI22_X1 U22879 ( .A1(n19690), .A2(n19766), .B1(n19726), .B2(n19711), .ZN(
        n19692) );
  AOI22_X1 U22880 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19728), .ZN(n19691) );
  OAI211_X1 U22881 ( .C1(n19693), .C2(n19710), .A(n19692), .B(n19691), .ZN(
        P3_U2981) );
  AOI22_X1 U22882 ( .A1(n19694), .A2(n19766), .B1(n19733), .B2(n19711), .ZN(
        n19696) );
  AOI22_X1 U22883 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19734), .ZN(n19695) );
  OAI211_X1 U22884 ( .C1(n19697), .C2(n19710), .A(n19696), .B(n19695), .ZN(
        P3_U2982) );
  AOI22_X1 U22885 ( .A1(n19698), .A2(n19766), .B1(n19739), .B2(n19711), .ZN(
        n19700) );
  AOI22_X1 U22886 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19740), .ZN(n19699) );
  OAI211_X1 U22887 ( .C1(n19701), .C2(n19710), .A(n19700), .B(n19699), .ZN(
        P3_U2983) );
  AOI22_X1 U22888 ( .A1(n19745), .A2(n19712), .B1(n19744), .B2(n19711), .ZN(
        n19703) );
  AOI22_X1 U22889 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19746), .ZN(n19702) );
  OAI211_X1 U22890 ( .C1(n19749), .C2(n19762), .A(n19703), .B(n19702), .ZN(
        P3_U2984) );
  AOI22_X1 U22891 ( .A1(n19704), .A2(n19766), .B1(n19751), .B2(n19711), .ZN(
        n19706) );
  AOI22_X1 U22892 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19752), .ZN(n19705) );
  OAI211_X1 U22893 ( .C1(n19707), .C2(n19710), .A(n19706), .B(n19705), .ZN(
        P3_U2985) );
  AOI22_X1 U22894 ( .A1(n19757), .A2(n19766), .B1(n19756), .B2(n19711), .ZN(
        n19709) );
  AOI22_X1 U22895 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19759), .ZN(n19708) );
  OAI211_X1 U22896 ( .C1(n19763), .C2(n19710), .A(n19709), .B(n19708), .ZN(
        P3_U2986) );
  AOI22_X1 U22897 ( .A1(n19767), .A2(n19712), .B1(n19765), .B2(n19711), .ZN(
        n19716) );
  AOI22_X1 U22898 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19714), .B1(
        n19713), .B2(n19768), .ZN(n19715) );
  OAI211_X1 U22899 ( .C1(n19773), .C2(n19762), .A(n19716), .B(n19715), .ZN(
        P3_U2987) );
  NOR2_X1 U22900 ( .A1(n19839), .A2(n19717), .ZN(n19764) );
  AOI22_X1 U22901 ( .A1(n19719), .A2(n19766), .B1(n19718), .B2(n19764), .ZN(
        n19724) );
  NAND2_X1 U22902 ( .A1(n19721), .A2(n19720), .ZN(n19770) );
  AOI22_X1 U22903 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19722), .ZN(n19723) );
  OAI211_X1 U22904 ( .C1(n19725), .C2(n19774), .A(n19724), .B(n19723), .ZN(
        P3_U2988) );
  AOI22_X1 U22905 ( .A1(n19727), .A2(n19766), .B1(n19726), .B2(n19764), .ZN(
        n19730) );
  AOI22_X1 U22906 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19728), .ZN(n19729) );
  OAI211_X1 U22907 ( .C1(n19774), .C2(n19731), .A(n19730), .B(n19729), .ZN(
        P3_U2989) );
  AOI22_X1 U22908 ( .A1(n19733), .A2(n19764), .B1(n19732), .B2(n19766), .ZN(
        n19736) );
  AOI22_X1 U22909 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19734), .ZN(n19735) );
  OAI211_X1 U22910 ( .C1(n19774), .C2(n19737), .A(n19736), .B(n19735), .ZN(
        P3_U2990) );
  AOI22_X1 U22911 ( .A1(n19739), .A2(n19764), .B1(n19738), .B2(n19766), .ZN(
        n19742) );
  AOI22_X1 U22912 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19740), .ZN(n19741) );
  OAI211_X1 U22913 ( .C1(n19774), .C2(n19743), .A(n19742), .B(n19741), .ZN(
        P3_U2991) );
  AOI22_X1 U22914 ( .A1(n19745), .A2(n19766), .B1(n19744), .B2(n19764), .ZN(
        n19748) );
  AOI22_X1 U22915 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19746), .ZN(n19747) );
  OAI211_X1 U22916 ( .C1(n19774), .C2(n19749), .A(n19748), .B(n19747), .ZN(
        P3_U2992) );
  AOI22_X1 U22917 ( .A1(n19751), .A2(n19764), .B1(n19750), .B2(n19766), .ZN(
        n19754) );
  AOI22_X1 U22918 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19752), .ZN(n19753) );
  OAI211_X1 U22919 ( .C1(n19774), .C2(n19755), .A(n19754), .B(n19753), .ZN(
        P3_U2993) );
  AOI22_X1 U22920 ( .A1(n19758), .A2(n19757), .B1(n19756), .B2(n19764), .ZN(
        n19761) );
  AOI22_X1 U22921 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19759), .ZN(n19760) );
  OAI211_X1 U22922 ( .C1(n19763), .C2(n19762), .A(n19761), .B(n19760), .ZN(
        P3_U2994) );
  AOI22_X1 U22923 ( .A1(n19767), .A2(n19766), .B1(n19765), .B2(n19764), .ZN(
        n19772) );
  AOI22_X1 U22924 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19768), .ZN(n19771) );
  OAI211_X1 U22925 ( .C1(n19774), .C2(n19773), .A(n19772), .B(n19771), .ZN(
        P3_U2995) );
  OAI21_X1 U22926 ( .B1(n19775), .B2(n19967), .A(n19794), .ZN(n19785) );
  AOI22_X1 U22927 ( .A1(n19812), .A2(n19776), .B1(n19786), .B2(n19785), .ZN(
        n19938) );
  NOR2_X1 U22928 ( .A1(n19802), .A2(n19938), .ZN(n19784) );
  INV_X1 U22929 ( .A(n19777), .ZN(n19781) );
  AOI21_X1 U22930 ( .B1(n19780), .B2(n19779), .A(n19778), .ZN(n19788) );
  OAI22_X1 U22931 ( .A1(n19794), .A2(n19786), .B1(n19781), .B2(n19788), .ZN(
        n19782) );
  AOI21_X1 U22932 ( .B1(n19787), .B2(n19953), .A(n19782), .ZN(n19941) );
  NAND2_X1 U22933 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19941), .ZN(
        n19783) );
  OAI22_X1 U22934 ( .A1(n19784), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19802), .B2(n19783), .ZN(n19807) );
  INV_X1 U22935 ( .A(n19785), .ZN(n19795) );
  AOI211_X1 U22936 ( .C1(n19961), .C2(n19953), .A(n19786), .B(n19795), .ZN(
        n19791) );
  INV_X1 U22937 ( .A(n19787), .ZN(n19789) );
  NOR3_X1 U22938 ( .A1(n19789), .A2(n19788), .A3(n19953), .ZN(n19790) );
  AOI211_X1 U22939 ( .C1(n19812), .C2(n19947), .A(n19791), .B(n19790), .ZN(
        n19950) );
  AOI22_X1 U22940 ( .A1(n19802), .A2(n19953), .B1(n19950), .B2(n19823), .ZN(
        n19804) );
  OAI22_X1 U22941 ( .A1(n19796), .A2(n19954), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19795), .ZN(n19959) );
  OR3_X1 U22942 ( .A1(n19963), .A2(n19799), .A3(n19797), .ZN(n19798) );
  AOI22_X1 U22943 ( .A1(n19963), .A2(n19799), .B1(n19959), .B2(n19798), .ZN(
        n19801) );
  INV_X1 U22944 ( .A(n19804), .ZN(n19809) );
  NAND2_X1 U22945 ( .A1(n19806), .A2(n19805), .ZN(n19808) );
  AOI21_X1 U22946 ( .B1(n19809), .B2(n19808), .A(n19807), .ZN(n19826) );
  INV_X1 U22947 ( .A(n19810), .ZN(n19818) );
  NOR2_X1 U22948 ( .A1(n19812), .A2(n19811), .ZN(n19815) );
  OAI222_X1 U22949 ( .A1(n19818), .A2(n19817), .B1(n19816), .B2(n19815), .C1(
        n19814), .C2(n19813), .ZN(n19980) );
  AOI221_X1 U22950 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n19820), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n19820), .A(n19819), .ZN(n19821) );
  OAI211_X1 U22951 ( .C1(n19824), .C2(n19823), .A(n19822), .B(n19821), .ZN(
        n19825) );
  AOI22_X1 U22952 ( .A1(n19962), .A2(n19995), .B1(n19990), .B2(n19982), .ZN(
        n19827) );
  INV_X1 U22953 ( .A(n19827), .ZN(n19832) );
  OAI211_X1 U22954 ( .C1(n19829), .C2(n19828), .A(n19985), .B(n19837), .ZN(
        n19936) );
  NAND2_X1 U22955 ( .A1(n19990), .A2(n20001), .ZN(n19838) );
  NAND2_X1 U22956 ( .A1(n19936), .A2(n19838), .ZN(n19840) );
  NOR2_X1 U22957 ( .A1(n19830), .A2(n19840), .ZN(n19831) );
  MUX2_X1 U22958 ( .A(n19832), .B(n19831), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19835) );
  INV_X1 U22959 ( .A(n19833), .ZN(n19834) );
  OAI211_X1 U22960 ( .C1(n19837), .C2(n19836), .A(n19835), .B(n19834), .ZN(
        P3_U2996) );
  NAND2_X1 U22961 ( .A1(n19990), .A2(n19982), .ZN(n19844) );
  NOR3_X1 U22962 ( .A1(n19946), .A2(n19992), .A3(n19838), .ZN(n19846) );
  INV_X1 U22963 ( .A(n19846), .ZN(n19843) );
  NAND4_X1 U22964 ( .A1(n10977), .A2(n19844), .A3(n19843), .A4(n19842), .ZN(
        P3_U2997) );
  OAI21_X1 U22965 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n19845), .ZN(n19847) );
  AOI21_X1 U22966 ( .B1(n19848), .B2(n19847), .A(n19846), .ZN(P3_U2998) );
  AND2_X1 U22967 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19931), .ZN(
        P3_U2999) );
  AND2_X1 U22968 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19931), .ZN(
        P3_U3000) );
  AND2_X1 U22969 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19931), .ZN(
        P3_U3001) );
  AND2_X1 U22970 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19931), .ZN(
        P3_U3002) );
  AND2_X1 U22971 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19931), .ZN(
        P3_U3003) );
  AND2_X1 U22972 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19931), .ZN(
        P3_U3004) );
  INV_X1 U22973 ( .A(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n21824) );
  NOR2_X1 U22974 ( .A1(n21824), .A2(n19934), .ZN(P3_U3005) );
  AND2_X1 U22975 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19931), .ZN(
        P3_U3006) );
  AND2_X1 U22976 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19931), .ZN(
        P3_U3007) );
  AND2_X1 U22977 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19931), .ZN(
        P3_U3008) );
  AND2_X1 U22978 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19931), .ZN(
        P3_U3009) );
  AND2_X1 U22979 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19931), .ZN(
        P3_U3010) );
  INV_X1 U22980 ( .A(P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21864) );
  NOR2_X1 U22981 ( .A1(n21864), .A2(n19934), .ZN(P3_U3011) );
  AND2_X1 U22982 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19931), .ZN(
        P3_U3012) );
  AND2_X1 U22983 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19931), .ZN(
        P3_U3013) );
  AND2_X1 U22984 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19931), .ZN(
        P3_U3014) );
  AND2_X1 U22985 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19931), .ZN(
        P3_U3015) );
  AND2_X1 U22986 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19931), .ZN(
        P3_U3016) );
  AND2_X1 U22987 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19931), .ZN(
        P3_U3017) );
  AND2_X1 U22988 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19931), .ZN(
        P3_U3018) );
  AND2_X1 U22989 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19931), .ZN(
        P3_U3019) );
  AND2_X1 U22990 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19931), .ZN(
        P3_U3020) );
  AND2_X1 U22991 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19931), .ZN(P3_U3021) );
  AND2_X1 U22992 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19931), .ZN(P3_U3022) );
  AND2_X1 U22993 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19931), .ZN(P3_U3023) );
  AND2_X1 U22994 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19931), .ZN(P3_U3024) );
  AND2_X1 U22995 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19931), .ZN(P3_U3025) );
  INV_X1 U22996 ( .A(P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n21813) );
  NOR2_X1 U22997 ( .A1(n21813), .A2(n19934), .ZN(P3_U3026) );
  AND2_X1 U22998 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19931), .ZN(P3_U3027) );
  AND2_X1 U22999 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19931), .ZN(P3_U3028) );
  OAI21_X1 U23000 ( .B1(n19849), .B2(n20723), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19850) );
  AOI22_X1 U23001 ( .A1(n19861), .A2(n19863), .B1(n19999), .B2(n19850), .ZN(
        n19851) );
  INV_X1 U23002 ( .A(NA), .ZN(n21656) );
  OR3_X1 U23003 ( .A1(n21656), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n19856) );
  OAI211_X1 U23004 ( .C1(n19852), .C2(n19981), .A(n19851), .B(n19856), .ZN(
        P3_U3029) );
  NOR2_X1 U23005 ( .A1(n19863), .A2(n20723), .ZN(n19859) );
  INV_X1 U23006 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19997) );
  OAI22_X1 U23007 ( .A1(n19859), .A2(n19997), .B1(n20723), .B2(n19852), .ZN(
        n19853) );
  AOI22_X1 U23008 ( .A1(n19990), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n19853), .ZN(n19854) );
  NAND2_X1 U23009 ( .A1(n19854), .A2(n19986), .ZN(P3_U3030) );
  NAND2_X1 U23010 ( .A1(n19990), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19857) );
  INV_X1 U23011 ( .A(n19857), .ZN(n19855) );
  AOI21_X1 U23012 ( .B1(n19861), .B2(n19856), .A(n19855), .ZN(n19862) );
  OAI22_X1 U23013 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19857), .ZN(n19858) );
  OAI22_X1 U23014 ( .A1(n19859), .A2(n19858), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19860) );
  OAI22_X1 U23015 ( .A1(n19862), .A2(n19863), .B1(n19861), .B2(n19860), .ZN(
        P3_U3031) );
  NAND2_X2 U23016 ( .A1(n19928), .A2(n19863), .ZN(n19908) );
  OAI222_X1 U23017 ( .A1(n19969), .A2(n19922), .B1(n19864), .B2(n19928), .C1(
        n19865), .C2(n19908), .ZN(P3_U3032) );
  OAI222_X1 U23018 ( .A1(n19908), .A2(n19867), .B1(n19866), .B2(n19928), .C1(
        n19865), .C2(n19922), .ZN(P3_U3033) );
  OAI222_X1 U23019 ( .A1(n19908), .A2(n19869), .B1(n19868), .B2(n19928), .C1(
        n19867), .C2(n19922), .ZN(P3_U3034) );
  OAI222_X1 U23020 ( .A1(n19908), .A2(n19872), .B1(n19870), .B2(n19928), .C1(
        n19869), .C2(n19922), .ZN(P3_U3035) );
  INV_X1 U23021 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19873) );
  OAI222_X1 U23022 ( .A1(n19872), .A2(n19922), .B1(n19871), .B2(n19928), .C1(
        n19873), .C2(n19908), .ZN(P3_U3036) );
  INV_X1 U23023 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19875) );
  OAI222_X1 U23024 ( .A1(n19908), .A2(n19875), .B1(n19874), .B2(n19928), .C1(
        n19873), .C2(n19922), .ZN(P3_U3037) );
  OAI222_X1 U23025 ( .A1(n19908), .A2(n19877), .B1(n19876), .B2(n19928), .C1(
        n19875), .C2(n19922), .ZN(P3_U3038) );
  OAI222_X1 U23026 ( .A1(n19877), .A2(n19922), .B1(n21953), .B2(n19928), .C1(
        n19878), .C2(n19908), .ZN(P3_U3039) );
  OAI222_X1 U23027 ( .A1(n19908), .A2(n19880), .B1(n19879), .B2(n19928), .C1(
        n19878), .C2(n19922), .ZN(P3_U3040) );
  OAI222_X1 U23028 ( .A1(n19908), .A2(n19882), .B1(n19881), .B2(n19928), .C1(
        n19880), .C2(n19922), .ZN(P3_U3041) );
  INV_X1 U23029 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n21826) );
  OAI222_X1 U23030 ( .A1(n19908), .A2(n21826), .B1(n19883), .B2(n19928), .C1(
        n19882), .C2(n19922), .ZN(P3_U3042) );
  OAI222_X1 U23031 ( .A1(n19908), .A2(n19885), .B1(n19884), .B2(n19928), .C1(
        n21826), .C2(n19922), .ZN(P3_U3043) );
  INV_X1 U23032 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19887) );
  OAI222_X1 U23033 ( .A1(n19908), .A2(n19887), .B1(n19886), .B2(n19928), .C1(
        n19885), .C2(n19922), .ZN(P3_U3044) );
  OAI222_X1 U23034 ( .A1(n19908), .A2(n19889), .B1(n19888), .B2(n19928), .C1(
        n19887), .C2(n19922), .ZN(P3_U3045) );
  OAI222_X1 U23035 ( .A1(n19908), .A2(n22035), .B1(n19890), .B2(n19928), .C1(
        n19889), .C2(n19922), .ZN(P3_U3046) );
  INV_X1 U23036 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19892) );
  OAI222_X1 U23037 ( .A1(n22035), .A2(n19922), .B1(n19891), .B2(n19928), .C1(
        n19892), .C2(n19908), .ZN(P3_U3047) );
  OAI222_X1 U23038 ( .A1(n19908), .A2(n19894), .B1(n19893), .B2(n19928), .C1(
        n19892), .C2(n19922), .ZN(P3_U3048) );
  OAI222_X1 U23039 ( .A1(n19908), .A2(n19896), .B1(n19895), .B2(n19928), .C1(
        n19894), .C2(n19922), .ZN(P3_U3049) );
  OAI222_X1 U23040 ( .A1(n19908), .A2(n19898), .B1(n19897), .B2(n19928), .C1(
        n19896), .C2(n19922), .ZN(P3_U3050) );
  OAI222_X1 U23041 ( .A1(n19908), .A2(n19900), .B1(n19899), .B2(n19928), .C1(
        n19898), .C2(n19922), .ZN(P3_U3051) );
  OAI222_X1 U23042 ( .A1(n19908), .A2(n19902), .B1(n19901), .B2(n19928), .C1(
        n19900), .C2(n19922), .ZN(P3_U3052) );
  OAI222_X1 U23043 ( .A1(n19908), .A2(n19904), .B1(n19903), .B2(n19928), .C1(
        n19902), .C2(n19922), .ZN(P3_U3053) );
  OAI222_X1 U23044 ( .A1(n19908), .A2(n19906), .B1(n19905), .B2(n19928), .C1(
        n19904), .C2(n19922), .ZN(P3_U3054) );
  OAI222_X1 U23045 ( .A1(n19908), .A2(n19909), .B1(n19907), .B2(n19928), .C1(
        n19906), .C2(n19922), .ZN(P3_U3055) );
  OAI222_X1 U23046 ( .A1(n19908), .A2(n19911), .B1(n19910), .B2(n19928), .C1(
        n19909), .C2(n19922), .ZN(P3_U3056) );
  OAI222_X1 U23047 ( .A1(n19908), .A2(n19913), .B1(n19912), .B2(n19928), .C1(
        n19911), .C2(n19922), .ZN(P3_U3057) );
  OAI222_X1 U23048 ( .A1(n19908), .A2(n19916), .B1(n19914), .B2(n19928), .C1(
        n19913), .C2(n19922), .ZN(P3_U3058) );
  OAI222_X1 U23049 ( .A1(n19916), .A2(n19922), .B1(n19915), .B2(n19928), .C1(
        n19917), .C2(n19908), .ZN(P3_U3059) );
  OAI222_X1 U23050 ( .A1(n19908), .A2(n19921), .B1(n19918), .B2(n19928), .C1(
        n19917), .C2(n19922), .ZN(P3_U3060) );
  OAI222_X1 U23051 ( .A1(n19922), .A2(n19921), .B1(n19920), .B2(n19928), .C1(
        n19919), .C2(n19908), .ZN(P3_U3061) );
  INV_X1 U23052 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19923) );
  AOI22_X1 U23053 ( .A1(n19928), .A2(n19924), .B1(n19923), .B2(n19999), .ZN(
        P3_U3274) );
  INV_X1 U23054 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19971) );
  INV_X1 U23055 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n21992) );
  AOI22_X1 U23056 ( .A1(n19928), .A2(n19971), .B1(n21992), .B2(n19999), .ZN(
        P3_U3275) );
  INV_X1 U23057 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19925) );
  AOI22_X1 U23058 ( .A1(n19928), .A2(n19926), .B1(n19925), .B2(n19999), .ZN(
        P3_U3276) );
  INV_X1 U23059 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19977) );
  INV_X1 U23060 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19927) );
  AOI22_X1 U23061 ( .A1(n19928), .A2(n19977), .B1(n19927), .B2(n19999), .ZN(
        P3_U3277) );
  INV_X1 U23062 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19930) );
  INV_X1 U23063 ( .A(n19932), .ZN(n19929) );
  AOI21_X1 U23064 ( .B1(n19931), .B2(n19930), .A(n19929), .ZN(P3_U3280) );
  OAI21_X1 U23065 ( .B1(n19934), .B2(n19933), .A(n19932), .ZN(P3_U3281) );
  OAI221_X1 U23066 ( .B1(n19937), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19937), 
        .C2(n19936), .A(n19935), .ZN(P3_U3282) );
  NOR2_X1 U23067 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19938), .ZN(
        n19940) );
  AOI22_X1 U23068 ( .A1(n20002), .A2(n19940), .B1(n19962), .B2(n19939), .ZN(
        n19944) );
  INV_X1 U23069 ( .A(n19941), .ZN(n19942) );
  AOI21_X1 U23070 ( .B1(n20002), .B2(n19942), .A(n19968), .ZN(n19943) );
  OAI22_X1 U23071 ( .A1(n19968), .A2(n19944), .B1(n19943), .B2(n10623), .ZN(
        P3_U3285) );
  AOI22_X1 U23072 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n10622), .B2(n19945), .ZN(
        n19955) );
  NOR2_X1 U23073 ( .A1(n19946), .A2(n19964), .ZN(n19956) );
  INV_X1 U23074 ( .A(n19962), .ZN(n19948) );
  OAI22_X1 U23075 ( .A1(n19950), .A2(n19949), .B1(n19948), .B2(n19947), .ZN(
        n19951) );
  AOI21_X1 U23076 ( .B1(n19955), .B2(n19956), .A(n19951), .ZN(n19952) );
  AOI22_X1 U23077 ( .A1(n19968), .A2(n19953), .B1(n19952), .B2(n19965), .ZN(
        P3_U3288) );
  INV_X1 U23078 ( .A(n19954), .ZN(n19958) );
  INV_X1 U23079 ( .A(n19955), .ZN(n19957) );
  AOI222_X1 U23080 ( .A1(n19959), .A2(n20002), .B1(n19962), .B2(n19958), .C1(
        n19957), .C2(n19956), .ZN(n19960) );
  AOI22_X1 U23081 ( .A1(n19968), .A2(n19961), .B1(n19960), .B2(n19965), .ZN(
        P3_U3289) );
  AOI222_X1 U23082 ( .A1(n19964), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n20002), 
        .B2(n19963), .C1(n19967), .C2(n19962), .ZN(n19966) );
  AOI22_X1 U23083 ( .A1(n19968), .A2(n19967), .B1(n19966), .B2(n19965), .ZN(
        P3_U3290) );
  AOI21_X1 U23084 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19970) );
  AOI22_X1 U23085 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19970), .B2(n19969), .ZN(n19972) );
  AOI22_X1 U23086 ( .A1(n19973), .A2(n19972), .B1(n19971), .B2(n19976), .ZN(
        P3_U3292) );
  NOR2_X1 U23087 ( .A1(n19976), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19974) );
  AOI22_X1 U23088 ( .A1(n19977), .A2(n19976), .B1(n19975), .B2(n19974), .ZN(
        P3_U3293) );
  INV_X1 U23089 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19978) );
  AOI22_X1 U23090 ( .A1(n19928), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19978), 
        .B2(n19999), .ZN(P3_U3294) );
  MUX2_X1 U23091 ( .A(P3_MORE_REG_SCAN_IN), .B(n19980), .S(n19979), .Z(
        P3_U3295) );
  AOI21_X1 U23092 ( .B1(n19982), .B2(n19981), .A(n20004), .ZN(n19983) );
  OAI21_X1 U23093 ( .B1(n19985), .B2(n19984), .A(n19983), .ZN(n19998) );
  AOI21_X1 U23094 ( .B1(n19988), .B2(n19987), .A(n19986), .ZN(n19989) );
  INV_X1 U23095 ( .A(n19989), .ZN(n19991) );
  AOI211_X1 U23096 ( .C1(n20003), .C2(n19991), .A(n19990), .B(n20001), .ZN(
        n19993) );
  NOR2_X1 U23097 ( .A1(n19993), .A2(n19992), .ZN(n19994) );
  OAI21_X1 U23098 ( .B1(n19995), .B2(n19994), .A(n19998), .ZN(n19996) );
  OAI21_X1 U23099 ( .B1(n19998), .B2(n19997), .A(n19996), .ZN(P3_U3296) );
  INV_X1 U23100 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n20006) );
  INV_X1 U23101 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n20000) );
  AOI22_X1 U23102 ( .A1(n19928), .A2(n20006), .B1(n20000), .B2(n19999), .ZN(
        P3_U3297) );
  AOI21_X1 U23103 ( .B1(n20002), .B2(n20001), .A(n20004), .ZN(n20007) );
  INV_X1 U23104 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n21931) );
  AOI22_X1 U23105 ( .A1(n20007), .A2(n21931), .B1(n20004), .B2(n20003), .ZN(
        P3_U3298) );
  AOI21_X1 U23106 ( .B1(n20007), .B2(n20006), .A(n20005), .ZN(P3_U3299) );
  INV_X1 U23107 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n20008) );
  INV_X1 U23108 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20731) );
  NAND2_X1 U23109 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20731), .ZN(n20722) );
  AOI22_X1 U23110 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20722), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n20728), .ZN(n20792) );
  OAI21_X1 U23111 ( .B1(n20728), .B2(n20008), .A(n20715), .ZN(P2_U2815) );
  AOI22_X1 U23112 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20009), .B1(n20847), 
        .B2(P2_CODEFETCH_REG_SCAN_IN), .ZN(n20010) );
  INV_X1 U23113 ( .A(n20010), .ZN(P2_U2816) );
  NAND2_X1 U23114 ( .A1(n20863), .A2(n20011), .ZN(n20718) );
  AOI21_X1 U23115 ( .B1(n20728), .B2(n20718), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n20012) );
  AOI21_X1 U23116 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n20862), .A(n20012), 
        .ZN(P2_U2817) );
  OAI21_X1 U23117 ( .B1(n20725), .B2(BS16), .A(n20792), .ZN(n20791) );
  OAI21_X1 U23118 ( .B1(n20792), .B2(n20481), .A(n20791), .ZN(P2_U2818) );
  NOR4_X1 U23119 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20016) );
  NOR4_X1 U23120 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20015) );
  NOR4_X1 U23121 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20014) );
  NOR4_X1 U23122 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20013) );
  NAND4_X1 U23123 ( .A1(n20016), .A2(n20015), .A3(n20014), .A4(n20013), .ZN(
        n20022) );
  NOR4_X1 U23124 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20020) );
  AOI211_X1 U23125 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_18__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20019) );
  NOR4_X1 U23126 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20018) );
  NOR4_X1 U23127 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20017) );
  NAND4_X1 U23128 ( .A1(n20020), .A2(n20019), .A3(n20018), .A4(n20017), .ZN(
        n20021) );
  NOR2_X1 U23129 ( .A1(n20022), .A2(n20021), .ZN(n20030) );
  INV_X1 U23130 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21816) );
  OAI21_X1 U23131 ( .B1(P2_REIP_REG_0__SCAN_IN), .B2(P2_REIP_REG_1__SCAN_IN), 
        .A(n20030), .ZN(n20023) );
  OAI21_X1 U23132 ( .B1(n20030), .B2(n21816), .A(n20023), .ZN(P2_U2820) );
  INV_X1 U23133 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20788) );
  NOR3_X1 U23134 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20027) );
  OAI21_X1 U23135 ( .B1(P2_REIP_REG_1__SCAN_IN), .B2(n20027), .A(n20030), .ZN(
        n20024) );
  OAI21_X1 U23136 ( .B1(n20030), .B2(n20788), .A(n20024), .ZN(P2_U2821) );
  AOI21_X1 U23137 ( .B1(P2_REIP_REG_0__SCAN_IN), .B2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20025) );
  OAI22_X1 U23138 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(n20732), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n20025), .ZN(n20026) );
  INV_X1 U23139 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20786) );
  INV_X1 U23140 ( .A(n20030), .ZN(n20028) );
  AOI22_X1 U23141 ( .A1(n20030), .A2(n20026), .B1(n20786), .B2(n20028), .ZN(
        P2_U2822) );
  INV_X1 U23142 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21862) );
  AOI21_X1 U23143 ( .B1(n20732), .B2(n21862), .A(n20027), .ZN(n20029) );
  INV_X1 U23144 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20784) );
  AOI22_X1 U23145 ( .A1(n20030), .A2(n20029), .B1(n20784), .B2(n20028), .ZN(
        P2_U2823) );
  AOI22_X1 U23146 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n20032), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20031), .ZN(n20050) );
  AOI21_X1 U23147 ( .B1(n20057), .B2(P2_REIP_REG_15__SCAN_IN), .A(n20033), 
        .ZN(n20034) );
  OAI21_X1 U23148 ( .B1(n20035), .B2(n20053), .A(n20034), .ZN(n20036) );
  AOI21_X1 U23149 ( .B1(n20038), .B2(n20037), .A(n20036), .ZN(n20049) );
  AOI22_X1 U23150 ( .A1(n20042), .A2(n20041), .B1(n20040), .B2(n20039), .ZN(
        n20048) );
  INV_X1 U23151 ( .A(n20043), .ZN(n20046) );
  OAI21_X1 U23152 ( .B1(n20046), .B2(n20045), .A(n20044), .ZN(n20047) );
  NAND4_X1 U23153 ( .A1(n20050), .A2(n20049), .A3(n20048), .A4(n20047), .ZN(
        P2_U2840) );
  OAI21_X1 U23154 ( .B1(n20052), .B2(n21970), .A(n20051), .ZN(n20056) );
  NOR2_X1 U23155 ( .A1(n20054), .A2(n20053), .ZN(n20055) );
  AOI211_X1 U23156 ( .C1(n20057), .C2(P2_REIP_REG_6__SCAN_IN), .A(n20056), .B(
        n20055), .ZN(n20072) );
  NAND2_X1 U23157 ( .A1(n20058), .A2(n20061), .ZN(n20060) );
  MUX2_X1 U23158 ( .A(n20061), .B(n20060), .S(n20059), .Z(n20070) );
  NOR2_X1 U23159 ( .A1(n20063), .A2(n20062), .ZN(n20069) );
  OAI22_X1 U23160 ( .A1(n20067), .A2(n20066), .B1(n20065), .B2(n20064), .ZN(
        n20068) );
  AOI21_X1 U23161 ( .B1(n20070), .B2(n20069), .A(n20068), .ZN(n20071) );
  OAI211_X1 U23162 ( .C1(n10665), .C2(n20073), .A(n20072), .B(n20071), .ZN(
        P2_U2849) );
  INV_X1 U23163 ( .A(n20074), .ZN(n20080) );
  AOI211_X1 U23164 ( .C1(n20078), .C2(n20077), .A(n20076), .B(n20075), .ZN(
        n20079) );
  AOI21_X1 U23165 ( .B1(n20080), .B2(n20082), .A(n20079), .ZN(n20081) );
  OAI21_X1 U23166 ( .B1(n20082), .B2(n11773), .A(n20081), .ZN(P2_U2877) );
  OAI22_X1 U23167 ( .A1(n20086), .A2(n20085), .B1(n20084), .B2(n20083), .ZN(
        n20087) );
  INV_X1 U23168 ( .A(n20087), .ZN(n20092) );
  XNOR2_X1 U23169 ( .A(n20089), .B(n20088), .ZN(n20090) );
  NAND2_X1 U23170 ( .A1(n20090), .A2(n22058), .ZN(n20091) );
  OAI211_X1 U23171 ( .C1(n20163), .C2(n22062), .A(n20092), .B(n20091), .ZN(
        P2_U2915) );
  AOI22_X1 U23172 ( .A1(n22053), .A2(n20828), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n20093), .ZN(n20099) );
  OAI21_X1 U23173 ( .B1(n20096), .B2(n20095), .A(n20094), .ZN(n20097) );
  NAND2_X1 U23174 ( .A1(n20097), .A2(n22058), .ZN(n20098) );
  OAI211_X1 U23175 ( .C1(n20148), .C2(n22062), .A(n20099), .B(n20098), .ZN(
        P2_U2918) );
  NOR2_X1 U23176 ( .A1(n20101), .A2(n20100), .ZN(P2_U2920) );
  AOI22_X1 U23177 ( .A1(n20130), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n20102) );
  OAI21_X1 U23178 ( .B1(n13856), .B2(n20132), .A(n20102), .ZN(P2_U2936) );
  AOI22_X1 U23179 ( .A1(n20130), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n20103) );
  OAI21_X1 U23180 ( .B1(n20104), .B2(n20132), .A(n20103), .ZN(P2_U2937) );
  AOI22_X1 U23181 ( .A1(n20130), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n20105) );
  OAI21_X1 U23182 ( .B1(n20106), .B2(n20132), .A(n20105), .ZN(P2_U2938) );
  AOI22_X1 U23183 ( .A1(n20130), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n20107) );
  OAI21_X1 U23184 ( .B1(n20108), .B2(n20132), .A(n20107), .ZN(P2_U2939) );
  AOI22_X1 U23185 ( .A1(n20130), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n20109) );
  OAI21_X1 U23186 ( .B1(n20110), .B2(n20132), .A(n20109), .ZN(P2_U2940) );
  AOI22_X1 U23187 ( .A1(n20130), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n20111) );
  OAI21_X1 U23188 ( .B1(n20112), .B2(n20132), .A(n20111), .ZN(P2_U2941) );
  AOI22_X1 U23189 ( .A1(n20130), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n20113) );
  OAI21_X1 U23190 ( .B1(n20114), .B2(n20132), .A(n20113), .ZN(P2_U2942) );
  AOI22_X1 U23191 ( .A1(n20130), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_8__SCAN_IN), .ZN(n20115) );
  OAI21_X1 U23192 ( .B1(n20116), .B2(n20132), .A(n20115), .ZN(P2_U2943) );
  AOI22_X1 U23193 ( .A1(n20130), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n20117) );
  OAI21_X1 U23194 ( .B1(n20118), .B2(n20132), .A(n20117), .ZN(P2_U2944) );
  AOI22_X1 U23195 ( .A1(n20130), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n20119) );
  OAI21_X1 U23196 ( .B1(n20120), .B2(n20132), .A(n20119), .ZN(P2_U2945) );
  INV_X1 U23197 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U23198 ( .A1(n20130), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_5__SCAN_IN), .ZN(n20121) );
  OAI21_X1 U23199 ( .B1(n20122), .B2(n20132), .A(n20121), .ZN(P2_U2946) );
  INV_X1 U23200 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n20124) );
  AOI22_X1 U23201 ( .A1(n20130), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_3__SCAN_IN), .ZN(n20123) );
  OAI21_X1 U23202 ( .B1(n20124), .B2(n20132), .A(n20123), .ZN(P2_U2948) );
  INV_X1 U23203 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20126) );
  AOI22_X1 U23204 ( .A1(n20130), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_2__SCAN_IN), .ZN(n20125) );
  OAI21_X1 U23205 ( .B1(n20126), .B2(n20132), .A(n20125), .ZN(P2_U2949) );
  AOI22_X1 U23206 ( .A1(n20130), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_1__SCAN_IN), .ZN(n20127) );
  OAI21_X1 U23207 ( .B1(n20128), .B2(n20132), .A(n20127), .ZN(P2_U2950) );
  AOI22_X1 U23208 ( .A1(n20130), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(n20129), 
        .B2(P2_LWORD_REG_0__SCAN_IN), .ZN(n20131) );
  OAI21_X1 U23209 ( .B1(n13924), .B2(n20132), .A(n20131), .ZN(P2_U2951) );
  AOI22_X1 U23210 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20175), .ZN(n20369) );
  NAND2_X1 U23211 ( .A1(n20812), .A2(n20821), .ZN(n20252) );
  NOR2_X1 U23212 ( .A1(n20416), .A2(n20252), .ZN(n20152) );
  INV_X1 U23213 ( .A(n20152), .ZN(n20182) );
  NAND2_X1 U23214 ( .A1(n20851), .A2(n20180), .ZN(n20257) );
  OAI22_X1 U23215 ( .A1(n20702), .A2(n20665), .B1(n20182), .B2(n20257), .ZN(
        n20135) );
  INV_X1 U23216 ( .A(n20135), .ZN(n20145) );
  AOI21_X1 U23217 ( .B1(n20702), .B2(n20220), .A(n20481), .ZN(n20136) );
  NOR2_X1 U23218 ( .A1(n20136), .A2(n20808), .ZN(n20140) );
  OAI21_X1 U23219 ( .B1(n20141), .B2(n20800), .A(n20814), .ZN(n20137) );
  AOI21_X1 U23220 ( .B1(n20140), .B2(n20657), .A(n20137), .ZN(n20138) );
  NOR2_X2 U23221 ( .A1(n20139), .A2(n20555), .ZN(n20653) );
  INV_X1 U23222 ( .A(n20657), .ZN(n20705) );
  OAI21_X1 U23223 ( .B1(n20705), .B2(n20152), .A(n20140), .ZN(n20143) );
  OAI21_X1 U23224 ( .B1(n20141), .B2(n20152), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20142) );
  AOI22_X1 U23225 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20186), .B1(
        n20653), .B2(n20185), .ZN(n20144) );
  OAI211_X1 U23226 ( .C1(n20369), .C2(n20220), .A(n20145), .B(n20144), .ZN(
        P2_U3048) );
  AOI22_X1 U23227 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20175), .ZN(n20589) );
  OAI22_X1 U23228 ( .A1(n22030), .A2(n20177), .B1(n21059), .B2(n20179), .ZN(
        n20586) );
  NAND2_X1 U23229 ( .A1(n20146), .A2(n20180), .ZN(n20267) );
  OAI22_X1 U23230 ( .A1(n20702), .A2(n20671), .B1(n20182), .B2(n20267), .ZN(
        n20147) );
  INV_X1 U23231 ( .A(n20147), .ZN(n20150) );
  NOR2_X2 U23232 ( .A1(n20148), .A2(n20555), .ZN(n20667) );
  AOI22_X1 U23233 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20186), .B1(
        n20667), .B2(n20185), .ZN(n20149) );
  OAI211_X1 U23234 ( .C1(n20589), .C2(n20220), .A(n20150), .B(n20149), .ZN(
        P2_U3049) );
  AOI22_X1 U23235 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20175), .ZN(n20677) );
  OAI22_X1 U23236 ( .A1(n21068), .A2(n20179), .B1(n21883), .B2(n20177), .ZN(
        n20674) );
  NOR2_X2 U23237 ( .A1(n11078), .A2(n20151), .ZN(n20672) );
  AOI22_X1 U23238 ( .A1(n20709), .A2(n20674), .B1(n20152), .B2(n20672), .ZN(
        n20155) );
  NOR2_X2 U23239 ( .A1(n20153), .A2(n20555), .ZN(n20673) );
  AOI22_X1 U23240 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20186), .B1(
        n20673), .B2(n20185), .ZN(n20154) );
  OAI211_X1 U23241 ( .C1(n20677), .C2(n20220), .A(n20155), .B(n20154), .ZN(
        P2_U3050) );
  AOI22_X1 U23242 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20175), .ZN(n20595) );
  AOI22_X1 U23243 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20175), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20176), .ZN(n20683) );
  NAND2_X1 U23244 ( .A1(n20156), .A2(n20180), .ZN(n20274) );
  OAI22_X1 U23245 ( .A1(n20702), .A2(n20683), .B1(n20182), .B2(n20274), .ZN(
        n20157) );
  INV_X1 U23246 ( .A(n20157), .ZN(n20159) );
  NOR2_X2 U23247 ( .A1(n22063), .A2(n20555), .ZN(n20679) );
  AOI22_X1 U23248 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20186), .B1(
        n20679), .B2(n20185), .ZN(n20158) );
  OAI211_X1 U23249 ( .C1(n20595), .C2(n20220), .A(n20159), .B(n20158), .ZN(
        P2_U3051) );
  AOI22_X1 U23250 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20175), .ZN(n20689) );
  OAI22_X1 U23251 ( .A1(n20160), .A2(n20177), .B1(n21082), .B2(n20179), .ZN(
        n20686) );
  NAND2_X1 U23252 ( .A1(n20161), .A2(n20180), .ZN(n20629) );
  OAI22_X1 U23253 ( .A1(n20702), .A2(n20630), .B1(n20182), .B2(n20629), .ZN(
        n20162) );
  INV_X1 U23254 ( .A(n20162), .ZN(n20165) );
  NOR2_X2 U23255 ( .A1(n20163), .A2(n20555), .ZN(n20685) );
  AOI22_X1 U23256 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20186), .B1(
        n20685), .B2(n20185), .ZN(n20164) );
  OAI211_X1 U23257 ( .C1(n20689), .C2(n20220), .A(n20165), .B(n20164), .ZN(
        P2_U3052) );
  AOI22_X1 U23258 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20175), .ZN(n20601) );
  AOI22_X1 U23259 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20175), .ZN(n20695) );
  NAND2_X1 U23260 ( .A1(n20166), .A2(n20180), .ZN(n20210) );
  OAI22_X1 U23261 ( .A1(n20702), .A2(n20695), .B1(n20182), .B2(n20210), .ZN(
        n20167) );
  INV_X1 U23262 ( .A(n20167), .ZN(n20171) );
  INV_X1 U23263 ( .A(n20168), .ZN(n20169) );
  NOR2_X2 U23264 ( .A1(n20169), .A2(n20555), .ZN(n20691) );
  AOI22_X1 U23265 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20186), .B1(
        n20691), .B2(n20185), .ZN(n20170) );
  OAI211_X1 U23266 ( .C1(n20601), .C2(n20220), .A(n20171), .B(n20170), .ZN(
        P2_U3053) );
  INV_X1 U23267 ( .A(n20696), .ZN(n20637) );
  OAI22_X1 U23268 ( .A1(n20702), .A2(n20638), .B1(n20637), .B2(n20182), .ZN(
        n20172) );
  INV_X1 U23269 ( .A(n20172), .ZN(n20174) );
  AOI22_X1 U23270 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20186), .B1(
        n20697), .B2(n20185), .ZN(n20173) );
  OAI211_X1 U23271 ( .C1(n20703), .C2(n20220), .A(n20174), .B(n20173), .ZN(
        P2_U3054) );
  AOI22_X1 U23272 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20176), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20175), .ZN(n20650) );
  OAI22_X1 U23273 ( .A1(n21103), .A2(n20179), .B1(n20178), .B2(n20177), .ZN(
        n20603) );
  INV_X1 U23274 ( .A(n20603), .ZN(n20714) );
  NAND2_X1 U23275 ( .A1(n20181), .A2(n20180), .ZN(n20643) );
  OAI22_X1 U23276 ( .A1(n20702), .A2(n20714), .B1(n20182), .B2(n20643), .ZN(
        n20183) );
  INV_X1 U23277 ( .A(n20183), .ZN(n20188) );
  NOR2_X2 U23278 ( .A1(n20184), .A2(n20555), .ZN(n20706) );
  AOI22_X1 U23279 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20186), .B1(
        n20706), .B2(n20185), .ZN(n20187) );
  OAI211_X1 U23280 ( .C1(n20650), .C2(n20220), .A(n20188), .B(n20187), .ZN(
        P2_U3055) );
  INV_X1 U23281 ( .A(n20252), .ZN(n20250) );
  NAND2_X1 U23282 ( .A1(n20250), .A2(n20831), .ZN(n20193) );
  INV_X1 U23283 ( .A(n20193), .ZN(n20189) );
  NAND2_X1 U23284 ( .A1(n20189), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20194) );
  INV_X1 U23285 ( .A(n20194), .ZN(n20215) );
  OAI21_X1 U23286 ( .B1(n20190), .B2(n20215), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20191) );
  AOI22_X1 U23287 ( .A1(n20216), .A2(n20653), .B1(n20652), .B2(n20215), .ZN(
        n20201) );
  NAND2_X1 U23288 ( .A1(n20199), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20392) );
  OAI21_X1 U23289 ( .B1(n20392), .B2(n20450), .A(n20193), .ZN(n20197) );
  OAI211_X1 U23290 ( .C1(n20195), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20194), 
        .B(n20808), .ZN(n20196) );
  NAND3_X1 U23291 ( .A1(n20197), .A2(n20660), .A3(n20196), .ZN(n20217) );
  AOI22_X1 U23292 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20217), .B1(
        n20246), .B2(n20662), .ZN(n20200) );
  OAI211_X1 U23293 ( .C1(n20665), .C2(n20220), .A(n20201), .B(n20200), .ZN(
        P2_U3056) );
  INV_X1 U23294 ( .A(n20267), .ZN(n20666) );
  AOI22_X1 U23295 ( .A1(n20216), .A2(n20667), .B1(n20666), .B2(n20215), .ZN(
        n20203) );
  INV_X1 U23296 ( .A(n20589), .ZN(n20668) );
  AOI22_X1 U23297 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20217), .B1(
        n20246), .B2(n20668), .ZN(n20202) );
  OAI211_X1 U23298 ( .C1(n20671), .C2(n20220), .A(n20203), .B(n20202), .ZN(
        P2_U3057) );
  AOI22_X1 U23299 ( .A1(n20216), .A2(n20673), .B1(n20672), .B2(n20215), .ZN(
        n20205) );
  INV_X1 U23300 ( .A(n20677), .ZN(n20623) );
  AOI22_X1 U23301 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20217), .B1(
        n20246), .B2(n20623), .ZN(n20204) );
  OAI211_X1 U23302 ( .C1(n20626), .C2(n20220), .A(n20205), .B(n20204), .ZN(
        P2_U3058) );
  INV_X1 U23303 ( .A(n20274), .ZN(n20678) );
  AOI22_X1 U23304 ( .A1(n20216), .A2(n20679), .B1(n20678), .B2(n20215), .ZN(
        n20207) );
  INV_X1 U23305 ( .A(n20595), .ZN(n20680) );
  AOI22_X1 U23306 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20217), .B1(
        n20246), .B2(n20680), .ZN(n20206) );
  OAI211_X1 U23307 ( .C1(n20683), .C2(n20220), .A(n20207), .B(n20206), .ZN(
        P2_U3059) );
  AOI22_X1 U23308 ( .A1(n20216), .A2(n20685), .B1(n20684), .B2(n20215), .ZN(
        n20209) );
  INV_X1 U23309 ( .A(n20689), .ZN(n20567) );
  AOI22_X1 U23310 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20217), .B1(
        n20246), .B2(n20567), .ZN(n20208) );
  OAI211_X1 U23311 ( .C1(n20630), .C2(n20220), .A(n20209), .B(n20208), .ZN(
        P2_U3060) );
  INV_X1 U23312 ( .A(n20210), .ZN(n20690) );
  AOI22_X1 U23313 ( .A1(n20216), .A2(n20691), .B1(n20690), .B2(n20215), .ZN(
        n20212) );
  INV_X1 U23314 ( .A(n20601), .ZN(n20692) );
  AOI22_X1 U23315 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20217), .B1(
        n20246), .B2(n20692), .ZN(n20211) );
  OAI211_X1 U23316 ( .C1(n20695), .C2(n20220), .A(n20212), .B(n20211), .ZN(
        P2_U3061) );
  AOI22_X1 U23317 ( .A1(n20216), .A2(n20697), .B1(n20696), .B2(n20215), .ZN(
        n20214) );
  AOI22_X1 U23318 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20217), .B1(
        n20246), .B2(n20572), .ZN(n20213) );
  OAI211_X1 U23319 ( .C1(n20638), .C2(n20220), .A(n20214), .B(n20213), .ZN(
        P2_U3062) );
  INV_X1 U23320 ( .A(n20643), .ZN(n20704) );
  AOI22_X1 U23321 ( .A1(n20216), .A2(n20706), .B1(n20704), .B2(n20215), .ZN(
        n20219) );
  INV_X1 U23322 ( .A(n20650), .ZN(n20708) );
  AOI22_X1 U23323 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20217), .B1(
        n20246), .B2(n20708), .ZN(n20218) );
  OAI211_X1 U23324 ( .C1(n20714), .C2(n20220), .A(n20219), .B(n20218), .ZN(
        P2_U3063) );
  NAND2_X1 U23325 ( .A1(n20296), .A2(n20250), .ZN(n20225) );
  NOR3_X2 U23326 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20831), .A3(
        n20252), .ZN(n20244) );
  OAI21_X1 U23327 ( .B1(n20221), .B2(n20244), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20222) );
  AOI22_X1 U23328 ( .A1(n20245), .A2(n20653), .B1(n20652), .B2(n20244), .ZN(
        n20231) );
  INV_X1 U23329 ( .A(n20287), .ZN(n20223) );
  OAI21_X1 U23330 ( .B1(n20223), .B2(n20246), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20224) );
  NAND2_X1 U23331 ( .A1(n20225), .A2(n20224), .ZN(n20229) );
  INV_X1 U23332 ( .A(n20244), .ZN(n20226) );
  OAI211_X1 U23333 ( .C1(n20227), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20226), 
        .B(n20808), .ZN(n20228) );
  NAND3_X1 U23334 ( .A1(n20229), .A2(n20660), .A3(n20228), .ZN(n20247) );
  INV_X1 U23335 ( .A(n20665), .ZN(n20582) );
  AOI22_X1 U23336 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20247), .B1(
        n20246), .B2(n20582), .ZN(n20230) );
  OAI211_X1 U23337 ( .C1(n20369), .C2(n20287), .A(n20231), .B(n20230), .ZN(
        P2_U3064) );
  AOI22_X1 U23338 ( .A1(n20245), .A2(n20667), .B1(n20666), .B2(n20244), .ZN(
        n20233) );
  AOI22_X1 U23339 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20247), .B1(
        n20246), .B2(n20586), .ZN(n20232) );
  OAI211_X1 U23340 ( .C1(n20589), .C2(n20287), .A(n20233), .B(n20232), .ZN(
        P2_U3065) );
  AOI22_X1 U23341 ( .A1(n20245), .A2(n20673), .B1(n20672), .B2(n20244), .ZN(
        n20235) );
  AOI22_X1 U23342 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20247), .B1(
        n20246), .B2(n20674), .ZN(n20234) );
  OAI211_X1 U23343 ( .C1(n20677), .C2(n20287), .A(n20235), .B(n20234), .ZN(
        P2_U3066) );
  AOI22_X1 U23344 ( .A1(n20245), .A2(n20679), .B1(n20678), .B2(n20244), .ZN(
        n20237) );
  INV_X1 U23345 ( .A(n20683), .ZN(n20592) );
  AOI22_X1 U23346 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20247), .B1(
        n20246), .B2(n20592), .ZN(n20236) );
  OAI211_X1 U23347 ( .C1(n20595), .C2(n20287), .A(n20237), .B(n20236), .ZN(
        P2_U3067) );
  AOI22_X1 U23348 ( .A1(n20245), .A2(n20685), .B1(n20684), .B2(n20244), .ZN(
        n20239) );
  AOI22_X1 U23349 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20247), .B1(
        n20246), .B2(n20686), .ZN(n20238) );
  OAI211_X1 U23350 ( .C1(n20689), .C2(n20287), .A(n20239), .B(n20238), .ZN(
        P2_U3068) );
  AOI22_X1 U23351 ( .A1(n20245), .A2(n20691), .B1(n20690), .B2(n20244), .ZN(
        n20241) );
  INV_X1 U23352 ( .A(n20695), .ZN(n20598) );
  AOI22_X1 U23353 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20247), .B1(
        n20246), .B2(n20598), .ZN(n20240) );
  OAI211_X1 U23354 ( .C1(n20601), .C2(n20287), .A(n20241), .B(n20240), .ZN(
        P2_U3069) );
  AOI22_X1 U23355 ( .A1(n20245), .A2(n20697), .B1(n20696), .B2(n20244), .ZN(
        n20243) );
  AOI22_X1 U23356 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20247), .B1(
        n20246), .B2(n20698), .ZN(n20242) );
  OAI211_X1 U23357 ( .C1(n20703), .C2(n20287), .A(n20243), .B(n20242), .ZN(
        P2_U3070) );
  AOI22_X1 U23358 ( .A1(n20245), .A2(n20706), .B1(n20704), .B2(n20244), .ZN(
        n20249) );
  AOI22_X1 U23359 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20247), .B1(
        n20246), .B2(n20603), .ZN(n20248) );
  OAI211_X1 U23360 ( .C1(n20650), .C2(n20287), .A(n20249), .B(n20248), .ZN(
        P2_U3071) );
  OR2_X1 U23361 ( .A1(n20392), .A2(n20264), .ZN(n20251) );
  NAND2_X1 U23362 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20250), .ZN(
        n20260) );
  NAND2_X1 U23363 ( .A1(n20251), .A2(n20260), .ZN(n20256) );
  OAI21_X1 U23364 ( .B1(n20259), .B2(n17300), .A(n20814), .ZN(n20254) );
  NOR2_X1 U23365 ( .A1(n20253), .A2(n20252), .ZN(n20283) );
  INV_X1 U23366 ( .A(n20283), .ZN(n20286) );
  AOI21_X1 U23367 ( .B1(n20254), .B2(n20286), .A(n20555), .ZN(n20255) );
  OAI22_X1 U23368 ( .A1(n20287), .A2(n20665), .B1(n20286), .B2(n20257), .ZN(
        n20258) );
  INV_X1 U23369 ( .A(n20258), .ZN(n20266) );
  NOR2_X1 U23370 ( .A1(n20259), .A2(n20283), .ZN(n20263) );
  INV_X1 U23371 ( .A(n20260), .ZN(n20261) );
  NAND2_X1 U23372 ( .A1(n20261), .A2(n20800), .ZN(n20262) );
  AOI22_X1 U23373 ( .A1(n20653), .A2(n20289), .B1(n20322), .B2(n20662), .ZN(
        n20265) );
  OAI211_X1 U23374 ( .C1(n20271), .C2(n21972), .A(n20266), .B(n20265), .ZN(
        P2_U3072) );
  OAI22_X1 U23375 ( .A1(n20287), .A2(n20671), .B1(n20286), .B2(n20267), .ZN(
        n20268) );
  INV_X1 U23376 ( .A(n20268), .ZN(n20270) );
  AOI22_X1 U23377 ( .A1(n20667), .A2(n20289), .B1(n20322), .B2(n20668), .ZN(
        n20269) );
  OAI211_X1 U23378 ( .C1(n20271), .C2(n11143), .A(n20270), .B(n20269), .ZN(
        P2_U3073) );
  AOI22_X1 U23379 ( .A1(n20322), .A2(n20623), .B1(n20283), .B2(n20672), .ZN(
        n20273) );
  AOI22_X1 U23380 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20290), .B1(
        n20673), .B2(n20289), .ZN(n20272) );
  OAI211_X1 U23381 ( .C1(n20626), .C2(n20287), .A(n20273), .B(n20272), .ZN(
        P2_U3074) );
  INV_X1 U23382 ( .A(n20322), .ZN(n20293) );
  OAI22_X1 U23383 ( .A1(n20287), .A2(n20683), .B1(n20286), .B2(n20274), .ZN(
        n20275) );
  INV_X1 U23384 ( .A(n20275), .ZN(n20277) );
  AOI22_X1 U23385 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20290), .B1(
        n20679), .B2(n20289), .ZN(n20276) );
  OAI211_X1 U23386 ( .C1(n20595), .C2(n20293), .A(n20277), .B(n20276), .ZN(
        P2_U3075) );
  OAI22_X1 U23387 ( .A1(n20287), .A2(n20630), .B1(n20286), .B2(n20629), .ZN(
        n20278) );
  INV_X1 U23388 ( .A(n20278), .ZN(n20280) );
  AOI22_X1 U23389 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20290), .B1(
        n20685), .B2(n20289), .ZN(n20279) );
  OAI211_X1 U23390 ( .C1(n20689), .C2(n20293), .A(n20280), .B(n20279), .ZN(
        P2_U3076) );
  AOI22_X1 U23391 ( .A1(n20322), .A2(n20692), .B1(n20283), .B2(n20690), .ZN(
        n20282) );
  AOI22_X1 U23392 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20290), .B1(
        n20691), .B2(n20289), .ZN(n20281) );
  OAI211_X1 U23393 ( .C1(n20695), .C2(n20287), .A(n20282), .B(n20281), .ZN(
        P2_U3077) );
  AOI22_X1 U23394 ( .A1(n20322), .A2(n20572), .B1(n20696), .B2(n20283), .ZN(
        n20285) );
  AOI22_X1 U23395 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20290), .B1(
        n20697), .B2(n20289), .ZN(n20284) );
  OAI211_X1 U23396 ( .C1(n20638), .C2(n20287), .A(n20285), .B(n20284), .ZN(
        P2_U3078) );
  OAI22_X1 U23397 ( .A1(n20287), .A2(n20714), .B1(n20286), .B2(n20643), .ZN(
        n20288) );
  INV_X1 U23398 ( .A(n20288), .ZN(n20292) );
  AOI22_X1 U23399 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20290), .B1(
        n20706), .B2(n20289), .ZN(n20291) );
  OAI211_X1 U23400 ( .C1(n20650), .C2(n20293), .A(n20292), .B(n20291), .ZN(
        P2_U3079) );
  NAND2_X1 U23401 ( .A1(n20812), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20388) );
  NOR2_X1 U23402 ( .A1(n20416), .A2(n20388), .ZN(n20320) );
  NOR2_X1 U23403 ( .A1(n20299), .A2(n20320), .ZN(n20298) );
  INV_X1 U23404 ( .A(n20295), .ZN(n20297) );
  INV_X1 U23405 ( .A(n20296), .ZN(n20549) );
  NAND2_X1 U23406 ( .A1(n20549), .A2(n20812), .ZN(n20303) );
  AOI22_X1 U23407 ( .A1(n20321), .A2(n20653), .B1(n20652), .B2(n20320), .ZN(
        n20307) );
  INV_X1 U23408 ( .A(n20299), .ZN(n20300) );
  AOI21_X1 U23409 ( .B1(n20300), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20305) );
  INV_X1 U23410 ( .A(n20548), .ZN(n20302) );
  OAI21_X1 U23411 ( .B1(n20322), .B2(n20351), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20301) );
  OAI21_X1 U23412 ( .B1(n20303), .B2(n20302), .A(n20301), .ZN(n20304) );
  AOI22_X1 U23413 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20582), .ZN(n20306) );
  OAI211_X1 U23414 ( .C1(n20369), .C2(n20347), .A(n20307), .B(n20306), .ZN(
        P2_U3080) );
  AOI22_X1 U23415 ( .A1(n20321), .A2(n20667), .B1(n20666), .B2(n20320), .ZN(
        n20309) );
  AOI22_X1 U23416 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20586), .ZN(n20308) );
  OAI211_X1 U23417 ( .C1(n20589), .C2(n20347), .A(n20309), .B(n20308), .ZN(
        P2_U3081) );
  AOI22_X1 U23418 ( .A1(n20321), .A2(n20673), .B1(n20672), .B2(n20320), .ZN(
        n20311) );
  AOI22_X1 U23419 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20674), .ZN(n20310) );
  OAI211_X1 U23420 ( .C1(n20677), .C2(n20347), .A(n20311), .B(n20310), .ZN(
        P2_U3082) );
  AOI22_X1 U23421 ( .A1(n20321), .A2(n20679), .B1(n20678), .B2(n20320), .ZN(
        n20313) );
  AOI22_X1 U23422 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20592), .ZN(n20312) );
  OAI211_X1 U23423 ( .C1(n20595), .C2(n20347), .A(n20313), .B(n20312), .ZN(
        P2_U3083) );
  AOI22_X1 U23424 ( .A1(n20321), .A2(n20685), .B1(n20684), .B2(n20320), .ZN(
        n20315) );
  AOI22_X1 U23425 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20686), .ZN(n20314) );
  OAI211_X1 U23426 ( .C1(n20689), .C2(n20347), .A(n20315), .B(n20314), .ZN(
        P2_U3084) );
  AOI22_X1 U23427 ( .A1(n20321), .A2(n20691), .B1(n20690), .B2(n20320), .ZN(
        n20317) );
  AOI22_X1 U23428 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20598), .ZN(n20316) );
  OAI211_X1 U23429 ( .C1(n20601), .C2(n20347), .A(n20317), .B(n20316), .ZN(
        P2_U3085) );
  AOI22_X1 U23430 ( .A1(n20321), .A2(n20697), .B1(n20696), .B2(n20320), .ZN(
        n20319) );
  AOI22_X1 U23431 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20698), .ZN(n20318) );
  OAI211_X1 U23432 ( .C1(n20703), .C2(n20347), .A(n20319), .B(n20318), .ZN(
        P2_U3086) );
  AOI22_X1 U23433 ( .A1(n20321), .A2(n20706), .B1(n20704), .B2(n20320), .ZN(
        n20325) );
  AOI22_X1 U23434 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20603), .ZN(n20324) );
  OAI211_X1 U23435 ( .C1(n20650), .C2(n20347), .A(n20325), .B(n20324), .ZN(
        P2_U3087) );
  NOR2_X1 U23436 ( .A1(n20388), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20330) );
  AOI22_X1 U23437 ( .A1(n20384), .A2(n20662), .B1(n20350), .B2(n20652), .ZN(
        n20336) );
  INV_X1 U23438 ( .A(n20331), .ZN(n20326) );
  AOI21_X1 U23439 ( .B1(n20326), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20329) );
  NOR2_X1 U23440 ( .A1(n20392), .A2(n20327), .ZN(n20334) );
  OR2_X1 U23441 ( .A1(n20330), .A2(n20334), .ZN(n20328) );
  NAND2_X1 U23442 ( .A1(n20800), .A2(n20330), .ZN(n20333) );
  NOR2_X1 U23443 ( .A1(n20331), .A2(n20350), .ZN(n20332) );
  AOI22_X1 U23444 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20353), .B1(
        n20653), .B2(n20352), .ZN(n20335) );
  OAI211_X1 U23445 ( .C1(n20665), .C2(n20347), .A(n20336), .B(n20335), .ZN(
        P2_U3088) );
  AOI22_X1 U23446 ( .A1(n20351), .A2(n20586), .B1(n20350), .B2(n20666), .ZN(
        n20338) );
  AOI22_X1 U23447 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20353), .B1(
        n20667), .B2(n20352), .ZN(n20337) );
  OAI211_X1 U23448 ( .C1(n20589), .C2(n20361), .A(n20338), .B(n20337), .ZN(
        P2_U3089) );
  AOI22_X1 U23449 ( .A1(n20384), .A2(n20623), .B1(n20350), .B2(n20672), .ZN(
        n20340) );
  AOI22_X1 U23450 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20353), .B1(
        n20673), .B2(n20352), .ZN(n20339) );
  OAI211_X1 U23451 ( .C1(n20626), .C2(n20347), .A(n20340), .B(n20339), .ZN(
        P2_U3090) );
  AOI22_X1 U23452 ( .A1(n20384), .A2(n20680), .B1(n20350), .B2(n20678), .ZN(
        n20342) );
  AOI22_X1 U23453 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20353), .B1(
        n20679), .B2(n20352), .ZN(n20341) );
  OAI211_X1 U23454 ( .C1(n20683), .C2(n20347), .A(n20342), .B(n20341), .ZN(
        P2_U3091) );
  AOI22_X1 U23455 ( .A1(n20351), .A2(n20686), .B1(n20350), .B2(n20684), .ZN(
        n20344) );
  AOI22_X1 U23456 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20353), .B1(
        n20685), .B2(n20352), .ZN(n20343) );
  OAI211_X1 U23457 ( .C1(n20689), .C2(n20361), .A(n20344), .B(n20343), .ZN(
        P2_U3092) );
  AOI22_X1 U23458 ( .A1(n20384), .A2(n20692), .B1(n20350), .B2(n20690), .ZN(
        n20346) );
  AOI22_X1 U23459 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20353), .B1(
        n20691), .B2(n20352), .ZN(n20345) );
  OAI211_X1 U23460 ( .C1(n20695), .C2(n20347), .A(n20346), .B(n20345), .ZN(
        P2_U3093) );
  AOI22_X1 U23461 ( .A1(n20351), .A2(n20698), .B1(n20696), .B2(n20350), .ZN(
        n20349) );
  AOI22_X1 U23462 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20353), .B1(
        n20697), .B2(n20352), .ZN(n20348) );
  OAI211_X1 U23463 ( .C1(n20703), .C2(n20361), .A(n20349), .B(n20348), .ZN(
        P2_U3094) );
  AOI22_X1 U23464 ( .A1(n20351), .A2(n20603), .B1(n20350), .B2(n20704), .ZN(
        n20355) );
  AOI22_X1 U23465 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20353), .B1(
        n20706), .B2(n20352), .ZN(n20354) );
  OAI211_X1 U23466 ( .C1(n20650), .C2(n20361), .A(n20355), .B(n20354), .ZN(
        P2_U3095) );
  INV_X1 U23467 ( .A(n20358), .ZN(n20489) );
  NAND2_X1 U23468 ( .A1(n20609), .A2(n20812), .ZN(n20393) );
  NOR2_X1 U23469 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20393), .ZN(
        n20382) );
  OAI21_X1 U23470 ( .B1(n20359), .B2(n20382), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20360) );
  AOI22_X1 U23471 ( .A1(n20383), .A2(n20653), .B1(n20652), .B2(n20382), .ZN(
        n20368) );
  AOI21_X1 U23472 ( .B1(n20361), .B2(n20415), .A(n20481), .ZN(n20366) );
  NOR2_X1 U23473 ( .A1(n20549), .A2(n20388), .ZN(n20365) );
  INV_X1 U23474 ( .A(n20382), .ZN(n20362) );
  OAI211_X1 U23475 ( .C1(n20363), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20362), 
        .B(n20808), .ZN(n20364) );
  AOI22_X1 U23476 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20582), .ZN(n20367) );
  OAI211_X1 U23477 ( .C1(n20369), .C2(n20415), .A(n20368), .B(n20367), .ZN(
        P2_U3096) );
  AOI22_X1 U23478 ( .A1(n20383), .A2(n20667), .B1(n20666), .B2(n20382), .ZN(
        n20371) );
  AOI22_X1 U23479 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20586), .ZN(n20370) );
  OAI211_X1 U23480 ( .C1(n20589), .C2(n20415), .A(n20371), .B(n20370), .ZN(
        P2_U3097) );
  AOI22_X1 U23481 ( .A1(n20383), .A2(n20673), .B1(n20672), .B2(n20382), .ZN(
        n20373) );
  AOI22_X1 U23482 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20674), .ZN(n20372) );
  OAI211_X1 U23483 ( .C1(n20677), .C2(n20415), .A(n20373), .B(n20372), .ZN(
        P2_U3098) );
  AOI22_X1 U23484 ( .A1(n20383), .A2(n20679), .B1(n20678), .B2(n20382), .ZN(
        n20375) );
  AOI22_X1 U23485 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20592), .ZN(n20374) );
  OAI211_X1 U23486 ( .C1(n20595), .C2(n20415), .A(n20375), .B(n20374), .ZN(
        P2_U3099) );
  AOI22_X1 U23487 ( .A1(n20383), .A2(n20685), .B1(n20684), .B2(n20382), .ZN(
        n20377) );
  AOI22_X1 U23488 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20686), .ZN(n20376) );
  OAI211_X1 U23489 ( .C1(n20689), .C2(n20415), .A(n20377), .B(n20376), .ZN(
        P2_U3100) );
  AOI22_X1 U23490 ( .A1(n20383), .A2(n20691), .B1(n20690), .B2(n20382), .ZN(
        n20379) );
  AOI22_X1 U23491 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20598), .ZN(n20378) );
  OAI211_X1 U23492 ( .C1(n20601), .C2(n20415), .A(n20379), .B(n20378), .ZN(
        P2_U3101) );
  AOI22_X1 U23493 ( .A1(n20383), .A2(n20697), .B1(n20696), .B2(n20382), .ZN(
        n20381) );
  AOI22_X1 U23494 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20698), .ZN(n20380) );
  OAI211_X1 U23495 ( .C1(n20703), .C2(n20415), .A(n20381), .B(n20380), .ZN(
        P2_U3102) );
  AOI22_X1 U23496 ( .A1(n20383), .A2(n20706), .B1(n20704), .B2(n20382), .ZN(
        n20387) );
  AOI22_X1 U23497 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20603), .ZN(n20386) );
  OAI211_X1 U23498 ( .C1(n20650), .C2(n20415), .A(n20387), .B(n20386), .ZN(
        P2_U3103) );
  INV_X1 U23499 ( .A(n20388), .ZN(n20389) );
  NAND2_X1 U23500 ( .A1(n20515), .A2(n20389), .ZN(n20425) );
  AOI22_X1 U23501 ( .A1(n20411), .A2(n20653), .B1(n20421), .B2(n20652), .ZN(
        n20398) );
  INV_X1 U23502 ( .A(n20391), .ZN(n20395) );
  OR2_X1 U23503 ( .A1(n20655), .A2(n20392), .ZN(n20809) );
  AOI22_X1 U23504 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20425), .B1(n20393), 
        .B2(n20809), .ZN(n20394) );
  NAND3_X1 U23505 ( .A1(n20395), .A2(n20394), .A3(n20660), .ZN(n20412) );
  AOI22_X1 U23506 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20412), .B1(
        n20417), .B2(n20662), .ZN(n20397) );
  OAI211_X1 U23507 ( .C1(n20665), .C2(n20415), .A(n20398), .B(n20397), .ZN(
        P2_U3104) );
  AOI22_X1 U23508 ( .A1(n20411), .A2(n20667), .B1(n20421), .B2(n20666), .ZN(
        n20400) );
  AOI22_X1 U23509 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20412), .B1(
        n20417), .B2(n20668), .ZN(n20399) );
  OAI211_X1 U23510 ( .C1(n20671), .C2(n20415), .A(n20400), .B(n20399), .ZN(
        P2_U3105) );
  AOI22_X1 U23511 ( .A1(n20411), .A2(n20673), .B1(n20421), .B2(n20672), .ZN(
        n20402) );
  AOI22_X1 U23512 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20412), .B1(
        n20417), .B2(n20623), .ZN(n20401) );
  OAI211_X1 U23513 ( .C1(n20626), .C2(n20415), .A(n20402), .B(n20401), .ZN(
        P2_U3106) );
  AOI22_X1 U23514 ( .A1(n20411), .A2(n20679), .B1(n20421), .B2(n20678), .ZN(
        n20404) );
  AOI22_X1 U23515 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20412), .B1(
        n20417), .B2(n20680), .ZN(n20403) );
  OAI211_X1 U23516 ( .C1(n20683), .C2(n20415), .A(n20404), .B(n20403), .ZN(
        P2_U3107) );
  AOI22_X1 U23517 ( .A1(n20411), .A2(n20685), .B1(n20421), .B2(n20684), .ZN(
        n20406) );
  AOI22_X1 U23518 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20412), .B1(
        n20417), .B2(n20567), .ZN(n20405) );
  OAI211_X1 U23519 ( .C1(n20630), .C2(n20415), .A(n20406), .B(n20405), .ZN(
        P2_U3108) );
  AOI22_X1 U23520 ( .A1(n20411), .A2(n20691), .B1(n20421), .B2(n20690), .ZN(
        n20408) );
  AOI22_X1 U23521 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20412), .B1(
        n20417), .B2(n20692), .ZN(n20407) );
  OAI211_X1 U23522 ( .C1(n20695), .C2(n20415), .A(n20408), .B(n20407), .ZN(
        P2_U3109) );
  AOI22_X1 U23523 ( .A1(n20411), .A2(n20697), .B1(n20696), .B2(n20421), .ZN(
        n20410) );
  AOI22_X1 U23524 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20412), .B1(
        n20417), .B2(n20572), .ZN(n20409) );
  OAI211_X1 U23525 ( .C1(n20638), .C2(n20415), .A(n20410), .B(n20409), .ZN(
        P2_U3110) );
  AOI22_X1 U23526 ( .A1(n20411), .A2(n20706), .B1(n20421), .B2(n20704), .ZN(
        n20414) );
  AOI22_X1 U23527 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20412), .B1(
        n20417), .B2(n20708), .ZN(n20413) );
  OAI211_X1 U23528 ( .C1(n20714), .C2(n20415), .A(n20414), .B(n20413), .ZN(
        P2_U3111) );
  NAND2_X1 U23529 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20821), .ZN(
        n20513) );
  NOR2_X1 U23530 ( .A1(n20416), .A2(n20513), .ZN(n20443) );
  AOI22_X1 U23531 ( .A1(n20470), .A2(n20662), .B1(n20443), .B2(n20652), .ZN(
        n20430) );
  INV_X1 U23532 ( .A(n20417), .ZN(n20418) );
  NAND2_X1 U23533 ( .A1(n20800), .A2(n20418), .ZN(n20419) );
  OR2_X1 U23534 ( .A1(n20470), .A2(n20419), .ZN(n20420) );
  NAND2_X1 U23535 ( .A1(n20800), .A2(n20481), .ZN(n20802) );
  NOR2_X1 U23536 ( .A1(n20428), .A2(n20421), .ZN(n20422) );
  OAI21_X1 U23537 ( .B1(n20424), .B2(n20443), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20427) );
  NOR2_X1 U23538 ( .A1(n20443), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20426) );
  AOI22_X1 U23539 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20445), .B1(
        n20653), .B2(n20444), .ZN(n20429) );
  OAI211_X1 U23540 ( .C1(n20665), .C2(n20448), .A(n20430), .B(n20429), .ZN(
        P2_U3112) );
  AOI22_X1 U23541 ( .A1(n20470), .A2(n20668), .B1(n20443), .B2(n20666), .ZN(
        n20432) );
  AOI22_X1 U23542 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20445), .B1(
        n20667), .B2(n20444), .ZN(n20431) );
  OAI211_X1 U23543 ( .C1(n20671), .C2(n20448), .A(n20432), .B(n20431), .ZN(
        P2_U3113) );
  AOI22_X1 U23544 ( .A1(n20470), .A2(n20623), .B1(n20443), .B2(n20672), .ZN(
        n20434) );
  AOI22_X1 U23545 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20445), .B1(
        n20673), .B2(n20444), .ZN(n20433) );
  OAI211_X1 U23546 ( .C1(n20626), .C2(n20448), .A(n20434), .B(n20433), .ZN(
        P2_U3114) );
  AOI22_X1 U23547 ( .A1(n20470), .A2(n20680), .B1(n20443), .B2(n20678), .ZN(
        n20436) );
  AOI22_X1 U23548 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20445), .B1(
        n20679), .B2(n20444), .ZN(n20435) );
  OAI211_X1 U23549 ( .C1(n20683), .C2(n20448), .A(n20436), .B(n20435), .ZN(
        P2_U3115) );
  AOI22_X1 U23550 ( .A1(n20470), .A2(n20567), .B1(n20443), .B2(n20684), .ZN(
        n20438) );
  AOI22_X1 U23551 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20445), .B1(
        n20685), .B2(n20444), .ZN(n20437) );
  OAI211_X1 U23552 ( .C1(n20630), .C2(n20448), .A(n20438), .B(n20437), .ZN(
        P2_U3116) );
  AOI22_X1 U23553 ( .A1(n20470), .A2(n20692), .B1(n20443), .B2(n20690), .ZN(
        n20440) );
  AOI22_X1 U23554 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20445), .B1(
        n20691), .B2(n20444), .ZN(n20439) );
  OAI211_X1 U23555 ( .C1(n20695), .C2(n20448), .A(n20440), .B(n20439), .ZN(
        P2_U3117) );
  AOI22_X1 U23556 ( .A1(n20470), .A2(n20572), .B1(n20696), .B2(n20443), .ZN(
        n20442) );
  AOI22_X1 U23557 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20445), .B1(
        n20697), .B2(n20444), .ZN(n20441) );
  OAI211_X1 U23558 ( .C1(n20638), .C2(n20448), .A(n20442), .B(n20441), .ZN(
        P2_U3118) );
  AOI22_X1 U23559 ( .A1(n20470), .A2(n20708), .B1(n20443), .B2(n20704), .ZN(
        n20447) );
  AOI22_X1 U23560 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20445), .B1(
        n20706), .B2(n20444), .ZN(n20446) );
  OAI211_X1 U23561 ( .C1(n20714), .C2(n20448), .A(n20447), .B(n20446), .ZN(
        P2_U3119) );
  NOR2_X1 U23562 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20513), .ZN(
        n20453) );
  NAND2_X1 U23563 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20453), .ZN(
        n20480) );
  INV_X1 U23564 ( .A(n20480), .ZN(n20473) );
  AOI22_X1 U23565 ( .A1(n20508), .A2(n20662), .B1(n20652), .B2(n20473), .ZN(
        n20459) );
  OAI21_X1 U23566 ( .B1(n20656), .B2(n20450), .A(n20800), .ZN(n20457) );
  OAI211_X1 U23567 ( .C1(n20451), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20480), 
        .B(n20808), .ZN(n20452) );
  INV_X1 U23568 ( .A(n20453), .ZN(n20456) );
  OAI21_X1 U23569 ( .B1(n20454), .B2(n20473), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20455) );
  AOI22_X1 U23570 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20475), .B1(
        n20653), .B2(n20474), .ZN(n20458) );
  OAI211_X1 U23571 ( .C1(n20665), .C2(n20478), .A(n20459), .B(n20458), .ZN(
        P2_U3120) );
  AOI22_X1 U23572 ( .A1(n20508), .A2(n20668), .B1(n20666), .B2(n20473), .ZN(
        n20461) );
  AOI22_X1 U23573 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20475), .B1(
        n20667), .B2(n20474), .ZN(n20460) );
  OAI211_X1 U23574 ( .C1(n20671), .C2(n20478), .A(n20461), .B(n20460), .ZN(
        P2_U3121) );
  AOI22_X1 U23575 ( .A1(n20470), .A2(n20674), .B1(n20672), .B2(n20473), .ZN(
        n20463) );
  AOI22_X1 U23576 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20475), .B1(
        n20673), .B2(n20474), .ZN(n20462) );
  OAI211_X1 U23577 ( .C1(n20677), .C2(n20505), .A(n20463), .B(n20462), .ZN(
        P2_U3122) );
  AOI22_X1 U23578 ( .A1(n20470), .A2(n20592), .B1(n20678), .B2(n20473), .ZN(
        n20465) );
  AOI22_X1 U23579 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20475), .B1(
        n20679), .B2(n20474), .ZN(n20464) );
  OAI211_X1 U23580 ( .C1(n20595), .C2(n20505), .A(n20465), .B(n20464), .ZN(
        P2_U3123) );
  AOI22_X1 U23581 ( .A1(n20508), .A2(n20567), .B1(n20684), .B2(n20473), .ZN(
        n20467) );
  AOI22_X1 U23582 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20475), .B1(
        n20685), .B2(n20474), .ZN(n20466) );
  OAI211_X1 U23583 ( .C1(n20630), .C2(n20478), .A(n20467), .B(n20466), .ZN(
        P2_U3124) );
  AOI22_X1 U23584 ( .A1(n20470), .A2(n20598), .B1(n20690), .B2(n20473), .ZN(
        n20469) );
  AOI22_X1 U23585 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20475), .B1(
        n20691), .B2(n20474), .ZN(n20468) );
  OAI211_X1 U23586 ( .C1(n20601), .C2(n20505), .A(n20469), .B(n20468), .ZN(
        P2_U3125) );
  AOI22_X1 U23587 ( .A1(n20470), .A2(n20698), .B1(n20696), .B2(n20473), .ZN(
        n20472) );
  AOI22_X1 U23588 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20475), .B1(
        n20697), .B2(n20474), .ZN(n20471) );
  OAI211_X1 U23589 ( .C1(n20703), .C2(n20505), .A(n20472), .B(n20471), .ZN(
        P2_U3126) );
  AOI22_X1 U23590 ( .A1(n20508), .A2(n20708), .B1(n20704), .B2(n20473), .ZN(
        n20477) );
  AOI22_X1 U23591 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20475), .B1(
        n20706), .B2(n20474), .ZN(n20476) );
  OAI211_X1 U23592 ( .C1(n20714), .C2(n20478), .A(n20477), .B(n20476), .ZN(
        P2_U3127) );
  INV_X1 U23593 ( .A(n20608), .ZN(n20479) );
  OAI221_X1 U23594 ( .B1(n20481), .B2(n20541), .C1(n20481), .C2(n20505), .A(
        n20480), .ZN(n20483) );
  OR2_X1 U23595 ( .A1(n20487), .A2(n17300), .ZN(n20482) );
  NAND3_X1 U23596 ( .A1(n20483), .A2(n20814), .A3(n20482), .ZN(n20485) );
  NOR2_X1 U23597 ( .A1(n20831), .A2(n20513), .ZN(n20525) );
  INV_X1 U23598 ( .A(n20525), .ZN(n20512) );
  NOR2_X1 U23599 ( .A1(n20512), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20506) );
  INV_X1 U23600 ( .A(n20506), .ZN(n20484) );
  NAND2_X1 U23601 ( .A1(n20485), .A2(n20484), .ZN(n20486) );
  OAI21_X1 U23602 ( .B1(n20487), .B2(n20506), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20488) );
  AOI22_X1 U23603 ( .A1(n20507), .A2(n20653), .B1(n20652), .B2(n20506), .ZN(
        n20491) );
  AOI22_X1 U23604 ( .A1(n20508), .A2(n20582), .B1(n20544), .B2(n20662), .ZN(
        n20490) );
  OAI211_X1 U23605 ( .C1(n20492), .C2(n16037), .A(n20491), .B(n20490), .ZN(
        P2_U3128) );
  AOI22_X1 U23606 ( .A1(n20507), .A2(n20667), .B1(n20666), .B2(n20506), .ZN(
        n20494) );
  AOI22_X1 U23607 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20509), .B1(
        n20544), .B2(n20668), .ZN(n20493) );
  OAI211_X1 U23608 ( .C1(n20671), .C2(n20505), .A(n20494), .B(n20493), .ZN(
        P2_U3129) );
  AOI22_X1 U23609 ( .A1(n20507), .A2(n20673), .B1(n20672), .B2(n20506), .ZN(
        n20496) );
  AOI22_X1 U23610 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20509), .B1(
        n20544), .B2(n20623), .ZN(n20495) );
  OAI211_X1 U23611 ( .C1(n20626), .C2(n20505), .A(n20496), .B(n20495), .ZN(
        P2_U3130) );
  AOI22_X1 U23612 ( .A1(n20507), .A2(n20679), .B1(n20678), .B2(n20506), .ZN(
        n20498) );
  AOI22_X1 U23613 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20592), .ZN(n20497) );
  OAI211_X1 U23614 ( .C1(n20595), .C2(n20541), .A(n20498), .B(n20497), .ZN(
        P2_U3131) );
  AOI22_X1 U23615 ( .A1(n20507), .A2(n20685), .B1(n20684), .B2(n20506), .ZN(
        n20500) );
  AOI22_X1 U23616 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20686), .ZN(n20499) );
  OAI211_X1 U23617 ( .C1(n20689), .C2(n20541), .A(n20500), .B(n20499), .ZN(
        P2_U3132) );
  AOI22_X1 U23618 ( .A1(n20507), .A2(n20691), .B1(n20690), .B2(n20506), .ZN(
        n20502) );
  AOI22_X1 U23619 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20509), .B1(
        n20544), .B2(n20692), .ZN(n20501) );
  OAI211_X1 U23620 ( .C1(n20695), .C2(n20505), .A(n20502), .B(n20501), .ZN(
        P2_U3133) );
  AOI22_X1 U23621 ( .A1(n20507), .A2(n20697), .B1(n20696), .B2(n20506), .ZN(
        n20504) );
  AOI22_X1 U23622 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20509), .B1(
        n20544), .B2(n20572), .ZN(n20503) );
  OAI211_X1 U23623 ( .C1(n20638), .C2(n20505), .A(n20504), .B(n20503), .ZN(
        P2_U3134) );
  AOI22_X1 U23624 ( .A1(n20507), .A2(n20706), .B1(n20704), .B2(n20506), .ZN(
        n20511) );
  AOI22_X1 U23625 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20603), .ZN(n20510) );
  OAI211_X1 U23626 ( .C1(n20650), .C2(n20541), .A(n20511), .B(n20510), .ZN(
        P2_U3135) );
  OR2_X1 U23627 ( .A1(n20512), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20518) );
  INV_X1 U23628 ( .A(n20513), .ZN(n20514) );
  NAND2_X1 U23629 ( .A1(n20515), .A2(n20514), .ZN(n20519) );
  NAND2_X1 U23630 ( .A1(n20519), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20516) );
  INV_X1 U23631 ( .A(n20519), .ZN(n20542) );
  AOI22_X1 U23632 ( .A1(n20543), .A2(n20653), .B1(n20652), .B2(n20542), .ZN(
        n20528) );
  INV_X1 U23633 ( .A(n20656), .ZN(n20524) );
  NAND2_X1 U23634 ( .A1(n20519), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20520) );
  NAND2_X1 U23635 ( .A1(n20660), .A2(n20520), .ZN(n20521) );
  NOR2_X1 U23636 ( .A1(n20522), .A2(n20521), .ZN(n20523) );
  OAI221_X1 U23637 ( .B1(n20525), .B2(n20801), .C1(n20525), .C2(n20524), .A(
        n20523), .ZN(n20545) );
  AOI22_X1 U23638 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20545), .B1(
        n20553), .B2(n20662), .ZN(n20527) );
  OAI211_X1 U23639 ( .C1(n20665), .C2(n20541), .A(n20528), .B(n20527), .ZN(
        P2_U3136) );
  AOI22_X1 U23640 ( .A1(n20543), .A2(n20667), .B1(n20666), .B2(n20542), .ZN(
        n20530) );
  AOI22_X1 U23641 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20545), .B1(
        n20553), .B2(n20668), .ZN(n20529) );
  OAI211_X1 U23642 ( .C1(n20671), .C2(n20541), .A(n20530), .B(n20529), .ZN(
        P2_U3137) );
  AOI22_X1 U23643 ( .A1(n20543), .A2(n20673), .B1(n20672), .B2(n20542), .ZN(
        n20532) );
  AOI22_X1 U23644 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20674), .ZN(n20531) );
  OAI211_X1 U23645 ( .C1(n20677), .C2(n20580), .A(n20532), .B(n20531), .ZN(
        P2_U3138) );
  AOI22_X1 U23646 ( .A1(n20543), .A2(n20679), .B1(n20678), .B2(n20542), .ZN(
        n20534) );
  AOI22_X1 U23647 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20545), .B1(
        n20553), .B2(n20680), .ZN(n20533) );
  OAI211_X1 U23648 ( .C1(n20683), .C2(n20541), .A(n20534), .B(n20533), .ZN(
        P2_U3139) );
  AOI22_X1 U23649 ( .A1(n20543), .A2(n20685), .B1(n20684), .B2(n20542), .ZN(
        n20536) );
  AOI22_X1 U23650 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20545), .B1(
        n20553), .B2(n20567), .ZN(n20535) );
  OAI211_X1 U23651 ( .C1(n20630), .C2(n20541), .A(n20536), .B(n20535), .ZN(
        P2_U3140) );
  AOI22_X1 U23652 ( .A1(n20543), .A2(n20691), .B1(n20690), .B2(n20542), .ZN(
        n20538) );
  AOI22_X1 U23653 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20598), .ZN(n20537) );
  OAI211_X1 U23654 ( .C1(n20601), .C2(n20580), .A(n20538), .B(n20537), .ZN(
        P2_U3141) );
  AOI22_X1 U23655 ( .A1(n20543), .A2(n20697), .B1(n20696), .B2(n20542), .ZN(
        n20540) );
  AOI22_X1 U23656 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20545), .B1(
        n20553), .B2(n20572), .ZN(n20539) );
  OAI211_X1 U23657 ( .C1(n20638), .C2(n20541), .A(n20540), .B(n20539), .ZN(
        P2_U3142) );
  AOI22_X1 U23658 ( .A1(n20543), .A2(n20706), .B1(n20704), .B2(n20542), .ZN(
        n20547) );
  AOI22_X1 U23659 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20603), .ZN(n20546) );
  OAI211_X1 U23660 ( .C1(n20650), .C2(n20580), .A(n20547), .B(n20546), .ZN(
        P2_U3143) );
  NAND3_X1 U23661 ( .A1(n20549), .A2(n20548), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20556) );
  NOR2_X1 U23662 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20550), .ZN(
        n20575) );
  AOI22_X1 U23663 ( .A1(n20576), .A2(n20653), .B1(n20652), .B2(n20575), .ZN(
        n20560) );
  OAI21_X1 U23664 ( .B1(n20553), .B2(n20604), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20557) );
  AOI211_X1 U23665 ( .C1(n20557), .C2(n20556), .A(n20555), .B(n20554), .ZN(
        n20558) );
  AOI22_X1 U23666 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20577), .B1(
        n20604), .B2(n20662), .ZN(n20559) );
  OAI211_X1 U23667 ( .C1(n20665), .C2(n20580), .A(n20560), .B(n20559), .ZN(
        P2_U3144) );
  AOI22_X1 U23668 ( .A1(n20576), .A2(n20667), .B1(n20666), .B2(n20575), .ZN(
        n20562) );
  AOI22_X1 U23669 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20577), .B1(
        n20604), .B2(n20668), .ZN(n20561) );
  OAI211_X1 U23670 ( .C1(n20671), .C2(n20580), .A(n20562), .B(n20561), .ZN(
        P2_U3145) );
  AOI22_X1 U23671 ( .A1(n20576), .A2(n20673), .B1(n20672), .B2(n20575), .ZN(
        n20564) );
  AOI22_X1 U23672 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20577), .B1(
        n20604), .B2(n20623), .ZN(n20563) );
  OAI211_X1 U23673 ( .C1(n20626), .C2(n20580), .A(n20564), .B(n20563), .ZN(
        P2_U3146) );
  AOI22_X1 U23674 ( .A1(n20576), .A2(n20679), .B1(n20678), .B2(n20575), .ZN(
        n20566) );
  AOI22_X1 U23675 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20577), .B1(
        n20604), .B2(n20680), .ZN(n20565) );
  OAI211_X1 U23676 ( .C1(n20683), .C2(n20580), .A(n20566), .B(n20565), .ZN(
        P2_U3147) );
  AOI22_X1 U23677 ( .A1(n20576), .A2(n20685), .B1(n20684), .B2(n20575), .ZN(
        n20569) );
  AOI22_X1 U23678 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20577), .B1(
        n20604), .B2(n20567), .ZN(n20568) );
  OAI211_X1 U23679 ( .C1(n20630), .C2(n20580), .A(n20569), .B(n20568), .ZN(
        P2_U3148) );
  AOI22_X1 U23680 ( .A1(n20576), .A2(n20691), .B1(n20690), .B2(n20575), .ZN(
        n20571) );
  AOI22_X1 U23681 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20577), .B1(
        n20604), .B2(n20692), .ZN(n20570) );
  OAI211_X1 U23682 ( .C1(n20695), .C2(n20580), .A(n20571), .B(n20570), .ZN(
        P2_U3149) );
  AOI22_X1 U23683 ( .A1(n20576), .A2(n20697), .B1(n20696), .B2(n20575), .ZN(
        n20574) );
  AOI22_X1 U23684 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20577), .B1(
        n20604), .B2(n20572), .ZN(n20573) );
  OAI211_X1 U23685 ( .C1(n20638), .C2(n20580), .A(n20574), .B(n20573), .ZN(
        P2_U3150) );
  AOI22_X1 U23686 ( .A1(n20576), .A2(n20706), .B1(n20704), .B2(n20575), .ZN(
        n20579) );
  AOI22_X1 U23687 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20577), .B1(
        n20604), .B2(n20708), .ZN(n20578) );
  OAI211_X1 U23688 ( .C1(n20714), .C2(n20580), .A(n20579), .B(n20578), .ZN(
        P2_U3151) );
  AOI22_X1 U23689 ( .A1(n20602), .A2(n20653), .B1(n20615), .B2(n20652), .ZN(
        n20584) );
  AOI22_X1 U23690 ( .A1(n20604), .A2(n20582), .B1(n20581), .B2(n20662), .ZN(
        n20583) );
  OAI211_X1 U23691 ( .C1(n20585), .C2(n16030), .A(n20584), .B(n20583), .ZN(
        P2_U3152) );
  AOI22_X1 U23692 ( .A1(n20602), .A2(n20667), .B1(n20615), .B2(n20666), .ZN(
        n20588) );
  AOI22_X1 U23693 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20586), .ZN(n20587) );
  OAI211_X1 U23694 ( .C1(n20589), .C2(n20644), .A(n20588), .B(n20587), .ZN(
        P2_U3153) );
  AOI22_X1 U23695 ( .A1(n20602), .A2(n20673), .B1(n20615), .B2(n20672), .ZN(
        n20591) );
  AOI22_X1 U23696 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20674), .ZN(n20590) );
  OAI211_X1 U23697 ( .C1(n20677), .C2(n20644), .A(n20591), .B(n20590), .ZN(
        P2_U3154) );
  AOI22_X1 U23698 ( .A1(n20602), .A2(n20679), .B1(n20615), .B2(n20678), .ZN(
        n20594) );
  AOI22_X1 U23699 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20592), .ZN(n20593) );
  OAI211_X1 U23700 ( .C1(n20595), .C2(n20644), .A(n20594), .B(n20593), .ZN(
        P2_U3155) );
  AOI22_X1 U23701 ( .A1(n20602), .A2(n20685), .B1(n20615), .B2(n20684), .ZN(
        n20597) );
  AOI22_X1 U23702 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20686), .ZN(n20596) );
  OAI211_X1 U23703 ( .C1(n20689), .C2(n20644), .A(n20597), .B(n20596), .ZN(
        P2_U3156) );
  AOI22_X1 U23704 ( .A1(n20602), .A2(n20691), .B1(n20615), .B2(n20690), .ZN(
        n20600) );
  AOI22_X1 U23705 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20598), .ZN(n20599) );
  OAI211_X1 U23706 ( .C1(n20601), .C2(n20644), .A(n20600), .B(n20599), .ZN(
        P2_U3157) );
  AOI22_X1 U23707 ( .A1(n20602), .A2(n20706), .B1(n20615), .B2(n20704), .ZN(
        n20607) );
  AOI22_X1 U23708 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20603), .ZN(n20606) );
  OAI211_X1 U23709 ( .C1(n20650), .C2(n20644), .A(n20607), .B(n20606), .ZN(
        P2_U3159) );
  NAND2_X1 U23710 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20609), .ZN(
        n20654) );
  NOR2_X1 U23711 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20654), .ZN(
        n20634) );
  AOI22_X1 U23712 ( .A1(n20699), .A2(n20662), .B1(n20652), .B2(n20634), .ZN(
        n20620) );
  NAND2_X1 U23713 ( .A1(n20644), .A2(n20800), .ZN(n20610) );
  OAI21_X1 U23714 ( .B1(n20610), .B2(n20699), .A(n20802), .ZN(n20614) );
  OAI21_X1 U23715 ( .B1(n20616), .B2(n20800), .A(n20814), .ZN(n20611) );
  AOI21_X1 U23716 ( .B1(n20614), .B2(n20612), .A(n20611), .ZN(n20613) );
  OAI21_X2 U23717 ( .B1(n20613), .B2(n20634), .A(n20660), .ZN(n20647) );
  OAI21_X1 U23718 ( .B1(n20615), .B2(n20634), .A(n20614), .ZN(n20618) );
  OAI21_X1 U23719 ( .B1(n20616), .B2(n20634), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20617) );
  AOI22_X1 U23720 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20647), .B1(
        n20653), .B2(n20646), .ZN(n20619) );
  OAI211_X1 U23721 ( .C1(n20665), .C2(n20644), .A(n20620), .B(n20619), .ZN(
        P2_U3160) );
  AOI22_X1 U23722 ( .A1(n20699), .A2(n20668), .B1(n20666), .B2(n20634), .ZN(
        n20622) );
  AOI22_X1 U23723 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20647), .B1(
        n20667), .B2(n20646), .ZN(n20621) );
  OAI211_X1 U23724 ( .C1(n20671), .C2(n20644), .A(n20622), .B(n20621), .ZN(
        P2_U3161) );
  AOI22_X1 U23725 ( .A1(n20699), .A2(n20623), .B1(n20672), .B2(n20634), .ZN(
        n20625) );
  AOI22_X1 U23726 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20647), .B1(
        n20673), .B2(n20646), .ZN(n20624) );
  OAI211_X1 U23727 ( .C1(n20626), .C2(n20644), .A(n20625), .B(n20624), .ZN(
        P2_U3162) );
  AOI22_X1 U23728 ( .A1(n20699), .A2(n20680), .B1(n20678), .B2(n20634), .ZN(
        n20628) );
  AOI22_X1 U23729 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20647), .B1(
        n20679), .B2(n20646), .ZN(n20627) );
  OAI211_X1 U23730 ( .C1(n20683), .C2(n20644), .A(n20628), .B(n20627), .ZN(
        P2_U3163) );
  INV_X1 U23731 ( .A(n20634), .ZN(n20642) );
  OAI22_X1 U23732 ( .A1(n20644), .A2(n20630), .B1(n20629), .B2(n20642), .ZN(
        n20631) );
  INV_X1 U23733 ( .A(n20631), .ZN(n20633) );
  AOI22_X1 U23734 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20647), .B1(
        n20685), .B2(n20646), .ZN(n20632) );
  OAI211_X1 U23735 ( .C1(n20689), .C2(n20713), .A(n20633), .B(n20632), .ZN(
        P2_U3164) );
  AOI22_X1 U23736 ( .A1(n20699), .A2(n20692), .B1(n20690), .B2(n20634), .ZN(
        n20636) );
  AOI22_X1 U23737 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20647), .B1(
        n20691), .B2(n20646), .ZN(n20635) );
  OAI211_X1 U23738 ( .C1(n20695), .C2(n20644), .A(n20636), .B(n20635), .ZN(
        P2_U3165) );
  OAI22_X1 U23739 ( .A1(n20644), .A2(n20638), .B1(n20637), .B2(n20642), .ZN(
        n20639) );
  INV_X1 U23740 ( .A(n20639), .ZN(n20641) );
  AOI22_X1 U23741 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20647), .B1(
        n20697), .B2(n20646), .ZN(n20640) );
  OAI211_X1 U23742 ( .C1(n20703), .C2(n20713), .A(n20641), .B(n20640), .ZN(
        P2_U3166) );
  OAI22_X1 U23743 ( .A1(n20644), .A2(n20714), .B1(n20643), .B2(n20642), .ZN(
        n20645) );
  INV_X1 U23744 ( .A(n20645), .ZN(n20649) );
  AOI22_X1 U23745 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20647), .B1(
        n20706), .B2(n20646), .ZN(n20648) );
  OAI211_X1 U23746 ( .C1(n20650), .C2(n20713), .A(n20649), .B(n20648), .ZN(
        P2_U3167) );
  OAI21_X1 U23747 ( .B1(n11271), .B2(n20705), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20651) );
  AOI22_X1 U23748 ( .A1(n20707), .A2(n20653), .B1(n20705), .B2(n20652), .ZN(
        n20664) );
  OAI21_X1 U23749 ( .B1(n20656), .B2(n20655), .A(n20654), .ZN(n20661) );
  OAI211_X1 U23750 ( .C1(n20658), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20657), 
        .B(n20808), .ZN(n20659) );
  NAND3_X1 U23751 ( .A1(n20661), .A2(n20660), .A3(n20659), .ZN(n20710) );
  AOI22_X1 U23752 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20710), .B1(
        n20709), .B2(n20662), .ZN(n20663) );
  OAI211_X1 U23753 ( .C1(n20665), .C2(n20713), .A(n20664), .B(n20663), .ZN(
        P2_U3168) );
  AOI22_X1 U23754 ( .A1(n20707), .A2(n20667), .B1(n20705), .B2(n20666), .ZN(
        n20670) );
  AOI22_X1 U23755 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20710), .B1(
        n20709), .B2(n20668), .ZN(n20669) );
  OAI211_X1 U23756 ( .C1(n20671), .C2(n20713), .A(n20670), .B(n20669), .ZN(
        P2_U3169) );
  AOI22_X1 U23757 ( .A1(n20707), .A2(n20673), .B1(n20705), .B2(n20672), .ZN(
        n20676) );
  AOI22_X1 U23758 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20710), .B1(
        n20699), .B2(n20674), .ZN(n20675) );
  OAI211_X1 U23759 ( .C1(n20677), .C2(n20702), .A(n20676), .B(n20675), .ZN(
        P2_U3170) );
  AOI22_X1 U23760 ( .A1(n20707), .A2(n20679), .B1(n20705), .B2(n20678), .ZN(
        n20682) );
  AOI22_X1 U23761 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20710), .B1(
        n20709), .B2(n20680), .ZN(n20681) );
  OAI211_X1 U23762 ( .C1(n20683), .C2(n20713), .A(n20682), .B(n20681), .ZN(
        P2_U3171) );
  AOI22_X1 U23763 ( .A1(n20707), .A2(n20685), .B1(n20705), .B2(n20684), .ZN(
        n20688) );
  AOI22_X1 U23764 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20710), .B1(
        n20699), .B2(n20686), .ZN(n20687) );
  OAI211_X1 U23765 ( .C1(n20689), .C2(n20702), .A(n20688), .B(n20687), .ZN(
        P2_U3172) );
  AOI22_X1 U23766 ( .A1(n20707), .A2(n20691), .B1(n20705), .B2(n20690), .ZN(
        n20694) );
  AOI22_X1 U23767 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20710), .B1(
        n20709), .B2(n20692), .ZN(n20693) );
  OAI211_X1 U23768 ( .C1(n20695), .C2(n20713), .A(n20694), .B(n20693), .ZN(
        P2_U3173) );
  AOI22_X1 U23769 ( .A1(n20707), .A2(n20697), .B1(n20705), .B2(n20696), .ZN(
        n20701) );
  AOI22_X1 U23770 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20710), .B1(
        n20699), .B2(n20698), .ZN(n20700) );
  OAI211_X1 U23771 ( .C1(n20703), .C2(n20702), .A(n20701), .B(n20700), .ZN(
        P2_U3174) );
  AOI22_X1 U23772 ( .A1(n20707), .A2(n20706), .B1(n20705), .B2(n20704), .ZN(
        n20712) );
  AOI22_X1 U23773 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20710), .B1(
        n20709), .B2(n20708), .ZN(n20711) );
  OAI211_X1 U23774 ( .C1(n20714), .C2(n20713), .A(n20712), .B(n20711), .ZN(
        P2_U3175) );
  AND2_X1 U23775 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20715), .ZN(
        P2_U3179) );
  AND2_X1 U23776 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20715), .ZN(
        P2_U3180) );
  AND2_X1 U23777 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20715), .ZN(
        P2_U3181) );
  AND2_X1 U23778 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20715), .ZN(
        P2_U3182) );
  AND2_X1 U23779 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20715), .ZN(
        P2_U3183) );
  AND2_X1 U23780 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20715), .ZN(
        P2_U3184) );
  AND2_X1 U23781 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20715), .ZN(
        P2_U3185) );
  AND2_X1 U23782 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20715), .ZN(
        P2_U3186) );
  AND2_X1 U23783 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20715), .ZN(
        P2_U3187) );
  AND2_X1 U23784 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20715), .ZN(
        P2_U3188) );
  AND2_X1 U23785 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20715), .ZN(
        P2_U3189) );
  AND2_X1 U23786 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20715), .ZN(
        P2_U3190) );
  AND2_X1 U23787 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20715), .ZN(
        P2_U3191) );
  INV_X1 U23788 ( .A(P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n21932) );
  NOR2_X1 U23789 ( .A1(n21932), .A2(n20792), .ZN(P2_U3192) );
  AND2_X1 U23790 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20715), .ZN(
        P2_U3193) );
  AND2_X1 U23791 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20715), .ZN(
        P2_U3194) );
  AND2_X1 U23792 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20715), .ZN(
        P2_U3195) );
  AND2_X1 U23793 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20715), .ZN(
        P2_U3196) );
  AND2_X1 U23794 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20715), .ZN(
        P2_U3197) );
  AND2_X1 U23795 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20715), .ZN(
        P2_U3198) );
  AND2_X1 U23796 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20715), .ZN(
        P2_U3199) );
  AND2_X1 U23797 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20715), .ZN(
        P2_U3200) );
  AND2_X1 U23798 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20715), .ZN(P2_U3201) );
  AND2_X1 U23799 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20715), .ZN(P2_U3202) );
  AND2_X1 U23800 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20715), .ZN(P2_U3203) );
  AND2_X1 U23801 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20715), .ZN(P2_U3204) );
  AND2_X1 U23802 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20715), .ZN(P2_U3205) );
  AND2_X1 U23803 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20715), .ZN(P2_U3206) );
  AND2_X1 U23804 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20715), .ZN(P2_U3207) );
  AND2_X1 U23805 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20715), .ZN(P2_U3208) );
  NAND2_X1 U23806 ( .A1(n20844), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20719) );
  NAND3_X1 U23807 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20719), .ZN(n20716) );
  NOR3_X1 U23808 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21656), .ZN(n20730) );
  AOI21_X1 U23809 ( .B1(n20731), .B2(n20716), .A(n20730), .ZN(n20717) );
  OAI221_X1 U23810 ( .B1(n20718), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20718), .C2(n20723), .A(n20717), .ZN(P2_U3209) );
  OAI22_X1 U23811 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20728), .B1(HOLD), .B2(
        n20728), .ZN(n20720) );
  INV_X1 U23812 ( .A(n20719), .ZN(n20724) );
  AOI211_X1 U23813 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20720), .A(
        n20853), .B(n20724), .ZN(n20721) );
  OAI21_X1 U23814 ( .B1(n20723), .B2(n20722), .A(n20721), .ZN(P2_U3210) );
  NOR3_X1 U23815 ( .A1(HOLD), .A2(n20724), .A3(n20728), .ZN(n20729) );
  NOR2_X1 U23816 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(HOLD), .ZN(n20727)
         );
  INV_X1 U23817 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20860) );
  AOI22_X1 U23818 ( .A1(n20725), .A2(n20860), .B1(n20724), .B2(n21656), .ZN(
        n20726) );
  OAI33_X1 U23819 ( .A1(n20731), .A2(n20730), .A3(n20729), .B1(n20728), .B2(
        n20727), .B3(n20726), .ZN(P2_U3211) );
  NAND2_X1 U23820 ( .A1(n20862), .A2(n20731), .ZN(n20782) );
  OAI222_X1 U23821 ( .A1(n20777), .A2(n20734), .B1(n20733), .B2(n20862), .C1(
        n20732), .C2(n20778), .ZN(P2_U3212) );
  OAI222_X1 U23822 ( .A1(n20782), .A2(n20736), .B1(n20735), .B2(n20862), .C1(
        n20734), .C2(n20778), .ZN(P2_U3213) );
  OAI222_X1 U23823 ( .A1(n20782), .A2(n20738), .B1(n20737), .B2(n20862), .C1(
        n20736), .C2(n20778), .ZN(P2_U3214) );
  OAI222_X1 U23824 ( .A1(n20782), .A2(n16904), .B1(n21832), .B2(n20862), .C1(
        n20738), .C2(n20778), .ZN(P2_U3215) );
  OAI222_X1 U23825 ( .A1(n20782), .A2(n21812), .B1(n20739), .B2(n20862), .C1(
        n16904), .C2(n20778), .ZN(P2_U3216) );
  OAI222_X1 U23826 ( .A1(n20782), .A2(n20741), .B1(n20740), .B2(n20862), .C1(
        n21812), .C2(n20778), .ZN(P2_U3217) );
  OAI222_X1 U23827 ( .A1(n20777), .A2(n20743), .B1(n20742), .B2(n20862), .C1(
        n20741), .C2(n20778), .ZN(P2_U3218) );
  OAI222_X1 U23828 ( .A1(n20777), .A2(n20745), .B1(n20744), .B2(n20862), .C1(
        n20743), .C2(n20778), .ZN(P2_U3219) );
  OAI222_X1 U23829 ( .A1(n20777), .A2(n16841), .B1(n20746), .B2(n20862), .C1(
        n20745), .C2(n20778), .ZN(P2_U3220) );
  OAI222_X1 U23830 ( .A1(n20777), .A2(n20748), .B1(n20747), .B2(n20862), .C1(
        n16841), .C2(n20778), .ZN(P2_U3221) );
  INV_X1 U23831 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20750) );
  OAI222_X1 U23832 ( .A1(n20777), .A2(n20750), .B1(n20749), .B2(n20862), .C1(
        n20748), .C2(n20778), .ZN(P2_U3222) );
  OAI222_X1 U23833 ( .A1(n20777), .A2(n16809), .B1(n20751), .B2(n20862), .C1(
        n20750), .C2(n20778), .ZN(P2_U3223) );
  OAI222_X1 U23834 ( .A1(n20782), .A2(n15813), .B1(n20752), .B2(n20862), .C1(
        n16809), .C2(n20778), .ZN(P2_U3224) );
  OAI222_X1 U23835 ( .A1(n20782), .A2(n16789), .B1(n20753), .B2(n20862), .C1(
        n15813), .C2(n20778), .ZN(P2_U3225) );
  OAI222_X1 U23836 ( .A1(n20782), .A2(n20755), .B1(n20754), .B2(n20862), .C1(
        n16789), .C2(n20778), .ZN(P2_U3226) );
  OAI222_X1 U23837 ( .A1(n20782), .A2(n20757), .B1(n20756), .B2(n20862), .C1(
        n20755), .C2(n20778), .ZN(P2_U3227) );
  OAI222_X1 U23838 ( .A1(n20782), .A2(n15772), .B1(n20758), .B2(n20862), .C1(
        n20757), .C2(n20778), .ZN(P2_U3228) );
  OAI222_X1 U23839 ( .A1(n20782), .A2(n20760), .B1(n20759), .B2(n20862), .C1(
        n15772), .C2(n20778), .ZN(P2_U3229) );
  OAI222_X1 U23840 ( .A1(n20777), .A2(n20762), .B1(n20761), .B2(n20862), .C1(
        n20760), .C2(n20778), .ZN(P2_U3230) );
  OAI222_X1 U23841 ( .A1(n20777), .A2(n20764), .B1(n20763), .B2(n20862), .C1(
        n20762), .C2(n20778), .ZN(P2_U3231) );
  OAI222_X1 U23842 ( .A1(n20777), .A2(n16717), .B1(n20765), .B2(n20862), .C1(
        n20764), .C2(n20778), .ZN(P2_U3232) );
  OAI222_X1 U23843 ( .A1(n20777), .A2(n20767), .B1(n20766), .B2(n20862), .C1(
        n16717), .C2(n20778), .ZN(P2_U3233) );
  OAI222_X1 U23844 ( .A1(n20777), .A2(n20769), .B1(n20768), .B2(n20862), .C1(
        n20767), .C2(n20778), .ZN(P2_U3234) );
  OAI222_X1 U23845 ( .A1(n20777), .A2(n21909), .B1(n20770), .B2(n20862), .C1(
        n20769), .C2(n20778), .ZN(P2_U3235) );
  OAI222_X1 U23846 ( .A1(n20777), .A2(n16677), .B1(n20771), .B2(n20862), .C1(
        n21909), .C2(n20778), .ZN(P2_U3236) );
  OAI222_X1 U23847 ( .A1(n20777), .A2(n20774), .B1(n20772), .B2(n20862), .C1(
        n16677), .C2(n20778), .ZN(P2_U3237) );
  OAI222_X1 U23848 ( .A1(n20778), .A2(n20774), .B1(n20773), .B2(n20862), .C1(
        n16654), .C2(n20777), .ZN(P2_U3238) );
  OAI222_X1 U23849 ( .A1(n20777), .A2(n20776), .B1(n20775), .B2(n20862), .C1(
        n16654), .C2(n20778), .ZN(P2_U3239) );
  INV_X1 U23850 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20779) );
  OAI222_X1 U23851 ( .A1(n20777), .A2(n20779), .B1(n21809), .B2(n20862), .C1(
        n20776), .C2(n20778), .ZN(P2_U3240) );
  OAI222_X1 U23852 ( .A1(n20782), .A2(n20781), .B1(n20780), .B2(n20862), .C1(
        n20779), .C2(n20778), .ZN(P2_U3241) );
  INV_X1 U23853 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20783) );
  AOI22_X1 U23854 ( .A1(n20862), .A2(n20784), .B1(n20783), .B2(n20863), .ZN(
        P2_U3585) );
  INV_X1 U23855 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n20785) );
  AOI22_X1 U23856 ( .A1(n20862), .A2(n20786), .B1(n20785), .B2(n20863), .ZN(
        P2_U3586) );
  INV_X1 U23857 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20787) );
  AOI22_X1 U23858 ( .A1(n20862), .A2(n20788), .B1(n20787), .B2(n20863), .ZN(
        P2_U3587) );
  INV_X1 U23859 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20789) );
  AOI22_X1 U23860 ( .A1(n20862), .A2(n21816), .B1(n20789), .B2(n20863), .ZN(
        P2_U3588) );
  OAI21_X1 U23861 ( .B1(n20792), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20791), 
        .ZN(n20790) );
  INV_X1 U23862 ( .A(n20790), .ZN(P2_U3591) );
  OAI21_X1 U23863 ( .B1(n20792), .B2(n21862), .A(n20791), .ZN(P2_U3592) );
  INV_X1 U23864 ( .A(n20793), .ZN(n20794) );
  OAI222_X1 U23865 ( .A1(n20817), .A2(n20797), .B1(n20796), .B2(n20803), .C1(
        n20795), .C2(n20794), .ZN(n20799) );
  MUX2_X1 U23866 ( .A(n20799), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n20798), .Z(P2_U3599) );
  AND2_X1 U23867 ( .A1(n20800), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20826) );
  NAND2_X1 U23868 ( .A1(n20801), .A2(n20826), .ZN(n20813) );
  OR2_X1 U23869 ( .A1(n20824), .A2(n20808), .ZN(n20804) );
  AND3_X1 U23870 ( .A1(n20804), .A2(n20803), .A3(n20802), .ZN(n20816) );
  NAND2_X1 U23871 ( .A1(n20813), .A2(n20816), .ZN(n20806) );
  AOI22_X1 U23872 ( .A1(n20806), .A2(n20805), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n22054), .ZN(n20807) );
  OAI21_X1 U23873 ( .B1(n20809), .B2(n20808), .A(n20807), .ZN(n20810) );
  INV_X1 U23874 ( .A(n20810), .ZN(n20811) );
  AOI22_X1 U23875 ( .A1(n20832), .A2(n20812), .B1(n20811), .B2(n20829), .ZN(
        P2_U3602) );
  INV_X1 U23876 ( .A(n20813), .ZN(n20819) );
  OAI22_X1 U23877 ( .A1(n20817), .A2(n20816), .B1(n20815), .B2(n20814), .ZN(
        n20818) );
  NOR2_X1 U23878 ( .A1(n20819), .A2(n20818), .ZN(n20820) );
  AOI22_X1 U23879 ( .A1(n20832), .A2(n20821), .B1(n20820), .B2(n20829), .ZN(
        P2_U3603) );
  AND2_X1 U23880 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20822) );
  NOR2_X1 U23881 ( .A1(n20823), .A2(n20822), .ZN(n20825) );
  MUX2_X1 U23882 ( .A(n20826), .B(n20825), .S(n20824), .Z(n20827) );
  AOI21_X1 U23883 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20828), .A(n20827), 
        .ZN(n20830) );
  AOI22_X1 U23884 ( .A1(n20832), .A2(n20831), .B1(n20830), .B2(n20829), .ZN(
        P2_U3604) );
  INV_X1 U23885 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20833) );
  AOI22_X1 U23886 ( .A1(n20862), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20833), 
        .B2(n20863), .ZN(P2_U3608) );
  INV_X1 U23887 ( .A(n20834), .ZN(n20839) );
  INV_X1 U23888 ( .A(n20835), .ZN(n20837) );
  NAND2_X1 U23889 ( .A1(n20837), .A2(n20836), .ZN(n20838) );
  OAI211_X1 U23890 ( .C1(n20841), .C2(n20840), .A(n20839), .B(n20838), .ZN(
        n20843) );
  MUX2_X1 U23891 ( .A(P2_MORE_REG_SCAN_IN), .B(n20843), .S(n20842), .Z(
        P2_U3609) );
  OR2_X1 U23892 ( .A1(n20845), .A2(n20844), .ZN(n20846) );
  OAI211_X1 U23893 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20848), .A(n20847), 
        .B(n20846), .ZN(n20861) );
  AOI21_X1 U23894 ( .B1(n20850), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n20849), 
        .ZN(n20858) );
  NOR3_X1 U23895 ( .A1(n20853), .A2(n20851), .A3(n10286), .ZN(n20856) );
  INV_X1 U23896 ( .A(n11084), .ZN(n20852) );
  AOI21_X1 U23897 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20853), .A(n20852), 
        .ZN(n20855) );
  MUX2_X1 U23898 ( .A(n20856), .B(n20855), .S(n20854), .Z(n20857) );
  OAI21_X1 U23899 ( .B1(n20858), .B2(n20857), .A(n20861), .ZN(n20859) );
  OAI21_X1 U23900 ( .B1(n20861), .B2(n20860), .A(n20859), .ZN(P2_U3610) );
  OAI22_X1 U23901 ( .A1(n20863), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20862), .ZN(n20864) );
  INV_X1 U23902 ( .A(n20864), .ZN(P2_U3611) );
  AOI21_X1 U23903 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21662), .A(n21661), 
        .ZN(n20871) );
  INV_X1 U23904 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20865) );
  AOI21_X1 U23905 ( .B1(n20871), .B2(n20865), .A(n21734), .ZN(P1_U2802) );
  OAI21_X1 U23906 ( .B1(n20867), .B2(n20866), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20868) );
  OAI21_X1 U23907 ( .B1(n20869), .B2(n21645), .A(n20868), .ZN(P1_U2803) );
  NOR2_X1 U23908 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20872) );
  OAI21_X1 U23909 ( .B1(n20872), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21746), .ZN(
        n20870) );
  OAI21_X1 U23910 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21746), .A(n20870), 
        .ZN(P1_U2804) );
  OAI21_X1 U23911 ( .B1(BS16), .B2(n20872), .A(n21724), .ZN(n21723) );
  OAI21_X1 U23912 ( .B1(n21724), .B2(n21880), .A(n21723), .ZN(P1_U2805) );
  INV_X1 U23913 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20874) );
  OAI21_X1 U23914 ( .B1(n20875), .B2(n20874), .A(n20873), .ZN(P1_U2806) );
  NOR4_X1 U23915 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20879) );
  NOR4_X1 U23916 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20878) );
  NOR4_X1 U23917 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20877) );
  NOR4_X1 U23918 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20876) );
  NAND4_X1 U23919 ( .A1(n20879), .A2(n20878), .A3(n20877), .A4(n20876), .ZN(
        n20885) );
  NOR4_X1 U23920 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20883) );
  AOI211_X1 U23921 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20882) );
  NOR4_X1 U23922 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20881) );
  NOR4_X1 U23923 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20880) );
  NAND4_X1 U23924 ( .A1(n20883), .A2(n20882), .A3(n20881), .A4(n20880), .ZN(
        n20884) );
  NOR2_X1 U23925 ( .A1(n20885), .A2(n20884), .ZN(n21732) );
  INV_X1 U23926 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21718) );
  NOR3_X1 U23927 ( .A1(P1_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P1_REIP_REG_0__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20887)
         );
  OAI21_X1 U23928 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20887), .A(n21732), .ZN(
        n20886) );
  OAI21_X1 U23929 ( .B1(n21732), .B2(n21718), .A(n20886), .ZN(P1_U2807) );
  INV_X1 U23930 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21725) );
  INV_X1 U23931 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21903) );
  AOI21_X1 U23932 ( .B1(n21725), .B2(n21903), .A(n20887), .ZN(n20888) );
  INV_X1 U23933 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21715) );
  INV_X1 U23934 ( .A(n21732), .ZN(n21727) );
  AOI22_X1 U23935 ( .A1(n21732), .A2(n20888), .B1(n21715), .B2(n21727), .ZN(
        P1_U2808) );
  NOR2_X1 U23936 ( .A1(n20938), .A2(n20889), .ZN(n20890) );
  AOI22_X1 U23937 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n20955), .B1(n20890), .B2(
        n21678), .ZN(n20899) );
  OAI22_X1 U23938 ( .A1(n20927), .A2(n20892), .B1(n21678), .B2(n20891), .ZN(
        n20893) );
  AOI211_X1 U23939 ( .C1(n20956), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20945), .B(n20893), .ZN(n20898) );
  INV_X1 U23940 ( .A(n20894), .ZN(n20895) );
  AOI22_X1 U23941 ( .A1(n20896), .A2(n20914), .B1(n20895), .B2(n20965), .ZN(
        n20897) );
  NAND3_X1 U23942 ( .A1(n20899), .A2(n20898), .A3(n20897), .ZN(P1_U2831) );
  NOR3_X1 U23943 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20905), .A3(n20923), .ZN(
        n20903) );
  OAI21_X1 U23944 ( .B1(n20901), .B2(n20900), .A(n20925), .ZN(n20902) );
  AOI211_X1 U23945 ( .C1(n20955), .C2(P1_EBX_REG_7__SCAN_IN), .A(n20903), .B(
        n20902), .ZN(n20911) );
  OAI21_X1 U23946 ( .B1(n20940), .B2(n20938), .A(n20904), .ZN(n20937) );
  AOI21_X1 U23947 ( .B1(n20959), .B2(n20905), .A(n20937), .ZN(n20922) );
  OAI222_X1 U23948 ( .A1(n20908), .A2(n20907), .B1(n21674), .B2(n20922), .C1(
        n20906), .C2(n20952), .ZN(n20909) );
  INV_X1 U23949 ( .A(n20909), .ZN(n20910) );
  OAI211_X1 U23950 ( .C1(n20927), .C2(n20912), .A(n20911), .B(n20910), .ZN(
        P1_U2833) );
  INV_X1 U23951 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21672) );
  INV_X1 U23952 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21670) );
  NOR3_X1 U23953 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n21670), .A3(n20923), .ZN(
        n20913) );
  AOI211_X1 U23954 ( .C1(n20956), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20945), .B(n20913), .ZN(n20920) );
  AOI22_X1 U23955 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n20955), .B1(n20954), .B2(
        n20970), .ZN(n20919) );
  NAND2_X1 U23956 ( .A1(n20971), .A2(n20914), .ZN(n20918) );
  INV_X1 U23957 ( .A(n20915), .ZN(n20916) );
  NAND2_X1 U23958 ( .A1(n20965), .A2(n20916), .ZN(n20917) );
  OAI21_X1 U23959 ( .B1(n20922), .B2(n21672), .A(n20921), .ZN(P1_U2834) );
  INV_X1 U23960 ( .A(n20923), .ZN(n20924) );
  AOI22_X1 U23961 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n20955), .B1(n20924), .B2(
        n21670), .ZN(n20933) );
  OAI21_X1 U23962 ( .B1(n20927), .B2(n20926), .A(n20925), .ZN(n20930) );
  AOI22_X1 U23963 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20956), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20937), .ZN(n20928) );
  INV_X1 U23964 ( .A(n20928), .ZN(n20929) );
  AOI211_X1 U23965 ( .C1(n20931), .C2(n20950), .A(n20930), .B(n20929), .ZN(
        n20932) );
  OAI211_X1 U23966 ( .C1(n20934), .C2(n20952), .A(n20933), .B(n20932), .ZN(
        P1_U2835) );
  OAI21_X1 U23967 ( .B1(n14450), .B2(n20935), .A(n14956), .ZN(n20936) );
  INV_X1 U23968 ( .A(n20936), .ZN(n21010) );
  AOI22_X1 U23969 ( .A1(n20954), .A2(n21010), .B1(P1_REIP_REG_4__SCAN_IN), 
        .B2(n20937), .ZN(n20947) );
  NOR3_X1 U23970 ( .A1(n20940), .A2(n20939), .A3(n20938), .ZN(n20941) );
  AOI21_X1 U23971 ( .B1(n20958), .B2(n20942), .A(n20941), .ZN(n20943) );
  INV_X1 U23972 ( .A(n20943), .ZN(n20944) );
  AOI211_X1 U23973 ( .C1(n20956), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20945), .B(n20944), .ZN(n20946) );
  OAI211_X1 U23974 ( .C1(n20977), .C2(n20948), .A(n20947), .B(n20946), .ZN(
        n20949) );
  AOI21_X1 U23975 ( .B1(n20999), .B2(n20950), .A(n20949), .ZN(n20951) );
  OAI21_X1 U23976 ( .B1(n21005), .B2(n20952), .A(n20951), .ZN(P1_U2836) );
  AOI21_X1 U23977 ( .B1(n20959), .B2(n21725), .A(n20953), .ZN(n20969) );
  INV_X1 U23978 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21665) );
  AOI22_X1 U23979 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(n20955), .B1(n20954), .B2(
        n21026), .ZN(n20968) );
  AOI22_X1 U23980 ( .A1(n20958), .A2(n20957), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20956), .ZN(n20961) );
  NAND3_X1 U23981 ( .A1(n20959), .A2(P1_REIP_REG_1__SCAN_IN), .A3(n21665), 
        .ZN(n20960) );
  OAI211_X1 U23982 ( .C1(n20963), .C2(n20962), .A(n20961), .B(n20960), .ZN(
        n20964) );
  AOI21_X1 U23983 ( .B1(n20966), .B2(n20965), .A(n20964), .ZN(n20967) );
  OAI211_X1 U23984 ( .C1(n20969), .C2(n21665), .A(n20968), .B(n20967), .ZN(
        P1_U2838) );
  AOI22_X1 U23985 ( .A1(n20971), .A2(n20975), .B1(n20974), .B2(n20970), .ZN(
        n20972) );
  OAI21_X1 U23986 ( .B1(n20978), .B2(n20973), .A(n20972), .ZN(P1_U2866) );
  AOI22_X1 U23987 ( .A1(n20999), .A2(n20975), .B1(n20974), .B2(n21010), .ZN(
        n20976) );
  OAI21_X1 U23988 ( .B1(n20978), .B2(n20977), .A(n20976), .ZN(P1_U2868) );
  AOI22_X1 U23989 ( .A1(n20980), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20979), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20981) );
  OAI21_X1 U23990 ( .B1(n21907), .B2(n20985), .A(n20981), .ZN(P1_U2923) );
  INV_X1 U23991 ( .A(P1_LWORD_REG_12__SCAN_IN), .ZN(n22002) );
  INV_X1 U23992 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n20984) );
  OAI22_X1 U23993 ( .A1(n20985), .A2(n20984), .B1(n20983), .B2(n20982), .ZN(
        n20986) );
  INV_X1 U23994 ( .A(n20986), .ZN(n20987) );
  OAI21_X1 U23995 ( .B1(n22002), .B2(n14160), .A(n20987), .ZN(P1_U2924) );
  AOI22_X1 U23996 ( .A1(n20989), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20988), .ZN(n20991) );
  NAND2_X1 U23997 ( .A1(n20991), .A2(n20990), .ZN(P1_U2965) );
  AOI22_X1 U23998 ( .A1(n20992), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n21051), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n21004) );
  INV_X1 U23999 ( .A(n20993), .ZN(n20996) );
  INV_X1 U24000 ( .A(n20994), .ZN(n20995) );
  NAND2_X1 U24001 ( .A1(n20996), .A2(n20995), .ZN(n20997) );
  NAND2_X1 U24002 ( .A1(n20998), .A2(n20997), .ZN(n21013) );
  INV_X1 U24003 ( .A(n21013), .ZN(n21002) );
  AOI22_X1 U24004 ( .A1(n21002), .A2(n21001), .B1(n21000), .B2(n20999), .ZN(
        n21003) );
  OAI211_X1 U24005 ( .C1(n21006), .C2(n21005), .A(n21004), .B(n21003), .ZN(
        P1_U2995) );
  NOR2_X1 U24006 ( .A1(n21008), .A2(n21007), .ZN(n21025) );
  NOR2_X1 U24007 ( .A1(n21025), .A2(n21009), .ZN(n21022) );
  AOI22_X1 U24008 ( .A1(n21051), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n21027), 
        .B2(n21010), .ZN(n21017) );
  AOI211_X1 U24009 ( .C1(n21018), .C2(n21023), .A(n21011), .B(n21024), .ZN(
        n21015) );
  NOR2_X1 U24010 ( .A1(n21013), .A2(n21012), .ZN(n21014) );
  NOR2_X1 U24011 ( .A1(n21015), .A2(n21014), .ZN(n21016) );
  OAI211_X1 U24012 ( .C1(n21022), .C2(n21018), .A(n21017), .B(n21016), .ZN(
        P1_U3027) );
  AOI222_X1 U24013 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n21051), .B1(n21027), 
        .B2(n21020), .C1(n21042), .C2(n21019), .ZN(n21021) );
  OAI221_X1 U24014 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21024), .C1(
        n21023), .C2(n21022), .A(n21021), .ZN(P1_U3028) );
  AOI21_X1 U24015 ( .B1(n21027), .B2(n21026), .A(n21025), .ZN(n21039) );
  NAND3_X1 U24016 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21028), .ZN(n21029) );
  OAI211_X1 U24017 ( .C1(n21031), .C2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n21030), .B(n21029), .ZN(n21032) );
  AOI22_X1 U24018 ( .A1(n21033), .A2(n21042), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21032), .ZN(n21038) );
  NAND2_X1 U24019 ( .A1(n21051), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n21037) );
  NAND3_X1 U24020 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21035), .A3(
        n21034), .ZN(n21036) );
  NAND4_X1 U24021 ( .A1(n21039), .A2(n21038), .A3(n21037), .A4(n21036), .ZN(
        P1_U3029) );
  NOR3_X1 U24022 ( .A1(n21041), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n21040), .ZN(n21050) );
  AND3_X1 U24023 ( .A1(n21044), .A2(n21043), .A3(n21042), .ZN(n21049) );
  AOI21_X1 U24024 ( .B1(n21047), .B2(n21046), .A(n21045), .ZN(n21048) );
  NOR3_X1 U24025 ( .A1(n21050), .A2(n21049), .A3(n21048), .ZN(n21053) );
  NAND2_X1 U24026 ( .A1(n21051), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21052) );
  OAI211_X1 U24027 ( .C1(n21055), .C2(n21054), .A(n21053), .B(n21052), .ZN(
        P1_U3030) );
  NOR2_X1 U24028 ( .A1(n21057), .A2(n21056), .ZN(P1_U3032) );
  INV_X1 U24029 ( .A(n21058), .ZN(n21071) );
  OAI22_X1 U24030 ( .A1(n21059), .A2(n21102), .B1(n14993), .B2(n21104), .ZN(
        n21597) );
  INV_X1 U24031 ( .A(n21597), .ZN(n21442) );
  INV_X1 U24032 ( .A(n21595), .ZN(n21267) );
  OAI22_X1 U24033 ( .A1(n21631), .A2(n21442), .B1(n21090), .B2(n21267), .ZN(
        n21061) );
  INV_X1 U24034 ( .A(n21061), .ZN(n21066) );
  INV_X1 U24035 ( .A(n21062), .ZN(n21063) );
  OAI22_X1 U24036 ( .A1(n21064), .A2(n21102), .B1(n15032), .B2(n21104), .ZN(
        n21478) );
  AOI22_X1 U24037 ( .A1(n21596), .A2(n21110), .B1(n21135), .B2(n21478), .ZN(
        n21065) );
  OAI211_X1 U24038 ( .C1(n21071), .C2(n13203), .A(n21066), .B(n21065), .ZN(
        P1_U3034) );
  OAI22_X1 U24039 ( .A1(n21067), .A2(n21102), .B1(n15024), .B2(n21104), .ZN(
        n21482) );
  INV_X1 U24040 ( .A(n21482), .ZN(n21606) );
  OAI22_X2 U24041 ( .A1(n21068), .A2(n21102), .B1(n14989), .B2(n21104), .ZN(
        n21603) );
  INV_X1 U24042 ( .A(n21603), .ZN(n21445) );
  INV_X1 U24043 ( .A(n21601), .ZN(n21069) );
  OAI22_X1 U24044 ( .A1(n21631), .A2(n21445), .B1(n21090), .B2(n21069), .ZN(
        n21070) );
  INV_X1 U24045 ( .A(n21070), .ZN(n21075) );
  INV_X1 U24046 ( .A(n21072), .ZN(n21073) );
  AOI22_X1 U24047 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n21058), .B1(
        n21602), .B2(n21110), .ZN(n21074) );
  OAI211_X1 U24048 ( .C1(n21606), .C2(n21132), .A(n21075), .B(n21074), .ZN(
        P1_U3035) );
  INV_X1 U24049 ( .A(DATAI_19_), .ZN(n21076) );
  OAI22_X1 U24050 ( .A1(n16594), .A2(n21102), .B1(n21076), .B2(n21104), .ZN(
        n21609) );
  INV_X1 U24051 ( .A(n21609), .ZN(n21560) );
  OAI22_X2 U24052 ( .A1(n21077), .A2(n21102), .B1(n14983), .B2(n21104), .ZN(
        n21557) );
  NAND2_X1 U24053 ( .A1(n12177), .A2(n21105), .ZN(n21402) );
  AOI22_X1 U24054 ( .A1(n21638), .A2(n21557), .B1(n21107), .B2(n21607), .ZN(
        n21080) );
  AOI22_X1 U24055 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n21058), .B1(
        n21608), .B2(n21110), .ZN(n21079) );
  OAI211_X1 U24056 ( .C1(n21560), .C2(n21132), .A(n21080), .B(n21079), .ZN(
        P1_U3036) );
  OAI22_X1 U24057 ( .A1(n15016), .A2(n21104), .B1(n21081), .B2(n21102), .ZN(
        n21489) );
  OAI22_X2 U24058 ( .A1(n21082), .A2(n21102), .B1(n14977), .B2(n21104), .ZN(
        n21615) );
  INV_X1 U24059 ( .A(n21615), .ZN(n21450) );
  INV_X1 U24060 ( .A(n21613), .ZN(n21275) );
  OAI22_X1 U24061 ( .A1(n21631), .A2(n21450), .B1(n21090), .B2(n21275), .ZN(
        n21083) );
  INV_X1 U24062 ( .A(n21083), .ZN(n21087) );
  INV_X1 U24063 ( .A(n21084), .ZN(n21085) );
  AOI22_X1 U24064 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n21058), .B1(
        n21614), .B2(n21110), .ZN(n21086) );
  OAI211_X1 U24065 ( .C1(n21618), .C2(n21132), .A(n21087), .B(n21086), .ZN(
        P1_U3037) );
  OAI22_X1 U24066 ( .A1(n15011), .A2(n21104), .B1(n21088), .B2(n21102), .ZN(
        n21621) );
  OAI22_X1 U24067 ( .A1(n21089), .A2(n21102), .B1(n14972), .B2(n21104), .ZN(
        n21563) );
  INV_X1 U24068 ( .A(n21563), .ZN(n21624) );
  NAND2_X1 U24069 ( .A1(n12186), .A2(n21105), .ZN(n21408) );
  OAI22_X1 U24070 ( .A1(n21631), .A2(n21624), .B1(n21090), .B2(n21408), .ZN(
        n21091) );
  INV_X1 U24071 ( .A(n21091), .ZN(n21095) );
  INV_X1 U24072 ( .A(n21092), .ZN(n21093) );
  AOI22_X1 U24073 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n21058), .B1(
        n21620), .B2(n21110), .ZN(n21094) );
  OAI211_X1 U24074 ( .C1(n21566), .C2(n21132), .A(n21095), .B(n21094), .ZN(
        P1_U3038) );
  OAI22_X1 U24075 ( .A1(n21096), .A2(n21102), .B1(n15007), .B2(n21104), .ZN(
        n21496) );
  OAI22_X2 U24076 ( .A1(n16509), .A2(n21102), .B1(n14967), .B2(n21104), .ZN(
        n21627) );
  AOI22_X1 U24077 ( .A1(n21638), .A2(n21627), .B1(n21107), .B2(n21625), .ZN(
        n21100) );
  INV_X1 U24078 ( .A(n21097), .ZN(n21098) );
  AOI22_X1 U24079 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n21058), .B1(
        n21626), .B2(n21110), .ZN(n21099) );
  OAI211_X1 U24080 ( .C1(n21632), .C2(n21132), .A(n21100), .B(n21099), .ZN(
        P1_U3039) );
  OAI22_X1 U24081 ( .A1(n21101), .A2(n21102), .B1(n15003), .B2(n21104), .ZN(
        n21637) );
  INV_X1 U24082 ( .A(n21637), .ZN(n21576) );
  INV_X1 U24083 ( .A(DATAI_31_), .ZN(n21928) );
  OAI22_X2 U24084 ( .A1(n21928), .A2(n21104), .B1(n21103), .B2(n21102), .ZN(
        n21571) );
  NAND2_X1 U24085 ( .A1(n21106), .A2(n21105), .ZN(n21417) );
  AOI22_X1 U24086 ( .A1(n21638), .A2(n21571), .B1(n21107), .B2(n21633), .ZN(
        n21112) );
  INV_X1 U24087 ( .A(n21108), .ZN(n21109) );
  AOI22_X1 U24088 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n21058), .B1(
        n21636), .B2(n21110), .ZN(n21111) );
  OAI211_X1 U24089 ( .C1(n21576), .C2(n21132), .A(n21112), .B(n21111), .ZN(
        P1_U3040) );
  NOR2_X1 U24090 ( .A1(n21509), .A2(n21113), .ZN(n21133) );
  AOI21_X1 U24091 ( .B1(n21173), .B2(n21510), .A(n21133), .ZN(n21115) );
  OAI22_X1 U24092 ( .A1(n21115), .A2(n21579), .B1(n21113), .B2(n21647), .ZN(
        n21134) );
  AOI22_X1 U24093 ( .A1(n21584), .A2(n21134), .B1(n21583), .B2(n21133), .ZN(
        n21119) );
  INV_X1 U24094 ( .A(n21113), .ZN(n21117) );
  OAI21_X1 U24095 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21474), .A(
        n21114), .ZN(n21431) );
  OAI211_X1 U24096 ( .C1(n21175), .C2(n21880), .A(n21517), .B(n21115), .ZN(
        n21116) );
  AOI22_X1 U24097 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n21136), .B1(
        n21135), .B2(n21549), .ZN(n21118) );
  OAI211_X1 U24098 ( .C1(n21552), .C2(n21160), .A(n21119), .B(n21118), .ZN(
        P1_U3041) );
  INV_X1 U24099 ( .A(n21478), .ZN(n21600) );
  AOI22_X1 U24100 ( .A1(n21596), .A2(n21134), .B1(n21595), .B2(n21133), .ZN(
        n21121) );
  AOI22_X1 U24101 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21136), .B1(
        n21135), .B2(n21597), .ZN(n21120) );
  OAI211_X1 U24102 ( .C1(n21600), .C2(n21160), .A(n21121), .B(n21120), .ZN(
        P1_U3042) );
  AOI22_X1 U24103 ( .A1(n21602), .A2(n21134), .B1(n21601), .B2(n21133), .ZN(
        n21123) );
  AOI22_X1 U24104 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n21136), .B1(
        n21135), .B2(n21603), .ZN(n21122) );
  OAI211_X1 U24105 ( .C1(n21606), .C2(n21160), .A(n21123), .B(n21122), .ZN(
        P1_U3043) );
  AOI22_X1 U24106 ( .A1(n21608), .A2(n21134), .B1(n21607), .B2(n21133), .ZN(
        n21125) );
  AOI22_X1 U24107 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n21136), .B1(
        n21135), .B2(n21557), .ZN(n21124) );
  OAI211_X1 U24108 ( .C1(n21560), .C2(n21160), .A(n21125), .B(n21124), .ZN(
        P1_U3044) );
  AOI22_X1 U24109 ( .A1(n21614), .A2(n21134), .B1(n21613), .B2(n21133), .ZN(
        n21127) );
  AOI22_X1 U24110 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n21136), .B1(
        n21135), .B2(n21615), .ZN(n21126) );
  OAI211_X1 U24111 ( .C1(n21618), .C2(n21160), .A(n21127), .B(n21126), .ZN(
        P1_U3045) );
  AOI22_X1 U24112 ( .A1(n21620), .A2(n21134), .B1(n21619), .B2(n21133), .ZN(
        n21129) );
  AOI22_X1 U24113 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n21136), .B1(
        n21135), .B2(n21563), .ZN(n21128) );
  OAI211_X1 U24114 ( .C1(n21566), .C2(n21160), .A(n21129), .B(n21128), .ZN(
        P1_U3046) );
  INV_X1 U24115 ( .A(n21627), .ZN(n21455) );
  AOI22_X1 U24116 ( .A1(n21626), .A2(n21134), .B1(n21625), .B2(n21133), .ZN(
        n21131) );
  AOI22_X1 U24117 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n21136), .B1(
        n21167), .B2(n21496), .ZN(n21130) );
  OAI211_X1 U24118 ( .C1(n21455), .C2(n21132), .A(n21131), .B(n21130), .ZN(
        P1_U3047) );
  AOI22_X1 U24119 ( .A1(n21636), .A2(n21134), .B1(n21633), .B2(n21133), .ZN(
        n21138) );
  AOI22_X1 U24120 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n21136), .B1(
        n21135), .B2(n21571), .ZN(n21137) );
  OAI211_X1 U24121 ( .C1(n21576), .C2(n21160), .A(n21138), .B(n21137), .ZN(
        P1_U3048) );
  INV_X1 U24122 ( .A(n21538), .ZN(n21140) );
  NAND2_X1 U24123 ( .A1(n21160), .A2(n21517), .ZN(n21141) );
  OAI21_X1 U24124 ( .B1(n21196), .B2(n21141), .A(n21464), .ZN(n21143) );
  NOR2_X1 U24125 ( .A1(n21142), .A2(n21384), .ZN(n21146) );
  OR2_X1 U24126 ( .A1(n21386), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21262) );
  INV_X1 U24127 ( .A(n21262), .ZN(n21144) );
  NAND3_X1 U24128 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21385), .A3(
        n21389), .ZN(n21177) );
  NOR2_X1 U24129 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21177), .ZN(
        n21166) );
  AOI22_X1 U24130 ( .A1(n21196), .A2(n21591), .B1(n21583), .B2(n21166), .ZN(
        n21149) );
  INV_X1 U24131 ( .A(n21143), .ZN(n21147) );
  INV_X1 U24132 ( .A(n21166), .ZN(n21159) );
  NOR2_X1 U24133 ( .A1(n21144), .A2(n21647), .ZN(n21259) );
  AOI211_X1 U24134 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n21159), .A(n21259), 
        .B(n21330), .ZN(n21145) );
  AOI22_X1 U24135 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21549), .ZN(n21148) );
  OAI211_X1 U24136 ( .C1(n21171), .C2(n21477), .A(n21149), .B(n21148), .ZN(
        P1_U3049) );
  INV_X1 U24137 ( .A(n21596), .ZN(n21481) );
  OAI22_X1 U24138 ( .A1(n21160), .A2(n21442), .B1(n21159), .B2(n21267), .ZN(
        n21150) );
  INV_X1 U24139 ( .A(n21150), .ZN(n21152) );
  AOI22_X1 U24140 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n21168), .B1(
        n21196), .B2(n21478), .ZN(n21151) );
  OAI211_X1 U24141 ( .C1(n21171), .C2(n21481), .A(n21152), .B(n21151), .ZN(
        P1_U3050) );
  AOI22_X1 U24142 ( .A1(n21196), .A2(n21482), .B1(n21166), .B2(n21601), .ZN(
        n21154) );
  AOI22_X1 U24143 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21603), .ZN(n21153) );
  OAI211_X1 U24144 ( .C1(n21171), .C2(n21485), .A(n21154), .B(n21153), .ZN(
        P1_U3051) );
  INV_X1 U24145 ( .A(n21608), .ZN(n21488) );
  AOI22_X1 U24146 ( .A1(n21196), .A2(n21609), .B1(n21166), .B2(n21607), .ZN(
        n21156) );
  AOI22_X1 U24147 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21557), .ZN(n21155) );
  OAI211_X1 U24148 ( .C1(n21171), .C2(n21488), .A(n21156), .B(n21155), .ZN(
        P1_U3052) );
  INV_X1 U24149 ( .A(n21614), .ZN(n21492) );
  AOI22_X1 U24150 ( .A1(n21196), .A2(n21489), .B1(n21166), .B2(n21613), .ZN(
        n21158) );
  AOI22_X1 U24151 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21615), .ZN(n21157) );
  OAI211_X1 U24152 ( .C1(n21171), .C2(n21492), .A(n21158), .B(n21157), .ZN(
        P1_U3053) );
  INV_X1 U24153 ( .A(n21620), .ZN(n21495) );
  OAI22_X1 U24154 ( .A1(n21160), .A2(n21624), .B1(n21159), .B2(n21408), .ZN(
        n21161) );
  INV_X1 U24155 ( .A(n21161), .ZN(n21163) );
  AOI22_X1 U24156 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n21168), .B1(
        n21196), .B2(n21621), .ZN(n21162) );
  OAI211_X1 U24157 ( .C1(n21171), .C2(n21495), .A(n21163), .B(n21162), .ZN(
        P1_U3054) );
  INV_X1 U24158 ( .A(n21626), .ZN(n21499) );
  AOI22_X1 U24159 ( .A1(n21196), .A2(n21496), .B1(n21166), .B2(n21625), .ZN(
        n21165) );
  AOI22_X1 U24160 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21627), .ZN(n21164) );
  OAI211_X1 U24161 ( .C1(n21171), .C2(n21499), .A(n21165), .B(n21164), .ZN(
        P1_U3055) );
  AOI22_X1 U24162 ( .A1(n21196), .A2(n21637), .B1(n21166), .B2(n21633), .ZN(
        n21170) );
  AOI22_X1 U24163 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n21168), .B1(
        n21167), .B2(n21571), .ZN(n21169) );
  OAI211_X1 U24164 ( .C1(n21171), .C2(n21505), .A(n21170), .B(n21169), .ZN(
        P1_U3056) );
  NAND2_X1 U24165 ( .A1(n13156), .A2(n21172), .ZN(n21426) );
  INV_X1 U24166 ( .A(n21426), .ZN(n21577) );
  NOR2_X1 U24167 ( .A1(n21424), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21195) );
  AOI21_X1 U24168 ( .B1(n21173), .B2(n21577), .A(n21195), .ZN(n21176) );
  AOI21_X1 U24169 ( .B1(n21175), .B2(n21517), .A(n21430), .ZN(n21180) );
  OAI22_X1 U24170 ( .A1(n21647), .A2(n21177), .B1(n21176), .B2(n21180), .ZN(
        n21174) );
  AOI22_X1 U24171 ( .A1(n21224), .A2(n21591), .B1(n21583), .B2(n21195), .ZN(
        n21182) );
  INV_X1 U24172 ( .A(n21176), .ZN(n21179) );
  AOI21_X1 U24173 ( .B1(n21579), .B2(n21177), .A(n21431), .ZN(n21178) );
  AOI22_X1 U24174 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n21197), .B1(
        n21196), .B2(n21549), .ZN(n21181) );
  OAI211_X1 U24175 ( .C1(n21200), .C2(n21477), .A(n21182), .B(n21181), .ZN(
        P1_U3057) );
  AOI22_X1 U24176 ( .A1(n21196), .A2(n21597), .B1(n21195), .B2(n21595), .ZN(
        n21184) );
  AOI22_X1 U24177 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n21197), .B1(
        n21224), .B2(n21478), .ZN(n21183) );
  OAI211_X1 U24178 ( .C1(n21200), .C2(n21481), .A(n21184), .B(n21183), .ZN(
        P1_U3058) );
  AOI22_X1 U24179 ( .A1(n21196), .A2(n21603), .B1(n21601), .B2(n21195), .ZN(
        n21186) );
  AOI22_X1 U24180 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n21197), .B1(
        n21224), .B2(n21482), .ZN(n21185) );
  OAI211_X1 U24181 ( .C1(n21200), .C2(n21485), .A(n21186), .B(n21185), .ZN(
        P1_U3059) );
  AOI22_X1 U24182 ( .A1(n21224), .A2(n21609), .B1(n21607), .B2(n21195), .ZN(
        n21188) );
  AOI22_X1 U24183 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n21197), .B1(
        n21196), .B2(n21557), .ZN(n21187) );
  OAI211_X1 U24184 ( .C1(n21200), .C2(n21488), .A(n21188), .B(n21187), .ZN(
        P1_U3060) );
  AOI22_X1 U24185 ( .A1(n21224), .A2(n21489), .B1(n21613), .B2(n21195), .ZN(
        n21190) );
  AOI22_X1 U24186 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n21197), .B1(
        n21196), .B2(n21615), .ZN(n21189) );
  OAI211_X1 U24187 ( .C1(n21200), .C2(n21492), .A(n21190), .B(n21189), .ZN(
        P1_U3061) );
  AOI22_X1 U24188 ( .A1(n21224), .A2(n21621), .B1(n21195), .B2(n21619), .ZN(
        n21192) );
  AOI22_X1 U24189 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n21197), .B1(
        n21196), .B2(n21563), .ZN(n21191) );
  OAI211_X1 U24190 ( .C1(n21200), .C2(n21495), .A(n21192), .B(n21191), .ZN(
        P1_U3062) );
  AOI22_X1 U24191 ( .A1(n21224), .A2(n21496), .B1(n21625), .B2(n21195), .ZN(
        n21194) );
  AOI22_X1 U24192 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n21197), .B1(
        n21196), .B2(n21627), .ZN(n21193) );
  OAI211_X1 U24193 ( .C1(n21200), .C2(n21499), .A(n21194), .B(n21193), .ZN(
        P1_U3063) );
  AOI22_X1 U24194 ( .A1(n21224), .A2(n21637), .B1(n21633), .B2(n21195), .ZN(
        n21199) );
  AOI22_X1 U24195 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n21197), .B1(
        n21196), .B2(n21571), .ZN(n21198) );
  OAI211_X1 U24196 ( .C1(n21200), .C2(n21505), .A(n21199), .B(n21198), .ZN(
        P1_U3064) );
  NOR2_X1 U24197 ( .A1(n15520), .A2(n21201), .ZN(n21295) );
  NAND3_X1 U24198 ( .A1(n21295), .A2(n21517), .A3(n21384), .ZN(n21202) );
  NAND3_X1 U24199 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21385), .A3(
        n21468), .ZN(n21231) );
  NOR2_X1 U24200 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21231), .ZN(
        n21222) );
  AOI22_X1 U24201 ( .A1(n21584), .A2(n21223), .B1(n21583), .B2(n21222), .ZN(
        n21209) );
  INV_X1 U24202 ( .A(n21245), .ZN(n21252) );
  OAI21_X1 U24203 ( .B1(n21224), .B2(n21252), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21205) );
  NAND2_X1 U24204 ( .A1(n21295), .A2(n21384), .ZN(n21204) );
  AOI21_X1 U24205 ( .B1(n21205), .B2(n21204), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21207) );
  AOI22_X1 U24206 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21549), .ZN(n21208) );
  OAI211_X1 U24207 ( .C1(n21552), .C2(n21245), .A(n21209), .B(n21208), .ZN(
        P1_U3065) );
  AOI22_X1 U24208 ( .A1(n21596), .A2(n21223), .B1(n21595), .B2(n21222), .ZN(
        n21211) );
  AOI22_X1 U24209 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21597), .ZN(n21210) );
  OAI211_X1 U24210 ( .C1(n21600), .C2(n21245), .A(n21211), .B(n21210), .ZN(
        P1_U3066) );
  AOI22_X1 U24211 ( .A1(n21602), .A2(n21223), .B1(n21601), .B2(n21222), .ZN(
        n21213) );
  AOI22_X1 U24212 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21603), .ZN(n21212) );
  OAI211_X1 U24213 ( .C1(n21606), .C2(n21245), .A(n21213), .B(n21212), .ZN(
        P1_U3067) );
  AOI22_X1 U24214 ( .A1(n21608), .A2(n21223), .B1(n21607), .B2(n21222), .ZN(
        n21215) );
  AOI22_X1 U24215 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21557), .ZN(n21214) );
  OAI211_X1 U24216 ( .C1(n21560), .C2(n21245), .A(n21215), .B(n21214), .ZN(
        P1_U3068) );
  AOI22_X1 U24217 ( .A1(n21614), .A2(n21223), .B1(n21613), .B2(n21222), .ZN(
        n21217) );
  AOI22_X1 U24218 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21615), .ZN(n21216) );
  OAI211_X1 U24219 ( .C1(n21618), .C2(n21245), .A(n21217), .B(n21216), .ZN(
        P1_U3069) );
  AOI22_X1 U24220 ( .A1(n21620), .A2(n21223), .B1(n21619), .B2(n21222), .ZN(
        n21219) );
  AOI22_X1 U24221 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21563), .ZN(n21218) );
  OAI211_X1 U24222 ( .C1(n21566), .C2(n21245), .A(n21219), .B(n21218), .ZN(
        P1_U3070) );
  AOI22_X1 U24223 ( .A1(n21626), .A2(n21223), .B1(n21625), .B2(n21222), .ZN(
        n21221) );
  AOI22_X1 U24224 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21627), .ZN(n21220) );
  OAI211_X1 U24225 ( .C1(n21632), .C2(n21245), .A(n21221), .B(n21220), .ZN(
        P1_U3071) );
  AOI22_X1 U24226 ( .A1(n21636), .A2(n21223), .B1(n21633), .B2(n21222), .ZN(
        n21227) );
  AOI22_X1 U24227 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n21225), .B1(
        n21224), .B2(n21571), .ZN(n21226) );
  OAI211_X1 U24228 ( .C1(n21576), .C2(n21245), .A(n21227), .B(n21226), .ZN(
        P1_U3072) );
  INV_X1 U24229 ( .A(n21549), .ZN(n21594) );
  NOR2_X1 U24230 ( .A1(n21509), .A2(n21231), .ZN(n21250) );
  AOI21_X1 U24231 ( .B1(n21295), .B2(n21510), .A(n21250), .ZN(n21232) );
  OAI22_X1 U24232 ( .A1(n21232), .A2(n21579), .B1(n21231), .B2(n21647), .ZN(
        n21251) );
  AOI22_X1 U24233 ( .A1(n21584), .A2(n21251), .B1(n21583), .B2(n21250), .ZN(
        n21236) );
  INV_X1 U24234 ( .A(n21228), .ZN(n21230) );
  NAND2_X1 U24235 ( .A1(n21229), .A2(n21517), .ZN(n21586) );
  NAND3_X1 U24236 ( .A1(n21230), .A2(n21464), .A3(n21586), .ZN(n21233) );
  AOI22_X1 U24237 ( .A1(n21233), .A2(n21232), .B1(n21231), .B2(n21579), .ZN(
        n21234) );
  NAND2_X1 U24238 ( .A1(n21588), .A2(n21234), .ZN(n21253) );
  AOI22_X1 U24239 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21253), .B1(
        n21289), .B2(n21591), .ZN(n21235) );
  OAI211_X1 U24240 ( .C1(n21594), .C2(n21245), .A(n21236), .B(n21235), .ZN(
        P1_U3073) );
  AOI22_X1 U24241 ( .A1(n21596), .A2(n21251), .B1(n21595), .B2(n21250), .ZN(
        n21238) );
  AOI22_X1 U24242 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21253), .B1(
        n21289), .B2(n21478), .ZN(n21237) );
  OAI211_X1 U24243 ( .C1(n21442), .C2(n21245), .A(n21238), .B(n21237), .ZN(
        P1_U3074) );
  AOI22_X1 U24244 ( .A1(n21602), .A2(n21251), .B1(n21601), .B2(n21250), .ZN(
        n21240) );
  AOI22_X1 U24245 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21253), .B1(
        n21289), .B2(n21482), .ZN(n21239) );
  OAI211_X1 U24246 ( .C1(n21445), .C2(n21245), .A(n21240), .B(n21239), .ZN(
        P1_U3075) );
  INV_X1 U24247 ( .A(n21557), .ZN(n21612) );
  AOI22_X1 U24248 ( .A1(n21608), .A2(n21251), .B1(n21607), .B2(n21250), .ZN(
        n21242) );
  AOI22_X1 U24249 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21253), .B1(
        n21289), .B2(n21609), .ZN(n21241) );
  OAI211_X1 U24250 ( .C1(n21612), .C2(n21245), .A(n21242), .B(n21241), .ZN(
        P1_U3076) );
  AOI22_X1 U24251 ( .A1(n21614), .A2(n21251), .B1(n21613), .B2(n21250), .ZN(
        n21244) );
  AOI22_X1 U24252 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21253), .B1(
        n21289), .B2(n21489), .ZN(n21243) );
  OAI211_X1 U24253 ( .C1(n21450), .C2(n21245), .A(n21244), .B(n21243), .ZN(
        P1_U3077) );
  AOI22_X1 U24254 ( .A1(n21620), .A2(n21251), .B1(n21619), .B2(n21250), .ZN(
        n21247) );
  AOI22_X1 U24255 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21563), .ZN(n21246) );
  OAI211_X1 U24256 ( .C1(n21566), .C2(n21287), .A(n21247), .B(n21246), .ZN(
        P1_U3078) );
  AOI22_X1 U24257 ( .A1(n21626), .A2(n21251), .B1(n21625), .B2(n21250), .ZN(
        n21249) );
  AOI22_X1 U24258 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21627), .ZN(n21248) );
  OAI211_X1 U24259 ( .C1(n21632), .C2(n21287), .A(n21249), .B(n21248), .ZN(
        P1_U3079) );
  AOI22_X1 U24260 ( .A1(n21636), .A2(n21251), .B1(n21633), .B2(n21250), .ZN(
        n21255) );
  AOI22_X1 U24261 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21571), .ZN(n21254) );
  OAI211_X1 U24262 ( .C1(n21576), .C2(n21287), .A(n21255), .B(n21254), .ZN(
        P1_U3080) );
  INV_X1 U24263 ( .A(n21583), .ZN(n21256) );
  INV_X1 U24264 ( .A(n21301), .ZN(n21296) );
  NOR2_X1 U24265 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21296), .ZN(
        n21288) );
  INV_X1 U24266 ( .A(n21288), .ZN(n21282) );
  OAI22_X1 U24267 ( .A1(n21287), .A2(n21594), .B1(n21256), .B2(n21282), .ZN(
        n21257) );
  INV_X1 U24268 ( .A(n21257), .ZN(n21266) );
  INV_X1 U24269 ( .A(n21325), .ZN(n21312) );
  NOR3_X1 U24270 ( .A1(n21312), .A2(n21289), .A3(n21579), .ZN(n21258) );
  INV_X1 U24271 ( .A(n21464), .ZN(n21513) );
  NOR2_X1 U24272 ( .A1(n21258), .A2(n21513), .ZN(n21264) );
  INV_X1 U24273 ( .A(n21264), .ZN(n21260) );
  NAND2_X1 U24274 ( .A1(n21295), .A2(n21540), .ZN(n21263) );
  AOI21_X1 U24275 ( .B1(n21260), .B2(n21263), .A(n21259), .ZN(n21261) );
  AOI22_X1 U24276 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n21291), .B1(
        n21584), .B2(n21290), .ZN(n21265) );
  OAI211_X1 U24277 ( .C1(n21552), .C2(n21325), .A(n21266), .B(n21265), .ZN(
        P1_U3081) );
  OAI22_X1 U24278 ( .A1(n21287), .A2(n21442), .B1(n21267), .B2(n21282), .ZN(
        n21268) );
  INV_X1 U24279 ( .A(n21268), .ZN(n21270) );
  AOI22_X1 U24280 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n21291), .B1(
        n21596), .B2(n21290), .ZN(n21269) );
  OAI211_X1 U24281 ( .C1(n21600), .C2(n21325), .A(n21270), .B(n21269), .ZN(
        P1_U3082) );
  AOI22_X1 U24282 ( .A1(n21312), .A2(n21482), .B1(n21601), .B2(n21288), .ZN(
        n21272) );
  AOI22_X1 U24283 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n21291), .B1(
        n21602), .B2(n21290), .ZN(n21271) );
  OAI211_X1 U24284 ( .C1(n21445), .C2(n21287), .A(n21272), .B(n21271), .ZN(
        P1_U3083) );
  AOI22_X1 U24285 ( .A1(n21289), .A2(n21557), .B1(n21607), .B2(n21288), .ZN(
        n21274) );
  AOI22_X1 U24286 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n21291), .B1(
        n21608), .B2(n21290), .ZN(n21273) );
  OAI211_X1 U24287 ( .C1(n21560), .C2(n21325), .A(n21274), .B(n21273), .ZN(
        P1_U3084) );
  OAI22_X1 U24288 ( .A1(n21287), .A2(n21450), .B1(n21275), .B2(n21282), .ZN(
        n21276) );
  INV_X1 U24289 ( .A(n21276), .ZN(n21278) );
  AOI22_X1 U24290 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n21291), .B1(
        n21614), .B2(n21290), .ZN(n21277) );
  OAI211_X1 U24291 ( .C1(n21618), .C2(n21325), .A(n21278), .B(n21277), .ZN(
        P1_U3085) );
  OAI22_X1 U24292 ( .A1(n21287), .A2(n21624), .B1(n21408), .B2(n21282), .ZN(
        n21279) );
  INV_X1 U24293 ( .A(n21279), .ZN(n21281) );
  AOI22_X1 U24294 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n21291), .B1(
        n21620), .B2(n21290), .ZN(n21280) );
  OAI211_X1 U24295 ( .C1(n21566), .C2(n21325), .A(n21281), .B(n21280), .ZN(
        P1_U3086) );
  INV_X1 U24296 ( .A(n21625), .ZN(n21283) );
  OAI22_X1 U24297 ( .A1(n21325), .A2(n21632), .B1(n21283), .B2(n21282), .ZN(
        n21284) );
  INV_X1 U24298 ( .A(n21284), .ZN(n21286) );
  AOI22_X1 U24299 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n21291), .B1(
        n21626), .B2(n21290), .ZN(n21285) );
  OAI211_X1 U24300 ( .C1(n21455), .C2(n21287), .A(n21286), .B(n21285), .ZN(
        P1_U3087) );
  AOI22_X1 U24301 ( .A1(n21289), .A2(n21571), .B1(n21633), .B2(n21288), .ZN(
        n21293) );
  AOI22_X1 U24302 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n21291), .B1(
        n21636), .B2(n21290), .ZN(n21292) );
  OAI211_X1 U24303 ( .C1(n21576), .C2(n21325), .A(n21293), .B(n21292), .ZN(
        P1_U3088) );
  INV_X1 U24304 ( .A(n21294), .ZN(n21320) );
  AOI21_X1 U24305 ( .B1(n21295), .B2(n21577), .A(n21320), .ZN(n21298) );
  OAI22_X1 U24306 ( .A1(n21298), .A2(n21579), .B1(n21647), .B2(n21296), .ZN(
        n21321) );
  AOI22_X1 U24307 ( .A1(n21584), .A2(n21321), .B1(n21320), .B2(n21583), .ZN(
        n21305) );
  INV_X1 U24308 ( .A(n21297), .ZN(n21585) );
  INV_X1 U24309 ( .A(n21586), .ZN(n21299) );
  OAI21_X1 U24310 ( .B1(n21585), .B2(n21299), .A(n21298), .ZN(n21300) );
  NAND2_X1 U24311 ( .A1(n21303), .A2(n21302), .ZN(n21315) );
  AOI22_X1 U24312 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n21322), .B1(
        n21351), .B2(n21591), .ZN(n21304) );
  OAI211_X1 U24313 ( .C1(n21594), .C2(n21325), .A(n21305), .B(n21304), .ZN(
        P1_U3089) );
  AOI22_X1 U24314 ( .A1(n21596), .A2(n21321), .B1(n21320), .B2(n21595), .ZN(
        n21307) );
  AOI22_X1 U24315 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n21322), .B1(
        n21351), .B2(n21478), .ZN(n21306) );
  OAI211_X1 U24316 ( .C1(n21442), .C2(n21325), .A(n21307), .B(n21306), .ZN(
        P1_U3090) );
  AOI22_X1 U24317 ( .A1(n21602), .A2(n21321), .B1(n21320), .B2(n21601), .ZN(
        n21309) );
  AOI22_X1 U24318 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n21322), .B1(
        n21351), .B2(n21482), .ZN(n21308) );
  OAI211_X1 U24319 ( .C1(n21445), .C2(n21325), .A(n21309), .B(n21308), .ZN(
        P1_U3091) );
  AOI22_X1 U24320 ( .A1(n21608), .A2(n21321), .B1(n21320), .B2(n21607), .ZN(
        n21311) );
  AOI22_X1 U24321 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n21322), .B1(
        n21351), .B2(n21609), .ZN(n21310) );
  OAI211_X1 U24322 ( .C1(n21612), .C2(n21325), .A(n21311), .B(n21310), .ZN(
        P1_U3092) );
  AOI22_X1 U24323 ( .A1(n21614), .A2(n21321), .B1(n21320), .B2(n21613), .ZN(
        n21314) );
  AOI22_X1 U24324 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n21322), .B1(
        n21312), .B2(n21615), .ZN(n21313) );
  OAI211_X1 U24325 ( .C1(n21618), .C2(n21315), .A(n21314), .B(n21313), .ZN(
        P1_U3093) );
  AOI22_X1 U24326 ( .A1(n21620), .A2(n21321), .B1(n21320), .B2(n21619), .ZN(
        n21317) );
  AOI22_X1 U24327 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n21322), .B1(
        n21351), .B2(n21621), .ZN(n21316) );
  OAI211_X1 U24328 ( .C1(n21624), .C2(n21325), .A(n21317), .B(n21316), .ZN(
        P1_U3094) );
  AOI22_X1 U24329 ( .A1(n21626), .A2(n21321), .B1(n21320), .B2(n21625), .ZN(
        n21319) );
  AOI22_X1 U24330 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n21322), .B1(
        n21351), .B2(n21496), .ZN(n21318) );
  OAI211_X1 U24331 ( .C1(n21455), .C2(n21325), .A(n21319), .B(n21318), .ZN(
        P1_U3095) );
  INV_X1 U24332 ( .A(n21571), .ZN(n21643) );
  AOI22_X1 U24333 ( .A1(n21636), .A2(n21321), .B1(n21320), .B2(n21633), .ZN(
        n21324) );
  AOI22_X1 U24334 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n21322), .B1(
        n21351), .B2(n21637), .ZN(n21323) );
  OAI211_X1 U24335 ( .C1(n21643), .C2(n21325), .A(n21324), .B(n21323), .ZN(
        P1_U3096) );
  NAND2_X1 U24336 ( .A1(n21327), .A2(n15520), .ZN(n21427) );
  INV_X1 U24337 ( .A(n21427), .ZN(n21355) );
  NAND3_X1 U24338 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21389), .A3(
        n21468), .ZN(n21356) );
  NOR2_X1 U24339 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21356), .ZN(
        n21349) );
  AOI21_X1 U24340 ( .B1(n21355), .B2(n21384), .A(n21349), .ZN(n21332) );
  AND2_X1 U24341 ( .A1(n21328), .A2(n21386), .ZN(n21466) );
  INV_X1 U24342 ( .A(n21466), .ZN(n21470) );
  OAI22_X1 U24343 ( .A1(n21332), .A2(n21579), .B1(n21329), .B2(n21470), .ZN(
        n21350) );
  AOI22_X1 U24344 ( .A1(n21584), .A2(n21350), .B1(n21583), .B2(n21349), .ZN(
        n21336) );
  INV_X1 U24345 ( .A(n21330), .ZN(n21391) );
  INV_X1 U24346 ( .A(n21380), .ZN(n21331) );
  OAI21_X1 U24347 ( .B1(n21331), .B2(n21351), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21333) );
  NAND2_X1 U24348 ( .A1(n21333), .A2(n21332), .ZN(n21334) );
  AOI22_X1 U24349 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21549), .ZN(n21335) );
  OAI211_X1 U24350 ( .C1(n21552), .C2(n21380), .A(n21336), .B(n21335), .ZN(
        P1_U3097) );
  AOI22_X1 U24351 ( .A1(n21596), .A2(n21350), .B1(n21595), .B2(n21349), .ZN(
        n21338) );
  AOI22_X1 U24352 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21597), .ZN(n21337) );
  OAI211_X1 U24353 ( .C1(n21600), .C2(n21380), .A(n21338), .B(n21337), .ZN(
        P1_U3098) );
  AOI22_X1 U24354 ( .A1(n21602), .A2(n21350), .B1(n21601), .B2(n21349), .ZN(
        n21340) );
  AOI22_X1 U24355 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21603), .ZN(n21339) );
  OAI211_X1 U24356 ( .C1(n21606), .C2(n21380), .A(n21340), .B(n21339), .ZN(
        P1_U3099) );
  AOI22_X1 U24357 ( .A1(n21608), .A2(n21350), .B1(n21607), .B2(n21349), .ZN(
        n21342) );
  AOI22_X1 U24358 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21557), .ZN(n21341) );
  OAI211_X1 U24359 ( .C1(n21560), .C2(n21380), .A(n21342), .B(n21341), .ZN(
        P1_U3100) );
  AOI22_X1 U24360 ( .A1(n21614), .A2(n21350), .B1(n21613), .B2(n21349), .ZN(
        n21344) );
  AOI22_X1 U24361 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21615), .ZN(n21343) );
  OAI211_X1 U24362 ( .C1(n21618), .C2(n21380), .A(n21344), .B(n21343), .ZN(
        P1_U3101) );
  AOI22_X1 U24363 ( .A1(n21620), .A2(n21350), .B1(n21619), .B2(n21349), .ZN(
        n21346) );
  AOI22_X1 U24364 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21563), .ZN(n21345) );
  OAI211_X1 U24365 ( .C1(n21566), .C2(n21380), .A(n21346), .B(n21345), .ZN(
        P1_U3102) );
  AOI22_X1 U24366 ( .A1(n21626), .A2(n21350), .B1(n21625), .B2(n21349), .ZN(
        n21348) );
  AOI22_X1 U24367 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21627), .ZN(n21347) );
  OAI211_X1 U24368 ( .C1(n21632), .C2(n21380), .A(n21348), .B(n21347), .ZN(
        P1_U3103) );
  AOI22_X1 U24369 ( .A1(n21636), .A2(n21350), .B1(n21633), .B2(n21349), .ZN(
        n21354) );
  AOI22_X1 U24370 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21571), .ZN(n21353) );
  OAI211_X1 U24371 ( .C1(n21576), .C2(n21380), .A(n21354), .B(n21353), .ZN(
        P1_U3104) );
  NOR2_X1 U24372 ( .A1(n21509), .A2(n21356), .ZN(n21375) );
  AOI21_X1 U24373 ( .B1(n21355), .B2(n21510), .A(n21375), .ZN(n21357) );
  OAI22_X1 U24374 ( .A1(n21357), .A2(n21579), .B1(n21356), .B2(n21647), .ZN(
        n21376) );
  AOI22_X1 U24375 ( .A1(n21584), .A2(n21376), .B1(n21583), .B2(n21375), .ZN(
        n21362) );
  INV_X1 U24376 ( .A(n21356), .ZN(n21359) );
  OAI211_X1 U24377 ( .C1(n21437), .C2(n21880), .A(n21517), .B(n21357), .ZN(
        n21358) );
  AOI22_X1 U24378 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21377), .B1(
        n21419), .B2(n21591), .ZN(n21361) );
  OAI211_X1 U24379 ( .C1(n21594), .C2(n21380), .A(n21362), .B(n21361), .ZN(
        P1_U3105) );
  AOI22_X1 U24380 ( .A1(n21596), .A2(n21376), .B1(n21595), .B2(n21375), .ZN(
        n21364) );
  AOI22_X1 U24381 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21377), .B1(
        n21419), .B2(n21478), .ZN(n21363) );
  OAI211_X1 U24382 ( .C1(n21442), .C2(n21380), .A(n21364), .B(n21363), .ZN(
        P1_U3106) );
  AOI22_X1 U24383 ( .A1(n21602), .A2(n21376), .B1(n21601), .B2(n21375), .ZN(
        n21366) );
  AOI22_X1 U24384 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21377), .B1(
        n21419), .B2(n21482), .ZN(n21365) );
  OAI211_X1 U24385 ( .C1(n21445), .C2(n21380), .A(n21366), .B(n21365), .ZN(
        P1_U3107) );
  AOI22_X1 U24386 ( .A1(n21608), .A2(n21376), .B1(n21607), .B2(n21375), .ZN(
        n21368) );
  AOI22_X1 U24387 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21377), .B1(
        n21419), .B2(n21609), .ZN(n21367) );
  OAI211_X1 U24388 ( .C1(n21612), .C2(n21380), .A(n21368), .B(n21367), .ZN(
        P1_U3108) );
  AOI22_X1 U24389 ( .A1(n21614), .A2(n21376), .B1(n21613), .B2(n21375), .ZN(
        n21370) );
  AOI22_X1 U24390 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21377), .B1(
        n21419), .B2(n21489), .ZN(n21369) );
  OAI211_X1 U24391 ( .C1(n21450), .C2(n21380), .A(n21370), .B(n21369), .ZN(
        P1_U3109) );
  AOI22_X1 U24392 ( .A1(n21620), .A2(n21376), .B1(n21619), .B2(n21375), .ZN(
        n21372) );
  AOI22_X1 U24393 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21377), .B1(
        n21419), .B2(n21621), .ZN(n21371) );
  OAI211_X1 U24394 ( .C1(n21624), .C2(n21380), .A(n21372), .B(n21371), .ZN(
        P1_U3110) );
  AOI22_X1 U24395 ( .A1(n21626), .A2(n21376), .B1(n21625), .B2(n21375), .ZN(
        n21374) );
  AOI22_X1 U24396 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21377), .B1(
        n21419), .B2(n21496), .ZN(n21373) );
  OAI211_X1 U24397 ( .C1(n21455), .C2(n21380), .A(n21374), .B(n21373), .ZN(
        P1_U3111) );
  AOI22_X1 U24398 ( .A1(n21636), .A2(n21376), .B1(n21633), .B2(n21375), .ZN(
        n21379) );
  AOI22_X1 U24399 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21377), .B1(
        n21419), .B2(n21637), .ZN(n21378) );
  OAI211_X1 U24400 ( .C1(n21643), .C2(n21380), .A(n21379), .B(n21378), .ZN(
        P1_U3112) );
  INV_X1 U24401 ( .A(n21419), .ZN(n21382) );
  NAND3_X1 U24402 ( .A1(n21382), .A2(n21517), .A3(n21461), .ZN(n21383) );
  NAND2_X1 U24403 ( .A1(n21383), .A2(n21464), .ZN(n21394) );
  NOR2_X1 U24404 ( .A1(n21427), .A2(n21384), .ZN(n21390) );
  OR2_X1 U24405 ( .A1(n21386), .A2(n21385), .ZN(n21542) );
  INV_X1 U24406 ( .A(n21542), .ZN(n21387) );
  NAND3_X1 U24407 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n21389), .ZN(n21432) );
  NOR2_X1 U24408 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21432), .ZN(
        n21412) );
  AOI22_X1 U24409 ( .A1(n21419), .A2(n21549), .B1(n21583), .B2(n21412), .ZN(
        n21397) );
  INV_X1 U24410 ( .A(n21390), .ZN(n21393) );
  NAND2_X1 U24411 ( .A1(n21542), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21546) );
  OAI211_X1 U24412 ( .C1(n21474), .C2(n21412), .A(n21546), .B(n21391), .ZN(
        n21392) );
  AOI21_X1 U24413 ( .B1(n21394), .B2(n21393), .A(n21392), .ZN(n21395) );
  INV_X1 U24414 ( .A(n21461), .ZN(n21413) );
  AOI22_X1 U24415 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21420), .B1(
        n21413), .B2(n21591), .ZN(n21396) );
  OAI211_X1 U24416 ( .C1(n21423), .C2(n21477), .A(n21397), .B(n21396), .ZN(
        P1_U3113) );
  AOI22_X1 U24417 ( .A1(n21413), .A2(n21478), .B1(n21595), .B2(n21412), .ZN(
        n21399) );
  AOI22_X1 U24418 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21420), .B1(
        n21419), .B2(n21597), .ZN(n21398) );
  OAI211_X1 U24419 ( .C1(n21423), .C2(n21481), .A(n21399), .B(n21398), .ZN(
        P1_U3114) );
  AOI22_X1 U24420 ( .A1(n21419), .A2(n21603), .B1(n21601), .B2(n21412), .ZN(
        n21401) );
  AOI22_X1 U24421 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21420), .B1(
        n21413), .B2(n21482), .ZN(n21400) );
  OAI211_X1 U24422 ( .C1(n21423), .C2(n21485), .A(n21401), .B(n21400), .ZN(
        P1_U3115) );
  INV_X1 U24423 ( .A(n21412), .ZN(n21416) );
  OAI22_X1 U24424 ( .A1(n21461), .A2(n21560), .B1(n21402), .B2(n21416), .ZN(
        n21403) );
  INV_X1 U24425 ( .A(n21403), .ZN(n21405) );
  AOI22_X1 U24426 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21420), .B1(
        n21419), .B2(n21557), .ZN(n21404) );
  OAI211_X1 U24427 ( .C1(n21423), .C2(n21488), .A(n21405), .B(n21404), .ZN(
        P1_U3116) );
  AOI22_X1 U24428 ( .A1(n21419), .A2(n21615), .B1(n21613), .B2(n21412), .ZN(
        n21407) );
  AOI22_X1 U24429 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21420), .B1(
        n21413), .B2(n21489), .ZN(n21406) );
  OAI211_X1 U24430 ( .C1(n21423), .C2(n21492), .A(n21407), .B(n21406), .ZN(
        P1_U3117) );
  OAI22_X1 U24431 ( .A1(n21461), .A2(n21566), .B1(n21408), .B2(n21416), .ZN(
        n21409) );
  INV_X1 U24432 ( .A(n21409), .ZN(n21411) );
  AOI22_X1 U24433 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21420), .B1(
        n21419), .B2(n21563), .ZN(n21410) );
  OAI211_X1 U24434 ( .C1(n21423), .C2(n21495), .A(n21411), .B(n21410), .ZN(
        P1_U3118) );
  AOI22_X1 U24435 ( .A1(n21419), .A2(n21627), .B1(n21625), .B2(n21412), .ZN(
        n21415) );
  AOI22_X1 U24436 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21420), .B1(
        n21413), .B2(n21496), .ZN(n21414) );
  OAI211_X1 U24437 ( .C1(n21423), .C2(n21499), .A(n21415), .B(n21414), .ZN(
        P1_U3119) );
  OAI22_X1 U24438 ( .A1(n21461), .A2(n21576), .B1(n21417), .B2(n21416), .ZN(
        n21418) );
  INV_X1 U24439 ( .A(n21418), .ZN(n21422) );
  AOI22_X1 U24440 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21420), .B1(
        n21419), .B2(n21571), .ZN(n21421) );
  OAI211_X1 U24441 ( .C1(n21423), .C2(n21505), .A(n21422), .B(n21421), .ZN(
        P1_U3120) );
  INV_X1 U24442 ( .A(n21424), .ZN(n21425) );
  NAND2_X1 U24443 ( .A1(n21425), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21429) );
  OAI21_X1 U24444 ( .B1(n21427), .B2(n21426), .A(n21429), .ZN(n21434) );
  INV_X1 U24445 ( .A(n21434), .ZN(n21428) );
  INV_X1 U24446 ( .A(n21429), .ZN(n21456) );
  AOI22_X1 U24447 ( .A1(n21584), .A2(n21457), .B1(n21583), .B2(n21456), .ZN(
        n21439) );
  AOI21_X1 U24448 ( .B1(n21437), .B2(n21517), .A(n21430), .ZN(n21435) );
  AOI21_X1 U24449 ( .B1(n21579), .B2(n21432), .A(n21431), .ZN(n21433) );
  NOR2_X4 U24450 ( .A1(n21437), .A2(n21436), .ZN(n21501) );
  AOI22_X1 U24451 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21458), .B1(
        n21501), .B2(n21591), .ZN(n21438) );
  OAI211_X1 U24452 ( .C1(n21594), .C2(n21461), .A(n21439), .B(n21438), .ZN(
        P1_U3121) );
  AOI22_X1 U24453 ( .A1(n21596), .A2(n21457), .B1(n21456), .B2(n21595), .ZN(
        n21441) );
  AOI22_X1 U24454 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21458), .B1(
        n21501), .B2(n21478), .ZN(n21440) );
  OAI211_X1 U24455 ( .C1(n21442), .C2(n21461), .A(n21441), .B(n21440), .ZN(
        P1_U3122) );
  AOI22_X1 U24456 ( .A1(n21602), .A2(n21457), .B1(n21456), .B2(n21601), .ZN(
        n21444) );
  AOI22_X1 U24457 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21458), .B1(
        n21501), .B2(n21482), .ZN(n21443) );
  OAI211_X1 U24458 ( .C1(n21445), .C2(n21461), .A(n21444), .B(n21443), .ZN(
        P1_U3123) );
  AOI22_X1 U24459 ( .A1(n21608), .A2(n21457), .B1(n21456), .B2(n21607), .ZN(
        n21447) );
  AOI22_X1 U24460 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21458), .B1(
        n21501), .B2(n21609), .ZN(n21446) );
  OAI211_X1 U24461 ( .C1(n21612), .C2(n21461), .A(n21447), .B(n21446), .ZN(
        P1_U3124) );
  AOI22_X1 U24462 ( .A1(n21614), .A2(n21457), .B1(n21456), .B2(n21613), .ZN(
        n21449) );
  AOI22_X1 U24463 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21458), .B1(
        n21501), .B2(n21489), .ZN(n21448) );
  OAI211_X1 U24464 ( .C1(n21450), .C2(n21461), .A(n21449), .B(n21448), .ZN(
        P1_U3125) );
  AOI22_X1 U24465 ( .A1(n21620), .A2(n21457), .B1(n21456), .B2(n21619), .ZN(
        n21452) );
  AOI22_X1 U24466 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21458), .B1(
        n21501), .B2(n21621), .ZN(n21451) );
  OAI211_X1 U24467 ( .C1(n21624), .C2(n21461), .A(n21452), .B(n21451), .ZN(
        P1_U3126) );
  AOI22_X1 U24468 ( .A1(n21626), .A2(n21457), .B1(n21456), .B2(n21625), .ZN(
        n21454) );
  AOI22_X1 U24469 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21458), .B1(
        n21501), .B2(n21496), .ZN(n21453) );
  OAI211_X1 U24470 ( .C1(n21455), .C2(n21461), .A(n21454), .B(n21453), .ZN(
        P1_U3127) );
  AOI22_X1 U24471 ( .A1(n21636), .A2(n21457), .B1(n21456), .B2(n21633), .ZN(
        n21460) );
  AOI22_X1 U24472 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21458), .B1(
        n21501), .B2(n21637), .ZN(n21459) );
  OAI211_X1 U24473 ( .C1(n21643), .C2(n21461), .A(n21460), .B(n21459), .ZN(
        P1_U3128) );
  INV_X1 U24474 ( .A(n21534), .ZN(n21463) );
  NAND2_X1 U24475 ( .A1(n21463), .A2(n21517), .ZN(n21465) );
  OAI21_X1 U24476 ( .B1(n21465), .B2(n21501), .A(n21464), .ZN(n21472) );
  OR2_X1 U24477 ( .A1(n15520), .A2(n10611), .ZN(n21508) );
  NOR2_X1 U24478 ( .A1(n21508), .A2(n21540), .ZN(n21469) );
  INV_X1 U24479 ( .A(n21541), .ZN(n21467) );
  NAND3_X1 U24480 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n21468), .ZN(n21511) );
  NOR2_X1 U24481 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21511), .ZN(
        n21500) );
  AOI22_X1 U24482 ( .A1(n21534), .A2(n21591), .B1(n21583), .B2(n21500), .ZN(
        n21476) );
  INV_X1 U24483 ( .A(n21469), .ZN(n21471) );
  AOI22_X1 U24484 ( .A1(n21472), .A2(n21471), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21470), .ZN(n21473) );
  AOI22_X1 U24485 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21502), .B1(
        n21501), .B2(n21549), .ZN(n21475) );
  OAI211_X1 U24486 ( .C1(n21506), .C2(n21477), .A(n21476), .B(n21475), .ZN(
        P1_U3129) );
  AOI22_X1 U24487 ( .A1(n21534), .A2(n21478), .B1(n21595), .B2(n21500), .ZN(
        n21480) );
  AOI22_X1 U24488 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21502), .B1(
        n21501), .B2(n21597), .ZN(n21479) );
  OAI211_X1 U24489 ( .C1(n21506), .C2(n21481), .A(n21480), .B(n21479), .ZN(
        P1_U3130) );
  AOI22_X1 U24490 ( .A1(n21534), .A2(n21482), .B1(n21601), .B2(n21500), .ZN(
        n21484) );
  AOI22_X1 U24491 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21502), .B1(
        n21501), .B2(n21603), .ZN(n21483) );
  OAI211_X1 U24492 ( .C1(n21506), .C2(n21485), .A(n21484), .B(n21483), .ZN(
        P1_U3131) );
  AOI22_X1 U24493 ( .A1(n21534), .A2(n21609), .B1(n21607), .B2(n21500), .ZN(
        n21487) );
  AOI22_X1 U24494 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21502), .B1(
        n21501), .B2(n21557), .ZN(n21486) );
  OAI211_X1 U24495 ( .C1(n21506), .C2(n21488), .A(n21487), .B(n21486), .ZN(
        P1_U3132) );
  AOI22_X1 U24496 ( .A1(n21534), .A2(n21489), .B1(n21613), .B2(n21500), .ZN(
        n21491) );
  AOI22_X1 U24497 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21502), .B1(
        n21501), .B2(n21615), .ZN(n21490) );
  OAI211_X1 U24498 ( .C1(n21506), .C2(n21492), .A(n21491), .B(n21490), .ZN(
        P1_U3133) );
  AOI22_X1 U24499 ( .A1(n21534), .A2(n21621), .B1(n21619), .B2(n21500), .ZN(
        n21494) );
  AOI22_X1 U24500 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21502), .B1(
        n21501), .B2(n21563), .ZN(n21493) );
  OAI211_X1 U24501 ( .C1(n21506), .C2(n21495), .A(n21494), .B(n21493), .ZN(
        P1_U3134) );
  AOI22_X1 U24502 ( .A1(n21534), .A2(n21496), .B1(n21625), .B2(n21500), .ZN(
        n21498) );
  AOI22_X1 U24503 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21502), .B1(
        n21501), .B2(n21627), .ZN(n21497) );
  OAI211_X1 U24504 ( .C1(n21506), .C2(n21499), .A(n21498), .B(n21497), .ZN(
        P1_U3135) );
  AOI22_X1 U24505 ( .A1(n21534), .A2(n21637), .B1(n21633), .B2(n21500), .ZN(
        n21504) );
  AOI22_X1 U24506 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21502), .B1(
        n21501), .B2(n21571), .ZN(n21503) );
  OAI211_X1 U24507 ( .C1(n21506), .C2(n21505), .A(n21504), .B(n21503), .ZN(
        P1_U3136) );
  NOR2_X1 U24508 ( .A1(n21509), .A2(n21511), .ZN(n21532) );
  AOI21_X1 U24509 ( .B1(n21578), .B2(n21510), .A(n21532), .ZN(n21512) );
  OAI22_X1 U24510 ( .A1(n21512), .A2(n21579), .B1(n21511), .B2(n21647), .ZN(
        n21533) );
  AOI22_X1 U24511 ( .A1(n21584), .A2(n21533), .B1(n21583), .B2(n21532), .ZN(
        n21519) );
  INV_X1 U24512 ( .A(n21511), .ZN(n21516) );
  OAI21_X1 U24513 ( .B1(n21514), .B2(n21513), .A(n21512), .ZN(n21515) );
  AOI22_X1 U24514 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21535), .B1(
        n21534), .B2(n21549), .ZN(n21518) );
  OAI211_X1 U24515 ( .C1(n21552), .C2(n21543), .A(n21519), .B(n21518), .ZN(
        P1_U3137) );
  AOI22_X1 U24516 ( .A1(n21596), .A2(n21533), .B1(n21595), .B2(n21532), .ZN(
        n21521) );
  AOI22_X1 U24517 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21535), .B1(
        n21534), .B2(n21597), .ZN(n21520) );
  OAI211_X1 U24518 ( .C1(n21600), .C2(n21543), .A(n21521), .B(n21520), .ZN(
        P1_U3138) );
  AOI22_X1 U24519 ( .A1(n21602), .A2(n21533), .B1(n21601), .B2(n21532), .ZN(
        n21523) );
  AOI22_X1 U24520 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21535), .B1(
        n21534), .B2(n21603), .ZN(n21522) );
  OAI211_X1 U24521 ( .C1(n21606), .C2(n21543), .A(n21523), .B(n21522), .ZN(
        P1_U3139) );
  AOI22_X1 U24522 ( .A1(n21608), .A2(n21533), .B1(n21607), .B2(n21532), .ZN(
        n21525) );
  AOI22_X1 U24523 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21535), .B1(
        n21534), .B2(n21557), .ZN(n21524) );
  OAI211_X1 U24524 ( .C1(n21560), .C2(n21543), .A(n21525), .B(n21524), .ZN(
        P1_U3140) );
  AOI22_X1 U24525 ( .A1(n21614), .A2(n21533), .B1(n21613), .B2(n21532), .ZN(
        n21527) );
  AOI22_X1 U24526 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21535), .B1(
        n21534), .B2(n21615), .ZN(n21526) );
  OAI211_X1 U24527 ( .C1(n21618), .C2(n21543), .A(n21527), .B(n21526), .ZN(
        P1_U3141) );
  AOI22_X1 U24528 ( .A1(n21620), .A2(n21533), .B1(n21619), .B2(n21532), .ZN(
        n21529) );
  AOI22_X1 U24529 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21535), .B1(
        n21534), .B2(n21563), .ZN(n21528) );
  OAI211_X1 U24530 ( .C1(n21566), .C2(n21543), .A(n21529), .B(n21528), .ZN(
        P1_U3142) );
  AOI22_X1 U24531 ( .A1(n21626), .A2(n21533), .B1(n21625), .B2(n21532), .ZN(
        n21531) );
  AOI22_X1 U24532 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21535), .B1(
        n21534), .B2(n21627), .ZN(n21530) );
  OAI211_X1 U24533 ( .C1(n21632), .C2(n21543), .A(n21531), .B(n21530), .ZN(
        P1_U3143) );
  AOI22_X1 U24534 ( .A1(n21636), .A2(n21533), .B1(n21633), .B2(n21532), .ZN(
        n21537) );
  AOI22_X1 U24535 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21535), .B1(
        n21534), .B2(n21571), .ZN(n21536) );
  OAI211_X1 U24536 ( .C1(n21576), .C2(n21543), .A(n21537), .B(n21536), .ZN(
        P1_U3144) );
  NAND2_X1 U24537 ( .A1(n21578), .A2(n21540), .ZN(n21544) );
  OAI22_X1 U24538 ( .A1(n21544), .A2(n21579), .B1(n21542), .B2(n21541), .ZN(
        n21570) );
  NOR2_X1 U24539 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21587), .ZN(
        n21569) );
  AOI22_X1 U24540 ( .A1(n21584), .A2(n21570), .B1(n21583), .B2(n21569), .ZN(
        n21551) );
  OAI21_X1 U24541 ( .B1(n21628), .B2(n21572), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21545) );
  AOI21_X1 U24542 ( .B1(n21545), .B2(n21544), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21548) );
  AOI22_X1 U24543 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21573), .B1(
        n21572), .B2(n21549), .ZN(n21550) );
  OAI211_X1 U24544 ( .C1(n21552), .C2(n21642), .A(n21551), .B(n21550), .ZN(
        P1_U3145) );
  AOI22_X1 U24545 ( .A1(n21596), .A2(n21570), .B1(n21595), .B2(n21569), .ZN(
        n21554) );
  AOI22_X1 U24546 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21573), .B1(
        n21572), .B2(n21597), .ZN(n21553) );
  OAI211_X1 U24547 ( .C1(n21600), .C2(n21642), .A(n21554), .B(n21553), .ZN(
        P1_U3146) );
  AOI22_X1 U24548 ( .A1(n21602), .A2(n21570), .B1(n21601), .B2(n21569), .ZN(
        n21556) );
  AOI22_X1 U24549 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21573), .B1(
        n21572), .B2(n21603), .ZN(n21555) );
  OAI211_X1 U24550 ( .C1(n21606), .C2(n21642), .A(n21556), .B(n21555), .ZN(
        P1_U3147) );
  AOI22_X1 U24551 ( .A1(n21608), .A2(n21570), .B1(n21607), .B2(n21569), .ZN(
        n21559) );
  AOI22_X1 U24552 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21573), .B1(
        n21572), .B2(n21557), .ZN(n21558) );
  OAI211_X1 U24553 ( .C1(n21560), .C2(n21642), .A(n21559), .B(n21558), .ZN(
        P1_U3148) );
  AOI22_X1 U24554 ( .A1(n21614), .A2(n21570), .B1(n21613), .B2(n21569), .ZN(
        n21562) );
  AOI22_X1 U24555 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21573), .B1(
        n21572), .B2(n21615), .ZN(n21561) );
  OAI211_X1 U24556 ( .C1(n21618), .C2(n21642), .A(n21562), .B(n21561), .ZN(
        P1_U3149) );
  AOI22_X1 U24557 ( .A1(n21620), .A2(n21570), .B1(n21619), .B2(n21569), .ZN(
        n21565) );
  AOI22_X1 U24558 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21573), .B1(
        n21572), .B2(n21563), .ZN(n21564) );
  OAI211_X1 U24559 ( .C1(n21566), .C2(n21642), .A(n21565), .B(n21564), .ZN(
        P1_U3150) );
  AOI22_X1 U24560 ( .A1(n21626), .A2(n21570), .B1(n21625), .B2(n21569), .ZN(
        n21568) );
  AOI22_X1 U24561 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21573), .B1(
        n21572), .B2(n21627), .ZN(n21567) );
  OAI211_X1 U24562 ( .C1(n21632), .C2(n21642), .A(n21568), .B(n21567), .ZN(
        P1_U3151) );
  AOI22_X1 U24563 ( .A1(n21636), .A2(n21570), .B1(n21633), .B2(n21569), .ZN(
        n21575) );
  AOI22_X1 U24564 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21573), .B1(
        n21572), .B2(n21571), .ZN(n21574) );
  OAI211_X1 U24565 ( .C1(n21576), .C2(n21642), .A(n21575), .B(n21574), .ZN(
        P1_U3152) );
  NAND2_X1 U24566 ( .A1(n21578), .A2(n21577), .ZN(n21580) );
  AOI21_X1 U24567 ( .B1(n21580), .B2(n21582), .A(n21579), .ZN(n21590) );
  INV_X1 U24568 ( .A(n21590), .ZN(n21581) );
  INV_X1 U24569 ( .A(n21582), .ZN(n21634) );
  AOI22_X1 U24570 ( .A1(n21584), .A2(n21635), .B1(n21634), .B2(n21583), .ZN(
        n21593) );
  AOI21_X1 U24571 ( .B1(n21587), .B2(n21586), .A(n21585), .ZN(n21589) );
  AOI22_X1 U24572 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21639), .B1(
        n21638), .B2(n21591), .ZN(n21592) );
  OAI211_X1 U24573 ( .C1(n21594), .C2(n21642), .A(n21593), .B(n21592), .ZN(
        P1_U3153) );
  AOI22_X1 U24574 ( .A1(n21596), .A2(n21635), .B1(n21634), .B2(n21595), .ZN(
        n21599) );
  AOI22_X1 U24575 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21639), .B1(
        n21628), .B2(n21597), .ZN(n21598) );
  OAI211_X1 U24576 ( .C1(n21600), .C2(n21631), .A(n21599), .B(n21598), .ZN(
        P1_U3154) );
  AOI22_X1 U24577 ( .A1(n21602), .A2(n21635), .B1(n21634), .B2(n21601), .ZN(
        n21605) );
  AOI22_X1 U24578 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21639), .B1(
        n21628), .B2(n21603), .ZN(n21604) );
  OAI211_X1 U24579 ( .C1(n21606), .C2(n21631), .A(n21605), .B(n21604), .ZN(
        P1_U3155) );
  AOI22_X1 U24580 ( .A1(n21608), .A2(n21635), .B1(n21634), .B2(n21607), .ZN(
        n21611) );
  AOI22_X1 U24581 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21639), .B1(
        n21638), .B2(n21609), .ZN(n21610) );
  OAI211_X1 U24582 ( .C1(n21612), .C2(n21642), .A(n21611), .B(n21610), .ZN(
        P1_U3156) );
  AOI22_X1 U24583 ( .A1(n21614), .A2(n21635), .B1(n21634), .B2(n21613), .ZN(
        n21617) );
  AOI22_X1 U24584 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21639), .B1(
        n21628), .B2(n21615), .ZN(n21616) );
  OAI211_X1 U24585 ( .C1(n21618), .C2(n21631), .A(n21617), .B(n21616), .ZN(
        P1_U3157) );
  AOI22_X1 U24586 ( .A1(n21620), .A2(n21635), .B1(n21634), .B2(n21619), .ZN(
        n21623) );
  AOI22_X1 U24587 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21639), .B1(
        n21638), .B2(n21621), .ZN(n21622) );
  OAI211_X1 U24588 ( .C1(n21624), .C2(n21642), .A(n21623), .B(n21622), .ZN(
        P1_U3158) );
  AOI22_X1 U24589 ( .A1(n21626), .A2(n21635), .B1(n21634), .B2(n21625), .ZN(
        n21630) );
  AOI22_X1 U24590 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21639), .B1(
        n21628), .B2(n21627), .ZN(n21629) );
  OAI211_X1 U24591 ( .C1(n21632), .C2(n21631), .A(n21630), .B(n21629), .ZN(
        P1_U3159) );
  AOI22_X1 U24592 ( .A1(n21636), .A2(n21635), .B1(n21634), .B2(n21633), .ZN(
        n21641) );
  AOI22_X1 U24593 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21639), .B1(
        n21638), .B2(n21637), .ZN(n21640) );
  OAI211_X1 U24594 ( .C1(n21643), .C2(n21642), .A(n21641), .B(n21640), .ZN(
        P1_U3160) );
  NOR2_X1 U24595 ( .A1(n21645), .A2(n21644), .ZN(n21648) );
  OAI21_X1 U24596 ( .B1(n21648), .B2(n21647), .A(n21646), .ZN(P1_U3163) );
  INV_X1 U24597 ( .A(n21724), .ZN(n21721) );
  AND2_X1 U24598 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21721), .ZN(
        P1_U3164) );
  AND2_X1 U24599 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21721), .ZN(
        P1_U3165) );
  AND2_X1 U24600 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21721), .ZN(
        P1_U3166) );
  AND2_X1 U24601 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21721), .ZN(
        P1_U3167) );
  AND2_X1 U24602 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21721), .ZN(
        P1_U3168) );
  AND2_X1 U24603 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21721), .ZN(
        P1_U3169) );
  AND2_X1 U24604 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21721), .ZN(
        P1_U3170) );
  AND2_X1 U24605 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21721), .ZN(
        P1_U3171) );
  AND2_X1 U24606 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21721), .ZN(
        P1_U3172) );
  AND2_X1 U24607 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21721), .ZN(
        P1_U3173) );
  INV_X1 U24608 ( .A(P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n22023) );
  NOR2_X1 U24609 ( .A1(n21724), .A2(n22023), .ZN(P1_U3174) );
  AND2_X1 U24610 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21721), .ZN(
        P1_U3175) );
  AND2_X1 U24611 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21721), .ZN(
        P1_U3176) );
  AND2_X1 U24612 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21721), .ZN(
        P1_U3177) );
  AND2_X1 U24613 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21721), .ZN(
        P1_U3178) );
  AND2_X1 U24614 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21721), .ZN(
        P1_U3179) );
  AND2_X1 U24615 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21721), .ZN(
        P1_U3180) );
  AND2_X1 U24616 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21721), .ZN(
        P1_U3181) );
  AND2_X1 U24617 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21721), .ZN(
        P1_U3182) );
  AND2_X1 U24618 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21721), .ZN(
        P1_U3183) );
  AND2_X1 U24619 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21721), .ZN(
        P1_U3184) );
  AND2_X1 U24620 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21721), .ZN(
        P1_U3185) );
  AND2_X1 U24621 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21721), .ZN(P1_U3186) );
  INV_X1 U24622 ( .A(P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21942) );
  NOR2_X1 U24623 ( .A1(n21724), .A2(n21942), .ZN(P1_U3187) );
  AND2_X1 U24624 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21721), .ZN(P1_U3188) );
  AND2_X1 U24625 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21721), .ZN(P1_U3189) );
  AND2_X1 U24626 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21721), .ZN(P1_U3190) );
  AND2_X1 U24627 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21721), .ZN(P1_U3191) );
  AND2_X1 U24628 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21721), .ZN(P1_U3192) );
  INV_X1 U24629 ( .A(P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21987) );
  NOR2_X1 U24630 ( .A1(n21724), .A2(n21987), .ZN(P1_U3193) );
  NAND2_X1 U24631 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21657), .ZN(n21655) );
  INV_X1 U24632 ( .A(n21655), .ZN(n21652) );
  OAI21_X1 U24633 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(HOLD), .ZN(n21649) );
  OAI211_X1 U24634 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n21656), .A(n21649), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21650) );
  INV_X1 U24635 ( .A(n21650), .ZN(n21651) );
  OAI22_X1 U24636 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21652), .B1(n21734), 
        .B2(n21651), .ZN(P1_U3194) );
  INV_X1 U24637 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21744) );
  OAI211_X1 U24638 ( .C1(NA), .C2(n21653), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n21662), .ZN(n21654) );
  OAI211_X1 U24639 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21744), .A(HOLD), .B(
        n21654), .ZN(n21660) );
  OAI211_X1 U24640 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21656), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21655), .ZN(n21659) );
  OR4_X1 U24641 ( .A1(n21744), .A2(n21661), .A3(n21657), .A4(NA), .ZN(n21658)
         );
  OAI211_X1 U24642 ( .C1(n21661), .C2(n21660), .A(n21659), .B(n21658), .ZN(
        P1_U3196) );
  NAND2_X1 U24643 ( .A1(n21734), .A2(n21662), .ZN(n21709) );
  INV_X1 U24644 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21663) );
  AND2_X1 U24645 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21734), .ZN(n21706) );
  INV_X1 U24646 ( .A(n21706), .ZN(n21713) );
  OAI222_X1 U24647 ( .A1(n21709), .A2(n21665), .B1(n21663), .B2(n21734), .C1(
        n21725), .C2(n21713), .ZN(P1_U3197) );
  INV_X1 U24648 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n21664) );
  OAI222_X1 U24649 ( .A1(n21713), .A2(n21665), .B1(n21664), .B2(n21734), .C1(
        n21989), .C2(n21709), .ZN(P1_U3198) );
  OAI222_X1 U24650 ( .A1(n21713), .A2(n21989), .B1(n21666), .B2(n21734), .C1(
        n21667), .C2(n21709), .ZN(P1_U3199) );
  INV_X1 U24651 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21668) );
  OAI222_X1 U24652 ( .A1(n21709), .A2(n21670), .B1(n21668), .B2(n21734), .C1(
        n21667), .C2(n21713), .ZN(P1_U3200) );
  INV_X1 U24653 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21669) );
  OAI222_X1 U24654 ( .A1(n21713), .A2(n21670), .B1(n21669), .B2(n21734), .C1(
        n21672), .C2(n21709), .ZN(P1_U3201) );
  INV_X1 U24655 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21671) );
  OAI222_X1 U24656 ( .A1(n21713), .A2(n21672), .B1(n21671), .B2(n21734), .C1(
        n21674), .C2(n21709), .ZN(P1_U3202) );
  INV_X1 U24657 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21673) );
  OAI222_X1 U24658 ( .A1(n21713), .A2(n21674), .B1(n21673), .B2(n21734), .C1(
        n21675), .C2(n21709), .ZN(P1_U3203) );
  INV_X1 U24659 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21676) );
  OAI222_X1 U24660 ( .A1(n21709), .A2(n21678), .B1(n21676), .B2(n21734), .C1(
        n21675), .C2(n21713), .ZN(P1_U3204) );
  INV_X1 U24661 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21677) );
  OAI222_X1 U24662 ( .A1(n21713), .A2(n21678), .B1(n21677), .B2(n21734), .C1(
        n21680), .C2(n21709), .ZN(P1_U3205) );
  INV_X1 U24663 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21679) );
  OAI222_X1 U24664 ( .A1(n21713), .A2(n21680), .B1(n21679), .B2(n21734), .C1(
        n21682), .C2(n21709), .ZN(P1_U3206) );
  AOI22_X1 U24665 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21746), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21705), .ZN(n21681) );
  OAI21_X1 U24666 ( .B1(n21682), .B2(n21713), .A(n21681), .ZN(P1_U3207) );
  AOI22_X1 U24667 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21746), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21706), .ZN(n21683) );
  OAI21_X1 U24668 ( .B1(n21685), .B2(n21709), .A(n21683), .ZN(P1_U3208) );
  INV_X1 U24669 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21684) );
  OAI222_X1 U24670 ( .A1(n21713), .A2(n21685), .B1(n21684), .B2(n21734), .C1(
        n21686), .C2(n21709), .ZN(P1_U3209) );
  INV_X1 U24671 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21687) );
  OAI222_X1 U24672 ( .A1(n21709), .A2(n21993), .B1(n21687), .B2(n21734), .C1(
        n21686), .C2(n21713), .ZN(P1_U3210) );
  INV_X1 U24673 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n22033) );
  OAI222_X1 U24674 ( .A1(n21709), .A2(n15207), .B1(n22033), .B2(n21734), .C1(
        n21993), .C2(n21713), .ZN(P1_U3211) );
  AOI222_X1 U24675 ( .A1(n21706), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n21746), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n21705), .ZN(n21688) );
  INV_X1 U24676 ( .A(n21688), .ZN(P1_U3212) );
  INV_X1 U24677 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21961) );
  OAI222_X1 U24678 ( .A1(n21709), .A2(n21690), .B1(n21961), .B2(n21734), .C1(
        n21799), .C2(n21713), .ZN(P1_U3213) );
  AOI22_X1 U24679 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21746), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21705), .ZN(n21689) );
  OAI21_X1 U24680 ( .B1(n21690), .B2(n21713), .A(n21689), .ZN(P1_U3214) );
  INV_X1 U24681 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21692) );
  AOI22_X1 U24682 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21746), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21705), .ZN(n21691) );
  OAI21_X1 U24683 ( .B1(n21692), .B2(n21713), .A(n21691), .ZN(P1_U3215) );
  AOI22_X1 U24684 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n21746), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21706), .ZN(n21693) );
  OAI21_X1 U24685 ( .B1(n21694), .B2(n21709), .A(n21693), .ZN(P1_U3216) );
  INV_X1 U24686 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21695) );
  OAI222_X1 U24687 ( .A1(n21709), .A2(n21696), .B1(n21695), .B2(n21734), .C1(
        n21694), .C2(n21713), .ZN(P1_U3217) );
  INV_X1 U24688 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21943) );
  OAI222_X1 U24689 ( .A1(n21713), .A2(n21696), .B1(n21943), .B2(n21734), .C1(
        n21698), .C2(n21709), .ZN(P1_U3218) );
  INV_X1 U24690 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n21697) );
  OAI222_X1 U24691 ( .A1(n21713), .A2(n21698), .B1(n21697), .B2(n21734), .C1(
        n21700), .C2(n21709), .ZN(P1_U3219) );
  INV_X1 U24692 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21699) );
  OAI222_X1 U24693 ( .A1(n21713), .A2(n21700), .B1(n21699), .B2(n21734), .C1(
        n21702), .C2(n21709), .ZN(P1_U3220) );
  AOI22_X1 U24694 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n21705), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21746), .ZN(n21701) );
  OAI21_X1 U24695 ( .B1(n21702), .B2(n21713), .A(n21701), .ZN(P1_U3221) );
  AOI22_X1 U24696 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n21706), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21746), .ZN(n21703) );
  OAI21_X1 U24697 ( .B1(n22020), .B2(n21709), .A(n21703), .ZN(P1_U3222) );
  AOI222_X1 U24698 ( .A1(n21706), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21746), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n21705), .ZN(n21704) );
  INV_X1 U24699 ( .A(n21704), .ZN(P1_U3223) );
  AOI222_X1 U24700 ( .A1(n21706), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21746), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21705), .ZN(n21707) );
  INV_X1 U24701 ( .A(n21707), .ZN(P1_U3224) );
  INV_X1 U24702 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n21998) );
  OAI222_X1 U24703 ( .A1(n21709), .A2(n21712), .B1(n21998), .B2(n21734), .C1(
        n21708), .C2(n21713), .ZN(P1_U3225) );
  INV_X1 U24704 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21711) );
  OAI222_X1 U24705 ( .A1(n21713), .A2(n21712), .B1(n21711), .B2(n21734), .C1(
        n21710), .C2(n21709), .ZN(P1_U3226) );
  INV_X1 U24706 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21714) );
  AOI22_X1 U24707 ( .A1(n21734), .A2(n21715), .B1(n21714), .B2(n21746), .ZN(
        P1_U3458) );
  INV_X1 U24708 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21728) );
  INV_X1 U24709 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21716) );
  AOI22_X1 U24710 ( .A1(n21734), .A2(n21728), .B1(n21716), .B2(n21746), .ZN(
        P1_U3459) );
  INV_X1 U24711 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21717) );
  AOI22_X1 U24712 ( .A1(n21734), .A2(n21718), .B1(n21717), .B2(n21746), .ZN(
        P1_U3460) );
  INV_X1 U24713 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21731) );
  INV_X1 U24714 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21719) );
  AOI22_X1 U24715 ( .A1(n21734), .A2(n21731), .B1(n21719), .B2(n21746), .ZN(
        P1_U3461) );
  INV_X1 U24716 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21722) );
  INV_X1 U24717 ( .A(n21723), .ZN(n21720) );
  AOI21_X1 U24718 ( .B1(n21722), .B2(n21721), .A(n21720), .ZN(P1_U3464) );
  OAI21_X1 U24719 ( .B1(n21724), .B2(n21903), .A(n21723), .ZN(P1_U3465) );
  AOI21_X1 U24720 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21726) );
  AOI22_X1 U24721 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21726), .B2(n21725), .ZN(n21729) );
  AOI22_X1 U24722 ( .A1(n21732), .A2(n21729), .B1(n21728), .B2(n21727), .ZN(
        P1_U3481) );
  OAI21_X1 U24723 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21732), .ZN(n21730) );
  OAI21_X1 U24724 ( .B1(n21732), .B2(n21731), .A(n21730), .ZN(P1_U3482) );
  INV_X1 U24725 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21733) );
  AOI22_X1 U24726 ( .A1(n21734), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21733), 
        .B2(n21746), .ZN(P1_U3483) );
  INV_X1 U24727 ( .A(n21735), .ZN(n21738) );
  INV_X1 U24728 ( .A(n21736), .ZN(n21737) );
  OAI211_X1 U24729 ( .C1(n21739), .C2(n14160), .A(n21738), .B(n21737), .ZN(
        n21745) );
  NAND3_X1 U24730 ( .A1(n21745), .A2(n21742), .A3(n21741), .ZN(n21743) );
  OAI21_X1 U24731 ( .B1(n21745), .B2(n21744), .A(n21743), .ZN(P1_U3485) );
  INV_X1 U24732 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21747) );
  AOI22_X1 U24733 ( .A1(n21734), .A2(n21747), .B1(n21968), .B2(n21746), .ZN(
        P1_U3486) );
  NOR4_X1 U24734 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .A4(n22000), .ZN(n21748) );
  NAND4_X1 U24735 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_3__6__SCAN_IN), .A3(P1_LWORD_REG_12__SCAN_IN), .A4(
        n21748), .ZN(n21756) );
  INV_X1 U24736 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21985) );
  NAND4_X1 U24737 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(n21985), .A4(n21993), .ZN(
        n21755) );
  NAND4_X1 U24738 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(BUF1_REG_16__SCAN_IN), 
        .A3(P1_DATAWIDTH_REG_2__SCAN_IN), .A4(n22005), .ZN(n21754) );
  NOR4_X1 U24739 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n22029), .A3(n22030), 
        .A4(n22038), .ZN(n21752) );
  NOR4_X1 U24740 ( .A1(P1_EAX_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(n22033), .A4(n21989), .ZN(n21751) );
  NOR4_X1 U24741 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_EAX_REG_18__SCAN_IN), .A3(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(
        n22023), .ZN(n21750) );
  NOR4_X1 U24742 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_12__5__SCAN_IN), .A3(P3_INSTQUEUE_REG_3__3__SCAN_IN), 
        .A4(n22035), .ZN(n21749) );
  NAND4_X1 U24743 ( .A1(n21752), .A2(n21751), .A3(n21750), .A4(n21749), .ZN(
        n21753) );
  NOR4_X1 U24744 ( .A1(n21756), .A2(n21755), .A3(n21754), .A4(n21753), .ZN(
        n21793) );
  NAND4_X1 U24745 ( .A1(P1_EAX_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .A3(n21956), .A4(n21757), .ZN(n21758) );
  OR4_X1 U24746 ( .A1(n21759), .A2(n21922), .A3(
        P1_INSTQUEUE_REG_11__4__SCAN_IN), .A4(n21758), .ZN(n21762) );
  NAND4_X1 U24747 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_16__SCAN_IN), .A3(P3_ADDRESS_REG_7__SCAN_IN), .A4(
        P3_UWORD_REG_4__SCAN_IN), .ZN(n21761) );
  NAND4_X1 U24748 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21929), .A3(n21928), 
        .A4(n21942), .ZN(n21760) );
  OR4_X1 U24749 ( .A1(n21762), .A2(n21761), .A3(n21760), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21791) );
  INV_X1 U24750 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21937) );
  NOR4_X1 U24751 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(P2_UWORD_REG_14__SCAN_IN), .A4(
        n21937), .ZN(n21766) );
  NOR4_X1 U24752 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_7__5__SCAN_IN), .A3(P1_REIP_REG_27__SCAN_IN), .A4(
        n22019), .ZN(n21765) );
  NOR4_X1 U24753 ( .A1(P2_EBX_REG_6__SCAN_IN), .A2(P1_EBX_REG_19__SCAN_IN), 
        .A3(n21972), .A4(n16052), .ZN(n21764) );
  NOR4_X1 U24754 ( .A1(BUF1_REG_13__SCAN_IN), .A2(P2_DATAWIDTH_REG_18__SCAN_IN), .A3(P3_READREQUEST_REG_SCAN_IN), .A4(n21968), .ZN(n21763) );
  NAND4_X1 U24755 ( .A1(n21766), .A2(n21765), .A3(n21764), .A4(n21763), .ZN(
        n21790) );
  NAND4_X1 U24756 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_1__3__SCAN_IN), .A3(P1_DATAO_REG_0__SCAN_IN), .A4(
        n21827), .ZN(n21767) );
  NOR3_X1 U24757 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(
        P2_BYTEENABLE_REG_0__SCAN_IN), .A3(n21767), .ZN(n21777) );
  INV_X1 U24758 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n21840) );
  NOR4_X1 U24759 ( .A1(P2_EBX_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n21840), .A4(n21843), .ZN(
        n21768) );
  NAND3_X1 U24760 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(n21768), .ZN(n21775) );
  NOR4_X1 U24761 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(P3_MORE_REG_SCAN_IN), .A4(n21959), .ZN(n21773) );
  NOR4_X1 U24762 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n16041), .A3(
        n11143), .A4(n21797), .ZN(n21772) );
  NOR4_X1 U24763 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(
        P2_LWORD_REG_4__SCAN_IN), .A3(n21812), .A4(n21813), .ZN(n21771) );
  NOR4_X1 U24764 ( .A1(n21809), .A2(n21769), .A3(P3_DATAO_REG_15__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21770) );
  NAND4_X1 U24765 ( .A1(n21773), .A2(n21772), .A3(n21771), .A4(n21770), .ZN(
        n21774) );
  NOR4_X1 U24766 ( .A1(P3_UWORD_REG_6__SCAN_IN), .A2(n11484), .A3(n21775), 
        .A4(n21774), .ZN(n21776) );
  NAND4_X1 U24767 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n21777), .A3(n21776), .A4(n21823), .ZN(n21789) );
  NAND4_X1 U24768 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_1__SCAN_IN), 
        .A4(n21904), .ZN(n21778) );
  NOR3_X1 U24769 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n21909), .A3(n21778), 
        .ZN(n21787) );
  NAND4_X1 U24770 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .A3(n21894), .A4(n21895), .ZN(n21785) );
  NAND4_X1 U24771 ( .A1(P2_EAX_REG_15__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .A3(P3_DATAO_REG_29__SCAN_IN), .A4(
        n21892), .ZN(n21784) );
  NOR4_X1 U24772 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_UWORD_REG_5__SCAN_IN), .A3(P3_DATAO_REG_26__SCAN_IN), .A4(n21861), 
        .ZN(n21782) );
  NOR4_X1 U24773 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21859), .A3(
        n21848), .A4(n21862), .ZN(n21781) );
  INV_X1 U24774 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n21876) );
  NOR4_X1 U24775 ( .A1(BUF2_REG_26__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .A3(P1_DATAO_REG_4__SCAN_IN), .A4(n21876), .ZN(n21780) );
  NOR4_X1 U24776 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21867), .A3(
        n21877), .A4(n15024), .ZN(n21779) );
  NAND4_X1 U24777 ( .A1(n21782), .A2(n21781), .A3(n21780), .A4(n21779), .ZN(
        n21783) );
  NOR3_X1 U24778 ( .A1(n21785), .A2(n21784), .A3(n21783), .ZN(n21786) );
  NAND4_X1 U24779 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(n21787), .A3(n21786), 
        .A4(n16037), .ZN(n21788) );
  NOR4_X1 U24780 ( .A1(n21791), .A2(n21790), .A3(n21789), .A4(n21788), .ZN(
        n21792) );
  AOI21_X1 U24781 ( .B1(n21793), .B2(n21792), .A(P1_ADDRESS_REG_28__SCAN_IN), 
        .ZN(n22052) );
  AOI22_X1 U24782 ( .A1(n16041), .A2(keyinput111), .B1(n11143), .B2(keyinput50), .ZN(n21794) );
  OAI221_X1 U24783 ( .B1(n16041), .B2(keyinput111), .C1(n11143), .C2(
        keyinput50), .A(n21794), .ZN(n21807) );
  INV_X1 U24784 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n21796) );
  AOI22_X1 U24785 ( .A1(n21797), .A2(keyinput9), .B1(n21796), .B2(keyinput43), 
        .ZN(n21795) );
  OAI221_X1 U24786 ( .B1(n21797), .B2(keyinput9), .C1(n21796), .C2(keyinput43), 
        .A(n21795), .ZN(n21806) );
  INV_X1 U24787 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n21800) );
  AOI22_X1 U24788 ( .A1(n21800), .A2(keyinput56), .B1(n21799), .B2(keyinput98), 
        .ZN(n21798) );
  OAI221_X1 U24789 ( .B1(n21800), .B2(keyinput56), .C1(n21799), .C2(keyinput98), .A(n21798), .ZN(n21805) );
  XOR2_X1 U24790 ( .A(n21801), .B(keyinput39), .Z(n21803) );
  XNOR2_X1 U24791 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput31), 
        .ZN(n21802) );
  NAND2_X1 U24792 ( .A1(n21803), .A2(n21802), .ZN(n21804) );
  NOR4_X1 U24793 ( .A1(n21807), .A2(n21806), .A3(n21805), .A4(n21804), .ZN(
        n21856) );
  AOI22_X1 U24794 ( .A1(n21810), .A2(keyinput52), .B1(n21809), .B2(keyinput42), 
        .ZN(n21808) );
  OAI221_X1 U24795 ( .B1(n21810), .B2(keyinput52), .C1(n21809), .C2(keyinput42), .A(n21808), .ZN(n21821) );
  AOI22_X1 U24796 ( .A1(n21813), .A2(keyinput122), .B1(n21812), .B2(
        keyinput112), .ZN(n21811) );
  OAI221_X1 U24797 ( .B1(n21813), .B2(keyinput122), .C1(n21812), .C2(
        keyinput112), .A(n21811), .ZN(n21820) );
  AOI22_X1 U24798 ( .A1(n13815), .A2(keyinput46), .B1(n16176), .B2(keyinput115), .ZN(n21814) );
  OAI221_X1 U24799 ( .B1(n13815), .B2(keyinput46), .C1(n16176), .C2(
        keyinput115), .A(n21814), .ZN(n21819) );
  AOI22_X1 U24800 ( .A1(n21817), .A2(keyinput78), .B1(keyinput38), .B2(n21816), 
        .ZN(n21815) );
  OAI221_X1 U24801 ( .B1(n21817), .B2(keyinput78), .C1(n21816), .C2(keyinput38), .A(n21815), .ZN(n21818) );
  NOR4_X1 U24802 ( .A1(n21821), .A2(n21820), .A3(n21819), .A4(n21818), .ZN(
        n21855) );
  AOI22_X1 U24803 ( .A1(n21824), .A2(keyinput58), .B1(n21823), .B2(keyinput81), 
        .ZN(n21822) );
  OAI221_X1 U24804 ( .B1(n21824), .B2(keyinput58), .C1(n21823), .C2(keyinput81), .A(n21822), .ZN(n21837) );
  AOI22_X1 U24805 ( .A1(n21827), .A2(keyinput72), .B1(n21826), .B2(keyinput87), 
        .ZN(n21825) );
  OAI221_X1 U24806 ( .B1(n21827), .B2(keyinput72), .C1(n21826), .C2(keyinput87), .A(n21825), .ZN(n21836) );
  INV_X1 U24807 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n21829) );
  AOI22_X1 U24808 ( .A1(n21830), .A2(keyinput82), .B1(n21829), .B2(keyinput17), 
        .ZN(n21828) );
  OAI221_X1 U24809 ( .B1(n21830), .B2(keyinput82), .C1(n21829), .C2(keyinput17), .A(n21828), .ZN(n21835) );
  AOI22_X1 U24810 ( .A1(n21833), .A2(keyinput13), .B1(n21832), .B2(keyinput99), 
        .ZN(n21831) );
  OAI221_X1 U24811 ( .B1(n21833), .B2(keyinput13), .C1(n21832), .C2(keyinput99), .A(n21831), .ZN(n21834) );
  NOR4_X1 U24812 ( .A1(n21837), .A2(n21836), .A3(n21835), .A4(n21834), .ZN(
        n21854) );
  AOI22_X1 U24813 ( .A1(n21840), .A2(keyinput121), .B1(keyinput16), .B2(n21839), .ZN(n21838) );
  OAI221_X1 U24814 ( .B1(n21840), .B2(keyinput121), .C1(n21839), .C2(
        keyinput16), .A(n21838), .ZN(n21852) );
  AOI22_X1 U24815 ( .A1(n21843), .A2(keyinput100), .B1(n21842), .B2(
        keyinput123), .ZN(n21841) );
  OAI221_X1 U24816 ( .B1(n21843), .B2(keyinput100), .C1(n21842), .C2(
        keyinput123), .A(n21841), .ZN(n21851) );
  AOI22_X1 U24817 ( .A1(n11484), .A2(keyinput33), .B1(keyinput24), .B2(n21845), 
        .ZN(n21844) );
  OAI221_X1 U24818 ( .B1(n11484), .B2(keyinput33), .C1(n21845), .C2(keyinput24), .A(n21844), .ZN(n21850) );
  INV_X1 U24819 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n21847) );
  AOI22_X1 U24820 ( .A1(n21848), .A2(keyinput36), .B1(n21847), .B2(keyinput65), 
        .ZN(n21846) );
  OAI221_X1 U24821 ( .B1(n21848), .B2(keyinput36), .C1(n21847), .C2(keyinput65), .A(n21846), .ZN(n21849) );
  NOR4_X1 U24822 ( .A1(n21852), .A2(n21851), .A3(n21850), .A4(n21849), .ZN(
        n21853) );
  NAND4_X1 U24823 ( .A1(n21856), .A2(n21855), .A3(n21854), .A4(n21853), .ZN(
        n22050) );
  AOI22_X1 U24824 ( .A1(n21859), .A2(keyinput89), .B1(n21858), .B2(keyinput101), .ZN(n21857) );
  OAI221_X1 U24825 ( .B1(n21859), .B2(keyinput89), .C1(n21858), .C2(
        keyinput101), .A(n21857), .ZN(n21872) );
  AOI22_X1 U24826 ( .A1(n21862), .A2(keyinput29), .B1(n21861), .B2(keyinput108), .ZN(n21860) );
  OAI221_X1 U24827 ( .B1(n21862), .B2(keyinput29), .C1(n21861), .C2(
        keyinput108), .A(n21860), .ZN(n21871) );
  AOI22_X1 U24828 ( .A1(n21865), .A2(keyinput8), .B1(keyinput11), .B2(n21864), 
        .ZN(n21863) );
  OAI221_X1 U24829 ( .B1(n21865), .B2(keyinput8), .C1(n21864), .C2(keyinput11), 
        .A(n21863), .ZN(n21870) );
  INV_X1 U24830 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n21868) );
  AOI22_X1 U24831 ( .A1(n21868), .A2(keyinput73), .B1(n21867), .B2(keyinput41), 
        .ZN(n21866) );
  OAI221_X1 U24832 ( .B1(n21868), .B2(keyinput73), .C1(n21867), .C2(keyinput41), .A(n21866), .ZN(n21869) );
  NOR4_X1 U24833 ( .A1(n21872), .A2(n21871), .A3(n21870), .A4(n21869), .ZN(
        n21920) );
  AOI22_X1 U24834 ( .A1(n21874), .A2(keyinput15), .B1(keyinput126), .B2(n15024), .ZN(n21873) );
  OAI221_X1 U24835 ( .B1(n21874), .B2(keyinput15), .C1(n15024), .C2(
        keyinput126), .A(n21873), .ZN(n21887) );
  AOI22_X1 U24836 ( .A1(n21877), .A2(keyinput68), .B1(n21876), .B2(keyinput44), 
        .ZN(n21875) );
  OAI221_X1 U24837 ( .B1(n21877), .B2(keyinput68), .C1(n21876), .C2(keyinput44), .A(n21875), .ZN(n21886) );
  AOI22_X1 U24838 ( .A1(n21880), .A2(keyinput109), .B1(keyinput61), .B2(n21879), .ZN(n21878) );
  OAI221_X1 U24839 ( .B1(n21880), .B2(keyinput109), .C1(n21879), .C2(
        keyinput61), .A(n21878), .ZN(n21885) );
  AOI22_X1 U24840 ( .A1(n21883), .A2(keyinput66), .B1(n21882), .B2(keyinput77), 
        .ZN(n21881) );
  OAI221_X1 U24841 ( .B1(n21883), .B2(keyinput66), .C1(n21882), .C2(keyinput77), .A(n21881), .ZN(n21884) );
  NOR4_X1 U24842 ( .A1(n21887), .A2(n21886), .A3(n21885), .A4(n21884), .ZN(
        n21919) );
  AOI22_X1 U24843 ( .A1(n21889), .A2(keyinput71), .B1(n13856), .B2(keyinput30), 
        .ZN(n21888) );
  OAI221_X1 U24844 ( .B1(n21889), .B2(keyinput71), .C1(n13856), .C2(keyinput30), .A(n21888), .ZN(n21901) );
  INV_X1 U24845 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n21891) );
  AOI22_X1 U24846 ( .A1(n21892), .A2(keyinput45), .B1(keyinput104), .B2(n21891), .ZN(n21890) );
  OAI221_X1 U24847 ( .B1(n21892), .B2(keyinput45), .C1(n21891), .C2(
        keyinput104), .A(n21890), .ZN(n21900) );
  AOI22_X1 U24848 ( .A1(n21895), .A2(keyinput110), .B1(n21894), .B2(keyinput67), .ZN(n21893) );
  OAI221_X1 U24849 ( .B1(n21895), .B2(keyinput110), .C1(n21894), .C2(
        keyinput67), .A(n21893), .ZN(n21899) );
  AOI22_X1 U24850 ( .A1(n21897), .A2(keyinput18), .B1(n16037), .B2(keyinput117), .ZN(n21896) );
  OAI221_X1 U24851 ( .B1(n21897), .B2(keyinput18), .C1(n16037), .C2(
        keyinput117), .A(n21896), .ZN(n21898) );
  NOR4_X1 U24852 ( .A1(n21901), .A2(n21900), .A3(n21899), .A4(n21898), .ZN(
        n21918) );
  AOI22_X1 U24853 ( .A1(n21904), .A2(keyinput32), .B1(keyinput116), .B2(n21903), .ZN(n21902) );
  OAI221_X1 U24854 ( .B1(n21904), .B2(keyinput32), .C1(n21903), .C2(
        keyinput116), .A(n21902), .ZN(n21916) );
  AOI22_X1 U24855 ( .A1(n21907), .A2(keyinput54), .B1(n21906), .B2(keyinput91), 
        .ZN(n21905) );
  OAI221_X1 U24856 ( .B1(n21907), .B2(keyinput54), .C1(n21906), .C2(keyinput91), .A(n21905), .ZN(n21915) );
  AOI22_X1 U24857 ( .A1(n21910), .A2(keyinput94), .B1(n21909), .B2(keyinput93), 
        .ZN(n21908) );
  OAI221_X1 U24858 ( .B1(n21910), .B2(keyinput94), .C1(n21909), .C2(keyinput93), .A(n21908), .ZN(n21914) );
  XOR2_X1 U24859 ( .A(n16175), .B(keyinput105), .Z(n21912) );
  XNOR2_X1 U24860 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B(keyinput63), .ZN(
        n21911) );
  NAND2_X1 U24861 ( .A1(n21912), .A2(n21911), .ZN(n21913) );
  NOR4_X1 U24862 ( .A1(n21916), .A2(n21915), .A3(n21914), .A4(n21913), .ZN(
        n21917) );
  NAND4_X1 U24863 ( .A1(n21920), .A2(n21919), .A3(n21918), .A4(n21917), .ZN(
        n22049) );
  AOI22_X1 U24864 ( .A1(n21922), .A2(keyinput25), .B1(n21759), .B2(keyinput119), .ZN(n21921) );
  OAI221_X1 U24865 ( .B1(n21922), .B2(keyinput25), .C1(n21759), .C2(
        keyinput119), .A(n21921), .ZN(n21926) );
  XOR2_X1 U24866 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B(keyinput97), .Z(
        n21925) );
  XNOR2_X1 U24867 ( .A(n21923), .B(keyinput102), .ZN(n21924) );
  OR3_X1 U24868 ( .A1(n21926), .A2(n21925), .A3(n21924), .ZN(n21935) );
  AOI22_X1 U24869 ( .A1(n21929), .A2(keyinput88), .B1(keyinput95), .B2(n21928), 
        .ZN(n21927) );
  OAI221_X1 U24870 ( .B1(n21929), .B2(keyinput88), .C1(n21928), .C2(keyinput95), .A(n21927), .ZN(n21934) );
  AOI22_X1 U24871 ( .A1(n21932), .A2(keyinput107), .B1(keyinput92), .B2(n21931), .ZN(n21930) );
  OAI221_X1 U24872 ( .B1(n21932), .B2(keyinput107), .C1(n21931), .C2(
        keyinput92), .A(n21930), .ZN(n21933) );
  NOR3_X1 U24873 ( .A1(n21935), .A2(n21934), .A3(n21933), .ZN(n21982) );
  AOI22_X1 U24874 ( .A1(n13203), .A2(keyinput57), .B1(keyinput1), .B2(n21937), 
        .ZN(n21936) );
  OAI221_X1 U24875 ( .B1(n13203), .B2(keyinput57), .C1(n21937), .C2(keyinput1), 
        .A(n21936), .ZN(n21950) );
  AOI22_X1 U24876 ( .A1(n21940), .A2(keyinput103), .B1(n21939), .B2(keyinput53), .ZN(n21938) );
  OAI221_X1 U24877 ( .B1(n21940), .B2(keyinput103), .C1(n21939), .C2(
        keyinput53), .A(n21938), .ZN(n21949) );
  AOI22_X1 U24878 ( .A1(n21943), .A2(keyinput55), .B1(keyinput49), .B2(n21942), 
        .ZN(n21941) );
  OAI221_X1 U24879 ( .B1(n21943), .B2(keyinput55), .C1(n21942), .C2(keyinput49), .A(n21941), .ZN(n21948) );
  AOI22_X1 U24880 ( .A1(n21946), .A2(keyinput83), .B1(n21945), .B2(keyinput21), 
        .ZN(n21944) );
  OAI221_X1 U24881 ( .B1(n21946), .B2(keyinput83), .C1(n21945), .C2(keyinput21), .A(n21944), .ZN(n21947) );
  NOR4_X1 U24882 ( .A1(n21950), .A2(n21949), .A3(n21948), .A4(n21947), .ZN(
        n21981) );
  AOI22_X1 U24883 ( .A1(n21953), .A2(keyinput127), .B1(keyinput120), .B2(
        n21952), .ZN(n21951) );
  OAI221_X1 U24884 ( .B1(n21953), .B2(keyinput127), .C1(n21952), .C2(
        keyinput120), .A(n21951), .ZN(n21966) );
  AOI22_X1 U24885 ( .A1(n21956), .A2(keyinput85), .B1(n21955), .B2(keyinput34), 
        .ZN(n21954) );
  OAI221_X1 U24886 ( .B1(n21956), .B2(keyinput85), .C1(n21955), .C2(keyinput34), .A(n21954), .ZN(n21965) );
  INV_X1 U24887 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n21958) );
  AOI22_X1 U24888 ( .A1(n21959), .A2(keyinput10), .B1(keyinput37), .B2(n21958), 
        .ZN(n21957) );
  OAI221_X1 U24889 ( .B1(n21959), .B2(keyinput10), .C1(n21958), .C2(keyinput37), .A(n21957), .ZN(n21964) );
  AOI22_X1 U24890 ( .A1(n21962), .A2(keyinput76), .B1(keyinput23), .B2(n21961), 
        .ZN(n21960) );
  OAI221_X1 U24891 ( .B1(n21962), .B2(keyinput76), .C1(n21961), .C2(keyinput23), .A(n21960), .ZN(n21963) );
  NOR4_X1 U24892 ( .A1(n21966), .A2(n21965), .A3(n21964), .A4(n21963), .ZN(
        n21980) );
  AOI22_X1 U24893 ( .A1(n14089), .A2(keyinput27), .B1(keyinput14), .B2(n21968), 
        .ZN(n21967) );
  OAI221_X1 U24894 ( .B1(n14089), .B2(keyinput27), .C1(n21968), .C2(keyinput14), .A(n21967), .ZN(n21978) );
  AOI22_X1 U24895 ( .A1(n21970), .A2(keyinput28), .B1(n16052), .B2(keyinput74), 
        .ZN(n21969) );
  OAI221_X1 U24896 ( .B1(n21970), .B2(keyinput28), .C1(n16052), .C2(keyinput74), .A(n21969), .ZN(n21977) );
  AOI22_X1 U24897 ( .A1(n21972), .A2(keyinput114), .B1(keyinput6), .B2(n12626), 
        .ZN(n21971) );
  OAI221_X1 U24898 ( .B1(n21972), .B2(keyinput114), .C1(n12626), .C2(keyinput6), .A(n21971), .ZN(n21976) );
  XNOR2_X1 U24899 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B(keyinput20), .ZN(
        n21974) );
  XNOR2_X1 U24900 ( .A(DATAI_11_), .B(keyinput0), .ZN(n21973) );
  NAND2_X1 U24901 ( .A1(n21974), .A2(n21973), .ZN(n21975) );
  NOR4_X1 U24902 ( .A1(n21978), .A2(n21977), .A3(n21976), .A4(n21975), .ZN(
        n21979) );
  NAND4_X1 U24903 ( .A1(n21982), .A2(n21981), .A3(n21980), .A4(n21979), .ZN(
        n22048) );
  AOI22_X1 U24904 ( .A1(n21985), .A2(keyinput5), .B1(keyinput47), .B2(n21984), 
        .ZN(n21983) );
  OAI221_X1 U24905 ( .B1(n21985), .B2(keyinput5), .C1(n21984), .C2(keyinput47), 
        .A(n21983), .ZN(n21997) );
  AOI22_X1 U24906 ( .A1(n21987), .A2(keyinput125), .B1(n17273), .B2(keyinput26), .ZN(n21986) );
  OAI221_X1 U24907 ( .B1(n21987), .B2(keyinput125), .C1(n17273), .C2(
        keyinput26), .A(n21986), .ZN(n21996) );
  AOI22_X1 U24908 ( .A1(n21990), .A2(keyinput48), .B1(keyinput75), .B2(n21989), 
        .ZN(n21988) );
  OAI221_X1 U24909 ( .B1(n21990), .B2(keyinput48), .C1(n21989), .C2(keyinput75), .A(n21988), .ZN(n21995) );
  AOI22_X1 U24910 ( .A1(n21993), .A2(keyinput4), .B1(keyinput40), .B2(n21992), 
        .ZN(n21991) );
  OAI221_X1 U24911 ( .B1(n21993), .B2(keyinput4), .C1(n21992), .C2(keyinput40), 
        .A(n21991), .ZN(n21994) );
  NOR4_X1 U24912 ( .A1(n21997), .A2(n21996), .A3(n21995), .A4(n21994), .ZN(
        n22046) );
  AOI22_X1 U24913 ( .A1(keyinput19), .A2(n22000), .B1(keyinput62), .B2(n21998), 
        .ZN(n21999) );
  OAI21_X1 U24914 ( .B1(n22000), .B2(keyinput19), .A(n21999), .ZN(n22011) );
  AOI22_X1 U24915 ( .A1(n12061), .A2(keyinput96), .B1(keyinput2), .B2(n22002), 
        .ZN(n22001) );
  OAI221_X1 U24916 ( .B1(n12061), .B2(keyinput96), .C1(n22002), .C2(keyinput2), 
        .A(n22001), .ZN(n22010) );
  AOI22_X1 U24917 ( .A1(n22005), .A2(keyinput79), .B1(n22004), .B2(keyinput12), 
        .ZN(n22003) );
  OAI221_X1 U24918 ( .B1(n22005), .B2(keyinput79), .C1(n22004), .C2(keyinput12), .A(n22003), .ZN(n22009) );
  INV_X1 U24919 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n22007) );
  AOI22_X1 U24920 ( .A1(n22007), .A2(keyinput69), .B1(keyinput64), .B2(n14112), 
        .ZN(n22006) );
  OAI221_X1 U24921 ( .B1(n22007), .B2(keyinput69), .C1(n14112), .C2(keyinput64), .A(n22006), .ZN(n22008) );
  NOR4_X1 U24922 ( .A1(n22011), .A2(n22010), .A3(n22009), .A4(n22008), .ZN(
        n22045) );
  AOI22_X1 U24923 ( .A1(n22014), .A2(keyinput60), .B1(n22013), .B2(keyinput70), 
        .ZN(n22012) );
  OAI221_X1 U24924 ( .B1(n22014), .B2(keyinput60), .C1(n22013), .C2(keyinput70), .A(n22012), .ZN(n22027) );
  INV_X1 U24925 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n22017) );
  AOI22_X1 U24926 ( .A1(n22017), .A2(keyinput35), .B1(keyinput113), .B2(n22016), .ZN(n22015) );
  OAI221_X1 U24927 ( .B1(n22017), .B2(keyinput35), .C1(n22016), .C2(
        keyinput113), .A(n22015), .ZN(n22026) );
  AOI22_X1 U24928 ( .A1(n22020), .A2(keyinput118), .B1(n22019), .B2(keyinput90), .ZN(n22018) );
  OAI221_X1 U24929 ( .B1(n22020), .B2(keyinput118), .C1(n22019), .C2(
        keyinput90), .A(n22018), .ZN(n22025) );
  INV_X1 U24930 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n22022) );
  AOI22_X1 U24931 ( .A1(n22023), .A2(keyinput22), .B1(n22022), .B2(keyinput124), .ZN(n22021) );
  OAI221_X1 U24932 ( .B1(n22023), .B2(keyinput22), .C1(n22022), .C2(
        keyinput124), .A(n22021), .ZN(n22024) );
  NOR4_X1 U24933 ( .A1(n22027), .A2(n22026), .A3(n22025), .A4(n22024), .ZN(
        n22044) );
  AOI22_X1 U24934 ( .A1(n22030), .A2(keyinput3), .B1(keyinput106), .B2(n22029), 
        .ZN(n22028) );
  OAI221_X1 U24935 ( .B1(n22030), .B2(keyinput3), .C1(n22029), .C2(keyinput106), .A(n22028), .ZN(n22042) );
  AOI22_X1 U24936 ( .A1(n22033), .A2(keyinput80), .B1(n22032), .B2(keyinput86), 
        .ZN(n22031) );
  OAI221_X1 U24937 ( .B1(n22033), .B2(keyinput80), .C1(n22032), .C2(keyinput86), .A(n22031), .ZN(n22041) );
  INV_X1 U24938 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n22036) );
  AOI22_X1 U24939 ( .A1(n22036), .A2(keyinput59), .B1(keyinput84), .B2(n22035), 
        .ZN(n22034) );
  OAI221_X1 U24940 ( .B1(n22036), .B2(keyinput59), .C1(n22035), .C2(keyinput84), .A(n22034), .ZN(n22040) );
  AOI22_X1 U24941 ( .A1(n22038), .A2(keyinput7), .B1(keyinput51), .B2(n14149), 
        .ZN(n22037) );
  OAI221_X1 U24942 ( .B1(n22038), .B2(keyinput7), .C1(n14149), .C2(keyinput51), 
        .A(n22037), .ZN(n22039) );
  NOR4_X1 U24943 ( .A1(n22042), .A2(n22041), .A3(n22040), .A4(n22039), .ZN(
        n22043) );
  NAND4_X1 U24944 ( .A1(n22046), .A2(n22045), .A3(n22044), .A4(n22043), .ZN(
        n22047) );
  NOR4_X1 U24945 ( .A1(n22050), .A2(n22049), .A3(n22048), .A4(n22047), .ZN(
        n22051) );
  OAI21_X1 U24946 ( .B1(keyinput62), .B2(n22052), .A(n22051), .ZN(n22065) );
  AOI22_X1 U24947 ( .A1(n22054), .A2(n22053), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20093), .ZN(n22061) );
  OAI21_X1 U24948 ( .B1(n22057), .B2(n22056), .A(n22055), .ZN(n22059) );
  NAND2_X1 U24949 ( .A1(n22059), .A2(n22058), .ZN(n22060) );
  OAI211_X1 U24950 ( .C1(n22063), .C2(n22062), .A(n22061), .B(n22060), .ZN(
        n22064) );
  XNOR2_X1 U24951 ( .A(n22065), .B(n22064), .ZN(P2_U2916) );
  NAND2_X1 U11199 ( .A1(n18088), .A2(n19961), .ZN(n18072) );
  NAND2_X2 U11277 ( .A1(n11066), .A2(n11417), .ZN(n11968) );
  BUF_X2 U11187 ( .A(n13322), .Z(n13724) );
  CLKBUF_X1 U11198 ( .A(n12132), .Z(n13645) );
  CLKBUF_X1 U11214 ( .A(n11113), .Z(n11114) );
  OR2_X1 U11258 ( .A1(n16289), .A2(n11015), .ZN(n16215) );
  CLKBUF_X1 U11274 ( .A(n12560), .Z(n9780) );
  CLKBUF_X2 U11275 ( .A(n11456), .Z(n11670) );
  INV_X2 U11276 ( .A(n21060), .ZN(n12185) );
  CLKBUF_X1 U11328 ( .A(n14455), .Z(n9763) );
  CLKBUF_X1 U11334 ( .A(n12562), .Z(n14392) );
  NAND2_X1 U11337 ( .A1(n18017), .A2(n10825), .ZN(n10566) );
endmodule

