

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900;

  INV_X1 U2291 ( .A(n2933), .ZN(n3664) );
  INV_X2 U2292 ( .A(n2720), .ZN(n3569) );
  XNOR2_X1 U2294 ( .A(n2766), .B(IR_REG_22__SCAN_IN), .ZN(n4038) );
  INV_X1 U2295 ( .A(n3664), .ZN(n3674) );
  OR2_X1 U2296 ( .A1(n3473), .A2(n3472), .ZN(n3476) );
  OAI22_X1 U2297 ( .A1(n3203), .A2(n3202), .B1(n3201), .B2(n3200), .ZN(n3227)
         );
  INV_X1 U2298 ( .A(n3720), .ZN(n3671) );
  AND2_X1 U2299 ( .A1(n2902), .A2(n2903), .ZN(n2921) );
  NOR2_X1 U2300 ( .A1(n3355), .A2(n3483), .ZN(n3356) );
  AND2_X1 U2301 ( .A1(n2768), .A2(n2942), .ZN(n4811) );
  AOI21_X2 U2302 ( .B1(n4167), .B2(n4807), .A(n4166), .ZN(n4343) );
  NOR2_X2 U2303 ( .A1(n3181), .A2(n3230), .ZN(n3238) );
  NAND4_X2 U2304 ( .A1(n2493), .A2(n2492), .A3(n2491), .A4(n2490), .ZN(n2912)
         );
  AND2_X2 U2305 ( .A1(n4214), .A2(n4011), .ZN(n4195) );
  NAND2_X2 U2306 ( .A1(n2457), .A2(IR_REG_31__SCAN_IN), .ZN(n2458) );
  AOI22_X2 U2307 ( .A1(n3556), .A2(n2703), .B1(n3828), .B2(n4321), .ZN(n4293)
         );
  AOI21_X2 U2308 ( .B1(n4311), .B2(n2694), .A(n2693), .ZN(n3556) );
  OAI21_X1 U2309 ( .B1(n3227), .B2(n3226), .A(n3225), .ZN(n3228) );
  INV_X2 U2310 ( .A(n4037), .ZN(n3719) );
  NAND2_X1 U2311 ( .A1(n2421), .A2(n2745), .ZN(n4153) );
  NAND2_X1 U2312 ( .A1(n2372), .A2(n2371), .ZN(n3865) );
  OR2_X1 U2313 ( .A1(n4295), .A2(n3924), .ZN(n2804) );
  OAI21_X1 U2314 ( .B1(n4231), .B2(n2284), .A(n2404), .ZN(n2403) );
  NAND2_X1 U2315 ( .A1(n3499), .A2(n2257), .ZN(n2389) );
  AND2_X1 U2316 ( .A1(n3473), .A2(n3472), .ZN(n3474) );
  NAND2_X1 U2317 ( .A1(n2369), .A2(n3321), .ZN(n3473) );
  OR2_X1 U2318 ( .A1(n3158), .A2(n3911), .ZN(n2784) );
  OAI21_X1 U2319 ( .B1(n4816), .B2(n2416), .A(n2414), .ZN(n3156) );
  NAND2_X2 U2320 ( .A1(n2957), .A2(n4863), .ZN(n4879) );
  OR2_X1 U2321 ( .A1(n3021), .A2(n3019), .ZN(n2368) );
  INV_X1 U2322 ( .A(n4805), .ZN(n4051) );
  NOR2_X1 U2323 ( .A1(n3147), .A2(n3148), .ZN(n4810) );
  BUF_X1 U2324 ( .A(n2923), .Z(n4056) );
  INV_X2 U2325 ( .A(n2921), .ZN(n4037) );
  NAND4_X2 U2326 ( .A1(n2509), .A2(n2508), .A3(n2507), .A4(n2506), .ZN(n4055)
         );
  NAND4_X1 U2327 ( .A1(n2502), .A2(n2501), .A3(n2500), .A4(n2499), .ZN(n2923)
         );
  NAND2_X2 U2328 ( .A1(n3044), .A2(n4033), .ZN(n3720) );
  OR2_X1 U2329 ( .A1(n3707), .A2(n2820), .ZN(n2456) );
  OR2_X1 U2330 ( .A1(n2821), .A2(n2820), .ZN(n2828) );
  AND2_X1 U2331 ( .A1(n2434), .A2(n2433), .ZN(n2432) );
  AND2_X1 U2332 ( .A1(n2437), .A2(n2293), .ZN(n2377) );
  AND2_X1 U2333 ( .A1(n2271), .A2(n2448), .ZN(n2434) );
  AND4_X1 U2334 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n2447)
         );
  AND2_X1 U2335 ( .A1(n2294), .A2(n2295), .ZN(n2293) );
  AND2_X1 U2336 ( .A1(n2407), .A2(n4617), .ZN(n2378) );
  NOR2_X1 U2337 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2665)
         );
  INV_X1 U2338 ( .A(IR_REG_4__SCAN_IN), .ZN(n2522) );
  NAND4_X2 U2339 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), .ZN(n4054)
         );
  INV_X2 U2340 ( .A(n2536), .ZN(n2720) );
  AND2_X1 U2341 ( .A1(n2465), .A2(n2464), .ZN(n2497) );
  AND2_X2 U2342 ( .A1(n2465), .A2(n2463), .ZN(n2498) );
  OAI22_X2 U2343 ( .A1(n3139), .A2(n2548), .B1(n3148), .B2(n4802), .ZN(n4816)
         );
  XNOR2_X2 U2344 ( .A(n2458), .B(IR_REG_29__SCAN_IN), .ZN(n2463) );
  AOI21_X1 U2345 ( .B1(n3497), .B2(n2399), .A(n2402), .ZN(n2401) );
  INV_X1 U2346 ( .A(n3579), .ZN(n2402) );
  AOI21_X1 U2347 ( .B1(n2279), .B2(n2401), .A(n2262), .ZN(n2395) );
  NAND2_X1 U2348 ( .A1(n3427), .A2(n2969), .ZN(n2364) );
  INV_X1 U2349 ( .A(n3980), .ZN(n2604) );
  NAND2_X1 U2350 ( .A1(n2768), .A2(n4023), .ZN(n3044) );
  OAI21_X1 U2351 ( .B1(n3239), .B2(n2591), .A(n2590), .ZN(n3295) );
  AND2_X1 U2352 ( .A1(n2374), .A2(n2449), .ZN(n2373) );
  INV_X1 U2353 ( .A(IR_REG_9__SCAN_IN), .ZN(n2443) );
  NOR2_X1 U2354 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2446)
         );
  NOR2_X1 U2355 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2445)
         );
  AND2_X1 U2356 ( .A1(n3745), .A2(n3743), .ZN(n3273) );
  OR2_X1 U2357 ( .A1(n3447), .A2(n3449), .ZN(n2323) );
  AOI21_X1 U2358 ( .B1(n2973), .B2(REG1_REG_3__SCAN_IN), .A(n2440), .ZN(n3448)
         );
  AND2_X1 U2359 ( .A1(n2972), .A2(n4431), .ZN(n2440) );
  INV_X1 U2360 ( .A(n4631), .ZN(n2365) );
  INV_X1 U2361 ( .A(n2403), .ZN(n4212) );
  NAND2_X1 U2362 ( .A1(n4222), .A2(n4241), .ZN(n2404) );
  NAND2_X1 U2363 ( .A1(n2998), .A2(n2511), .ZN(n2426) );
  NAND2_X1 U2364 ( .A1(n2809), .A2(n2808), .ZN(n4807) );
  NAND2_X1 U2365 ( .A1(n2764), .A2(n2455), .ZN(n2470) );
  INV_X1 U2366 ( .A(n2510), .ZN(n2406) );
  NOR2_X1 U2367 ( .A1(n2314), .A2(n2313), .ZN(n2312) );
  NOR2_X1 U2368 ( .A1(n4747), .A2(n4814), .ZN(n2313) );
  INV_X1 U2369 ( .A(n4746), .ZN(n2314) );
  NOR2_X1 U2370 ( .A1(n3497), .A2(n2399), .ZN(n2398) );
  INV_X1 U2371 ( .A(IR_REG_1__SCAN_IN), .ZN(n2294) );
  NAND2_X1 U2372 ( .A1(n2349), .A2(REG2_REG_2__SCAN_IN), .ZN(n2348) );
  INV_X1 U2373 ( .A(n4082), .ZN(n2346) );
  NOR2_X1 U2374 ( .A1(n2348), .A2(n2347), .ZN(n2344) );
  NOR2_X1 U2375 ( .A1(n4714), .A2(REG2_REG_12__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U2376 ( .A1(n2264), .A2(REG1_REG_12__SCAN_IN), .ZN(n2309) );
  AND2_X1 U2377 ( .A1(n2677), .A2(n3531), .ZN(n2678) );
  OAI21_X1 U2378 ( .B1(n2604), .B2(n2412), .A(n2618), .ZN(n2411) );
  AND2_X1 U2379 ( .A1(n2569), .A2(n2418), .ZN(n2417) );
  NAND2_X1 U2380 ( .A1(n4815), .A2(n2559), .ZN(n2418) );
  AND2_X1 U2381 ( .A1(n4038), .A2(n4023), .ZN(n2941) );
  INV_X1 U2382 ( .A(n3048), .ZN(n2297) );
  NOR2_X1 U2383 ( .A1(n3702), .A2(n3074), .ZN(n2296) );
  INV_X1 U2384 ( .A(IR_REG_22__SCAN_IN), .ZN(n2819) );
  INV_X1 U2385 ( .A(n2381), .ZN(n2380) );
  AOI21_X1 U2386 ( .B1(n2387), .B2(n2381), .A(n2261), .ZN(n2379) );
  NAND2_X1 U2387 ( .A1(n3718), .A2(n3047), .ZN(n2913) );
  INV_X1 U2388 ( .A(n3598), .ZN(n2392) );
  INV_X1 U2389 ( .A(n2282), .ZN(n2391) );
  AND2_X1 U2390 ( .A1(n3481), .A2(n3480), .ZN(n3497) );
  NAND2_X1 U2391 ( .A1(n2388), .A2(n2385), .ZN(n2384) );
  INV_X1 U2392 ( .A(n3826), .ZN(n2385) );
  NAND2_X1 U2393 ( .A1(n3757), .A2(n2386), .ZN(n2383) );
  XNOR2_X1 U2394 ( .A(n2906), .B(n3671), .ZN(n2916) );
  AND2_X1 U2395 ( .A1(n2737), .A2(n2462), .ZN(n3866) );
  NAND2_X1 U2397 ( .A1(n4081), .A2(n4082), .ZN(n4080) );
  XNOR2_X1 U2398 ( .A(n4087), .B(REG1_REG_2__SCAN_IN), .ZN(n2890) );
  INV_X1 U2399 ( .A(n2293), .ZN(n2488) );
  OAI21_X1 U2400 ( .B1(n3448), .B2(n2320), .A(n2318), .ZN(n3454) );
  INV_X1 U2401 ( .A(n2321), .ZN(n2320) );
  AOI21_X1 U2402 ( .B1(n2321), .B2(n2319), .A(n2283), .ZN(n2318) );
  OAI21_X1 U2403 ( .B1(n4653), .B2(n4795), .A(n2333), .ZN(n3433) );
  OR2_X1 U2404 ( .A1(n4640), .A2(n2332), .ZN(n2331) );
  NAND2_X1 U2405 ( .A1(n2334), .A2(n4795), .ZN(n2332) );
  XNOR2_X1 U2406 ( .A(n3437), .B(n3436), .ZN(n4684) );
  NAND2_X1 U2407 ( .A1(n3460), .A2(n3459), .ZN(n3461) );
  OR2_X1 U2408 ( .A1(n3457), .A2(n4846), .ZN(n3460) );
  AND2_X1 U2409 ( .A1(n2317), .A2(n2281), .ZN(n3457) );
  OR2_X1 U2410 ( .A1(n4705), .A2(n4706), .ZN(n2310) );
  XNOR2_X1 U2411 ( .A(n4094), .B(n4093), .ZN(n3466) );
  INV_X1 U2412 ( .A(n2341), .ZN(n2338) );
  AND2_X1 U2413 ( .A1(n4118), .A2(n4111), .ZN(n2340) );
  OR2_X1 U2414 ( .A1(n4102), .A2(n4101), .ZN(n4119) );
  OR2_X1 U2415 ( .A1(n4118), .A2(n4111), .ZN(n2341) );
  AND2_X1 U2416 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2689)
         );
  NOR2_X1 U2417 ( .A1(n2352), .A2(n2355), .ZN(n2351) );
  INV_X1 U2418 ( .A(n2354), .ZN(n2352) );
  OAI21_X1 U2419 ( .B1(n4195), .B2(n3995), .A(n3992), .ZN(n4174) );
  NAND2_X1 U2420 ( .A1(n4219), .A2(n4207), .ZN(n2423) );
  AND2_X1 U2421 ( .A1(n2734), .A2(n4201), .ZN(n2422) );
  INV_X1 U2422 ( .A(n4192), .ZN(n2424) );
  AND2_X1 U2423 ( .A1(n2479), .A2(n2478), .ZN(n4244) );
  OR2_X1 U2424 ( .A1(n2731), .A2(n4266), .ZN(n2732) );
  OAI22_X1 U2425 ( .A1(n2730), .A2(n4251), .B1(n4259), .B2(n4277), .ZN(n2405)
         );
  AND2_X1 U2426 ( .A1(n2724), .A2(n2723), .ZN(n4267) );
  NAND2_X1 U2427 ( .A1(n2413), .A2(n2604), .ZN(n3297) );
  OAI21_X1 U2428 ( .B1(n3156), .B2(n2581), .A(n2580), .ZN(n3239) );
  NAND2_X1 U2429 ( .A1(n2986), .A2(n2505), .ZN(n2998) );
  NAND2_X1 U2430 ( .A1(n3030), .A2(n3029), .ZN(n3028) );
  AND2_X1 U2431 ( .A1(n2812), .A2(n2955), .ZN(n2942) );
  AND2_X1 U2432 ( .A1(n4183), .A2(n4157), .ZN(n4155) );
  OR2_X1 U2433 ( .A1(n4752), .A2(n4038), .ZN(n4760) );
  NAND2_X1 U2434 ( .A1(n2773), .A2(n2431), .ZN(n2430) );
  INV_X1 U2435 ( .A(IR_REG_27__SCAN_IN), .ZN(n2431) );
  INV_X1 U2436 ( .A(IR_REG_28__SCAN_IN), .ZN(n2773) );
  INV_X1 U2437 ( .A(IR_REG_21__SCAN_IN), .ZN(n2433) );
  INV_X1 U2438 ( .A(IR_REG_20__SCAN_IN), .ZN(n2760) );
  NAND2_X1 U2439 ( .A1(n2269), .A2(IR_REG_31__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U2440 ( .A1(n3320), .A2(n2291), .ZN(n2369) );
  AND2_X1 U2441 ( .A1(n2272), .A2(n4637), .ZN(n2321) );
  INV_X1 U2442 ( .A(n2366), .ZN(n4632) );
  OR2_X1 U2443 ( .A1(n3426), .A2(n2367), .ZN(n2366) );
  XNOR2_X1 U2444 ( .A(n3433), .B(n4837), .ZN(n4668) );
  NAND2_X1 U2445 ( .A1(n4668), .A2(REG2_REG_8__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U2446 ( .A1(n4678), .A2(n4679), .ZN(n4677) );
  XNOR2_X1 U2447 ( .A(n3461), .B(n3436), .ZN(n4686) );
  OAI21_X1 U2448 ( .B1(n4731), .B2(n2325), .A(n2324), .ZN(n4139) );
  NAND2_X1 U2449 ( .A1(n2327), .A2(n2326), .ZN(n2325) );
  INV_X1 U2450 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2326) );
  OAI211_X1 U2451 ( .C1(n4134), .C2(n2353), .A(n2350), .B(n4710), .ZN(n2358)
         );
  NAND2_X1 U2452 ( .A1(n2356), .A2(n2354), .ZN(n2353) );
  NAND2_X1 U2453 ( .A1(n4134), .A2(n2351), .ZN(n2350) );
  NAND2_X1 U2454 ( .A1(n2357), .A2(n4735), .ZN(n2356) );
  AND2_X1 U2455 ( .A1(n4062), .A2(n2980), .ZN(n4744) );
  AOI22_X1 U2456 ( .A1(n4153), .A2(n4160), .B1(n4175), .B2(n4162), .ZN(n2758)
         );
  OR2_X1 U2457 ( .A1(n2759), .A2(IR_REG_19__SCAN_IN), .ZN(n2691) );
  AND2_X1 U2458 ( .A1(n2695), .A2(REG3_REG_21__SCAN_IN), .ZN(n2704) );
  AND2_X1 U2459 ( .A1(n2682), .A2(REG3_REG_20__SCAN_IN), .ZN(n2695) );
  NOR2_X1 U2460 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2444)
         );
  NAND2_X1 U2461 ( .A1(n4080), .A2(n2348), .ZN(n2968) );
  INV_X1 U2462 ( .A(n2323), .ZN(n2319) );
  INV_X1 U2463 ( .A(IR_REG_5__SCAN_IN), .ZN(n2407) );
  NOR2_X1 U2464 ( .A1(n4144), .A2(n4131), .ZN(n2359) );
  NOR2_X1 U2465 ( .A1(n2359), .A2(n4735), .ZN(n2355) );
  OR2_X1 U2466 ( .A1(n4198), .A2(n4185), .ZN(n4158) );
  INV_X1 U2467 ( .A(n4237), .ZN(n3665) );
  NAND2_X1 U2468 ( .A1(n2704), .A2(REG3_REG_22__SCAN_IN), .ZN(n2722) );
  AND2_X1 U2469 ( .A1(REG3_REG_19__SCAN_IN), .A2(n2683), .ZN(n2682) );
  NAND2_X1 U2470 ( .A1(n2299), .A2(n4185), .ZN(n2298) );
  NOR2_X1 U2471 ( .A1(n4162), .A2(n2300), .ZN(n2299) );
  INV_X1 U2472 ( .A(n3938), .ZN(n2300) );
  AND2_X1 U2473 ( .A1(n4328), .A2(n4327), .ZN(n3561) );
  AND2_X1 U2474 ( .A1(n3256), .A2(n3258), .ZN(n3980) );
  INV_X1 U2475 ( .A(IR_REG_6__SCAN_IN), .ZN(n2557) );
  OR3_X1 U2476 ( .A1(n2578), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2588) );
  AND2_X2 U2477 ( .A1(n2519), .A2(n2522), .ZN(n2437) );
  AOI22_X1 U2478 ( .A1(n4054), .A2(n2921), .B1(n3718), .B2(n3074), .ZN(n3014)
         );
  NOR2_X1 U2479 ( .A1(n3646), .A2(n2382), .ZN(n2381) );
  INV_X1 U2480 ( .A(n2384), .ZN(n2382) );
  NOR2_X1 U2481 ( .A1(n2925), .A2(n2924), .ZN(n2926) );
  AND2_X1 U2482 ( .A1(n2933), .A2(n2923), .ZN(n2924) );
  INV_X1 U2483 ( .A(n3516), .ZN(n3854) );
  AOI22_X1 U2484 ( .A1(n4802), .A2(n3674), .B1(n3719), .B2(n3148), .ZN(n3190)
         );
  INV_X1 U2485 ( .A(n4201), .ZN(n4207) );
  NAND2_X1 U2486 ( .A1(n2631), .A2(REG3_REG_14__SCAN_IN), .ZN(n2640) );
  OR2_X1 U2487 ( .A1(n2640), .A2(n2639), .ZN(n2653) );
  NAND2_X1 U2488 ( .A1(n2394), .A2(n2282), .ZN(n2393) );
  INV_X1 U2489 ( .A(n3499), .ZN(n2394) );
  NAND4_X2 U2490 ( .A1(n2487), .A2(n2485), .A3(n2484), .A4(n2486), .ZN(n2909)
         );
  NAND2_X1 U2491 ( .A1(n2495), .A2(REG3_REG_1__SCAN_IN), .ZN(n2487) );
  AOI22_X1 U2492 ( .A1(n2890), .A2(n4083), .B1(n2349), .B2(REG1_REG_2__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U2493 ( .A1(n2343), .A2(n2342), .ZN(n2894) );
  NAND2_X1 U2494 ( .A1(n4080), .A2(n2260), .ZN(n2342) );
  AOI21_X1 U2495 ( .B1(n4081), .B2(n2345), .A(n2344), .ZN(n2343) );
  NOR2_X1 U2496 ( .A1(n2894), .A2(n2895), .ZN(n2967) );
  INV_X1 U2497 ( .A(n2364), .ZN(n2367) );
  OAI21_X1 U2498 ( .B1(n3426), .B2(n2259), .A(n2268), .ZN(n3430) );
  NAND2_X1 U2499 ( .A1(n4677), .A2(n3435), .ZN(n3437) );
  NAND2_X1 U2500 ( .A1(n4684), .A2(REG2_REG_10__SCAN_IN), .ZN(n4683) );
  NAND2_X1 U2501 ( .A1(n3441), .A2(n2363), .ZN(n2362) );
  AOI21_X1 U2502 ( .B1(n3441), .B2(n2361), .A(n2288), .ZN(n2360) );
  NOR2_X1 U2503 ( .A1(n3442), .A2(n4093), .ZN(n4098) );
  NAND2_X1 U2504 ( .A1(n2308), .A2(n2264), .ZN(n2307) );
  NAND2_X1 U2505 ( .A1(n2270), .A2(n4717), .ZN(n2308) );
  INV_X1 U2506 ( .A(n4116), .ZN(n2327) );
  NAND2_X1 U2507 ( .A1(n2667), .A2(n2441), .ZN(n2688) );
  INV_X1 U2508 ( .A(n4133), .ZN(n2357) );
  AOI21_X1 U2509 ( .B1(n4133), .B2(n2355), .A(n2290), .ZN(n2354) );
  NAND2_X1 U2510 ( .A1(n4198), .A2(n2744), .ZN(n2745) );
  NAND2_X1 U2511 ( .A1(n4181), .A2(n2743), .ZN(n2421) );
  INV_X1 U2512 ( .A(n4180), .ZN(n4173) );
  AND2_X1 U2513 ( .A1(n4158), .A2(n3932), .ZN(n4180) );
  NOR2_X1 U2514 ( .A1(n2669), .A2(n3855), .ZN(n2683) );
  AND2_X1 U2515 ( .A1(n3366), .A2(n2678), .ZN(n2681) );
  NOR2_X1 U2516 ( .A1(n2653), .A2(n4529), .ZN(n2670) );
  INV_X1 U2517 ( .A(n2411), .ZN(n2410) );
  AND2_X1 U2518 ( .A1(n2608), .A2(REG3_REG_12__SCAN_IN), .ZN(n2621) );
  OR2_X1 U2519 ( .A1(n2582), .A2(n4582), .ZN(n2593) );
  INV_X1 U2520 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4582) );
  AOI21_X1 U2521 ( .B1(n2417), .B2(n2415), .A(n2278), .ZN(n2414) );
  INV_X1 U2522 ( .A(n2417), .ZN(n2416) );
  INV_X1 U2523 ( .A(n2559), .ZN(n2415) );
  NAND2_X1 U2524 ( .A1(n2420), .A2(n2419), .ZN(n4818) );
  INV_X1 U2525 ( .A(n4815), .ZN(n2419) );
  NAND2_X1 U2526 ( .A1(n2525), .A2(REG3_REG_6__SCAN_IN), .ZN(n2550) );
  AND4_X1 U2527 ( .A1(n2533), .A2(n2532), .A3(n2531), .A4(n2530), .ZN(n3144)
         );
  NOR3_X1 U2528 ( .A1(n4350), .A2(n4339), .A3(n2298), .ZN(n4337) );
  INV_X1 U2529 ( .A(n4282), .ZN(n4800) );
  NOR2_X1 U2530 ( .A1(n4350), .A2(n2744), .ZN(n4183) );
  OR2_X1 U2531 ( .A1(n4225), .A2(n4207), .ZN(n4350) );
  NAND2_X1 U2532 ( .A1(n4243), .A2(n4226), .ZN(n4225) );
  AND2_X1 U2533 ( .A1(n4264), .A2(n4241), .ZN(n4243) );
  NOR2_X1 U2534 ( .A1(n4302), .A2(n2303), .ZN(n4264) );
  OR2_X1 U2535 ( .A1(n4288), .A2(n4259), .ZN(n2303) );
  AND2_X1 U2536 ( .A1(n3561), .A2(n3630), .ZN(n4304) );
  NAND2_X1 U2537 ( .A1(n4304), .A2(n4303), .ZN(n4302) );
  NOR2_X1 U2538 ( .A1(n3513), .A2(n3854), .ZN(n4328) );
  OR2_X1 U2539 ( .A1(n4388), .A2(n3806), .ZN(n3513) );
  NAND2_X1 U2540 ( .A1(n3389), .A2(n2302), .ZN(n4388) );
  AND2_X1 U2541 ( .A1(n3589), .A2(n3388), .ZN(n2302) );
  NAND2_X1 U2542 ( .A1(n3389), .A2(n3388), .ZN(n3387) );
  INV_X1 U2543 ( .A(n4878), .ZN(n3388) );
  AND2_X1 U2544 ( .A1(n3356), .A2(n3501), .ZN(n3389) );
  NAND2_X1 U2545 ( .A1(n3238), .A2(n2285), .ZN(n3355) );
  NAND2_X1 U2546 ( .A1(n3238), .A2(n2263), .ZN(n3293) );
  INV_X1 U2547 ( .A(n3747), .ZN(n3244) );
  AND2_X1 U2548 ( .A1(n3238), .A2(n3244), .ZN(n3294) );
  INV_X1 U2549 ( .A(n3204), .ZN(n3212) );
  OR2_X1 U2550 ( .A1(n4813), .A2(n3212), .ZN(n3181) );
  NAND2_X1 U2551 ( .A1(n2258), .A2(n2275), .ZN(n3147) );
  NAND2_X1 U2552 ( .A1(n2258), .A2(n2297), .ZN(n3067) );
  AND2_X1 U2553 ( .A1(n3009), .A2(n3008), .ZN(n3069) );
  NOR2_X1 U2554 ( .A1(n3048), .A2(n3702), .ZN(n3009) );
  INV_X1 U2555 ( .A(n2838), .ZN(n2847) );
  AND2_X1 U2556 ( .A1(n2903), .A2(n2872), .ZN(n3087) );
  NAND2_X1 U2557 ( .A1(n2470), .A2(IR_REG_31__SCAN_IN), .ZN(n2775) );
  AND2_X1 U2558 ( .A1(n2453), .A2(n2824), .ZN(n2816) );
  AND2_X1 U2559 ( .A1(n2452), .A2(n2819), .ZN(n2824) );
  NOR2_X1 U2560 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2452)
         );
  NOR2_X1 U2561 ( .A1(n2375), .A2(n2277), .ZN(n2374) );
  INV_X1 U2562 ( .A(n2441), .ZN(n2375) );
  AND2_X1 U2563 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2438)
         );
  NAND2_X1 U2564 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2646) );
  NOR2_X1 U2565 ( .A1(n2588), .A2(IR_REG_9__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U2566 ( .A1(n2488), .A2(n2328), .ZN(n4068) );
  INV_X1 U2567 ( .A(n2329), .ZN(n2328) );
  INV_X1 U2568 ( .A(n3863), .ZN(n2370) );
  INV_X1 U2569 ( .A(n3497), .ZN(n2397) );
  NAND2_X1 U2570 ( .A1(n3499), .A2(n3498), .ZN(n2400) );
  AOI21_X1 U2571 ( .B1(n2257), .B2(n2391), .A(n2286), .ZN(n2390) );
  INV_X1 U2572 ( .A(n3047), .ZN(n3698) );
  CLKBUF_X1 U2573 ( .A(n3840), .Z(n4877) );
  NAND2_X1 U2574 ( .A1(n2383), .A2(n2384), .ZN(n3836) );
  NAND2_X1 U2575 ( .A1(n3278), .A2(n3277), .ZN(n3279) );
  INV_X1 U2576 ( .A(n3275), .ZN(n3278) );
  NOR2_X1 U2577 ( .A1(n2960), .A2(n2978), .ZN(n3840) );
  INV_X1 U2578 ( .A(n2922), .ZN(n3702) );
  OR2_X1 U2579 ( .A1(n2945), .A2(n2944), .ZN(n3871) );
  NAND4_X1 U2580 ( .A1(n2469), .A2(n2468), .A3(n2467), .A4(n2466), .ZN(n4219)
         );
  NAND4_X1 U2581 ( .A1(n2483), .A2(n2482), .A3(n2481), .A4(n2480), .ZN(n4260)
         );
  NAND4_X1 U2582 ( .A1(n2729), .A2(n2728), .A3(n2727), .A4(n2726), .ZN(n4277)
         );
  NAND4_X1 U2583 ( .A1(n2711), .A2(n2710), .A3(n2709), .A4(n2708), .ZN(n4278)
         );
  NAND4_X1 U2584 ( .A1(n2701), .A2(n2700), .A3(n2699), .A4(n2698), .ZN(n4321)
         );
  NAND4_X1 U2585 ( .A1(n2599), .A2(n2598), .A3(n2597), .A4(n2596), .ZN(n4048)
         );
  INV_X1 U2586 ( .A(n3144), .ZN(n4053) );
  NAND2_X1 U2587 ( .A1(n2495), .A2(REG3_REG_0__SCAN_IN), .ZN(n2493) );
  AND2_X1 U2588 ( .A1(n2887), .A2(n2886), .ZN(n4062) );
  XNOR2_X1 U2589 ( .A(n4068), .B(REG2_REG_1__SCAN_IN), .ZN(n4075) );
  XNOR2_X1 U2590 ( .A(n4083), .B(n2305), .ZN(n4084) );
  INV_X1 U2591 ( .A(n2890), .ZN(n2305) );
  XNOR2_X1 U2592 ( .A(n3448), .B(n3447), .ZN(n3450) );
  AND2_X1 U2593 ( .A1(n2970), .A2(REG2_REG_4__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U2594 ( .A1(n3448), .A2(n2323), .ZN(n2322) );
  AND2_X1 U2595 ( .A1(n2322), .A2(n2272), .ZN(n4636) );
  XNOR2_X1 U2596 ( .A(n3430), .B(n4787), .ZN(n4641) );
  NAND2_X1 U2597 ( .A1(n3455), .A2(n4645), .ZN(n4658) );
  INV_X1 U2598 ( .A(n2317), .ZN(n4662) );
  AND2_X1 U2599 ( .A1(n2317), .A2(n2265), .ZN(n4674) );
  NAND2_X1 U2600 ( .A1(n4667), .A2(n3434), .ZN(n4678) );
  NAND2_X1 U2601 ( .A1(n4685), .A2(n3462), .ZN(n4695) );
  NAND2_X1 U2602 ( .A1(n4711), .A2(REG2_REG_12__SCAN_IN), .ZN(n4709) );
  AND2_X1 U2603 ( .A1(n2310), .A2(n2270), .ZN(n4719) );
  NAND2_X1 U2604 ( .A1(n4709), .A2(n3441), .ZN(n4716) );
  XNOR2_X1 U2605 ( .A(n4112), .B(n4111), .ZN(n4731) );
  OAI211_X1 U2606 ( .C1(n4119), .C2(n2339), .A(n3373), .B(n2335), .ZN(n4727)
         );
  NAND2_X1 U2607 ( .A1(n2341), .A2(n4111), .ZN(n2339) );
  NOR2_X1 U2608 ( .A1(n2338), .A2(n2340), .ZN(n2337) );
  OAI211_X1 U2609 ( .C1(n4119), .C2(n4111), .A(n2341), .B(n2336), .ZN(n4728)
         );
  NAND2_X1 U2610 ( .A1(n4119), .A2(n2340), .ZN(n2336) );
  NOR2_X1 U2611 ( .A1(n4731), .A2(REG1_REG_16__SCAN_IN), .ZN(n4732) );
  AND2_X1 U2612 ( .A1(n2746), .A2(n2738), .ZN(n4179) );
  NAND2_X1 U2613 ( .A1(n3297), .A2(n2606), .ZN(n3255) );
  NAND2_X1 U2614 ( .A1(n4333), .A2(n3046), .ZN(n4859) );
  INV_X1 U2615 ( .A(n4814), .ZN(n4168) );
  NAND2_X1 U2616 ( .A1(n2426), .A2(n2512), .ZN(n3072) );
  INV_X1 U2617 ( .A(n4863), .ZN(n4847) );
  AND2_X1 U2618 ( .A1(n4333), .A2(n3045), .ZN(n4851) );
  XOR2_X1 U2619 ( .A(n4022), .B(n4337), .Z(n3578) );
  AND2_X1 U2620 ( .A1(n2848), .A2(n2847), .ZN(n2873) );
  NAND2_X1 U2621 ( .A1(n2429), .A2(n2428), .ZN(n2427) );
  INV_X1 U2622 ( .A(IR_REG_29__SCAN_IN), .ZN(n2428) );
  INV_X1 U2623 ( .A(n2430), .ZN(n2429) );
  INV_X1 U2624 ( .A(IR_REG_30__SCAN_IN), .ZN(n3708) );
  NOR2_X1 U2625 ( .A1(n2470), .A2(IR_REG_27__SCAN_IN), .ZN(n2772) );
  XNOR2_X1 U2626 ( .A(n2763), .B(IR_REG_21__SCAN_IN), .ZN(n4023) );
  INV_X1 U2627 ( .A(n4068), .ZN(n4432) );
  NAND2_X1 U2628 ( .A1(n2322), .A2(n2321), .ZN(n4635) );
  AOI21_X1 U2629 ( .B1(n2267), .B2(n4138), .A(n4137), .ZN(n4143) );
  NAND2_X1 U2630 ( .A1(n2315), .A2(n2311), .ZN(U3259) );
  NAND2_X1 U2631 ( .A1(n4745), .A2(n4744), .ZN(n2315) );
  AND2_X1 U2632 ( .A1(n2358), .A2(n2312), .ZN(n2311) );
  AND2_X1 U2633 ( .A1(n2854), .A2(n2853), .ZN(n2855) );
  OR2_X1 U2634 ( .A1(n4147), .A2(n4383), .ZN(n2854) );
  AND2_X1 U2635 ( .A1(n2395), .A2(n2392), .ZN(n2257) );
  XNOR2_X1 U2636 ( .A(n2503), .B(n4617), .ZN(n4087) );
  INV_X1 U2637 ( .A(n4087), .ZN(n2349) );
  AND2_X1 U2638 ( .A1(n3008), .A2(n2296), .ZN(n2258) );
  NAND2_X1 U2639 ( .A1(n2364), .A2(n3428), .ZN(n2259) );
  NAND2_X1 U2640 ( .A1(n2406), .A2(n2437), .ZN(n2534) );
  AND2_X1 U2641 ( .A1(n2348), .A2(n2347), .ZN(n2260) );
  OR2_X1 U2642 ( .A1(n3735), .A2(n3734), .ZN(n2261) );
  AND2_X1 U2643 ( .A1(n2398), .A2(n2396), .ZN(n2262) );
  INV_X1 U2644 ( .A(n3428), .ZN(n3429) );
  AND2_X1 U2645 ( .A1(n3244), .A2(n3302), .ZN(n2263) );
  INV_X1 U2646 ( .A(n4714), .ZN(n2363) );
  OR2_X1 U2647 ( .A1(n4871), .A2(REG1_REG_13__SCAN_IN), .ZN(n2264) );
  INV_X1 U2648 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2316) );
  NAND2_X1 U2649 ( .A1(n2393), .A2(n2395), .ZN(n3792) );
  NOR2_X4 U2650 ( .A1(n2465), .A2(n2463), .ZN(n2496) );
  OR2_X1 U2651 ( .A1(n4837), .A2(n3456), .ZN(n2265) );
  NAND2_X1 U2652 ( .A1(n3757), .A2(n3626), .ZN(n3768) );
  AND2_X1 U2653 ( .A1(n2383), .A2(n2381), .ZN(n2266) );
  MUX2_X1 U2654 ( .A(n2489), .B(n4068), .S(n2536), .Z(n3034) );
  OR2_X1 U2655 ( .A1(n4134), .A2(n4133), .ZN(n2267) );
  XNOR2_X1 U2656 ( .A(n2761), .B(n2760), .ZN(n2768) );
  OR2_X1 U2657 ( .A1(n2365), .A2(n3429), .ZN(n2268) );
  NAND2_X1 U2658 ( .A1(n2667), .A2(n2373), .ZN(n2269) );
  OR2_X1 U2659 ( .A1(n3465), .A2(n4870), .ZN(n2270) );
  AND2_X1 U2660 ( .A1(n2628), .A2(n2432), .ZN(n2764) );
  INV_X1 U2661 ( .A(IR_REG_2__SCAN_IN), .ZN(n4617) );
  AND4_X1 U2662 ( .A1(n2665), .A2(n2451), .A3(n2450), .A4(n2449), .ZN(n2271)
         );
  NAND2_X1 U2663 ( .A1(n3447), .A2(n3449), .ZN(n2272) );
  OR2_X1 U2664 ( .A1(n4350), .A2(n2298), .ZN(n2273) );
  INV_X1 U2665 ( .A(n3108), .ZN(n3118) );
  NAND2_X1 U2666 ( .A1(n2628), .A2(n2434), .ZN(n2762) );
  NOR2_X1 U2667 ( .A1(n4732), .A2(n4113), .ZN(n2274) );
  AND2_X1 U2668 ( .A1(n2297), .A2(n3108), .ZN(n2275) );
  NAND2_X1 U2669 ( .A1(n3757), .A2(n3756), .ZN(n2276) );
  OR2_X1 U2670 ( .A1(n2438), .A2(n2689), .ZN(n2277) );
  AND2_X1 U2671 ( .A1(n4051), .A2(n3212), .ZN(n2278) );
  INV_X1 U2672 ( .A(n2387), .ZN(n2386) );
  NAND2_X1 U2673 ( .A1(n3626), .A2(n2388), .ZN(n2387) );
  NAND2_X1 U2674 ( .A1(n3498), .A2(n2399), .ZN(n2279) );
  AND2_X1 U2675 ( .A1(n4119), .A2(n4118), .ZN(n2280) );
  INV_X1 U2676 ( .A(n3431), .ZN(n2334) );
  AND2_X1 U2677 ( .A1(n2265), .A2(n2316), .ZN(n2281) );
  INV_X1 U2678 ( .A(IR_REG_13__SCAN_IN), .ZN(n2448) );
  INV_X1 U2679 ( .A(n3580), .ZN(n2399) );
  OR2_X1 U2680 ( .A1(n2401), .A2(n2398), .ZN(n2282) );
  AND2_X1 U2681 ( .A1(n2377), .A2(n2378), .ZN(n2546) );
  INV_X1 U2682 ( .A(n3324), .ZN(n2301) );
  AND2_X1 U2683 ( .A1(n3452), .A2(REG1_REG_5__SCAN_IN), .ZN(n2283) );
  INV_X1 U2684 ( .A(n2304), .ZN(n4367) );
  NOR2_X1 U2685 ( .A1(n4302), .A2(n4288), .ZN(n2304) );
  AND2_X1 U2686 ( .A1(n4260), .A2(n4236), .ZN(n2284) );
  AND2_X1 U2687 ( .A1(n2263), .A2(n2301), .ZN(n2285) );
  OR2_X1 U2688 ( .A1(n3597), .A2(n3790), .ZN(n2286) );
  AND2_X1 U2689 ( .A1(n2400), .A2(n2397), .ZN(n2287) );
  INV_X1 U2690 ( .A(n3589), .ZN(n3798) );
  INV_X1 U2691 ( .A(n2606), .ZN(n2412) );
  INV_X1 U2692 ( .A(IR_REG_31__SCAN_IN), .ZN(n2820) );
  AOI21_X1 U2693 ( .B1(n3055), .B2(n2539), .A(n2442), .ZN(n3139) );
  NAND2_X1 U2694 ( .A1(n4818), .A2(n2559), .ZN(n3173) );
  NAND2_X1 U2695 ( .A1(n2915), .A2(n2436), .ZN(n2976) );
  INV_X1 U2696 ( .A(n3498), .ZN(n2396) );
  NOR2_X1 U2697 ( .A1(n3018), .A2(n2368), .ZN(n3105) );
  AND2_X1 U2698 ( .A1(n4722), .A2(n3360), .ZN(n2288) );
  OR2_X1 U2699 ( .A1(n4663), .A2(n4664), .ZN(n2317) );
  CLKBUF_X1 U2700 ( .A(n2909), .Z(n4057) );
  INV_X1 U2701 ( .A(n2909), .ZN(n2425) );
  INV_X1 U2702 ( .A(n4710), .ZN(n4748) );
  AND2_X1 U2703 ( .A1(n4062), .A2(n2893), .ZN(n4710) );
  AND2_X1 U2704 ( .A1(n2366), .A2(n2365), .ZN(n2289) );
  AND2_X1 U2705 ( .A1(n2359), .A2(n4735), .ZN(n2290) );
  NAND2_X1 U2706 ( .A1(n3285), .A2(n3284), .ZN(n2291) );
  AND2_X1 U2707 ( .A1(n3028), .A2(n2494), .ZN(n2292) );
  NOR2_X1 U2708 ( .A1(n2470), .A2(n2427), .ZN(n3707) );
  INV_X1 U2709 ( .A(n4431), .ZN(n2347) );
  INV_X1 U2710 ( .A(IR_REG_3__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U2711 ( .A1(n2293), .A2(n4617), .ZN(n2510) );
  NOR2_X1 U2712 ( .A1(n2488), .A2(IR_REG_13__SCAN_IN), .ZN(n2376) );
  NAND2_X1 U2713 ( .A1(IR_REG_31__SCAN_IN), .A2(n2488), .ZN(n2503) );
  INV_X1 U2714 ( .A(IR_REG_0__SCAN_IN), .ZN(n2295) );
  MUX2_X1 U2715 ( .A(n2472), .B(n2471), .S(n2775), .Z(n2536) );
  OR2_X1 U2716 ( .A1(n4705), .A2(n2309), .ZN(n2306) );
  NAND2_X1 U2717 ( .A1(n2307), .A2(n2306), .ZN(n4094) );
  INV_X1 U2718 ( .A(n2310), .ZN(n4704) );
  XNOR2_X1 U2719 ( .A(n3456), .B(n4837), .ZN(n4663) );
  NAND2_X1 U2720 ( .A1(n4113), .A2(n2327), .ZN(n2324) );
  OAI21_X1 U2721 ( .B1(IR_REG_31__SCAN_IN), .B2(IR_REG_1__SCAN_IN), .A(n2330), 
        .ZN(n2329) );
  NAND3_X1 U2722 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .A3(
        IR_REG_31__SCAN_IN), .ZN(n2330) );
  NAND2_X1 U2723 ( .A1(n2331), .A2(REG2_REG_7__SCAN_IN), .ZN(n2333) );
  NOR2_X1 U2724 ( .A1(n4640), .A2(n3431), .ZN(n4653) );
  NAND2_X1 U2725 ( .A1(n4119), .A2(n2337), .ZN(n2335) );
  NAND2_X1 U2726 ( .A1(n4120), .A2(n4727), .ZN(n4121) );
  NOR2_X1 U2727 ( .A1(n2346), .A2(n2347), .ZN(n2345) );
  OAI21_X1 U2728 ( .B1(n4711), .B2(n2362), .A(n2360), .ZN(n3442) );
  NOR2_X2 U2729 ( .A1(n2936), .A2(n2935), .ZN(n3018) );
  NAND2_X1 U2730 ( .A1(n3668), .A2(n3667), .ZN(n2371) );
  NAND2_X1 U2731 ( .A1(n3666), .A2(n3781), .ZN(n2372) );
  NAND3_X1 U2732 ( .A1(n2372), .A2(n2371), .A3(n2370), .ZN(n3687) );
  NAND2_X1 U2733 ( .A1(n2667), .A2(n2374), .ZN(n2759) );
  NAND4_X1 U2734 ( .A1(n2447), .A2(n2378), .A3(n2437), .A4(n2376), .ZN(n2637)
         );
  AND2_X2 U2735 ( .A1(n2546), .A2(n2447), .ZN(n2628) );
  OAI21_X2 U2736 ( .B1(n3757), .B2(n2380), .A(n2379), .ZN(n3736) );
  INV_X1 U2737 ( .A(n3641), .ZN(n2388) );
  NAND2_X2 U2738 ( .A1(n2389), .A2(n2390), .ZN(n3847) );
  NAND2_X2 U2739 ( .A1(n2405), .A2(n2732), .ZN(n4231) );
  NAND2_X1 U2740 ( .A1(n3028), .A2(n2408), .ZN(n2986) );
  AND2_X1 U2741 ( .A1(n2987), .A2(n2494), .ZN(n2408) );
  OAI21_X1 U2742 ( .B1(n2987), .B2(n2292), .A(n2986), .ZN(n4768) );
  INV_X1 U2743 ( .A(n3295), .ZN(n2413) );
  NAND2_X1 U2744 ( .A1(n2409), .A2(n2410), .ZN(n2620) );
  NAND2_X1 U2745 ( .A1(n3295), .A2(n2606), .ZN(n2409) );
  INV_X1 U2746 ( .A(n4816), .ZN(n2420) );
  AOI21_X2 U2747 ( .B1(n2424), .B2(n2423), .A(n2422), .ZN(n4181) );
  NAND2_X1 U2748 ( .A1(n2425), .A2(n3089), .ZN(n3895) );
  NAND3_X1 U2749 ( .A1(n2426), .A2(n2512), .A3(n3071), .ZN(n3055) );
  OR2_X2 U2750 ( .A1(n2470), .A2(n2430), .ZN(n2457) );
  AOI21_X2 U2751 ( .B1(n3107), .B2(n3106), .A(n3105), .ZN(n3126) );
  INV_X1 U2752 ( .A(n2463), .ZN(n2464) );
  NOR2_X2 U2753 ( .A1(n3701), .A2(n3700), .ZN(n3699) );
  AOI21_X4 U2754 ( .B1(n3476), .B2(n3475), .A(n3474), .ZN(n3499) );
  NOR2_X1 U2755 ( .A1(n2680), .A2(n3529), .ZN(n2435) );
  AND2_X2 U2756 ( .A1(n2852), .A2(n3042), .ZN(n4835) );
  INV_X1 U2757 ( .A(n4831), .ZN(n2856) );
  OR2_X1 U2758 ( .A1(n2903), .A2(n4059), .ZN(n2436) );
  INV_X1 U2759 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2570) );
  OR2_X1 U2760 ( .A1(n4046), .A2(n3483), .ZN(n2439) );
  INV_X1 U2761 ( .A(n4682), .ZN(n3436) );
  NAND2_X1 U2762 ( .A1(n2666), .A2(IR_REG_31__SCAN_IN), .ZN(n2441) );
  INV_X1 U2763 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2549) );
  INV_X1 U2764 ( .A(n3432), .ZN(n4837) );
  AND2_X1 U2765 ( .A1(n3144), .A2(n3108), .ZN(n2442) );
  INV_X1 U2766 ( .A(IR_REG_19__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U2767 ( .A1(n3458), .A2(REG1_REG_9__SCAN_IN), .ZN(n3459) );
  AND2_X1 U2768 ( .A1(n4213), .A2(n3964), .ZN(n4011) );
  INV_X1 U2769 ( .A(IR_REG_26__SCAN_IN), .ZN(n2454) );
  INV_X1 U2770 ( .A(n3276), .ZN(n3277) );
  INV_X1 U2771 ( .A(n3127), .ZN(n3128) );
  AND2_X1 U2772 ( .A1(n2459), .A2(REG3_REG_23__SCAN_IN), .ZN(n2477) );
  INV_X1 U2773 ( .A(n3447), .ZN(n2969) );
  INV_X1 U2774 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2592) );
  INV_X1 U2775 ( .A(n4799), .ZN(n4809) );
  NAND2_X1 U2776 ( .A1(n2909), .A2(n3034), .ZN(n3892) );
  AND2_X1 U2777 ( .A1(n2816), .A2(n2454), .ZN(n2455) );
  AND2_X1 U2778 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2472)
         );
  NOR2_X1 U2779 ( .A1(n3034), .A2(n2907), .ZN(n2908) );
  NAND2_X1 U2780 ( .A1(n2477), .A2(REG3_REG_24__SCAN_IN), .ZN(n2479) );
  INV_X1 U2781 ( .A(n2498), .ZN(n2607) );
  OAI22_X1 U2782 ( .A1(n4695), .A2(n3463), .B1(REG1_REG_11__SCAN_IN), .B2(
        n4693), .ZN(n3465) );
  INV_X1 U2783 ( .A(n4185), .ZN(n2744) );
  NOR2_X1 U2784 ( .A1(n2479), .A2(n2460), .ZN(n2735) );
  INV_X1 U2785 ( .A(n4303), .ZN(n4296) );
  NAND2_X1 U2786 ( .A1(n2670), .A2(REG3_REG_17__SCAN_IN), .ZN(n2669) );
  AND2_X1 U2787 ( .A1(n2621), .A2(REG3_REG_13__SCAN_IN), .ZN(n2631) );
  NOR2_X1 U2788 ( .A1(n2593), .A2(n2592), .ZN(n2608) );
  OR2_X1 U2789 ( .A1(n2571), .A2(n2570), .ZN(n2582) );
  AND3_X1 U2790 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2525) );
  OR2_X1 U2791 ( .A1(n3535), .A2(n3527), .ZN(n3531) );
  INV_X1 U2792 ( .A(n3002), .ZN(n3008) );
  AOI21_X1 U2793 ( .B1(n3736), .B2(n3660), .A(n3661), .ZN(n3814) );
  INV_X1 U2794 ( .A(n2607), .ZN(n2878) );
  NOR2_X1 U2795 ( .A1(n4642), .A2(n4641), .ZN(n4640) );
  AOI21_X1 U2796 ( .B1(n4737), .B2(ADDR_REG_18__SCAN_IN), .A(n4135), .ZN(n4136) );
  OR2_X1 U2797 ( .A1(n2746), .A2(n3726), .ZN(n4146) );
  INV_X1 U2798 ( .A(n4260), .ZN(n4222) );
  OR2_X1 U2799 ( .A1(n4297), .A2(n4281), .ZN(n4256) );
  AND2_X1 U2800 ( .A1(n4003), .A2(n3999), .ZN(n3952) );
  INV_X1 U2801 ( .A(n4801), .ZN(n4324) );
  INV_X1 U2802 ( .A(n3417), .ZN(n3806) );
  INV_X1 U2803 ( .A(n4807), .ZN(n4300) );
  AND2_X1 U2804 ( .A1(n2840), .A2(n4428), .ZN(n2870) );
  OR2_X1 U2805 ( .A1(n3087), .A2(n2876), .ZN(n2886) );
  INV_X1 U2806 ( .A(n4266), .ZN(n4259) );
  INV_X1 U2807 ( .A(n3760), .ZN(n4875) );
  INV_X1 U2808 ( .A(n3871), .ZN(n4886) );
  AND4_X1 U2809 ( .A1(n2565), .A2(n2564), .A3(n2563), .A4(n2562), .ZN(n4805)
         );
  NAND2_X1 U2810 ( .A1(n3444), .A2(n3443), .ZN(n3445) );
  AOI21_X1 U2811 ( .B1(n4134), .B2(n4133), .A(n4748), .ZN(n4138) );
  AND2_X1 U2812 ( .A1(n4146), .A2(n2747), .ZN(n4154) );
  INV_X1 U2813 ( .A(n3952), .ZN(n3366) );
  NOR2_X1 U2814 ( .A1(n2550), .A2(n2549), .ZN(n2560) );
  INV_X1 U2815 ( .A(n4859), .ZN(n4896) );
  NAND2_X1 U2816 ( .A1(n2856), .A2(REG1_REG_29__SCAN_IN), .ZN(n2853) );
  AOI21_X1 U2817 ( .B1(n2870), .B2(n2874), .A(n2873), .ZN(n2939) );
  AND3_X1 U2818 ( .A1(n2846), .A2(n2938), .A3(n2845), .ZN(n2852) );
  XNOR2_X1 U2819 ( .A(n2823), .B(IR_REG_24__SCAN_IN), .ZN(n2838) );
  AND2_X1 U2820 ( .A1(n2658), .A2(n2648), .ZN(n4107) );
  AND2_X1 U2821 ( .A1(n2877), .A2(n2886), .ZN(n4737) );
  NAND4_X1 U2822 ( .A1(n2742), .A2(n2741), .A3(n2740), .A4(n2739), .ZN(n4198)
         );
  NAND4_X1 U2823 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .ZN(n4237)
         );
  NAND4_X1 U2824 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n4046)
         );
  NAND4_X1 U2825 ( .A1(n2587), .A2(n2586), .A3(n2585), .A4(n2584), .ZN(n4049)
         );
  AND2_X1 U2826 ( .A1(n3306), .A2(n3305), .ZN(n4868) );
  OR2_X1 U2827 ( .A1(n2956), .A2(n4760), .ZN(n4863) );
  NAND2_X1 U2828 ( .A1(n4333), .A2(n4819), .ZN(n4335) );
  AND2_X2 U2829 ( .A1(n3043), .A2(n4863), .ZN(n4900) );
  NAND2_X1 U2830 ( .A1(n4831), .A2(n4811), .ZN(n4383) );
  AND2_X2 U2831 ( .A1(n2852), .A2(n2939), .ZN(n4831) );
  AND2_X1 U2832 ( .A1(n2850), .A2(n2849), .ZN(n2851) );
  NAND2_X1 U2833 ( .A1(n4835), .A2(n4811), .ZN(n4423) );
  INV_X1 U2834 ( .A(n4835), .ZN(n4832) );
  AND2_X1 U2835 ( .A1(n4034), .A2(STATE_REG_SCAN_IN), .ZN(n2872) );
  XNOR2_X1 U2836 ( .A(n2818), .B(IR_REG_26__SCAN_IN), .ZN(n4428) );
  INV_X1 U2837 ( .A(n4111), .ZN(n4893) );
  INV_X1 U2838 ( .A(n4693), .ZN(n4856) );
  INV_X1 U2839 ( .A(n4650), .ZN(n4795) );
  NOR2_X1 U2840 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2451)
         );
  NOR2_X1 U2841 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2450)
         );
  INV_X1 U2842 ( .A(IR_REG_25__SCAN_IN), .ZN(n2453) );
  XNOR2_X2 U2843 ( .A(n2456), .B(n3708), .ZN(n2465) );
  NAND2_X1 U2844 ( .A1(n2513), .A2(REG2_REG_26__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U2845 ( .A1(n2878), .A2(REG1_REG_26__SCAN_IN), .ZN(n2468) );
  INV_X1 U2846 ( .A(n2465), .ZN(n4427) );
  AND2_X2 U2847 ( .A1(n4427), .A2(n2463), .ZN(n2495) );
  NAND2_X1 U2848 ( .A1(n2560), .A2(REG3_REG_8__SCAN_IN), .ZN(n2571) );
  INV_X1 U2849 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2639) );
  INV_X1 U2850 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4529) );
  INV_X1 U2851 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3855) );
  INV_X1 U2852 ( .A(n2722), .ZN(n2459) );
  NAND2_X1 U2853 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2460) );
  INV_X1 U2854 ( .A(n2735), .ZN(n2737) );
  INV_X1 U2855 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4598) );
  INV_X1 U2856 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2461) );
  OAI21_X1 U2857 ( .B1(n2479), .B2(n4598), .A(n2461), .ZN(n2462) );
  NAND2_X1 U2858 ( .A1(n2753), .A2(n3866), .ZN(n2467) );
  BUF_X4 U2859 ( .A(n2497), .Z(n2725) );
  NAND2_X1 U2860 ( .A1(n2725), .A2(REG0_REG_26__SCAN_IN), .ZN(n2466) );
  INV_X1 U2861 ( .A(n4219), .ZN(n2734) );
  NOR2_X1 U2862 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2471)
         );
  NAND2_X1 U2863 ( .A1(n2720), .A2(DATAI_26_), .ZN(n4201) );
  NAND2_X1 U2864 ( .A1(n2513), .A2(REG2_REG_25__SCAN_IN), .ZN(n2476) );
  NAND2_X1 U2865 ( .A1(n2878), .A2(REG1_REG_25__SCAN_IN), .ZN(n2475) );
  XNOR2_X1 U2866 ( .A(n2479), .B(REG3_REG_25__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U2867 ( .A1(n2753), .A2(n3784), .ZN(n2474) );
  NAND2_X1 U2868 ( .A1(n2725), .A2(REG0_REG_25__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U2869 ( .A1(n2720), .A2(DATAI_25_), .ZN(n4226) );
  INV_X1 U2870 ( .A(n4226), .ZN(n4218) );
  NAND2_X1 U2871 ( .A1(n2513), .A2(REG2_REG_24__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U2872 ( .A1(n2878), .A2(REG1_REG_24__SCAN_IN), .ZN(n2482) );
  INV_X1 U2873 ( .A(n2477), .ZN(n2724) );
  INV_X1 U2874 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U2875 ( .A1(n2724), .A2(n4436), .ZN(n2478) );
  NAND2_X1 U2876 ( .A1(n2753), .A2(n4244), .ZN(n2481) );
  NAND2_X1 U2877 ( .A1(n2725), .A2(REG0_REG_24__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U2878 ( .A1(n2720), .A2(DATAI_24_), .ZN(n4241) );
  INV_X1 U2879 ( .A(n4241), .ZN(n4236) );
  NAND2_X1 U2880 ( .A1(n2496), .A2(REG2_REG_1__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U2881 ( .A1(n2497), .A2(REG0_REG_1__SCAN_IN), .ZN(n2485) );
  NAND2_X1 U2882 ( .A1(n2498), .A2(REG1_REG_1__SCAN_IN), .ZN(n2484) );
  INV_X1 U2883 ( .A(DATAI_1_), .ZN(n2489) );
  NAND2_X1 U2884 ( .A1(n3895), .A2(n3892), .ZN(n3030) );
  NAND2_X1 U2885 ( .A1(n2496), .A2(REG2_REG_0__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U2886 ( .A1(n2497), .A2(REG0_REG_0__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U2887 ( .A1(n2498), .A2(REG1_REG_0__SCAN_IN), .ZN(n2490) );
  MUX2_X1 U2888 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(n2536), .Z(n3047) );
  AND2_X1 U2889 ( .A1(n2912), .A2(n3047), .ZN(n3029) );
  INV_X1 U2890 ( .A(n3034), .ZN(n3089) );
  NAND2_X1 U2891 ( .A1(n4057), .A2(n3089), .ZN(n2494) );
  NAND2_X1 U2892 ( .A1(n2495), .A2(REG3_REG_2__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U2893 ( .A1(n2496), .A2(REG2_REG_2__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U2894 ( .A1(n2497), .A2(REG0_REG_2__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U2895 ( .A1(n2498), .A2(REG1_REG_2__SCAN_IN), .ZN(n2499) );
  INV_X1 U2896 ( .A(DATAI_2_), .ZN(n2504) );
  MUX2_X1 U2897 ( .A(n2504), .B(n4087), .S(n2536), .Z(n2922) );
  OR2_X1 U2898 ( .A1(n2923), .A2(n2922), .ZN(n3896) );
  NAND2_X1 U2899 ( .A1(n4056), .A2(n2922), .ZN(n3899) );
  NAND2_X1 U2900 ( .A1(n3896), .A2(n3899), .ZN(n2987) );
  INV_X1 U2901 ( .A(n4056), .ZN(n3005) );
  NAND2_X1 U2902 ( .A1(n3005), .A2(n2922), .ZN(n2505) );
  NAND2_X1 U2903 ( .A1(n2498), .A2(REG1_REG_3__SCAN_IN), .ZN(n2509) );
  NAND2_X1 U2904 ( .A1(n2495), .A2(n4772), .ZN(n2508) );
  NAND2_X1 U2905 ( .A1(n2725), .A2(REG0_REG_3__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U2906 ( .A1(n2513), .A2(REG2_REG_3__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U2907 ( .A1(n2510), .A2(IR_REG_31__SCAN_IN), .ZN(n2520) );
  XNOR2_X1 U2908 ( .A(n2520), .B(IR_REG_3__SCAN_IN), .ZN(n4431) );
  MUX2_X1 U2909 ( .A(DATAI_3_), .B(n4431), .S(n2536), .Z(n3002) );
  NAND2_X1 U2910 ( .A1(n4055), .A2(n3002), .ZN(n2511) );
  INV_X1 U2911 ( .A(n4055), .ZN(n2934) );
  NAND2_X1 U2912 ( .A1(n2934), .A2(n3008), .ZN(n2512) );
  NAND2_X1 U2913 ( .A1(n2513), .A2(REG2_REG_4__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U2914 ( .A1(n2498), .A2(REG1_REG_4__SCAN_IN), .ZN(n2517) );
  INV_X1 U2915 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2514) );
  XNOR2_X1 U2916 ( .A(n2514), .B(REG3_REG_3__SCAN_IN), .ZN(n3080) );
  NAND2_X1 U2917 ( .A1(n2495), .A2(n3080), .ZN(n2516) );
  NAND2_X1 U2918 ( .A1(n2725), .A2(REG0_REG_4__SCAN_IN), .ZN(n2515) );
  INV_X1 U2919 ( .A(DATAI_4_), .ZN(n2524) );
  NAND2_X1 U2920 ( .A1(n2520), .A2(n2519), .ZN(n2521) );
  NAND2_X1 U2921 ( .A1(n2521), .A2(IR_REG_31__SCAN_IN), .ZN(n2523) );
  XNOR2_X1 U2922 ( .A(n2523), .B(n2522), .ZN(n3447) );
  MUX2_X1 U2923 ( .A(n2524), .B(n3447), .S(n2536), .Z(n3068) );
  OR2_X1 U2924 ( .A1(n4054), .A2(n3068), .ZN(n3902) );
  NAND2_X1 U2925 ( .A1(n4054), .A2(n3068), .ZN(n3906) );
  NAND2_X1 U2926 ( .A1(n3902), .A2(n3906), .ZN(n3071) );
  INV_X1 U2927 ( .A(n3068), .ZN(n3074) );
  NAND2_X1 U2928 ( .A1(n4054), .A2(n3074), .ZN(n3056) );
  INV_X1 U2929 ( .A(n2525), .ZN(n2540) );
  INV_X1 U2930 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2527) );
  NAND2_X1 U2931 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2526) );
  NAND2_X1 U2932 ( .A1(n2527), .A2(n2526), .ZN(n2528) );
  NAND2_X1 U2933 ( .A1(n2540), .A2(n2528), .ZN(n3121) );
  INV_X1 U2934 ( .A(n3121), .ZN(n2529) );
  NAND2_X1 U2935 ( .A1(n2495), .A2(n2529), .ZN(n2533) );
  NAND2_X1 U2936 ( .A1(n2513), .A2(REG2_REG_5__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U2937 ( .A1(n2725), .A2(REG0_REG_5__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U2938 ( .A1(n2498), .A2(REG1_REG_5__SCAN_IN), .ZN(n2530) );
  INV_X1 U2939 ( .A(DATAI_5_), .ZN(n2537) );
  NAND2_X1 U2940 ( .A1(n2534), .A2(IR_REG_31__SCAN_IN), .ZN(n2535) );
  XNOR2_X1 U2941 ( .A(n2535), .B(IR_REG_5__SCAN_IN), .ZN(n3452) );
  INV_X1 U2942 ( .A(n3452), .ZN(n4785) );
  MUX2_X1 U2943 ( .A(n2537), .B(n4785), .S(n3569), .Z(n3108) );
  NAND2_X1 U2944 ( .A1(n4053), .A2(n3118), .ZN(n2538) );
  AND2_X1 U2945 ( .A1(n3056), .A2(n2538), .ZN(n2539) );
  NAND2_X1 U2946 ( .A1(n2498), .A2(REG1_REG_6__SCAN_IN), .ZN(n2545) );
  INV_X1 U2947 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U2948 ( .A1(n2540), .A2(n3132), .ZN(n2541) );
  AND2_X1 U2949 ( .A1(n2541), .A2(n2550), .ZN(n4788) );
  NAND2_X1 U2950 ( .A1(n2495), .A2(n4788), .ZN(n2544) );
  NAND2_X1 U2951 ( .A1(n2725), .A2(REG0_REG_6__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U2952 ( .A1(n2513), .A2(REG2_REG_6__SCAN_IN), .ZN(n2542) );
  NAND4_X1 U2953 ( .A1(n2545), .A2(n2544), .A3(n2543), .A4(n2542), .ZN(n4802)
         );
  OR2_X1 U2954 ( .A1(n2546), .A2(n2820), .ZN(n2547) );
  XNOR2_X1 U2955 ( .A(n2547), .B(IR_REG_6__SCAN_IN), .ZN(n3453) );
  MUX2_X1 U2956 ( .A(DATAI_6_), .B(n3453), .S(n3569), .Z(n3148) );
  AND2_X1 U2957 ( .A1(n4802), .A2(n3148), .ZN(n2548) );
  NAND2_X1 U2958 ( .A1(n2498), .A2(REG1_REG_7__SCAN_IN), .ZN(n2556) );
  AND2_X1 U2959 ( .A1(n2550), .A2(n2549), .ZN(n2551) );
  OR2_X1 U2960 ( .A1(n2551), .A2(n2560), .ZN(n4824) );
  INV_X1 U2961 ( .A(n4824), .ZN(n2552) );
  NAND2_X1 U2962 ( .A1(n2495), .A2(n2552), .ZN(n2555) );
  NAND2_X1 U2963 ( .A1(n2725), .A2(REG0_REG_7__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U2964 ( .A1(n2513), .A2(REG2_REG_7__SCAN_IN), .ZN(n2553) );
  NAND4_X1 U2965 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n4052)
         );
  NAND2_X1 U2966 ( .A1(n2546), .A2(n2557), .ZN(n2578) );
  NAND2_X1 U2967 ( .A1(n2578), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  XNOR2_X1 U2968 ( .A(n2566), .B(IR_REG_7__SCAN_IN), .ZN(n4650) );
  MUX2_X1 U2969 ( .A(DATAI_7_), .B(n4650), .S(n3569), .Z(n4799) );
  OR2_X1 U2970 ( .A1(n4052), .A2(n4799), .ZN(n2558) );
  NAND2_X1 U2971 ( .A1(n4052), .A2(n4799), .ZN(n2559) );
  NAND2_X1 U2972 ( .A1(n2558), .A2(n2559), .ZN(n4815) );
  OR2_X1 U2973 ( .A1(n2560), .A2(REG3_REG_8__SCAN_IN), .ZN(n2561) );
  AND2_X1 U2974 ( .A1(n2571), .A2(n2561), .ZN(n4838) );
  NAND2_X1 U2975 ( .A1(n2495), .A2(n4838), .ZN(n2565) );
  NAND2_X1 U2976 ( .A1(n2513), .A2(REG2_REG_8__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U2977 ( .A1(n2725), .A2(REG0_REG_8__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U2978 ( .A1(n2878), .A2(REG1_REG_8__SCAN_IN), .ZN(n2562) );
  INV_X1 U2979 ( .A(DATAI_8_), .ZN(n4836) );
  INV_X1 U2980 ( .A(IR_REG_7__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U2981 ( .A1(n2566), .A2(n4521), .ZN(n2567) );
  NAND2_X1 U2982 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2568) );
  XNOR2_X1 U2983 ( .A(n2568), .B(IR_REG_8__SCAN_IN), .ZN(n3432) );
  MUX2_X1 U2984 ( .A(n4836), .B(n4837), .S(n3569), .Z(n3204) );
  NAND2_X1 U2985 ( .A1(n4805), .A2(n3204), .ZN(n2569) );
  NAND2_X1 U2986 ( .A1(n2878), .A2(REG1_REG_9__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U2987 ( .A1(n2571), .A2(n2570), .ZN(n2572) );
  NAND2_X1 U2988 ( .A1(n2582), .A2(n2572), .ZN(n3233) );
  INV_X1 U2989 ( .A(n3233), .ZN(n2573) );
  NAND2_X1 U2990 ( .A1(n2495), .A2(n2573), .ZN(n2576) );
  NAND2_X1 U2991 ( .A1(n2725), .A2(REG0_REG_9__SCAN_IN), .ZN(n2575) );
  NAND2_X1 U2992 ( .A1(n2513), .A2(REG2_REG_9__SCAN_IN), .ZN(n2574) );
  NAND4_X1 U2993 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n4050)
         );
  NAND2_X1 U2994 ( .A1(n2588), .A2(IR_REG_31__SCAN_IN), .ZN(n2579) );
  XNOR2_X1 U2995 ( .A(n2579), .B(IR_REG_9__SCAN_IN), .ZN(n4671) );
  MUX2_X1 U2996 ( .A(DATAI_9_), .B(n4671), .S(n3569), .Z(n3230) );
  AND2_X1 U2997 ( .A1(n4050), .A2(n3230), .ZN(n2581) );
  INV_X1 U2998 ( .A(n4050), .ZN(n3221) );
  INV_X1 U2999 ( .A(n3230), .ZN(n3220) );
  NAND2_X1 U3000 ( .A1(n3221), .A2(n3220), .ZN(n2580) );
  NAND2_X1 U3001 ( .A1(n2582), .A2(n4582), .ZN(n2583) );
  AND2_X1 U3002 ( .A1(n2593), .A2(n2583), .ZN(n4848) );
  NAND2_X1 U3003 ( .A1(n2753), .A2(n4848), .ZN(n2587) );
  NAND2_X1 U3004 ( .A1(n2513), .A2(REG2_REG_10__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U3005 ( .A1(n2725), .A2(REG0_REG_10__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U3006 ( .A1(n2878), .A2(REG1_REG_10__SCAN_IN), .ZN(n2584) );
  OR2_X1 U3007 ( .A1(n2601), .A2(n2820), .ZN(n2589) );
  XNOR2_X1 U3008 ( .A(n2589), .B(IR_REG_10__SCAN_IN), .ZN(n4682) );
  MUX2_X1 U3009 ( .A(DATAI_10_), .B(n4682), .S(n3569), .Z(n3747) );
  NOR2_X1 U3010 ( .A1(n4049), .A2(n3747), .ZN(n2591) );
  NAND2_X1 U3011 ( .A1(n4049), .A2(n3747), .ZN(n2590) );
  AND2_X1 U3012 ( .A1(n2593), .A2(n2592), .ZN(n2594) );
  OR2_X1 U3013 ( .A1(n2594), .A2(n2608), .ZN(n4864) );
  INV_X1 U3014 ( .A(n4864), .ZN(n2595) );
  NAND2_X1 U3015 ( .A1(n2495), .A2(n2595), .ZN(n2599) );
  NAND2_X1 U3016 ( .A1(n2513), .A2(REG2_REG_11__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U3017 ( .A1(n2725), .A2(REG0_REG_11__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U3018 ( .A1(n2878), .A2(REG1_REG_11__SCAN_IN), .ZN(n2596) );
  INV_X1 U3019 ( .A(DATAI_11_), .ZN(n2603) );
  INV_X1 U3020 ( .A(IR_REG_10__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U3021 ( .A1(n2601), .A2(n2600), .ZN(n2602) );
  NAND2_X1 U3022 ( .A1(n2602), .A2(IR_REG_31__SCAN_IN), .ZN(n2615) );
  XNOR2_X1 U3023 ( .A(n2615), .B(IR_REG_11__SCAN_IN), .ZN(n4693) );
  MUX2_X1 U3024 ( .A(n2603), .B(n4856), .S(n3569), .Z(n3302) );
  OR2_X1 U3025 ( .A1(n4048), .A2(n3302), .ZN(n3256) );
  NAND2_X1 U3026 ( .A1(n4048), .A2(n3302), .ZN(n3258) );
  INV_X1 U3027 ( .A(n4048), .ZN(n2605) );
  NAND2_X1 U3028 ( .A1(n2605), .A2(n3302), .ZN(n2606) );
  NAND2_X1 U3029 ( .A1(n2496), .A2(REG2_REG_12__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U3030 ( .A1(n2878), .A2(REG1_REG_12__SCAN_IN), .ZN(n2612) );
  NOR2_X1 U3031 ( .A1(n2608), .A2(REG3_REG_12__SCAN_IN), .ZN(n2609) );
  OR2_X1 U3032 ( .A1(n2621), .A2(n2609), .ZN(n3327) );
  INV_X1 U3033 ( .A(n3327), .ZN(n3263) );
  NAND2_X1 U3034 ( .A1(n2753), .A2(n3263), .ZN(n2611) );
  NAND2_X1 U3035 ( .A1(n2725), .A2(REG0_REG_12__SCAN_IN), .ZN(n2610) );
  NAND4_X1 U3036 ( .A1(n2613), .A2(n2612), .A3(n2611), .A4(n2610), .ZN(n4047)
         );
  INV_X1 U3037 ( .A(IR_REG_11__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U3038 ( .A1(n2615), .A2(n2614), .ZN(n2616) );
  NAND2_X1 U3039 ( .A1(n2616), .A2(IR_REG_31__SCAN_IN), .ZN(n2617) );
  XNOR2_X1 U3040 ( .A(n2617), .B(IR_REG_12__SCAN_IN), .ZN(n3464) );
  MUX2_X1 U3041 ( .A(DATAI_12_), .B(n3464), .S(n3569), .Z(n3324) );
  NAND2_X1 U3042 ( .A1(n4047), .A2(n3324), .ZN(n2618) );
  INV_X1 U3043 ( .A(n4047), .ZN(n3351) );
  NAND2_X1 U3044 ( .A1(n3351), .A2(n2301), .ZN(n2619) );
  NAND2_X1 U3045 ( .A1(n2620), .A2(n2619), .ZN(n3344) );
  INV_X1 U3046 ( .A(n3344), .ZN(n2630) );
  NAND2_X1 U3047 ( .A1(n2496), .A2(REG2_REG_13__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U3048 ( .A1(n2878), .A2(REG1_REG_13__SCAN_IN), .ZN(n2626) );
  NOR2_X1 U3049 ( .A1(n2621), .A2(REG3_REG_13__SCAN_IN), .ZN(n2622) );
  OR2_X1 U3050 ( .A1(n2631), .A2(n2622), .ZN(n3486) );
  INV_X1 U3051 ( .A(n3486), .ZN(n2623) );
  NAND2_X1 U3052 ( .A1(n2753), .A2(n2623), .ZN(n2625) );
  NAND2_X1 U3053 ( .A1(n2725), .A2(REG0_REG_13__SCAN_IN), .ZN(n2624) );
  OR2_X1 U3054 ( .A1(n2628), .A2(n2820), .ZN(n2629) );
  XNOR2_X1 U3055 ( .A(n2629), .B(IR_REG_13__SCAN_IN), .ZN(n4871) );
  MUX2_X1 U3056 ( .A(DATAI_13_), .B(n4871), .S(n3569), .Z(n3483) );
  NAND2_X1 U3057 ( .A1(n2630), .A2(n2439), .ZN(n3332) );
  NAND2_X1 U3058 ( .A1(n2878), .A2(REG1_REG_14__SCAN_IN), .ZN(n2636) );
  NAND2_X1 U3059 ( .A1(n2513), .A2(REG2_REG_14__SCAN_IN), .ZN(n2635) );
  OR2_X1 U3060 ( .A1(n2631), .A2(REG3_REG_14__SCAN_IN), .ZN(n2632) );
  AND2_X1 U3061 ( .A1(n2632), .A2(n2640), .ZN(n3504) );
  NAND2_X1 U3062 ( .A1(n2753), .A2(n3504), .ZN(n2634) );
  NAND2_X1 U3063 ( .A1(n2725), .A2(REG0_REG_14__SCAN_IN), .ZN(n2633) );
  NAND4_X1 U3064 ( .A1(n2636), .A2(n2635), .A3(n2634), .A4(n2633), .ZN(n4874)
         );
  INV_X1 U3065 ( .A(DATAI_14_), .ZN(n4535) );
  NAND2_X1 U3066 ( .A1(n2637), .A2(IR_REG_31__SCAN_IN), .ZN(n2647) );
  INV_X1 U3067 ( .A(IR_REG_14__SCAN_IN), .ZN(n2638) );
  XNOR2_X1 U3068 ( .A(n2647), .B(n2638), .ZN(n4093) );
  MUX2_X1 U3069 ( .A(n4535), .B(n4093), .S(n3569), .Z(n3501) );
  OR2_X1 U3070 ( .A1(n4874), .A2(n3501), .ZN(n3887) );
  NAND2_X1 U3071 ( .A1(n4874), .A2(n3501), .ZN(n3875) );
  NAND2_X1 U3072 ( .A1(n3887), .A2(n3875), .ZN(n3945) );
  NAND2_X1 U3073 ( .A1(n2878), .A2(REG1_REG_15__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U3074 ( .A1(n2640), .A2(n2639), .ZN(n2641) );
  NAND2_X1 U3075 ( .A1(n2653), .A2(n2641), .ZN(n4890) );
  INV_X1 U3076 ( .A(n4890), .ZN(n3390) );
  NAND2_X1 U3077 ( .A1(n2753), .A2(n3390), .ZN(n2644) );
  NAND2_X1 U3078 ( .A1(n2725), .A2(REG0_REG_15__SCAN_IN), .ZN(n2643) );
  NAND2_X1 U3079 ( .A1(n2496), .A2(REG2_REG_15__SCAN_IN), .ZN(n2642) );
  NAND4_X1 U3080 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .ZN(n4045)
         );
  NAND2_X1 U3081 ( .A1(n2647), .A2(n2646), .ZN(n2664) );
  OR2_X1 U3082 ( .A1(n2664), .A2(IR_REG_15__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3083 ( .A1(n2664), .A2(IR_REG_15__SCAN_IN), .ZN(n2648) );
  MUX2_X1 U3084 ( .A(DATAI_15_), .B(n4107), .S(n3569), .Z(n4878) );
  NAND2_X1 U3085 ( .A1(n4045), .A2(n4878), .ZN(n2649) );
  NAND2_X1 U3086 ( .A1(n4046), .A2(n3483), .ZN(n3331) );
  AND3_X1 U3087 ( .A1(n3945), .A2(n2649), .A3(n3331), .ZN(n2652) );
  INV_X1 U3088 ( .A(n2649), .ZN(n2650) );
  INV_X1 U3089 ( .A(n3501), .ZN(n3505) );
  OR2_X1 U3090 ( .A1(n4874), .A2(n3505), .ZN(n3379) );
  OAI22_X1 U3091 ( .A1(n2650), .A2(n3379), .B1(n4878), .B2(n4045), .ZN(n2651)
         );
  AOI21_X2 U3092 ( .B1(n3332), .B2(n2652), .A(n2651), .ZN(n3365) );
  NAND2_X1 U3093 ( .A1(n2496), .A2(REG2_REG_16__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U3094 ( .A1(n2878), .A2(REG1_REG_16__SCAN_IN), .ZN(n2656) );
  AOI21_X1 U3095 ( .B1(n2653), .B2(n4529), .A(n2670), .ZN(n3372) );
  NAND2_X1 U3096 ( .A1(n2753), .A2(n3372), .ZN(n2655) );
  NAND2_X1 U3097 ( .A1(n2725), .A2(REG0_REG_16__SCAN_IN), .ZN(n2654) );
  NAND4_X1 U3098 ( .A1(n2657), .A2(n2656), .A3(n2655), .A4(n2654), .ZN(n4876)
         );
  INV_X1 U3099 ( .A(DATAI_16_), .ZN(n4892) );
  NAND2_X1 U3100 ( .A1(n2658), .A2(IR_REG_31__SCAN_IN), .ZN(n2659) );
  XNOR2_X1 U3101 ( .A(n2659), .B(IR_REG_16__SCAN_IN), .ZN(n4111) );
  MUX2_X1 U3102 ( .A(n4892), .B(n4893), .S(n3569), .Z(n3589) );
  OR2_X1 U3103 ( .A1(n4876), .A2(n3589), .ZN(n4003) );
  NAND2_X1 U3104 ( .A1(n4876), .A2(n3589), .ZN(n3999) );
  NAND2_X1 U3105 ( .A1(n2878), .A2(REG1_REG_18__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3106 ( .A1(n2513), .A2(REG2_REG_18__SCAN_IN), .ZN(n2662) );
  AOI21_X1 U3107 ( .B1(n3855), .B2(n2669), .A(n2683), .ZN(n3525) );
  NAND2_X1 U3108 ( .A1(n2495), .A2(n3525), .ZN(n2661) );
  NAND2_X1 U3109 ( .A1(n2725), .A2(REG0_REG_18__SCAN_IN), .ZN(n2660) );
  NAND4_X1 U3110 ( .A1(n2663), .A2(n2662), .A3(n2661), .A4(n2660), .ZN(n4043)
         );
  INV_X1 U3111 ( .A(n4043), .ZN(n4325) );
  INV_X1 U3112 ( .A(DATAI_18_), .ZN(n4456) );
  INV_X1 U3113 ( .A(n2664), .ZN(n2667) );
  INV_X1 U3114 ( .A(n2665), .ZN(n2666) );
  OR2_X1 U3115 ( .A1(n2688), .A2(n2689), .ZN(n2668) );
  XNOR2_X1 U3116 ( .A(n2668), .B(IR_REG_18__SCAN_IN), .ZN(n4144) );
  MUX2_X1 U3117 ( .A(n4456), .B(n4144), .S(n3569), .Z(n3516) );
  NAND2_X1 U3118 ( .A1(n4325), .A2(n3516), .ZN(n2677) );
  OR2_X1 U3119 ( .A1(n4043), .A2(n3516), .ZN(n4312) );
  NAND2_X1 U3120 ( .A1(n4043), .A2(n3516), .ZN(n4313) );
  NAND2_X1 U3121 ( .A1(n4312), .A2(n4313), .ZN(n3948) );
  INV_X1 U3122 ( .A(n3948), .ZN(n3535) );
  NAND2_X1 U3123 ( .A1(n2878), .A2(REG1_REG_17__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3124 ( .A1(n2513), .A2(REG2_REG_17__SCAN_IN), .ZN(n2674) );
  OAI21_X1 U3125 ( .B1(REG3_REG_17__SCAN_IN), .B2(n2670), .A(n2669), .ZN(n3809) );
  INV_X1 U3126 ( .A(n3809), .ZN(n2671) );
  NAND2_X1 U3127 ( .A1(n2753), .A2(n2671), .ZN(n2673) );
  NAND2_X1 U3128 ( .A1(n2725), .A2(REG0_REG_17__SCAN_IN), .ZN(n2672) );
  NAND4_X1 U3129 ( .A1(n2675), .A2(n2674), .A3(n2673), .A4(n2672), .ZN(n4044)
         );
  INV_X1 U3130 ( .A(n4044), .ZN(n3522) );
  INV_X1 U3131 ( .A(DATAI_17_), .ZN(n2676) );
  XNOR2_X1 U3132 ( .A(n2688), .B(IR_REG_17__SCAN_IN), .ZN(n4117) );
  MUX2_X1 U3133 ( .A(n2676), .B(n4117), .S(n3569), .Z(n3417) );
  NAND2_X1 U3134 ( .A1(n3522), .A2(n3417), .ZN(n3527) );
  INV_X1 U3135 ( .A(n2678), .ZN(n2680) );
  NAND2_X1 U3136 ( .A1(n4876), .A2(n3798), .ZN(n3412) );
  NAND2_X1 U3137 ( .A1(n4044), .A2(n3806), .ZN(n2679) );
  AND2_X1 U3138 ( .A1(n3412), .A2(n2679), .ZN(n3526) );
  AND2_X1 U3139 ( .A1(n3526), .A2(n3948), .ZN(n3529) );
  AOI21_X1 U3140 ( .B1(n3365), .B2(n2681), .A(n2435), .ZN(n4311) );
  NAND2_X1 U3141 ( .A1(n2496), .A2(REG2_REG_19__SCAN_IN), .ZN(n2687) );
  NAND2_X1 U3142 ( .A1(n2878), .A2(REG1_REG_19__SCAN_IN), .ZN(n2686) );
  INV_X1 U3143 ( .A(n2682), .ZN(n2696) );
  OAI21_X1 U3144 ( .B1(REG3_REG_19__SCAN_IN), .B2(n2683), .A(n2696), .ZN(n4329) );
  INV_X1 U3145 ( .A(n4329), .ZN(n3763) );
  NAND2_X1 U3146 ( .A1(n2753), .A2(n3763), .ZN(n2685) );
  NAND2_X1 U3147 ( .A1(n2725), .A2(REG0_REG_19__SCAN_IN), .ZN(n2684) );
  NAND4_X1 U31480 ( .A1(n2687), .A2(n2686), .A3(n2685), .A4(n2684), .ZN(n4042)
         );
  INV_X1 U31490 ( .A(DATAI_19_), .ZN(n2692) );
  NAND2_X1 U3150 ( .A1(n2759), .A2(IR_REG_19__SCAN_IN), .ZN(n2690) );
  NAND2_X2 U3151 ( .A1(n2691), .A2(n2690), .ZN(n4814) );
  MUX2_X1 U3152 ( .A(n2692), .B(n4814), .S(n3569), .Z(n4327) );
  INV_X1 U3153 ( .A(n4327), .ZN(n4319) );
  NAND2_X1 U3154 ( .A1(n4042), .A2(n4319), .ZN(n2694) );
  NOR2_X1 U3155 ( .A1(n4042), .A2(n4319), .ZN(n2693) );
  NAND2_X1 U3156 ( .A1(n2878), .A2(REG1_REG_20__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U3157 ( .A1(n2496), .A2(REG2_REG_20__SCAN_IN), .ZN(n2700) );
  INV_X1 U3158 ( .A(n2695), .ZN(n2706) );
  INV_X1 U3159 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U3160 ( .A1(n2696), .A2(n4605), .ZN(n2697) );
  AND2_X1 U3161 ( .A1(n2706), .A2(n2697), .ZN(n3562) );
  NAND2_X1 U3162 ( .A1(n2753), .A2(n3562), .ZN(n2699) );
  NAND2_X1 U3163 ( .A1(n2725), .A2(REG0_REG_20__SCAN_IN), .ZN(n2698) );
  INV_X1 U3164 ( .A(n4321), .ZN(n2702) );
  NAND2_X1 U3165 ( .A1(n2720), .A2(DATAI_20_), .ZN(n3630) );
  NAND2_X1 U3166 ( .A1(n2702), .A2(n3630), .ZN(n2703) );
  INV_X1 U3167 ( .A(n3630), .ZN(n3828) );
  NAND2_X1 U3168 ( .A1(n2878), .A2(REG1_REG_21__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3169 ( .A1(n2496), .A2(REG2_REG_21__SCAN_IN), .ZN(n2710) );
  INV_X1 U3170 ( .A(n2704), .ZN(n2713) );
  INV_X1 U3171 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U3172 ( .A1(n2706), .A2(n2705), .ZN(n2707) );
  AND2_X1 U3173 ( .A1(n2713), .A2(n2707), .ZN(n3774) );
  NAND2_X1 U3174 ( .A1(n2753), .A2(n3774), .ZN(n2709) );
  NAND2_X1 U3175 ( .A1(n2725), .A2(REG0_REG_21__SCAN_IN), .ZN(n2708) );
  NAND2_X1 U3176 ( .A1(n2720), .A2(DATAI_21_), .ZN(n4303) );
  NAND2_X1 U3177 ( .A1(n4278), .A2(n4296), .ZN(n4249) );
  NAND2_X1 U3178 ( .A1(n2496), .A2(REG2_REG_22__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U3179 ( .A1(n2878), .A2(REG1_REG_22__SCAN_IN), .ZN(n2717) );
  INV_X1 U3180 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2712) );
  NAND2_X1 U3181 ( .A1(n2713), .A2(n2712), .ZN(n2714) );
  AND2_X1 U3182 ( .A1(n2722), .A2(n2714), .ZN(n3839) );
  NAND2_X1 U3183 ( .A1(n2753), .A2(n3839), .ZN(n2716) );
  NAND2_X1 U3184 ( .A1(n2725), .A2(REG0_REG_22__SCAN_IN), .ZN(n2715) );
  NAND4_X1 U3185 ( .A1(n2718), .A2(n2717), .A3(n2716), .A4(n2715), .ZN(n4297)
         );
  NAND2_X1 U3186 ( .A1(n2720), .A2(DATAI_22_), .ZN(n4281) );
  NAND2_X1 U3187 ( .A1(n4297), .A2(n4281), .ZN(n2801) );
  NAND2_X1 U3188 ( .A1(n4256), .A2(n2801), .ZN(n4275) );
  INV_X1 U3189 ( .A(n4275), .ZN(n2719) );
  NOR2_X1 U3190 ( .A1(n4278), .A2(n4296), .ZN(n4250) );
  AOI211_X1 U3191 ( .C1(n4293), .C2(n4249), .A(n2719), .B(n4250), .ZN(n2730)
         );
  INV_X1 U3192 ( .A(n4297), .ZN(n3645) );
  NOR2_X1 U3193 ( .A1(n3645), .A2(n4281), .ZN(n4251) );
  NAND2_X1 U3194 ( .A1(n2720), .A2(DATAI_23_), .ZN(n4266) );
  NAND2_X1 U3195 ( .A1(n2513), .A2(REG2_REG_23__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U3196 ( .A1(n2878), .A2(REG1_REG_23__SCAN_IN), .ZN(n2728) );
  INV_X1 U3197 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U3198 ( .A1(n2722), .A2(n2721), .ZN(n2723) );
  NAND2_X1 U3199 ( .A1(n2753), .A2(n4267), .ZN(n2727) );
  NAND2_X1 U3200 ( .A1(n2725), .A2(REG0_REG_23__SCAN_IN), .ZN(n2726) );
  INV_X1 U3201 ( .A(n4277), .ZN(n2731) );
  OAI21_X1 U3202 ( .B1(n4218), .B2(n4237), .A(n4212), .ZN(n2733) );
  OAI21_X1 U3203 ( .B1(n3665), .B2(n4226), .A(n2733), .ZN(n4192) );
  NAND2_X1 U3204 ( .A1(n2513), .A2(REG2_REG_27__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U3205 ( .A1(n2878), .A2(REG1_REG_27__SCAN_IN), .ZN(n2741) );
  NAND2_X1 U3206 ( .A1(n2735), .A2(REG3_REG_27__SCAN_IN), .ZN(n2746) );
  INV_X1 U3207 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2736) );
  NAND2_X1 U3208 ( .A1(n2737), .A2(n2736), .ZN(n2738) );
  NAND2_X1 U3209 ( .A1(n2753), .A2(n4179), .ZN(n2740) );
  NAND2_X1 U32100 ( .A1(n2725), .A2(REG0_REG_27__SCAN_IN), .ZN(n2739) );
  NAND2_X1 U32110 ( .A1(n2720), .A2(DATAI_27_), .ZN(n4185) );
  NAND2_X1 U32120 ( .A1(n4165), .A2(n4185), .ZN(n2743) );
  INV_X1 U32130 ( .A(n4198), .ZN(n4165) );
  NAND2_X1 U32140 ( .A1(n2513), .A2(REG2_REG_28__SCAN_IN), .ZN(n2751) );
  NAND2_X1 U32150 ( .A1(n2878), .A2(REG1_REG_28__SCAN_IN), .ZN(n2750) );
  INV_X1 U32160 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U32170 ( .A1(n2746), .A2(n3726), .ZN(n2747) );
  NAND2_X1 U32180 ( .A1(n2753), .A2(n4154), .ZN(n2749) );
  NAND2_X1 U32190 ( .A1(n2725), .A2(REG0_REG_28__SCAN_IN), .ZN(n2748) );
  NAND4_X1 U32200 ( .A1(n2751), .A2(n2750), .A3(n2749), .A4(n2748), .ZN(n4175)
         );
  NAND2_X1 U32210 ( .A1(n2720), .A2(DATAI_28_), .ZN(n4157) );
  OR2_X1 U32220 ( .A1(n4175), .A2(n4157), .ZN(n2806) );
  NAND2_X1 U32230 ( .A1(n4175), .A2(n4157), .ZN(n3934) );
  NAND2_X1 U32240 ( .A1(n2806), .A2(n3934), .ZN(n4160) );
  INV_X1 U32250 ( .A(n4157), .ZN(n4162) );
  NAND2_X1 U32260 ( .A1(n2513), .A2(REG2_REG_29__SCAN_IN), .ZN(n2757) );
  NAND2_X1 U32270 ( .A1(n2878), .A2(REG1_REG_29__SCAN_IN), .ZN(n2756) );
  INV_X1 U32280 ( .A(n4146), .ZN(n2752) );
  NAND2_X1 U32290 ( .A1(n2753), .A2(n2752), .ZN(n2755) );
  NAND2_X1 U32300 ( .A1(n2725), .A2(REG0_REG_29__SCAN_IN), .ZN(n2754) );
  NAND4_X1 U32310 ( .A1(n2757), .A2(n2756), .A3(n2755), .A4(n2754), .ZN(n4163)
         );
  NAND2_X1 U32320 ( .A1(n2720), .A2(DATAI_29_), .ZN(n3938) );
  XNOR2_X1 U32330 ( .A(n4163), .B(n3938), .ZN(n3984) );
  XNOR2_X1 U32340 ( .A(n2758), .B(n3984), .ZN(n4145) );
  NAND2_X1 U32350 ( .A1(n2762), .A2(IR_REG_31__SCAN_IN), .ZN(n2763) );
  INV_X1 U32360 ( .A(n2764), .ZN(n2765) );
  NAND2_X1 U32370 ( .A1(n2765), .A2(IR_REG_31__SCAN_IN), .ZN(n2766) );
  XNOR2_X1 U32380 ( .A(n3044), .B(n4038), .ZN(n2767) );
  NAND2_X1 U32390 ( .A1(n2767), .A2(n4814), .ZN(n3557) );
  NAND2_X1 U32400 ( .A1(n2768), .A2(n4168), .ZN(n4752) );
  NAND2_X1 U32410 ( .A1(n3557), .A2(n4760), .ZN(n4826) );
  NAND2_X1 U32420 ( .A1(n2878), .A2(REG1_REG_30__SCAN_IN), .ZN(n2771) );
  NAND2_X1 U32430 ( .A1(n2513), .A2(REG2_REG_30__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U32440 ( .A1(n2725), .A2(REG0_REG_30__SCAN_IN), .ZN(n2769) );
  AND3_X1 U32450 ( .A1(n2771), .A2(n2770), .A3(n2769), .ZN(n3935) );
  OR2_X1 U32460 ( .A1(n2772), .A2(n2820), .ZN(n2774) );
  XNOR2_X1 U32470 ( .A(n2774), .B(n2773), .ZN(n4895) );
  AND2_X2 U32480 ( .A1(n4895), .A2(n2941), .ZN(n4320) );
  XNOR2_X1 U32490 ( .A(n2775), .B(IR_REG_27__SCAN_IN), .ZN(n4060) );
  NAND2_X1 U32500 ( .A1(n4060), .A2(B_REG_SCAN_IN), .ZN(n2776) );
  NAND2_X1 U32510 ( .A1(n4320), .A2(n2776), .ZN(n3570) );
  INV_X1 U32520 ( .A(n3030), .ZN(n3959) );
  NOR2_X1 U32530 ( .A1(n2912), .A2(n3698), .ZN(n3894) );
  NAND2_X1 U32540 ( .A1(n3959), .A2(n3894), .ZN(n3031) );
  NAND2_X1 U32550 ( .A1(n3031), .A2(n3895), .ZN(n2988) );
  INV_X1 U32560 ( .A(n2987), .ZN(n3960) );
  NAND2_X1 U32570 ( .A1(n2988), .A2(n3960), .ZN(n2777) );
  NAND2_X1 U32580 ( .A1(n2777), .A2(n3896), .ZN(n3000) );
  OR2_X1 U32590 ( .A1(n4055), .A2(n3008), .ZN(n3901) );
  NAND2_X1 U32600 ( .A1(n4055), .A2(n3008), .ZN(n3898) );
  NAND2_X1 U32610 ( .A1(n3901), .A2(n3898), .ZN(n2997) );
  INV_X1 U32620 ( .A(n2997), .ZN(n3958) );
  NAND2_X1 U32630 ( .A1(n3000), .A2(n3958), .ZN(n2999) );
  NAND2_X1 U32640 ( .A1(n2999), .A2(n3901), .ZN(n3070) );
  INV_X1 U32650 ( .A(n3902), .ZN(n2778) );
  OR2_X1 U32660 ( .A1(n3070), .A2(n2778), .ZN(n2779) );
  NAND2_X1 U32670 ( .A1(n2779), .A2(n3906), .ZN(n3059) );
  AND2_X1 U32680 ( .A1(n4053), .A2(n3108), .ZN(n3057) );
  OR2_X1 U32690 ( .A1(n4053), .A2(n3108), .ZN(n3881) );
  OAI21_X1 U32700 ( .B1(n3059), .B2(n3057), .A(n3881), .ZN(n3140) );
  INV_X1 U32710 ( .A(n3148), .ZN(n2780) );
  NAND2_X1 U32720 ( .A1(n4802), .A2(n2780), .ZN(n3905) );
  NAND2_X1 U32730 ( .A1(n3140), .A2(n3905), .ZN(n4797) );
  OR2_X1 U32740 ( .A1(n4802), .A2(n2780), .ZN(n4796) );
  OR2_X1 U32750 ( .A1(n4052), .A2(n4809), .ZN(n2781) );
  AND2_X1 U32760 ( .A1(n4796), .A2(n2781), .ZN(n3909) );
  NAND2_X1 U32770 ( .A1(n4797), .A2(n3909), .ZN(n2782) );
  NAND2_X1 U32780 ( .A1(n4052), .A2(n4809), .ZN(n3877) );
  NAND2_X1 U32790 ( .A1(n2782), .A2(n3877), .ZN(n3174) );
  OR2_X1 U32800 ( .A1(n4051), .A2(n3204), .ZN(n3912) );
  NAND2_X1 U32810 ( .A1(n3174), .A2(n3912), .ZN(n2783) );
  NAND2_X1 U32820 ( .A1(n4051), .A2(n3204), .ZN(n3878) );
  NAND2_X1 U32830 ( .A1(n2783), .A2(n3878), .ZN(n3158) );
  AND2_X1 U32840 ( .A1(n4050), .A2(n3220), .ZN(n3911) );
  OR2_X1 U32850 ( .A1(n4050), .A2(n3220), .ZN(n3913) );
  NAND2_X1 U32860 ( .A1(n2784), .A2(n3913), .ZN(n3241) );
  NAND2_X1 U32870 ( .A1(n4049), .A2(n3244), .ZN(n3882) );
  NAND2_X1 U32880 ( .A1(n3241), .A2(n3882), .ZN(n2785) );
  OR2_X1 U32890 ( .A1(n4049), .A2(n3244), .ZN(n3885) );
  NAND2_X1 U32900 ( .A1(n2785), .A2(n3885), .ZN(n3299) );
  NAND2_X1 U32910 ( .A1(n4047), .A2(n2301), .ZN(n3345) );
  INV_X1 U32920 ( .A(n3483), .ZN(n3358) );
  NAND2_X1 U32930 ( .A1(n4046), .A2(n3358), .ZN(n2786) );
  NAND2_X1 U32940 ( .A1(n3345), .A2(n2786), .ZN(n2788) );
  INV_X1 U32950 ( .A(n3258), .ZN(n2787) );
  NOR2_X1 U32960 ( .A1(n2788), .A2(n2787), .ZN(n3883) );
  NAND2_X1 U32970 ( .A1(n3299), .A2(n3883), .ZN(n2792) );
  INV_X1 U32980 ( .A(n2788), .ZN(n2791) );
  OR2_X1 U32990 ( .A1(n4047), .A2(n2301), .ZN(n3347) );
  NAND2_X1 U33000 ( .A1(n3256), .A2(n3347), .ZN(n2790) );
  NOR2_X1 U33010 ( .A1(n4046), .A2(n3358), .ZN(n2789) );
  AOI21_X1 U33020 ( .B1(n2791), .B2(n2790), .A(n2789), .ZN(n3888) );
  NAND2_X1 U33030 ( .A1(n2792), .A2(n3888), .ZN(n4001) );
  INV_X1 U33040 ( .A(n3945), .ZN(n3334) );
  NAND2_X1 U33050 ( .A1(n4001), .A2(n3334), .ZN(n3382) );
  OR2_X1 U33060 ( .A1(n4045), .A2(n3388), .ZN(n3886) );
  NAND2_X1 U33070 ( .A1(n4045), .A2(n3388), .ZN(n3876) );
  NAND2_X1 U33080 ( .A1(n3886), .A2(n3876), .ZN(n3953) );
  INV_X1 U33090 ( .A(n3887), .ZN(n2793) );
  NOR2_X1 U33100 ( .A1(n3953), .A2(n2793), .ZN(n2794) );
  NAND2_X1 U33110 ( .A1(n3382), .A2(n2794), .ZN(n2795) );
  NAND2_X1 U33120 ( .A1(n2795), .A2(n3876), .ZN(n3367) );
  NAND2_X1 U33130 ( .A1(n3367), .A2(n3952), .ZN(n2796) );
  NAND2_X1 U33140 ( .A1(n2796), .A2(n3999), .ZN(n3520) );
  NAND2_X1 U33150 ( .A1(n4042), .A2(n4327), .ZN(n3942) );
  AND2_X1 U33160 ( .A1(n4313), .A2(n3942), .ZN(n2798) );
  NAND2_X1 U33170 ( .A1(n4044), .A2(n3417), .ZN(n3517) );
  AND2_X1 U33180 ( .A1(n2798), .A2(n3517), .ZN(n3548) );
  NAND2_X1 U33190 ( .A1(n4321), .A2(n3630), .ZN(n3550) );
  AND2_X1 U33200 ( .A1(n3548), .A2(n3550), .ZN(n3921) );
  INV_X1 U33210 ( .A(n3921), .ZN(n4002) );
  OR2_X2 U33220 ( .A1(n3520), .A2(n4002), .ZN(n2800) );
  OR2_X1 U33230 ( .A1(n4044), .A2(n3417), .ZN(n3518) );
  NAND2_X1 U33240 ( .A1(n4312), .A2(n3518), .ZN(n2797) );
  NAND2_X1 U33250 ( .A1(n2798), .A2(n2797), .ZN(n2799) );
  OR2_X1 U33260 ( .A1(n4042), .A2(n4327), .ZN(n3943) );
  NAND2_X1 U33270 ( .A1(n2799), .A2(n3943), .ZN(n3547) );
  NOR2_X1 U33280 ( .A1(n4321), .A2(n3630), .ZN(n3551) );
  OAI21_X1 U33290 ( .B1(n3547), .B2(n3551), .A(n3550), .ZN(n4005) );
  NAND2_X2 U33300 ( .A1(n2800), .A2(n4005), .ZN(n4295) );
  OR2_X1 U33310 ( .A1(n4278), .A2(n4303), .ZN(n4253) );
  NAND2_X1 U33320 ( .A1(n4256), .A2(n4253), .ZN(n3924) );
  NAND2_X1 U33330 ( .A1(n4277), .A2(n4266), .ZN(n3966) );
  AND2_X1 U33340 ( .A1(n2801), .A2(n3966), .ZN(n3927) );
  AND2_X1 U33350 ( .A1(n4278), .A2(n4303), .ZN(n3946) );
  NAND2_X1 U33360 ( .A1(n3946), .A2(n4256), .ZN(n2802) );
  NAND2_X1 U33370 ( .A1(n3927), .A2(n2802), .ZN(n4008) );
  INV_X1 U33380 ( .A(n4008), .ZN(n2803) );
  NAND2_X1 U33390 ( .A1(n2804), .A2(n2803), .ZN(n4233) );
  OR2_X1 U33400 ( .A1(n4277), .A2(n4266), .ZN(n4232) );
  OR2_X1 U33410 ( .A1(n4260), .A2(n4241), .ZN(n3965) );
  NAND2_X1 U33420 ( .A1(n4232), .A2(n3965), .ZN(n4012) );
  INV_X1 U33430 ( .A(n4012), .ZN(n2805) );
  NAND2_X1 U33440 ( .A1(n4233), .A2(n2805), .ZN(n4214) );
  NAND2_X1 U33450 ( .A1(n4260), .A2(n4241), .ZN(n4213) );
  NAND2_X1 U33460 ( .A1(n4237), .A2(n4226), .ZN(n3964) );
  OR2_X1 U33470 ( .A1(n4237), .A2(n4226), .ZN(n4193) );
  OR2_X1 U33480 ( .A1(n4219), .A2(n4201), .ZN(n3970) );
  NAND2_X1 U33490 ( .A1(n4193), .A2(n3970), .ZN(n3995) );
  NAND2_X1 U33500 ( .A1(n4219), .A2(n4201), .ZN(n3992) );
  NAND2_X1 U33510 ( .A1(n4198), .A2(n4185), .ZN(n3932) );
  NOR2_X2 U33520 ( .A1(n4174), .A2(n4173), .ZN(n4172) );
  NAND2_X1 U3353 ( .A1(n4158), .A2(n2806), .ZN(n3996) );
  OAI21_X1 U33540 ( .B1(n4172), .B2(n3996), .A(n3934), .ZN(n2807) );
  XNOR2_X1 U3355 ( .A(n2807), .B(n3984), .ZN(n2810) );
  INV_X1 U3356 ( .A(n2768), .ZN(n4027) );
  NAND2_X1 U3357 ( .A1(n4027), .A2(n4023), .ZN(n2809) );
  INV_X1 U3358 ( .A(n4038), .ZN(n2812) );
  OR2_X1 U3359 ( .A1(n4814), .A2(n2812), .ZN(n2808) );
  NAND2_X1 U3360 ( .A1(n2810), .A2(n4807), .ZN(n2815) );
  INV_X1 U3361 ( .A(n2941), .ZN(n2811) );
  NOR2_X2 U3362 ( .A1(n4895), .A2(n2811), .ZN(n4801) );
  INV_X1 U3363 ( .A(n4023), .ZN(n2955) );
  NAND2_X1 U3364 ( .A1(n4027), .A2(n2942), .ZN(n4282) );
  NOR2_X1 U3365 ( .A1(n3938), .A2(n4282), .ZN(n2813) );
  AOI21_X1 U3366 ( .B1(n4175), .B2(n4801), .A(n2813), .ZN(n2814) );
  OAI211_X1 U3367 ( .C1(n3935), .C2(n3570), .A(n2815), .B(n2814), .ZN(n4149)
         );
  AOI21_X1 U3368 ( .B1(n4145), .B2(n4826), .A(n4149), .ZN(n2857) );
  NOR2_X1 U3369 ( .A1(n4760), .A2(n4023), .ZN(n2829) );
  NAND2_X1 U3370 ( .A1(n2764), .A2(n2816), .ZN(n2817) );
  NAND2_X1 U3371 ( .A1(n2817), .A2(IR_REG_31__SCAN_IN), .ZN(n2818) );
  AND2_X1 U3372 ( .A1(n2764), .A2(n2819), .ZN(n2821) );
  INV_X1 U3373 ( .A(IR_REG_23__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U3374 ( .A1(n2828), .A2(n2827), .ZN(n2822) );
  NAND2_X1 U3375 ( .A1(n2822), .A2(IR_REG_31__SCAN_IN), .ZN(n2823) );
  NAND2_X1 U3376 ( .A1(n2764), .A2(n2824), .ZN(n2825) );
  NAND2_X1 U3377 ( .A1(n2825), .A2(IR_REG_31__SCAN_IN), .ZN(n2826) );
  XNOR2_X1 U3378 ( .A(n2826), .B(IR_REG_25__SCAN_IN), .ZN(n4429) );
  NAND3_X1 U3379 ( .A1(n4428), .A2(n2838), .A3(n4429), .ZN(n2903) );
  INV_X1 U3380 ( .A(n2903), .ZN(n2949) );
  XNOR2_X1 U3381 ( .A(n2828), .B(n2827), .ZN(n4034) );
  NAND2_X1 U3382 ( .A1(n2768), .A2(n4814), .ZN(n2943) );
  NAND2_X1 U3383 ( .A1(n2943), .A2(n2941), .ZN(n2947) );
  NAND2_X1 U3384 ( .A1(n3087), .A2(n2947), .ZN(n3038) );
  NOR2_X1 U3385 ( .A1(n2829), .A2(n3038), .ZN(n2846) );
  NOR4_X1 U3386 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2833) );
  NOR4_X1 U3387 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2832) );
  NOR4_X1 U3388 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2831) );
  NOR4_X1 U3389 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2830) );
  NAND4_X1 U3390 ( .A1(n2833), .A2(n2832), .A3(n2831), .A4(n2830), .ZN(n2842)
         );
  NOR2_X1 U3391 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_31__SCAN_IN), .ZN(n2837)
         );
  NOR4_X1 U3392 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2836) );
  NOR4_X1 U3393 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2835) );
  NOR4_X1 U3394 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2834) );
  NAND4_X1 U3395 ( .A1(n2837), .A2(n2836), .A3(n2835), .A4(n2834), .ZN(n2841)
         );
  INV_X1 U3396 ( .A(n4429), .ZN(n2844) );
  NAND2_X1 U3397 ( .A1(n2847), .A2(n2844), .ZN(n2839) );
  MUX2_X1 U3398 ( .A(n2847), .B(n2839), .S(B_REG_SCAN_IN), .Z(n2840) );
  OAI21_X1 U3399 ( .B1(n2842), .B2(n2841), .A(n2870), .ZN(n2938) );
  INV_X1 U3400 ( .A(D_REG_1__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U3401 ( .A1(n2870), .A2(n2843), .ZN(n3039) );
  INV_X1 U3402 ( .A(n4428), .ZN(n2848) );
  NAND2_X1 U3403 ( .A1(n2848), .A2(n2844), .ZN(n2937) );
  NAND2_X1 U3404 ( .A1(n3039), .A2(n2937), .ZN(n2845) );
  INV_X1 U3405 ( .A(D_REG_0__SCAN_IN), .ZN(n2874) );
  INV_X1 U3406 ( .A(n2939), .ZN(n3042) );
  NAND2_X1 U3407 ( .A1(n3698), .A2(n3034), .ZN(n3048) );
  NAND2_X1 U3408 ( .A1(n4810), .A2(n4809), .ZN(n4813) );
  INV_X1 U3409 ( .A(n4281), .ZN(n4288) );
  OAI21_X1 U3410 ( .B1(n4155), .B2(n3938), .A(n2273), .ZN(n4147) );
  OR2_X1 U3411 ( .A1(n4147), .A2(n4423), .ZN(n2850) );
  NAND2_X1 U3412 ( .A1(n4832), .A2(REG0_REG_29__SCAN_IN), .ZN(n2849) );
  OAI21_X1 U3413 ( .B1(n2857), .B2(n4832), .A(n2851), .ZN(U3515) );
  OAI21_X1 U3414 ( .B1(n2857), .B2(n2856), .A(n2855), .ZN(U3547) );
  INV_X2 U3415 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3416 ( .A(n2872), .ZN(n2858) );
  OR2_X2 U3417 ( .A1(n2903), .A2(n2858), .ZN(n4058) );
  INV_X1 U3418 ( .A(n4058), .ZN(U4043) );
  MUX2_X1 U3419 ( .A(n2524), .B(n3447), .S(STATE_REG_SCAN_IN), .Z(n2859) );
  INV_X1 U3420 ( .A(n2859), .ZN(U3348) );
  INV_X1 U3421 ( .A(DATAI_15_), .ZN(n4537) );
  NAND2_X1 U3422 ( .A1(n4107), .A2(STATE_REG_SCAN_IN), .ZN(n2860) );
  OAI21_X1 U3423 ( .B1(STATE_REG_SCAN_IN), .B2(n4537), .A(n2860), .ZN(U3337)
         );
  INV_X1 U3424 ( .A(DATAI_21_), .ZN(n4553) );
  NAND2_X1 U3425 ( .A1(n4023), .A2(STATE_REG_SCAN_IN), .ZN(n2861) );
  OAI21_X1 U3426 ( .B1(STATE_REG_SCAN_IN), .B2(n4553), .A(n2861), .ZN(U3331)
         );
  INV_X1 U3427 ( .A(n4117), .ZN(n4130) );
  NAND2_X1 U3428 ( .A1(n4130), .A2(STATE_REG_SCAN_IN), .ZN(n2862) );
  OAI21_X1 U3429 ( .B1(STATE_REG_SCAN_IN), .B2(n2676), .A(n2862), .ZN(U3335)
         );
  INV_X1 U3430 ( .A(DATAI_22_), .ZN(n2864) );
  NAND2_X1 U3431 ( .A1(n4038), .A2(STATE_REG_SCAN_IN), .ZN(n2863) );
  OAI21_X1 U3432 ( .B1(STATE_REG_SCAN_IN), .B2(n2864), .A(n2863), .ZN(U3330)
         );
  INV_X1 U3433 ( .A(DATAI_27_), .ZN(n4541) );
  NAND2_X1 U3434 ( .A1(n4060), .A2(STATE_REG_SCAN_IN), .ZN(n2865) );
  OAI21_X1 U3435 ( .B1(STATE_REG_SCAN_IN), .B2(n4541), .A(n2865), .ZN(U3325)
         );
  MUX2_X1 U3436 ( .A(n2692), .B(n4814), .S(STATE_REG_SCAN_IN), .Z(n2866) );
  INV_X1 U3437 ( .A(n2866), .ZN(U3333) );
  INV_X1 U3438 ( .A(DATAI_29_), .ZN(n4444) );
  NAND2_X1 U3439 ( .A1(n2463), .A2(STATE_REG_SCAN_IN), .ZN(n2867) );
  OAI21_X1 U3440 ( .B1(STATE_REG_SCAN_IN), .B2(n4444), .A(n2867), .ZN(U3323)
         );
  INV_X1 U3441 ( .A(DATAI_20_), .ZN(n2869) );
  NAND2_X1 U3442 ( .A1(n4027), .A2(STATE_REG_SCAN_IN), .ZN(n2868) );
  OAI21_X1 U3443 ( .B1(STATE_REG_SCAN_IN), .B2(n2869), .A(n2868), .ZN(U3332)
         );
  INV_X1 U3444 ( .A(n2870), .ZN(n2871) );
  NAND2_X2 U3445 ( .A1(n2871), .A2(n3087), .ZN(n4434) );
  AOI22_X1 U3446 ( .A1(n4434), .A2(n2874), .B1(n2873), .B2(n2872), .ZN(U3458)
         );
  AND2_X1 U3447 ( .A1(n4034), .A2(n2941), .ZN(n2875) );
  NOR2_X1 U3448 ( .A1(n3569), .A2(n2875), .ZN(n2887) );
  INV_X1 U3449 ( .A(n2887), .ZN(n2877) );
  OR2_X1 U3450 ( .A1(n4034), .A2(U3149), .ZN(n4433) );
  INV_X1 U3451 ( .A(n4433), .ZN(n2876) );
  NOR2_X1 U3452 ( .A1(n4737), .A2(U4043), .ZN(U3148) );
  NAND2_X1 U3453 ( .A1(n2878), .A2(REG1_REG_31__SCAN_IN), .ZN(n2881) );
  NAND2_X1 U3454 ( .A1(n2513), .A2(REG2_REG_31__SCAN_IN), .ZN(n2880) );
  NAND2_X1 U3455 ( .A1(n2725), .A2(REG0_REG_31__SCAN_IN), .ZN(n2879) );
  AND3_X1 U3456 ( .A1(n2881), .A2(n2880), .A3(n2879), .ZN(n4019) );
  NAND2_X1 U3457 ( .A1(n4058), .A2(DATAO_REG_31__SCAN_IN), .ZN(n2882) );
  OAI21_X1 U34580 ( .B1(n4019), .B2(n4058), .A(n2882), .ZN(U3581) );
  NAND2_X1 U34590 ( .A1(n4058), .A2(DATAO_REG_30__SCAN_IN), .ZN(n2883) );
  OAI21_X1 U3460 ( .B1(n3935), .B2(n4058), .A(n2883), .ZN(U3580) );
  INV_X1 U3461 ( .A(n4434), .ZN(n2885) );
  NAND2_X1 U3462 ( .A1(n2885), .A2(n2937), .ZN(n2884) );
  OAI21_X1 U3463 ( .B1(n2885), .B2(n2843), .A(n2884), .ZN(U3459) );
  NAND2_X1 U3464 ( .A1(n4062), .A2(n4895), .ZN(n4747) );
  INV_X1 U3465 ( .A(n4060), .ZN(n2980) );
  NAND2_X1 U3466 ( .A1(n4432), .A2(REG1_REG_1__SCAN_IN), .ZN(n2889) );
  INV_X1 U34670 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4764) );
  NAND2_X1 U3468 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n4069) );
  AOI21_X1 U34690 ( .B1(n4068), .B2(n4764), .A(n4069), .ZN(n2888) );
  NAND2_X1 U3470 ( .A1(n2889), .A2(n2888), .ZN(n4072) );
  NAND2_X1 U34710 ( .A1(n4072), .A2(n2889), .ZN(n4083) );
  XNOR2_X1 U3472 ( .A(n2971), .B(n4431), .ZN(n2973) );
  XOR2_X1 U34730 ( .A(REG1_REG_3__SCAN_IN), .B(n2973), .Z(n2897) );
  INV_X1 U3474 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2895) );
  INV_X1 U34750 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2892) );
  AND2_X1 U3476 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4074)
         );
  NAND2_X1 U34770 ( .A1(n4075), .A2(n4074), .ZN(n4073) );
  NAND2_X1 U3478 ( .A1(n4432), .A2(REG2_REG_1__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U34790 ( .A1(n4073), .A2(n2891), .ZN(n4081) );
  MUX2_X1 U3480 ( .A(n2892), .B(REG2_REG_2__SCAN_IN), .S(n4087), .Z(n4082) );
  NOR2_X1 U34810 ( .A1(n4895), .A2(n2980), .ZN(n2893) );
  AOI211_X1 U3482 ( .C1(n2895), .C2(n2894), .A(n2967), .B(n4748), .ZN(n2896)
         );
  AOI21_X1 U34830 ( .B1(n4744), .B2(n2897), .A(n2896), .ZN(n2899) );
  INV_X1 U3484 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4772) );
  NOR2_X1 U34850 ( .A1(STATE_REG_SCAN_IN), .A2(n4772), .ZN(n2961) );
  AOI21_X1 U3486 ( .B1(n4737), .B2(ADDR_REG_3__SCAN_IN), .A(n2961), .ZN(n2898)
         );
  OAI211_X1 U34870 ( .C1(n2347), .C2(n4747), .A(n2899), .B(n2898), .ZN(U3243)
         );
  INV_X1 U3488 ( .A(n4760), .ZN(n4781) );
  AND2_X1 U34890 ( .A1(n2912), .A2(n3698), .ZN(n3891) );
  OR2_X1 U3490 ( .A1(n3891), .A2(n3894), .ZN(n4754) );
  AND2_X1 U34910 ( .A1(n3047), .A2(n2942), .ZN(n4753) );
  INV_X1 U3492 ( .A(n4320), .ZN(n4804) );
  INV_X1 U34930 ( .A(n3557), .ZN(n3298) );
  OAI21_X1 U3494 ( .B1(n3298), .B2(n4807), .A(n4754), .ZN(n2900) );
  OAI21_X1 U34950 ( .B1(n2425), .B2(n4804), .A(n2900), .ZN(n4751) );
  AOI211_X1 U3496 ( .C1(n4781), .C2(n4754), .A(n4753), .B(n4751), .ZN(n4750)
         );
  NAND2_X1 U34970 ( .A1(n2856), .A2(REG1_REG_0__SCAN_IN), .ZN(n2901) );
  OAI21_X1 U3498 ( .B1(n4750), .B2(n2856), .A(n2901), .ZN(U3518) );
  INV_X1 U34990 ( .A(n3044), .ZN(n2902) );
  NAND2_X1 U3500 ( .A1(n2909), .A2(n2921), .ZN(n2905) );
  AND2_X4 U35010 ( .A1(n3044), .A2(n2903), .ZN(n3718) );
  NAND2_X1 U3502 ( .A1(n3089), .A2(n3718), .ZN(n2904) );
  NAND2_X1 U35030 ( .A1(n2905), .A2(n2904), .ZN(n2906) );
  NAND2_X1 U3504 ( .A1(n4814), .A2(n4038), .ZN(n4033) );
  INV_X1 U35050 ( .A(n4811), .ZN(n4759) );
  AND2_X2 U35060 ( .A1(n3718), .A2(n4759), .ZN(n2933) );
  INV_X1 U35070 ( .A(n2921), .ZN(n2907) );
  AOI21_X1 U35080 ( .B1(n2909), .B2(n2933), .A(n2908), .ZN(n2917) );
  XNOR2_X1 U35090 ( .A(n2916), .B(n2917), .ZN(n3083) );
  NAND2_X1 U35100 ( .A1(n2912), .A2(n2933), .ZN(n2911) );
  AOI22_X1 U35110 ( .A1(n3047), .A2(n2921), .B1(n2949), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2910) );
  NAND2_X1 U35120 ( .A1(n2911), .A2(n2910), .ZN(n2977) );
  NAND2_X1 U35130 ( .A1(n2921), .A2(n2912), .ZN(n2914) );
  AND2_X1 U35140 ( .A1(n2914), .A2(n2913), .ZN(n2915) );
  INV_X1 U35150 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U35160 ( .A1(n2977), .A2(n2976), .B1(n3671), .B2(n2915), .ZN(n3084)
         );
  OAI22_X1 U35170 ( .A1(n3083), .A2(n3084), .B1(n2917), .B2(n2916), .ZN(n3701)
         );
  NAND2_X1 U35180 ( .A1(n2923), .A2(n2921), .ZN(n2919) );
  NAND2_X1 U35190 ( .A1(n3702), .A2(n3718), .ZN(n2918) );
  NAND2_X1 U35200 ( .A1(n2919), .A2(n2918), .ZN(n2920) );
  XNOR2_X1 U35210 ( .A(n2920), .B(n3671), .ZN(n2927) );
  NOR2_X1 U35220 ( .A1(n2922), .A2(n4037), .ZN(n2925) );
  NAND2_X1 U35230 ( .A1(n2927), .A2(n2926), .ZN(n2928) );
  OAI21_X1 U35240 ( .B1(n2927), .B2(n2926), .A(n2928), .ZN(n3700) );
  INV_X1 U35250 ( .A(n2928), .ZN(n2929) );
  NOR2_X1 U35260 ( .A1(n3699), .A2(n2929), .ZN(n2936) );
  NAND2_X1 U35270 ( .A1(n4055), .A2(n2921), .ZN(n2931) );
  NAND2_X1 U35280 ( .A1(n3002), .A2(n3718), .ZN(n2930) );
  NAND2_X1 U35290 ( .A1(n2931), .A2(n2930), .ZN(n2932) );
  XNOR2_X1 U35300 ( .A(n2932), .B(n3720), .ZN(n3017) );
  OAI22_X1 U35310 ( .A1(n2934), .A2(n3664), .B1(n4037), .B2(n3008), .ZN(n3016)
         );
  XNOR2_X1 U35320 ( .A(n3017), .B(n3016), .ZN(n2935) );
  AOI21_X1 U35330 ( .B1(n2936), .B2(n2935), .A(n3018), .ZN(n2966) );
  AND2_X1 U35340 ( .A1(n2938), .A2(n2937), .ZN(n3041) );
  NAND3_X1 U35350 ( .A1(n3041), .A2(n2939), .A3(n3039), .ZN(n2959) );
  INV_X1 U35360 ( .A(n3087), .ZN(n2940) );
  NOR2_X1 U35370 ( .A1(n2959), .A2(n2940), .ZN(n2954) );
  INV_X1 U35380 ( .A(n2954), .ZN(n2945) );
  AOI21_X1 U35390 ( .B1(n2943), .B2(n2942), .A(n2941), .ZN(n2946) );
  INV_X1 U35400 ( .A(n2946), .ZN(n2944) );
  NAND2_X1 U35410 ( .A1(n2959), .A2(n2946), .ZN(n2948) );
  NAND2_X1 U35420 ( .A1(n2948), .A2(n2947), .ZN(n3085) );
  OAI21_X1 U35430 ( .B1(n3085), .B2(n2949), .A(STATE_REG_SCAN_IN), .ZN(n2953)
         );
  NOR2_X1 U35440 ( .A1(n3044), .A2(n4033), .ZN(n2950) );
  NAND2_X1 U35450 ( .A1(n2950), .A2(n3087), .ZN(n2958) );
  OAI21_X1 U35460 ( .B1(U3149), .B2(n4282), .A(n2958), .ZN(n2951) );
  NAND2_X1 U35470 ( .A1(n2959), .A2(n2951), .ZN(n3086) );
  AND2_X1 U35480 ( .A1(n3086), .A2(n4433), .ZN(n2952) );
  AND2_X2 U35490 ( .A1(n2953), .A2(n2952), .ZN(n4891) );
  NAND2_X1 U35500 ( .A1(n2954), .A2(n4800), .ZN(n2957) );
  NAND2_X1 U35510 ( .A1(n3087), .A2(n2955), .ZN(n2956) );
  OR2_X1 U35520 ( .A1(n2959), .A2(n2958), .ZN(n2960) );
  INV_X1 U35530 ( .A(n4895), .ZN(n2978) );
  AOI22_X1 U35540 ( .A1(n4879), .A2(n3002), .B1(n3840), .B2(n4054), .ZN(n2963)
         );
  OR2_X1 U35550 ( .A1(n2960), .A2(n4895), .ZN(n3760) );
  AOI21_X1 U35560 ( .B1(n4875), .B2(n4056), .A(n2961), .ZN(n2962) );
  OAI211_X1 U35570 ( .C1(n4891), .C2(REG3_REG_3__SCAN_IN), .A(n2963), .B(n2962), .ZN(n2964) );
  INV_X1 U35580 ( .A(n2964), .ZN(n2965) );
  OAI21_X1 U35590 ( .B1(n2966), .B2(n3871), .A(n2965), .ZN(U3215) );
  AND2_X1 U35600 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3022) );
  AOI21_X1 U35610 ( .B1(n4431), .B2(n2968), .A(n2967), .ZN(n3425) );
  XNOR2_X1 U35620 ( .A(n3425), .B(n2969), .ZN(n2970) );
  OAI21_X1 U35630 ( .B1(REG2_REG_4__SCAN_IN), .B2(n2970), .A(n4710), .ZN(n2983) );
  INV_X1 U35640 ( .A(n2971), .ZN(n2972) );
  XNOR2_X1 U35650 ( .A(REG1_REG_4__SCAN_IN), .B(n3450), .ZN(n2974) );
  NAND2_X1 U35660 ( .A1(n4744), .A2(n2974), .ZN(n2982) );
  INV_X1 U35670 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4756) );
  AND2_X1 U35680 ( .A1(n4060), .A2(n4756), .ZN(n2975) );
  NOR2_X1 U35690 ( .A1(n4895), .A2(n2975), .ZN(n4064) );
  XOR2_X1 U35700 ( .A(n2976), .B(n2977), .Z(n3695) );
  NAND2_X1 U35710 ( .A1(n3695), .A2(n2980), .ZN(n2979) );
  OAI211_X1 U35720 ( .C1(n4074), .C2(n2980), .A(n2979), .B(n2978), .ZN(n2981)
         );
  OAI211_X1 U35730 ( .C1(IR_REG_0__SCAN_IN), .C2(n4064), .A(n2981), .B(U4043), 
        .ZN(n4091) );
  OAI211_X1 U35740 ( .C1(n3426), .C2(n2983), .A(n2982), .B(n4091), .ZN(n2984)
         );
  AOI211_X1 U35750 ( .C1(n4737), .C2(ADDR_REG_4__SCAN_IN), .A(n3022), .B(n2984), .ZN(n2985) );
  OAI21_X1 U35760 ( .B1(n3447), .B2(n4747), .A(n2985), .ZN(U3244) );
  XNOR2_X1 U35770 ( .A(n2988), .B(n3960), .ZN(n2992) );
  NAND2_X1 U35780 ( .A1(n4768), .A2(n3298), .ZN(n2990) );
  AOI22_X1 U35790 ( .A1(n4055), .A2(n4320), .B1(n3702), .B2(n4800), .ZN(n2989)
         );
  OAI211_X1 U35800 ( .C1(n2425), .C2(n4324), .A(n2990), .B(n2989), .ZN(n2991)
         );
  AOI21_X1 U35810 ( .B1(n2992), .B2(n4807), .A(n2991), .ZN(n4771) );
  INV_X1 U3582 ( .A(n4771), .ZN(n2993) );
  AOI21_X1 U3583 ( .B1(n4781), .B2(n4768), .A(n2993), .ZN(n2996) );
  AOI21_X1 U3584 ( .B1(n3702), .B2(n3048), .A(n3009), .ZN(n4767) );
  INV_X1 U3585 ( .A(n4383), .ZN(n3169) );
  AOI22_X1 U3586 ( .A1(n4767), .A2(n3169), .B1(REG1_REG_2__SCAN_IN), .B2(n2856), .ZN(n2994) );
  OAI21_X1 U3587 ( .B1(n2996), .B2(n2856), .A(n2994), .ZN(U3520) );
  INV_X1 U3588 ( .A(n4423), .ZN(n3167) );
  AOI22_X1 U3589 ( .A1(n4767), .A2(n3167), .B1(REG0_REG_2__SCAN_IN), .B2(n4832), .ZN(n2995) );
  OAI21_X1 U3590 ( .B1(n2996), .B2(n4832), .A(n2995), .ZN(U3471) );
  XNOR2_X1 U3591 ( .A(n2998), .B(n2997), .ZN(n4774) );
  OAI21_X1 U3592 ( .B1(n3958), .B2(n3000), .A(n2999), .ZN(n3001) );
  NAND2_X1 U3593 ( .A1(n3001), .A2(n4807), .ZN(n3004) );
  AOI22_X1 U3594 ( .A1(n4054), .A2(n4320), .B1(n4800), .B2(n3002), .ZN(n3003)
         );
  OAI211_X1 U3595 ( .C1(n3005), .C2(n4324), .A(n3004), .B(n3003), .ZN(n3006)
         );
  AOI21_X1 U3596 ( .B1(n3298), .B2(n4774), .A(n3006), .ZN(n4777) );
  INV_X1 U3597 ( .A(n4777), .ZN(n3007) );
  AOI21_X1 U3598 ( .B1(n4781), .B2(n4774), .A(n3007), .ZN(n3013) );
  NOR2_X1 U3599 ( .A1(n3009), .A2(n3008), .ZN(n3010) );
  NOR2_X1 U3600 ( .A1(n3010), .A2(n3069), .ZN(n4773) );
  AOI22_X1 U3601 ( .A1(n4773), .A2(n3169), .B1(REG1_REG_3__SCAN_IN), .B2(n2856), .ZN(n3011) );
  OAI21_X1 U3602 ( .B1(n3013), .B2(n2856), .A(n3011), .ZN(U3521) );
  AOI22_X1 U3603 ( .A1(n4773), .A2(n3167), .B1(REG0_REG_3__SCAN_IN), .B2(n4832), .ZN(n3012) );
  OAI21_X1 U3604 ( .B1(n3013), .B2(n4832), .A(n3012), .ZN(U3473) );
  XNOR2_X1 U3605 ( .A(n3014), .B(n3720), .ZN(n3104) );
  NOR2_X1 U3606 ( .A1(n3068), .A2(n4037), .ZN(n3015) );
  AOI21_X1 U3607 ( .B1(n4054), .B2(n3674), .A(n3015), .ZN(n3103) );
  XNOR2_X1 U3608 ( .A(n3104), .B(n3103), .ZN(n3021) );
  NOR2_X1 U3609 ( .A1(n3017), .A2(n3016), .ZN(n3019) );
  OR2_X1 U3610 ( .A1(n3018), .A2(n3019), .ZN(n3020) );
  AOI211_X1 U3611 ( .C1(n3021), .C2(n3020), .A(n3871), .B(n3105), .ZN(n3027)
         );
  INV_X1 U3612 ( .A(n3080), .ZN(n3025) );
  AOI22_X1 U3613 ( .A1(n3074), .A2(n4879), .B1(n4053), .B2(n3840), .ZN(n3024)
         );
  AOI21_X1 U3614 ( .B1(n4875), .B2(n4055), .A(n3022), .ZN(n3023) );
  OAI211_X1 U3615 ( .C1(n4891), .C2(n3025), .A(n3024), .B(n3023), .ZN(n3026)
         );
  OR2_X1 U3616 ( .A1(n3027), .A2(n3026), .ZN(U3227) );
  OAI21_X1 U3617 ( .B1(n3030), .B2(n3029), .A(n3028), .ZN(n4761) );
  OAI21_X1 U3618 ( .B1(n3959), .B2(n3894), .A(n3031), .ZN(n3036) );
  NAND2_X1 U3619 ( .A1(n2912), .A2(n4801), .ZN(n3033) );
  NAND2_X1 U3620 ( .A1(n4056), .A2(n4320), .ZN(n3032) );
  OAI211_X1 U3621 ( .C1(n4282), .C2(n3034), .A(n3033), .B(n3032), .ZN(n3035)
         );
  AOI21_X1 U3622 ( .B1(n3036), .B2(n4807), .A(n3035), .ZN(n3037) );
  OAI21_X1 U3623 ( .B1(n3557), .B2(n4761), .A(n3037), .ZN(n4763) );
  INV_X1 U3624 ( .A(n4763), .ZN(n3054) );
  INV_X1 U3625 ( .A(n3038), .ZN(n3040) );
  NAND4_X1 U3626 ( .A1(n3042), .A2(n3041), .A3(n3040), .A4(n3039), .ZN(n3043)
         );
  INV_X1 U3627 ( .A(n4761), .ZN(n3052) );
  OR2_X1 U3628 ( .A1(n3044), .A2(n4814), .ZN(n3094) );
  INV_X1 U3629 ( .A(n3094), .ZN(n3045) );
  INV_X2 U3630 ( .A(n4900), .ZN(n4333) );
  AND2_X1 U3631 ( .A1(n4811), .A2(n4814), .ZN(n3046) );
  NAND2_X1 U3632 ( .A1(n3089), .A2(n3047), .ZN(n3049) );
  NAND2_X1 U3633 ( .A1(n3049), .A2(n3048), .ZN(n4758) );
  AOI22_X1 U3634 ( .A1(n4900), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4847), .ZN(n3050) );
  OAI21_X1 U3635 ( .B1(n4859), .B2(n4758), .A(n3050), .ZN(n3051) );
  AOI21_X1 U3636 ( .B1(n3052), .B2(n4851), .A(n3051), .ZN(n3053) );
  OAI21_X1 U3637 ( .B1(n3054), .B2(n4900), .A(n3053), .ZN(U3289) );
  NAND2_X1 U3638 ( .A1(n3055), .A2(n3056), .ZN(n3058) );
  INV_X1 U3639 ( .A(n3057), .ZN(n3904) );
  AND2_X1 U3640 ( .A1(n3904), .A2(n3881), .ZN(n3977) );
  XNOR2_X1 U3641 ( .A(n3058), .B(n3977), .ZN(n3093) );
  XNOR2_X1 U3642 ( .A(n3059), .B(n3977), .ZN(n3062) );
  AOI22_X1 U3643 ( .A1(n4054), .A2(n4801), .B1(n3118), .B2(n4800), .ZN(n3061)
         );
  NAND2_X1 U3644 ( .A1(n4802), .A2(n4320), .ZN(n3060) );
  OAI211_X1 U3645 ( .C1(n3062), .C2(n4300), .A(n3061), .B(n3060), .ZN(n3095)
         );
  AOI21_X1 U3646 ( .B1(n3093), .B2(n4826), .A(n3095), .ZN(n3066) );
  INV_X1 U3647 ( .A(n3147), .ZN(n3063) );
  AOI21_X1 U3648 ( .B1(n3118), .B2(n3067), .A(n3063), .ZN(n3099) );
  AOI22_X1 U3649 ( .A1(n3099), .A2(n3169), .B1(REG1_REG_5__SCAN_IN), .B2(n2856), .ZN(n3064) );
  OAI21_X1 U3650 ( .B1(n3066), .B2(n2856), .A(n3064), .ZN(U3523) );
  AOI22_X1 U3651 ( .A1(n3099), .A2(n3167), .B1(REG0_REG_5__SCAN_IN), .B2(n4832), .ZN(n3065) );
  OAI21_X1 U3652 ( .B1(n3066), .B2(n4832), .A(n3065), .ZN(U3477) );
  OAI211_X1 U3653 ( .C1(n3069), .C2(n3068), .A(n4811), .B(n3067), .ZN(n4778)
         );
  NOR2_X1 U3654 ( .A1(n4778), .A2(n4168), .ZN(n3079) );
  XNOR2_X1 U3655 ( .A(n3070), .B(n3071), .ZN(n3078) );
  INV_X1 U3656 ( .A(n3071), .ZN(n3978) );
  NAND2_X1 U3657 ( .A1(n3072), .A2(n3978), .ZN(n3073) );
  AND2_X1 U3658 ( .A1(n3055), .A2(n3073), .ZN(n4782) );
  AOI22_X1 U3659 ( .A1(n4055), .A2(n4801), .B1(n3074), .B2(n4800), .ZN(n3075)
         );
  OAI21_X1 U3660 ( .B1(n3144), .B2(n4804), .A(n3075), .ZN(n3076) );
  AOI21_X1 U3661 ( .B1(n4782), .B2(n3298), .A(n3076), .ZN(n3077) );
  OAI21_X1 U3662 ( .B1(n4300), .B2(n3078), .A(n3077), .ZN(n4779) );
  AOI211_X1 U3663 ( .C1(n4847), .C2(n3080), .A(n3079), .B(n4779), .ZN(n3082)
         );
  AOI22_X1 U3664 ( .A1(n4782), .A2(n4851), .B1(REG2_REG_4__SCAN_IN), .B2(n4900), .ZN(n3081) );
  OAI21_X1 U3665 ( .B1(n3082), .B2(n4900), .A(n3081), .ZN(U3286) );
  XNOR2_X1 U3666 ( .A(n3083), .B(n3084), .ZN(n3092) );
  AOI22_X1 U3667 ( .A1(n4875), .A2(n2912), .B1(n4877), .B2(n4056), .ZN(n3091)
         );
  INV_X1 U3668 ( .A(n3085), .ZN(n3088) );
  NAND3_X1 U3669 ( .A1(n3088), .A2(n3087), .A3(n3086), .ZN(n3703) );
  AOI22_X1 U3670 ( .A1(REG3_REG_1__SCAN_IN), .A2(n3703), .B1(n4879), .B2(n3089), .ZN(n3090) );
  OAI211_X1 U3671 ( .C1(n3092), .C2(n3871), .A(n3091), .B(n3090), .ZN(U3219)
         );
  INV_X1 U3672 ( .A(n3093), .ZN(n3102) );
  NAND2_X1 U3673 ( .A1(n3557), .A2(n3094), .ZN(n4819) );
  NAND2_X1 U3674 ( .A1(n3095), .A2(n4333), .ZN(n3101) );
  NOR2_X1 U3675 ( .A1(n3121), .A2(n4863), .ZN(n3098) );
  INV_X1 U3676 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3096) );
  NOR2_X1 U3677 ( .A1(n4333), .A2(n3096), .ZN(n3097) );
  AOI211_X1 U3678 ( .C1(n3099), .C2(n4896), .A(n3098), .B(n3097), .ZN(n3100)
         );
  OAI211_X1 U3679 ( .C1(n3102), .C2(n4335), .A(n3101), .B(n3100), .ZN(U3285)
         );
  INV_X1 U3680 ( .A(n3103), .ZN(n3107) );
  INV_X1 U3681 ( .A(n3104), .ZN(n3106) );
  INV_X1 U3682 ( .A(n3718), .ZN(n3662) );
  OAI22_X1 U3683 ( .A1(n3144), .A2(n4037), .B1(n3662), .B2(n3108), .ZN(n3109)
         );
  XNOR2_X1 U3684 ( .A(n3109), .B(n3671), .ZN(n3115) );
  INV_X1 U3685 ( .A(n3115), .ZN(n3113) );
  OR2_X1 U3686 ( .A1(n3144), .A2(n3664), .ZN(n3111) );
  NAND2_X1 U3687 ( .A1(n3118), .A2(n3719), .ZN(n3110) );
  AND2_X1 U3688 ( .A1(n3111), .A2(n3110), .ZN(n3114) );
  INV_X1 U3689 ( .A(n3114), .ZN(n3112) );
  NAND2_X1 U3690 ( .A1(n3113), .A2(n3112), .ZN(n3125) );
  INV_X1 U3691 ( .A(n3125), .ZN(n3116) );
  AND2_X1 U3692 ( .A1(n3115), .A2(n3114), .ZN(n3127) );
  NOR2_X1 U3693 ( .A1(n3116), .A2(n3127), .ZN(n3117) );
  XNOR2_X1 U3694 ( .A(n3126), .B(n3117), .ZN(n3123) );
  INV_X1 U3695 ( .A(n3760), .ZN(n3818) );
  AOI22_X1 U3696 ( .A1(n4879), .A2(n3118), .B1(n3818), .B2(n4054), .ZN(n3120)
         );
  NOR2_X1 U3697 ( .A1(STATE_REG_SCAN_IN), .A2(n2527), .ZN(n4633) );
  AOI21_X1 U3698 ( .B1(n4877), .B2(n4802), .A(n4633), .ZN(n3119) );
  OAI211_X1 U3699 ( .C1(n4891), .C2(n3121), .A(n3120), .B(n3119), .ZN(n3122)
         );
  AOI21_X1 U3700 ( .B1(n3123), .B2(n4886), .A(n3122), .ZN(n3124) );
  INV_X1 U3701 ( .A(n3124), .ZN(U3224) );
  NAND2_X1 U3702 ( .A1(n3126), .A2(n3125), .ZN(n3129) );
  NAND2_X1 U3703 ( .A1(n3129), .A2(n3128), .ZN(n3191) );
  INV_X1 U3704 ( .A(n3191), .ZN(n3194) );
  AOI22_X1 U3705 ( .A1(n4802), .A2(n3719), .B1(n3718), .B2(n3148), .ZN(n3130)
         );
  XNOR2_X1 U3706 ( .A(n3130), .B(n3720), .ZN(n3189) );
  XNOR2_X1 U3707 ( .A(n3189), .B(n3190), .ZN(n3131) );
  XNOR2_X1 U3708 ( .A(n3194), .B(n3131), .ZN(n3137) );
  INV_X1 U3709 ( .A(n4788), .ZN(n3135) );
  AOI22_X1 U3710 ( .A1(n3148), .A2(n4879), .B1(n4053), .B2(n4875), .ZN(n3134)
         );
  NOR2_X1 U3711 ( .A1(STATE_REG_SCAN_IN), .A2(n3132), .ZN(n4643) );
  AOI21_X1 U3712 ( .B1(n4877), .B2(n4052), .A(n4643), .ZN(n3133) );
  OAI211_X1 U3713 ( .C1(n4891), .C2(n3135), .A(n3134), .B(n3133), .ZN(n3136)
         );
  AOI21_X1 U3714 ( .B1(n3137), .B2(n4886), .A(n3136), .ZN(n3138) );
  INV_X1 U3715 ( .A(n3138), .ZN(U3236) );
  INV_X1 U3716 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3151) );
  AND2_X1 U3717 ( .A1(n4796), .A2(n3905), .ZN(n3954) );
  XNOR2_X1 U3718 ( .A(n3139), .B(n3954), .ZN(n4790) );
  INV_X1 U3719 ( .A(n4790), .ZN(n3146) );
  XNOR2_X1 U3720 ( .A(n3140), .B(n3954), .ZN(n3141) );
  NAND2_X1 U3721 ( .A1(n3141), .A2(n4807), .ZN(n3143) );
  AOI22_X1 U3722 ( .A1(n4052), .A2(n4320), .B1(n3148), .B2(n4800), .ZN(n3142)
         );
  OAI211_X1 U3723 ( .C1(n3144), .C2(n4324), .A(n3143), .B(n3142), .ZN(n3145)
         );
  AOI21_X1 U3724 ( .B1(n3298), .B2(n4790), .A(n3145), .ZN(n4793) );
  OAI21_X1 U3725 ( .B1(n4760), .B2(n3146), .A(n4793), .ZN(n3152) );
  NAND2_X1 U3726 ( .A1(n3152), .A2(n4835), .ZN(n3150) );
  AOI21_X1 U3727 ( .B1(n3148), .B2(n3147), .A(n4810), .ZN(n4789) );
  NAND2_X1 U3728 ( .A1(n4789), .A2(n3167), .ZN(n3149) );
  OAI211_X1 U3729 ( .C1(n4835), .C2(n3151), .A(n3150), .B(n3149), .ZN(U3479)
         );
  INV_X1 U3730 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U3731 ( .A1(n3152), .A2(n4831), .ZN(n3154) );
  NAND2_X1 U3732 ( .A1(n4789), .A2(n3169), .ZN(n3153) );
  OAI211_X1 U3733 ( .C1(n4831), .C2(n3155), .A(n3154), .B(n3153), .ZN(U3524)
         );
  INV_X1 U3734 ( .A(n3911), .ZN(n3879) );
  AND2_X1 U3735 ( .A1(n3879), .A2(n3913), .ZN(n3961) );
  XNOR2_X1 U3736 ( .A(n3156), .B(n3961), .ZN(n3166) );
  INV_X1 U3737 ( .A(n3166), .ZN(n3164) );
  AOI21_X1 U3738 ( .B1(n3230), .B2(n3181), .A(n3238), .ZN(n3170) );
  INV_X1 U3739 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3424) );
  OAI22_X1 U3740 ( .A1(n3233), .A2(n4863), .B1(n3424), .B2(n4333), .ZN(n3157)
         );
  AOI21_X1 U3741 ( .B1(n3170), .B2(n4896), .A(n3157), .ZN(n3163) );
  XNOR2_X1 U3742 ( .A(n3158), .B(n3961), .ZN(n3161) );
  OAI22_X1 U3743 ( .A1(n4805), .A2(n4324), .B1(n4282), .B2(n3220), .ZN(n3159)
         );
  AOI21_X1 U3744 ( .B1(n4320), .B2(n4049), .A(n3159), .ZN(n3160) );
  OAI21_X1 U3745 ( .B1(n3161), .B2(n4300), .A(n3160), .ZN(n3165) );
  NAND2_X1 U3746 ( .A1(n3165), .A2(n4333), .ZN(n3162) );
  OAI211_X1 U3747 ( .C1(n3164), .C2(n4335), .A(n3163), .B(n3162), .ZN(U3281)
         );
  AOI21_X1 U3748 ( .B1(n3166), .B2(n4826), .A(n3165), .ZN(n3172) );
  AOI22_X1 U3749 ( .A1(n3170), .A2(n3167), .B1(REG0_REG_9__SCAN_IN), .B2(n4832), .ZN(n3168) );
  OAI21_X1 U3750 ( .B1(n3172), .B2(n4832), .A(n3168), .ZN(U3485) );
  AOI22_X1 U3751 ( .A1(n3170), .A2(n3169), .B1(REG1_REG_9__SCAN_IN), .B2(n2856), .ZN(n3171) );
  OAI21_X1 U3752 ( .B1(n3172), .B2(n2856), .A(n3171), .ZN(U3527) );
  AND2_X1 U3753 ( .A1(n3912), .A2(n3878), .ZN(n3975) );
  XNOR2_X1 U3754 ( .A(n3173), .B(n3975), .ZN(n4841) );
  INV_X1 U3755 ( .A(n4841), .ZN(n3179) );
  XNOR2_X1 U3756 ( .A(n3174), .B(n3975), .ZN(n3177) );
  OAI22_X1 U3757 ( .A1(n3221), .A2(n4804), .B1(n3204), .B2(n4282), .ZN(n3175)
         );
  AOI21_X1 U3758 ( .B1(n4801), .B2(n4052), .A(n3175), .ZN(n3176) );
  OAI21_X1 U3759 ( .B1(n3177), .B2(n4300), .A(n3176), .ZN(n3178) );
  AOI21_X1 U3760 ( .B1(n3298), .B2(n4841), .A(n3178), .ZN(n4844) );
  OAI21_X1 U3761 ( .B1(n4760), .B2(n3179), .A(n4844), .ZN(n3186) );
  NAND2_X1 U3762 ( .A1(n4813), .A2(n3212), .ZN(n3180) );
  NAND2_X1 U3763 ( .A1(n3181), .A2(n3180), .ZN(n4839) );
  INV_X1 U3764 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4664) );
  OAI22_X1 U3765 ( .A1(n4839), .A2(n4383), .B1(n4831), .B2(n4664), .ZN(n3182)
         );
  AOI21_X1 U3766 ( .B1(n3186), .B2(n4831), .A(n3182), .ZN(n3183) );
  INV_X1 U3767 ( .A(n3183), .ZN(U3526) );
  INV_X1 U3768 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3184) );
  OAI22_X1 U3769 ( .A1(n4839), .A2(n4423), .B1(n4835), .B2(n3184), .ZN(n3185)
         );
  AOI21_X1 U3770 ( .B1(n3186), .B2(n4835), .A(n3185), .ZN(n3187) );
  INV_X1 U3771 ( .A(n3187), .ZN(U3483) );
  AOI22_X1 U3772 ( .A1(n4052), .A2(n3719), .B1(n3718), .B2(n4799), .ZN(n3188)
         );
  XNOR2_X1 U3773 ( .A(n3188), .B(n3720), .ZN(n3200) );
  AOI22_X1 U3774 ( .A1(n4052), .A2(n2933), .B1(n3719), .B2(n4799), .ZN(n3201)
         );
  XNOR2_X1 U3775 ( .A(n3200), .B(n3201), .ZN(n3202) );
  INV_X1 U3776 ( .A(n3190), .ZN(n3193) );
  AOI21_X1 U3777 ( .B1(n3191), .B2(n3190), .A(n3189), .ZN(n3192) );
  AOI21_X2 U3778 ( .B1(n3194), .B2(n3193), .A(n3192), .ZN(n3203) );
  XOR2_X1 U3779 ( .A(n3202), .B(n3203), .Z(n3198) );
  AOI22_X1 U3780 ( .A1(n4879), .A2(n4799), .B1(n3818), .B2(n4802), .ZN(n3196)
         );
  NOR2_X1 U3781 ( .A1(STATE_REG_SCAN_IN), .A2(n2549), .ZN(n4654) );
  AOI21_X1 U3782 ( .B1(n4051), .B2(n3840), .A(n4654), .ZN(n3195) );
  OAI211_X1 U3783 ( .C1(n4891), .C2(n4824), .A(n3196), .B(n3195), .ZN(n3197)
         );
  AOI21_X1 U3784 ( .B1(n3198), .B2(n4886), .A(n3197), .ZN(n3199) );
  INV_X1 U3785 ( .A(n3199), .ZN(U3210) );
  OAI22_X1 U3786 ( .A1(n4805), .A2(n4037), .B1(n3662), .B2(n3204), .ZN(n3205)
         );
  XNOR2_X1 U3787 ( .A(n3205), .B(n3671), .ZN(n3209) );
  OR2_X1 U3788 ( .A1(n4805), .A2(n3664), .ZN(n3207) );
  NAND2_X1 U3789 ( .A1(n3212), .A2(n3719), .ZN(n3206) );
  AND2_X1 U3790 ( .A1(n3207), .A2(n3206), .ZN(n3208) );
  NOR2_X1 U3791 ( .A1(n3209), .A2(n3208), .ZN(n3226) );
  INV_X1 U3792 ( .A(n3226), .ZN(n3210) );
  NAND2_X1 U3793 ( .A1(n3209), .A2(n3208), .ZN(n3225) );
  NAND2_X1 U3794 ( .A1(n3210), .A2(n3225), .ZN(n3211) );
  XNOR2_X1 U3795 ( .A(n3227), .B(n3211), .ZN(n3218) );
  INV_X1 U3796 ( .A(n4838), .ZN(n3216) );
  AOI22_X1 U3797 ( .A1(n4879), .A2(n3212), .B1(n3818), .B2(n4052), .ZN(n3215)
         );
  INV_X1 U3798 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3213) );
  NOR2_X1 U3799 ( .A1(STATE_REG_SCAN_IN), .A2(n3213), .ZN(n4665) );
  AOI21_X1 U3800 ( .B1(n4877), .B2(n4050), .A(n4665), .ZN(n3214) );
  OAI211_X1 U3801 ( .C1(n4891), .C2(n3216), .A(n3215), .B(n3214), .ZN(n3217)
         );
  AOI21_X1 U3802 ( .B1(n3218), .B2(n4886), .A(n3217), .ZN(n3219) );
  INV_X1 U3803 ( .A(n3219), .ZN(U3218) );
  OAI22_X1 U3804 ( .A1(n3221), .A2(n3664), .B1(n4037), .B2(n3220), .ZN(n3270)
         );
  NAND2_X1 U3805 ( .A1(n4050), .A2(n3719), .ZN(n3223) );
  NAND2_X1 U3806 ( .A1(n3230), .A2(n3718), .ZN(n3222) );
  NAND2_X1 U3807 ( .A1(n3223), .A2(n3222), .ZN(n3224) );
  XNOR2_X1 U3808 ( .A(n3224), .B(n3720), .ZN(n3269) );
  XOR2_X1 U3809 ( .A(n3270), .B(n3269), .Z(n3229) );
  NAND2_X1 U3810 ( .A1(n3228), .A2(n3229), .ZN(n3274) );
  OAI21_X1 U3811 ( .B1(n3229), .B2(n3228), .A(n3274), .ZN(n3235) );
  AOI22_X1 U3812 ( .A1(n3230), .A2(n4879), .B1(n4051), .B2(n4875), .ZN(n3232)
         );
  NOR2_X1 U3813 ( .A1(STATE_REG_SCAN_IN), .A2(n2570), .ZN(n4675) );
  AOI21_X1 U3814 ( .B1(n4877), .B2(n4049), .A(n4675), .ZN(n3231) );
  OAI211_X1 U3815 ( .C1(n4891), .C2(n3233), .A(n3232), .B(n3231), .ZN(n3234)
         );
  AOI21_X1 U3816 ( .B1(n3235), .B2(n4886), .A(n3234), .ZN(n3236) );
  INV_X1 U3817 ( .A(n3236), .ZN(U3228) );
  INV_X1 U3818 ( .A(n3294), .ZN(n3237) );
  OAI21_X1 U3819 ( .B1(n3238), .B2(n3244), .A(n3237), .ZN(n4849) );
  NAND2_X1 U3820 ( .A1(n3885), .A2(n3882), .ZN(n3973) );
  XNOR2_X1 U3821 ( .A(n3239), .B(n3973), .ZN(n4852) );
  NAND2_X1 U3822 ( .A1(n4852), .A2(n3298), .ZN(n3248) );
  INV_X1 U3823 ( .A(n3973), .ZN(n3240) );
  XNOR2_X1 U3824 ( .A(n3241), .B(n3240), .ZN(n3246) );
  NAND2_X1 U3825 ( .A1(n4050), .A2(n4801), .ZN(n3243) );
  NAND2_X1 U3826 ( .A1(n4048), .A2(n4320), .ZN(n3242) );
  OAI211_X1 U3827 ( .C1(n4282), .C2(n3244), .A(n3243), .B(n3242), .ZN(n3245)
         );
  AOI21_X1 U3828 ( .B1(n3246), .B2(n4807), .A(n3245), .ZN(n3247) );
  AND2_X1 U3829 ( .A1(n3248), .A2(n3247), .ZN(n4855) );
  NAND2_X1 U3830 ( .A1(n4852), .A2(n4781), .ZN(n3249) );
  AND2_X1 U3831 ( .A1(n4855), .A2(n3249), .ZN(n3252) );
  INV_X1 U3832 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3250) );
  MUX2_X1 U3833 ( .A(n3252), .B(n3250), .S(n4832), .Z(n3251) );
  OAI21_X1 U3834 ( .B1(n4849), .B2(n4423), .A(n3251), .ZN(U3487) );
  INV_X1 U3835 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3253) );
  MUX2_X1 U3836 ( .A(n3253), .B(n3252), .S(n4831), .Z(n3254) );
  OAI21_X1 U3837 ( .B1(n4849), .B2(n4383), .A(n3254), .ZN(U3528) );
  NAND2_X1 U3838 ( .A1(n3347), .A2(n3345), .ZN(n3944) );
  XNOR2_X1 U3839 ( .A(n3255), .B(n3944), .ZN(n3314) );
  INV_X1 U3840 ( .A(n3314), .ZN(n3267) );
  INV_X1 U3841 ( .A(n3256), .ZN(n3257) );
  AOI21_X1 U3842 ( .B1(n3299), .B2(n3258), .A(n3257), .ZN(n3348) );
  XOR2_X1 U3843 ( .A(n3944), .B(n3348), .Z(n3261) );
  AOI22_X1 U3844 ( .A1(n4048), .A2(n4801), .B1(n3324), .B2(n4800), .ZN(n3260)
         );
  NAND2_X1 U3845 ( .A1(n4046), .A2(n4320), .ZN(n3259) );
  OAI211_X1 U3846 ( .C1(n3261), .C2(n4300), .A(n3260), .B(n3259), .ZN(n3313)
         );
  NAND2_X1 U3847 ( .A1(n3293), .A2(n3324), .ZN(n3262) );
  NAND2_X1 U3848 ( .A1(n3355), .A2(n3262), .ZN(n3319) );
  AOI22_X1 U3849 ( .A1(n4900), .A2(REG2_REG_12__SCAN_IN), .B1(n3263), .B2(
        n4847), .ZN(n3264) );
  OAI21_X1 U3850 ( .B1(n3319), .B2(n4859), .A(n3264), .ZN(n3265) );
  AOI21_X1 U3851 ( .B1(n3313), .B2(n4333), .A(n3265), .ZN(n3266) );
  OAI21_X1 U3852 ( .B1(n3267), .B2(n4335), .A(n3266), .ZN(U3278) );
  AOI22_X1 U3853 ( .A1(n4049), .A2(n2933), .B1(n3719), .B2(n3747), .ZN(n3276)
         );
  AOI22_X1 U3854 ( .A1(n4049), .A2(n3719), .B1(n3718), .B2(n3747), .ZN(n3268)
         );
  XNOR2_X1 U3855 ( .A(n3268), .B(n3720), .ZN(n3275) );
  XOR2_X1 U3856 ( .A(n3276), .B(n3275), .Z(n3745) );
  INV_X1 U3857 ( .A(n3269), .ZN(n3272) );
  INV_X1 U3858 ( .A(n3270), .ZN(n3271) );
  NAND2_X1 U3859 ( .A1(n3272), .A2(n3271), .ZN(n3743) );
  NAND2_X1 U3860 ( .A1(n3274), .A2(n3273), .ZN(n3744) );
  NAND2_X1 U3861 ( .A1(n3744), .A2(n3279), .ZN(n3320) );
  NAND2_X1 U3862 ( .A1(n4048), .A2(n3719), .ZN(n3281) );
  INV_X1 U3863 ( .A(n3302), .ZN(n3287) );
  NAND2_X1 U3864 ( .A1(n3287), .A2(n3718), .ZN(n3280) );
  NAND2_X1 U3865 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  XNOR2_X1 U3866 ( .A(n3282), .B(n3671), .ZN(n3285) );
  NOR2_X1 U3867 ( .A1(n3302), .A2(n4037), .ZN(n3283) );
  AOI21_X1 U3868 ( .B1(n4048), .B2(n2933), .A(n3283), .ZN(n3284) );
  OR2_X1 U3869 ( .A1(n3285), .A2(n3284), .ZN(n3321) );
  NAND2_X1 U3870 ( .A1(n2291), .A2(n3321), .ZN(n3286) );
  XNOR2_X1 U3871 ( .A(n3320), .B(n3286), .ZN(n3291) );
  AOI22_X1 U3872 ( .A1(n4879), .A2(n3287), .B1(n4875), .B2(n4049), .ZN(n3289)
         );
  AND2_X1 U3873 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4697) );
  AOI21_X1 U3874 ( .B1(n4877), .B2(n4047), .A(n4697), .ZN(n3288) );
  OAI211_X1 U3875 ( .C1(n4891), .C2(n4864), .A(n3289), .B(n3288), .ZN(n3290)
         );
  AOI21_X1 U3876 ( .B1(n3291), .B2(n4886), .A(n3290), .ZN(n3292) );
  INV_X1 U3877 ( .A(n3292), .ZN(U3233) );
  OAI21_X1 U3878 ( .B1(n3294), .B2(n3302), .A(n3293), .ZN(n4858) );
  NAND2_X1 U3879 ( .A1(n3295), .A2(n3980), .ZN(n3296) );
  NAND2_X1 U3880 ( .A1(n3297), .A2(n3296), .ZN(n4857) );
  NAND2_X1 U3881 ( .A1(n4857), .A2(n3298), .ZN(n3306) );
  XNOR2_X1 U3882 ( .A(n3299), .B(n3980), .ZN(n3304) );
  NAND2_X1 U3883 ( .A1(n4049), .A2(n4801), .ZN(n3301) );
  NAND2_X1 U3884 ( .A1(n4047), .A2(n4320), .ZN(n3300) );
  OAI211_X1 U3885 ( .C1(n4282), .C2(n3302), .A(n3301), .B(n3300), .ZN(n3303)
         );
  AOI21_X1 U3886 ( .B1(n3304), .B2(n4807), .A(n3303), .ZN(n3305) );
  NAND2_X1 U3887 ( .A1(n4857), .A2(n4781), .ZN(n3307) );
  NAND2_X1 U3888 ( .A1(n4868), .A2(n3307), .ZN(n3310) );
  MUX2_X1 U3889 ( .A(REG0_REG_11__SCAN_IN), .B(n3310), .S(n4835), .Z(n3308) );
  INV_X1 U3890 ( .A(n3308), .ZN(n3309) );
  OAI21_X1 U3891 ( .B1(n4858), .B2(n4423), .A(n3309), .ZN(U3489) );
  MUX2_X1 U3892 ( .A(REG1_REG_11__SCAN_IN), .B(n3310), .S(n4831), .Z(n3311) );
  INV_X1 U3893 ( .A(n3311), .ZN(n3312) );
  OAI21_X1 U3894 ( .B1(n4383), .B2(n4858), .A(n3312), .ZN(U3529) );
  INV_X1 U3895 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4706) );
  AOI21_X1 U3896 ( .B1(n4826), .B2(n3314), .A(n3313), .ZN(n3316) );
  MUX2_X1 U3897 ( .A(n4706), .B(n3316), .S(n4831), .Z(n3315) );
  OAI21_X1 U3898 ( .B1(n3319), .B2(n4383), .A(n3315), .ZN(U3530) );
  INV_X1 U3899 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3317) );
  MUX2_X1 U3900 ( .A(n3317), .B(n3316), .S(n4835), .Z(n3318) );
  OAI21_X1 U3901 ( .B1(n3319), .B2(n4423), .A(n3318), .ZN(U3491) );
  OAI22_X1 U3902 ( .A1(n3351), .A2(n4037), .B1(n3662), .B2(n2301), .ZN(n3322)
         );
  XNOR2_X1 U3903 ( .A(n3322), .B(n3720), .ZN(n3475) );
  AOI22_X1 U3904 ( .A1(n4047), .A2(n2933), .B1(n3719), .B2(n3324), .ZN(n3471)
         );
  INV_X1 U3905 ( .A(n3471), .ZN(n3472) );
  XNOR2_X1 U3906 ( .A(n3475), .B(n3472), .ZN(n3323) );
  XNOR2_X1 U3907 ( .A(n3473), .B(n3323), .ZN(n3329) );
  AOI22_X1 U3908 ( .A1(n4879), .A2(n3324), .B1(n4877), .B2(n4046), .ZN(n3326)
         );
  INV_X1 U3909 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4490) );
  NOR2_X1 U3910 ( .A1(STATE_REG_SCAN_IN), .A2(n4490), .ZN(n4707) );
  AOI21_X1 U3911 ( .B1(n4875), .B2(n4048), .A(n4707), .ZN(n3325) );
  OAI211_X1 U3912 ( .C1(n4891), .C2(n3327), .A(n3326), .B(n3325), .ZN(n3328)
         );
  AOI21_X1 U3913 ( .B1(n3329), .B2(n4886), .A(n3328), .ZN(n3330) );
  INV_X1 U3914 ( .A(n3330), .ZN(U3221) );
  AND2_X1 U3915 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  NAND2_X1 U3916 ( .A1(n3333), .A2(n3945), .ZN(n3380) );
  OAI21_X1 U3917 ( .B1(n3333), .B2(n3945), .A(n3380), .ZN(n3405) );
  INV_X1 U3918 ( .A(n3405), .ZN(n3343) );
  INV_X1 U3919 ( .A(n4045), .ZN(n3338) );
  OAI21_X1 U3920 ( .B1(n3334), .B2(n4001), .A(n3382), .ZN(n3335) );
  NAND2_X1 U3921 ( .A1(n3335), .A2(n4807), .ZN(n3337) );
  AOI22_X1 U3922 ( .A1(n4046), .A2(n4801), .B1(n4800), .B2(n3505), .ZN(n3336)
         );
  OAI211_X1 U3923 ( .C1(n3338), .C2(n4804), .A(n3337), .B(n3336), .ZN(n3404)
         );
  NOR2_X1 U3924 ( .A1(n3356), .A2(n3501), .ZN(n3339) );
  OR2_X1 U3925 ( .A1(n3389), .A2(n3339), .ZN(n3411) );
  AOI22_X1 U3926 ( .A1(n4900), .A2(REG2_REG_14__SCAN_IN), .B1(n3504), .B2(
        n4847), .ZN(n3340) );
  OAI21_X1 U3927 ( .B1(n3411), .B2(n4859), .A(n3340), .ZN(n3341) );
  AOI21_X1 U3928 ( .B1(n3404), .B2(n4333), .A(n3341), .ZN(n3342) );
  OAI21_X1 U3929 ( .B1(n3343), .B2(n4335), .A(n3342), .ZN(U3276) );
  XNOR2_X1 U3930 ( .A(n4046), .B(n3358), .ZN(n3983) );
  XOR2_X1 U3931 ( .A(n3983), .B(n3344), .Z(n3395) );
  INV_X1 U3932 ( .A(n4851), .ZN(n4860) );
  INV_X1 U3933 ( .A(n3345), .ZN(n3346) );
  AOI21_X1 U3934 ( .B1(n3348), .B2(n3347), .A(n3346), .ZN(n3349) );
  XOR2_X1 U3935 ( .A(n3983), .B(n3349), .Z(n3353) );
  AOI22_X1 U3936 ( .A1(n4874), .A2(n4320), .B1(n3483), .B2(n4800), .ZN(n3350)
         );
  OAI21_X1 U3937 ( .B1(n3351), .B2(n4324), .A(n3350), .ZN(n3352) );
  AOI21_X1 U3938 ( .B1(n3353), .B2(n4807), .A(n3352), .ZN(n3354) );
  OAI21_X1 U3939 ( .B1(n3395), .B2(n3557), .A(n3354), .ZN(n3396) );
  NAND2_X1 U3940 ( .A1(n3396), .A2(n4333), .ZN(n3364) );
  INV_X1 U3941 ( .A(n3355), .ZN(n3359) );
  INV_X1 U3942 ( .A(n3356), .ZN(n3357) );
  OAI21_X1 U3943 ( .B1(n3359), .B2(n3358), .A(n3357), .ZN(n3403) );
  INV_X1 U3944 ( .A(n3403), .ZN(n3362) );
  INV_X1 U3945 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3360) );
  OAI22_X1 U3946 ( .A1(n4333), .A2(n3360), .B1(n3486), .B2(n4863), .ZN(n3361)
         );
  AOI21_X1 U3947 ( .B1(n3362), .B2(n4896), .A(n3361), .ZN(n3363) );
  OAI211_X1 U3948 ( .C1(n3395), .C2(n4860), .A(n3364), .B(n3363), .ZN(U3277)
         );
  NAND2_X1 U3949 ( .A1(n3365), .A2(n3366), .ZN(n3530) );
  OAI21_X1 U3950 ( .B1(n3365), .B2(n3366), .A(n3530), .ZN(n4392) );
  XNOR2_X1 U3951 ( .A(n3367), .B(n3366), .ZN(n3371) );
  NAND2_X1 U3952 ( .A1(n4044), .A2(n4320), .ZN(n3369) );
  NAND2_X1 U3953 ( .A1(n4045), .A2(n4801), .ZN(n3368) );
  OAI211_X1 U3954 ( .C1(n4282), .C2(n3589), .A(n3369), .B(n3368), .ZN(n3370)
         );
  AOI21_X1 U3955 ( .B1(n3371), .B2(n4807), .A(n3370), .ZN(n4390) );
  INV_X1 U3956 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3373) );
  INV_X1 U3957 ( .A(n3372), .ZN(n3801) );
  OAI22_X1 U3958 ( .A1(n4333), .A2(n3373), .B1(n3801), .B2(n4863), .ZN(n3374)
         );
  INV_X1 U3959 ( .A(n3374), .ZN(n3376) );
  NAND2_X1 U3960 ( .A1(n3387), .A2(n3798), .ZN(n4387) );
  NAND3_X1 U3961 ( .A1(n4388), .A2(n4896), .A3(n4387), .ZN(n3375) );
  OAI211_X1 U3962 ( .C1(n4390), .C2(n4900), .A(n3376), .B(n3375), .ZN(n3377)
         );
  INV_X1 U3963 ( .A(n3377), .ZN(n3378) );
  OAI21_X1 U3964 ( .B1(n4392), .B2(n4335), .A(n3378), .ZN(U3274) );
  NAND2_X1 U3965 ( .A1(n3380), .A2(n3379), .ZN(n3381) );
  XNOR2_X1 U3966 ( .A(n3381), .B(n3953), .ZN(n3491) );
  INV_X1 U3967 ( .A(n3491), .ZN(n3394) );
  NAND2_X1 U3968 ( .A1(n3382), .A2(n3887), .ZN(n3383) );
  XNOR2_X1 U3969 ( .A(n3383), .B(n3953), .ZN(n3386) );
  INV_X1 U3970 ( .A(n4874), .ZN(n3502) );
  OAI22_X1 U3971 ( .A1(n3502), .A2(n4324), .B1(n4282), .B2(n3388), .ZN(n3384)
         );
  AOI21_X1 U3972 ( .B1(n4320), .B2(n4876), .A(n3384), .ZN(n3385) );
  OAI21_X1 U3973 ( .B1(n3386), .B2(n4300), .A(n3385), .ZN(n3490) );
  OAI21_X1 U3974 ( .B1(n3389), .B2(n3388), .A(n3387), .ZN(n3496) );
  AOI22_X1 U3975 ( .A1(n4900), .A2(REG2_REG_15__SCAN_IN), .B1(n3390), .B2(
        n4847), .ZN(n3391) );
  OAI21_X1 U3976 ( .B1(n3496), .B2(n4859), .A(n3391), .ZN(n3392) );
  AOI21_X1 U3977 ( .B1(n3490), .B2(n4333), .A(n3392), .ZN(n3393) );
  OAI21_X1 U3978 ( .B1(n3394), .B2(n4335), .A(n3393), .ZN(U3275) );
  INV_X1 U3979 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3398) );
  INV_X1 U3980 ( .A(n3395), .ZN(n3397) );
  AOI21_X1 U3981 ( .B1(n4781), .B2(n3397), .A(n3396), .ZN(n3400) );
  MUX2_X1 U3982 ( .A(n3398), .B(n3400), .S(n4835), .Z(n3399) );
  OAI21_X1 U3983 ( .B1(n3403), .B2(n4423), .A(n3399), .ZN(U3493) );
  INV_X1 U3984 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3401) );
  MUX2_X1 U3985 ( .A(n3401), .B(n3400), .S(n4831), .Z(n3402) );
  OAI21_X1 U3986 ( .B1(n4383), .B2(n3403), .A(n3402), .ZN(U3531) );
  AOI21_X1 U3987 ( .B1(n3405), .B2(n4826), .A(n3404), .ZN(n3409) );
  INV_X1 U3988 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3406) );
  MUX2_X1 U3989 ( .A(n3409), .B(n3406), .S(n4832), .Z(n3407) );
  OAI21_X1 U3990 ( .B1(n3411), .B2(n4423), .A(n3407), .ZN(U3495) );
  INV_X1 U3991 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3408) );
  MUX2_X1 U3992 ( .A(n3409), .B(n3408), .S(n2856), .Z(n3410) );
  OAI21_X1 U3993 ( .B1(n4383), .B2(n3411), .A(n3410), .ZN(U3532) );
  NAND2_X1 U3994 ( .A1(n3518), .A2(n3517), .ZN(n3974) );
  NAND2_X1 U3995 ( .A1(n3530), .A2(n3412), .ZN(n3413) );
  XOR2_X1 U3996 ( .A(n3974), .B(n3413), .Z(n3541) );
  INV_X1 U3997 ( .A(n3541), .ZN(n3423) );
  INV_X1 U3998 ( .A(n3520), .ZN(n3549) );
  XNOR2_X1 U3999 ( .A(n3549), .B(n3974), .ZN(n3416) );
  AOI22_X1 U4000 ( .A1(n4876), .A2(n4801), .B1(n3806), .B2(n4800), .ZN(n3415)
         );
  NAND2_X1 U4001 ( .A1(n4043), .A2(n4320), .ZN(n3414) );
  OAI211_X1 U4002 ( .C1(n3416), .C2(n4300), .A(n3415), .B(n3414), .ZN(n3540)
         );
  INV_X1 U4003 ( .A(n4388), .ZN(n3418) );
  OAI21_X1 U4004 ( .B1(n3418), .B2(n3417), .A(n3513), .ZN(n3546) );
  NOR2_X1 U4005 ( .A1(n3546), .A2(n4859), .ZN(n3421) );
  INV_X1 U4006 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3419) );
  OAI22_X1 U4007 ( .A1(n4333), .A2(n3419), .B1(n3809), .B2(n4863), .ZN(n3420)
         );
  AOI211_X1 U4008 ( .C1(n3540), .C2(n4333), .A(n3421), .B(n3420), .ZN(n3422)
         );
  OAI21_X1 U4009 ( .B1(n3423), .B2(n4335), .A(n3422), .ZN(U3273) );
  INV_X1 U4010 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3446) );
  NAND2_X1 U4011 ( .A1(n4693), .A2(REG2_REG_11__SCAN_IN), .ZN(n3439) );
  INV_X1 U4012 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4862) );
  AOI22_X1 U4013 ( .A1(n4693), .A2(REG2_REG_11__SCAN_IN), .B1(n4862), .B2(
        n4856), .ZN(n4701) );
  NAND2_X1 U4014 ( .A1(n4671), .A2(REG2_REG_9__SCAN_IN), .ZN(n3435) );
  INV_X1 U4015 ( .A(n4671), .ZN(n4846) );
  AOI22_X1 U4016 ( .A1(n4671), .A2(REG2_REG_9__SCAN_IN), .B1(n3424), .B2(n4846), .ZN(n4679) );
  INV_X1 U4017 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4642) );
  INV_X1 U4018 ( .A(n3425), .ZN(n3427) );
  NAND2_X1 U4019 ( .A1(n3452), .A2(REG2_REG_5__SCAN_IN), .ZN(n3428) );
  OAI21_X1 U4020 ( .B1(n3452), .B2(REG2_REG_5__SCAN_IN), .A(n3428), .ZN(n4631)
         );
  INV_X1 U4021 ( .A(n3453), .ZN(n4787) );
  NOR2_X1 U4022 ( .A1(n3430), .A2(n4787), .ZN(n3431) );
  INV_X1 U4023 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4649) );
  NAND2_X1 U4024 ( .A1(n3432), .A2(n3433), .ZN(n3434) );
  NAND2_X1 U4025 ( .A1(n3437), .A2(n4682), .ZN(n3438) );
  NAND2_X1 U4026 ( .A1(n3438), .A2(n4683), .ZN(n4700) );
  NAND2_X1 U4027 ( .A1(n4701), .A2(n4700), .ZN(n4699) );
  NAND2_X1 U4028 ( .A1(n3439), .A2(n4699), .ZN(n3440) );
  NAND2_X1 U4029 ( .A1(n3464), .A2(n3440), .ZN(n3441) );
  XOR2_X1 U4030 ( .A(n3440), .B(n3464), .Z(n4711) );
  INV_X1 U4031 ( .A(n4871), .ZN(n4722) );
  NOR2_X1 U4032 ( .A1(n4722), .A2(n3360), .ZN(n4714) );
  INV_X1 U4033 ( .A(n4098), .ZN(n3444) );
  NAND2_X1 U4034 ( .A1(n3442), .A2(n4093), .ZN(n3443) );
  NOR2_X1 U4035 ( .A1(n3445), .A2(n3446), .ZN(n4097) );
  AOI211_X1 U4036 ( .C1(n3446), .C2(n3445), .A(n4097), .B(n4748), .ZN(n3470)
         );
  INV_X1 U4037 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4830) );
  NOR2_X1 U4038 ( .A1(n4795), .A2(n4830), .ZN(n4656) );
  INV_X1 U4039 ( .A(REG1_REG_4__SCAN_IN), .ZN(n3449) );
  INV_X1 U4040 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4041 ( .A1(n3452), .A2(REG1_REG_5__SCAN_IN), .B1(n3451), .B2(n4785), .ZN(n4637) );
  NAND2_X1 U4042 ( .A1(n3453), .A2(n3454), .ZN(n3455) );
  XOR2_X1 U40430 ( .A(n3454), .B(n3453), .Z(n4646) );
  NAND2_X1 U4044 ( .A1(REG1_REG_6__SCAN_IN), .A2(n4646), .ZN(n4645) );
  OAI22_X1 U4045 ( .A1(n4656), .A2(n4658), .B1(n4650), .B2(REG1_REG_7__SCAN_IN), .ZN(n3456) );
  INV_X1 U4046 ( .A(n4674), .ZN(n3458) );
  NAND2_X1 U4047 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4686), .ZN(n4685) );
  NAND2_X1 U4048 ( .A1(n3461), .A2(n4682), .ZN(n3462) );
  AND2_X1 U4049 ( .A1(n4693), .A2(REG1_REG_11__SCAN_IN), .ZN(n3463) );
  INV_X1 U4050 ( .A(n3464), .ZN(n4870) );
  XNOR2_X1 U4051 ( .A(n3465), .B(n4870), .ZN(n4705) );
  NAND2_X1 U4052 ( .A1(n4871), .A2(REG1_REG_13__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U4053 ( .A1(REG1_REG_14__SCAN_IN), .A2(n3466), .ZN(n4095) );
  OAI211_X1 U4054 ( .C1(n3466), .C2(REG1_REG_14__SCAN_IN), .A(n4744), .B(n4095), .ZN(n3468) );
  AND2_X1 U4055 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n3506) );
  AOI21_X1 U4056 ( .B1(n4737), .B2(ADDR_REG_14__SCAN_IN), .A(n3506), .ZN(n3467) );
  OAI211_X1 U4057 ( .C1(n4747), .C2(n4093), .A(n3468), .B(n3467), .ZN(n3469)
         );
  OR2_X1 U4058 ( .A1(n3470), .A2(n3469), .ZN(U3254) );
  NAND2_X1 U4059 ( .A1(n4046), .A2(n3719), .ZN(n3478) );
  NAND2_X1 U4060 ( .A1(n3483), .A2(n3718), .ZN(n3477) );
  NAND2_X1 U4061 ( .A1(n3478), .A2(n3477), .ZN(n3479) );
  XNOR2_X1 U4062 ( .A(n3479), .B(n3671), .ZN(n3481) );
  AOI22_X1 U4063 ( .A1(n4046), .A2(n2933), .B1(n3719), .B2(n3483), .ZN(n3480)
         );
  OR2_X1 U4064 ( .A1(n3481), .A2(n3480), .ZN(n3498) );
  NOR2_X1 U4065 ( .A1(n2396), .A2(n3497), .ZN(n3482) );
  XNOR2_X1 U4066 ( .A(n3499), .B(n3482), .ZN(n3488) );
  AOI22_X1 U4067 ( .A1(n4879), .A2(n3483), .B1(n3840), .B2(n4874), .ZN(n3485)
         );
  INV_X1 U4068 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4609) );
  NOR2_X1 U4069 ( .A1(STATE_REG_SCAN_IN), .A2(n4609), .ZN(n4724) );
  AOI21_X1 U4070 ( .B1(n4875), .B2(n4047), .A(n4724), .ZN(n3484) );
  OAI211_X1 U4071 ( .C1(n4891), .C2(n3486), .A(n3485), .B(n3484), .ZN(n3487)
         );
  AOI21_X1 U4072 ( .B1(n3488), .B2(n4886), .A(n3487), .ZN(n3489) );
  INV_X1 U4073 ( .A(n3489), .ZN(U3231) );
  AOI21_X1 U4074 ( .B1(n3491), .B2(n4826), .A(n3490), .ZN(n3494) );
  INV_X1 U4075 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3492) );
  MUX2_X1 U4076 ( .A(n3494), .B(n3492), .S(n4832), .Z(n3493) );
  OAI21_X1 U4077 ( .B1(n3496), .B2(n4423), .A(n3493), .ZN(U3497) );
  INV_X1 U4078 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4092) );
  MUX2_X1 U4079 ( .A(n3494), .B(n4092), .S(n2856), .Z(n3495) );
  OAI21_X1 U4080 ( .B1(n4383), .B2(n3496), .A(n3495), .ZN(U3533) );
  AOI22_X1 U4081 ( .A1(n4874), .A2(n3719), .B1(n3718), .B2(n3505), .ZN(n3500)
         );
  XOR2_X1 U4082 ( .A(n3720), .B(n3500), .Z(n3579) );
  OAI22_X1 U4083 ( .A1(n3502), .A2(n3664), .B1(n4037), .B2(n3501), .ZN(n3580)
         );
  XNOR2_X1 U4084 ( .A(n3579), .B(n3580), .ZN(n3503) );
  XNOR2_X1 U4085 ( .A(n2287), .B(n3503), .ZN(n3511) );
  INV_X1 U4086 ( .A(n3504), .ZN(n3509) );
  AOI22_X1 U4087 ( .A1(n4879), .A2(n3505), .B1(n4877), .B2(n4045), .ZN(n3508)
         );
  AOI21_X1 U4088 ( .B1(n4875), .B2(n4046), .A(n3506), .ZN(n3507) );
  OAI211_X1 U4089 ( .C1(n4891), .C2(n3509), .A(n3508), .B(n3507), .ZN(n3510)
         );
  AOI21_X1 U4090 ( .B1(n3511), .B2(n4886), .A(n3510), .ZN(n3512) );
  INV_X1 U4091 ( .A(n3512), .ZN(U3212) );
  INV_X1 U4092 ( .A(n3513), .ZN(n3515) );
  INV_X1 U4093 ( .A(n4328), .ZN(n3514) );
  OAI211_X1 U4094 ( .C1(n3516), .C2(n3515), .A(n3514), .B(n4811), .ZN(n4384)
         );
  INV_X1 U4095 ( .A(n3517), .ZN(n3519) );
  OAI21_X1 U4096 ( .B1(n3520), .B2(n3519), .A(n3518), .ZN(n4315) );
  XNOR2_X1 U4097 ( .A(n4315), .B(n3535), .ZN(n3524) );
  AOI22_X1 U4098 ( .A1(n4042), .A2(n4320), .B1(n4800), .B2(n3854), .ZN(n3521)
         );
  OAI21_X1 U4099 ( .B1(n3522), .B2(n4324), .A(n3521), .ZN(n3523) );
  AOI21_X1 U4100 ( .B1(n3524), .B2(n4807), .A(n3523), .ZN(n4385) );
  OAI21_X1 U4101 ( .B1(n4168), .B2(n4384), .A(n4385), .ZN(n3538) );
  INV_X1 U4102 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4131) );
  INV_X1 U4103 ( .A(n3525), .ZN(n3858) );
  OAI22_X1 U4104 ( .A1(n4333), .A2(n4131), .B1(n3858), .B2(n4863), .ZN(n3537)
         );
  NAND2_X1 U4105 ( .A1(n3530), .A2(n3526), .ZN(n3528) );
  AND2_X1 U4106 ( .A1(n3528), .A2(n3527), .ZN(n3534) );
  NAND2_X1 U4107 ( .A1(n3530), .A2(n3529), .ZN(n3532) );
  NAND2_X1 U4108 ( .A1(n3532), .A2(n3531), .ZN(n3533) );
  AOI21_X1 U4109 ( .B1(n3535), .B2(n3534), .A(n3533), .ZN(n4386) );
  NOR2_X1 U4110 ( .A1(n4386), .A2(n4335), .ZN(n3536) );
  AOI211_X1 U4111 ( .C1(n4333), .C2(n3538), .A(n3537), .B(n3536), .ZN(n3539)
         );
  INV_X1 U4112 ( .A(n3539), .ZN(U3272) );
  AOI21_X1 U4113 ( .B1(n3541), .B2(n4826), .A(n3540), .ZN(n3543) );
  MUX2_X1 U4114 ( .A(n4115), .B(n3543), .S(n4831), .Z(n3542) );
  OAI21_X1 U4115 ( .B1(n4383), .B2(n3546), .A(n3542), .ZN(U3535) );
  INV_X1 U4116 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3544) );
  MUX2_X1 U4117 ( .A(n3544), .B(n3543), .S(n4835), .Z(n3545) );
  OAI21_X1 U4118 ( .B1(n3546), .B2(n4423), .A(n3545), .ZN(U3501) );
  AOI21_X1 U4119 ( .B1(n3549), .B2(n3548), .A(n3547), .ZN(n3553) );
  INV_X1 U4120 ( .A(n3550), .ZN(n3552) );
  OR2_X1 U4121 ( .A1(n3552), .A2(n3551), .ZN(n3947) );
  XNOR2_X1 U4122 ( .A(n3553), .B(n3947), .ZN(n3560) );
  INV_X1 U4123 ( .A(n4042), .ZN(n3555) );
  AOI22_X1 U4124 ( .A1(n4278), .A2(n4320), .B1(n3828), .B2(n4800), .ZN(n3554)
         );
  OAI21_X1 U4125 ( .B1(n3555), .B2(n4324), .A(n3554), .ZN(n3559) );
  XNOR2_X1 U4126 ( .A(n3556), .B(n3947), .ZN(n4379) );
  NOR2_X1 U4127 ( .A1(n4379), .A2(n3557), .ZN(n3558) );
  AOI211_X1 U4128 ( .C1(n3560), .C2(n4807), .A(n3559), .B(n3558), .ZN(n4378)
         );
  INV_X1 U4129 ( .A(n4379), .ZN(n3566) );
  INV_X1 U4130 ( .A(n4304), .ZN(n4376) );
  INV_X1 U4131 ( .A(n3561), .ZN(n4326) );
  NAND2_X1 U4132 ( .A1(n4326), .A2(n3828), .ZN(n4375) );
  AND3_X1 U4133 ( .A1(n4376), .A2(n4896), .A3(n4375), .ZN(n3565) );
  INV_X1 U4134 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3563) );
  INV_X1 U4135 ( .A(n3562), .ZN(n3831) );
  OAI22_X1 U4136 ( .A1(n4333), .A2(n3563), .B1(n3831), .B2(n4863), .ZN(n3564)
         );
  AOI211_X1 U4137 ( .C1(n3566), .C2(n4851), .A(n3565), .B(n3564), .ZN(n3567)
         );
  OAI21_X1 U4138 ( .B1(n4378), .B2(n4900), .A(n3567), .ZN(U3270) );
  INV_X1 U4139 ( .A(DATAI_31_), .ZN(n3709) );
  NOR2_X1 U4140 ( .A1(n3569), .A2(n3709), .ZN(n4022) );
  INV_X1 U4141 ( .A(DATAI_30_), .ZN(n3568) );
  NOR2_X1 U4142 ( .A1(n3569), .A2(n3568), .ZN(n4339) );
  NOR2_X1 U4143 ( .A1(n4019), .A2(n3570), .ZN(n4338) );
  AOI21_X1 U4144 ( .B1(n4022), .B2(n4800), .A(n4338), .ZN(n3575) );
  NOR2_X1 U4145 ( .A1(n3575), .A2(n4832), .ZN(n3571) );
  AOI21_X1 U4146 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4832), .A(n3571), .ZN(n3572) );
  OAI21_X1 U4147 ( .B1(n3578), .B2(n4423), .A(n3572), .ZN(U3517) );
  NOR2_X1 U4148 ( .A1(n3575), .A2(n2856), .ZN(n3573) );
  AOI21_X1 U4149 ( .B1(REG1_REG_31__SCAN_IN), .B2(n2856), .A(n3573), .ZN(n3574) );
  OAI21_X1 U4150 ( .B1(n3578), .B2(n4383), .A(n3574), .ZN(U3549) );
  NOR2_X1 U4151 ( .A1(n3575), .A2(n4900), .ZN(n3576) );
  AOI21_X1 U4152 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4900), .A(n3576), .ZN(n3577) );
  OAI21_X1 U4153 ( .B1(n3578), .B2(n4859), .A(n3577), .ZN(U3260) );
  NAND2_X1 U4154 ( .A1(n4045), .A2(n3719), .ZN(n3582) );
  NAND2_X1 U4155 ( .A1(n4878), .A2(n3718), .ZN(n3581) );
  NAND2_X1 U4156 ( .A1(n3582), .A2(n3581), .ZN(n3583) );
  XNOR2_X1 U4157 ( .A(n3583), .B(n3720), .ZN(n4884) );
  INV_X1 U4158 ( .A(n4884), .ZN(n3592) );
  NAND2_X1 U4159 ( .A1(n4045), .A2(n3674), .ZN(n3585) );
  NAND2_X1 U4160 ( .A1(n4878), .A2(n3719), .ZN(n3584) );
  NAND2_X1 U4161 ( .A1(n3585), .A2(n3584), .ZN(n4883) );
  INV_X1 U4162 ( .A(n4883), .ZN(n3794) );
  NAND2_X1 U4163 ( .A1(n4876), .A2(n3719), .ZN(n3587) );
  NAND2_X1 U4164 ( .A1(n3798), .A2(n3718), .ZN(n3586) );
  NAND2_X1 U4165 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  XNOR2_X1 U4166 ( .A(n3588), .B(n3671), .ZN(n3593) );
  NOR2_X1 U4167 ( .A1(n3589), .A2(n4037), .ZN(n3590) );
  AOI21_X1 U4168 ( .B1(n4876), .B2(n2933), .A(n3590), .ZN(n3594) );
  NOR2_X1 U4169 ( .A1(n3593), .A2(n3594), .ZN(n3791) );
  INV_X1 U4170 ( .A(n3791), .ZN(n3591) );
  OAI21_X1 U4171 ( .B1(n3592), .B2(n3794), .A(n3591), .ZN(n3598) );
  NOR3_X1 U4172 ( .A1(n3791), .A2(n4883), .A3(n4884), .ZN(n3597) );
  INV_X1 U4173 ( .A(n3593), .ZN(n3596) );
  INV_X1 U4174 ( .A(n3594), .ZN(n3595) );
  NOR2_X1 U4175 ( .A1(n3596), .A2(n3595), .ZN(n3790) );
  NAND2_X1 U4176 ( .A1(n4044), .A2(n3719), .ZN(n3600) );
  NAND2_X1 U4177 ( .A1(n3806), .A2(n3718), .ZN(n3599) );
  NAND2_X1 U4178 ( .A1(n3600), .A2(n3599), .ZN(n3601) );
  XNOR2_X1 U4179 ( .A(n3601), .B(n3720), .ZN(n3618) );
  NAND2_X1 U4180 ( .A1(n4044), .A2(n3674), .ZN(n3603) );
  NAND2_X1 U4181 ( .A1(n3806), .A2(n3719), .ZN(n3602) );
  NAND2_X1 U4182 ( .A1(n3603), .A2(n3602), .ZN(n3619) );
  NAND2_X1 U4183 ( .A1(n3618), .A2(n3619), .ZN(n3846) );
  NAND2_X1 U4184 ( .A1(n4043), .A2(n3719), .ZN(n3605) );
  NAND2_X1 U4185 ( .A1(n3854), .A2(n3718), .ZN(n3604) );
  NAND2_X1 U4186 ( .A1(n3605), .A2(n3604), .ZN(n3606) );
  XNOR2_X1 U4187 ( .A(n3606), .B(n3720), .ZN(n3850) );
  NAND2_X1 U4188 ( .A1(n4043), .A2(n3674), .ZN(n3608) );
  NAND2_X1 U4189 ( .A1(n3854), .A2(n3719), .ZN(n3607) );
  NAND2_X1 U4190 ( .A1(n3608), .A2(n3607), .ZN(n3851) );
  NAND2_X1 U4191 ( .A1(n3850), .A2(n3851), .ZN(n3617) );
  AND2_X1 U4192 ( .A1(n3846), .A2(n3617), .ZN(n3753) );
  NAND2_X1 U4193 ( .A1(n4042), .A2(n3719), .ZN(n3610) );
  NAND2_X1 U4194 ( .A1(n4319), .A2(n3718), .ZN(n3609) );
  NAND2_X1 U4195 ( .A1(n3610), .A2(n3609), .ZN(n3611) );
  XNOR2_X1 U4196 ( .A(n3611), .B(n3671), .ZN(n3614) );
  NOR2_X1 U4197 ( .A1(n4327), .A2(n4037), .ZN(n3612) );
  AOI21_X1 U4198 ( .B1(n4042), .B2(n2933), .A(n3612), .ZN(n3613) );
  NAND2_X1 U4199 ( .A1(n3614), .A2(n3613), .ZN(n3625) );
  OAI21_X1 U4200 ( .B1(n3614), .B2(n3613), .A(n3625), .ZN(n3758) );
  INV_X1 U4201 ( .A(n3758), .ZN(n3615) );
  AND2_X1 U4202 ( .A1(n3753), .A2(n3615), .ZN(n3616) );
  NAND2_X1 U4203 ( .A1(n3847), .A2(n3616), .ZN(n3757) );
  INV_X1 U4204 ( .A(n3617), .ZN(n3624) );
  OR2_X1 U4205 ( .A1(n3850), .A2(n3851), .ZN(n3622) );
  INV_X1 U4206 ( .A(n3618), .ZN(n3621) );
  INV_X1 U4207 ( .A(n3619), .ZN(n3620) );
  NAND2_X1 U4208 ( .A1(n3621), .A2(n3620), .ZN(n3848) );
  AND2_X1 U4209 ( .A1(n3622), .A2(n3848), .ZN(n3623) );
  OR2_X1 U4210 ( .A1(n3624), .A2(n3623), .ZN(n3754) );
  OR2_X1 U4211 ( .A1(n3758), .A2(n3754), .ZN(n3756) );
  AND2_X1 U4212 ( .A1(n3625), .A2(n3756), .ZN(n3626) );
  NAND2_X1 U4213 ( .A1(n4321), .A2(n3719), .ZN(n3628) );
  NAND2_X1 U4214 ( .A1(n3828), .A2(n3718), .ZN(n3627) );
  NAND2_X1 U4215 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  XNOR2_X1 U4216 ( .A(n3629), .B(n3671), .ZN(n3640) );
  INV_X1 U4217 ( .A(n3640), .ZN(n3633) );
  NOR2_X1 U4218 ( .A1(n4037), .A2(n3630), .ZN(n3631) );
  AOI21_X1 U4219 ( .B1(n4321), .B2(n3674), .A(n3631), .ZN(n3639) );
  INV_X1 U4220 ( .A(n3639), .ZN(n3632) );
  NAND2_X1 U4221 ( .A1(n3633), .A2(n3632), .ZN(n3826) );
  NAND2_X1 U4222 ( .A1(n4278), .A2(n3719), .ZN(n3635) );
  NAND2_X1 U4223 ( .A1(n4296), .A2(n3718), .ZN(n3634) );
  NAND2_X1 U4224 ( .A1(n3635), .A2(n3634), .ZN(n3636) );
  XNOR2_X1 U4225 ( .A(n3636), .B(n3720), .ZN(n3771) );
  NAND2_X1 U4226 ( .A1(n4278), .A2(n2933), .ZN(n3638) );
  NAND2_X1 U4227 ( .A1(n4296), .A2(n3719), .ZN(n3637) );
  NAND2_X1 U4228 ( .A1(n3638), .A2(n3637), .ZN(n3770) );
  NAND2_X1 U4229 ( .A1(n3640), .A2(n3639), .ZN(n3825) );
  OAI21_X1 U4230 ( .B1(n3771), .B2(n3770), .A(n3825), .ZN(n3641) );
  INV_X1 U4231 ( .A(n3771), .ZN(n3643) );
  INV_X1 U4232 ( .A(n3770), .ZN(n3642) );
  NOR2_X1 U4233 ( .A1(n3643), .A2(n3642), .ZN(n3835) );
  OAI22_X1 U4234 ( .A1(n3645), .A2(n4037), .B1(n3662), .B2(n4281), .ZN(n3644)
         );
  XNOR2_X1 U4235 ( .A(n3644), .B(n3720), .ZN(n3648) );
  OAI22_X1 U4236 ( .A1(n3645), .A2(n3664), .B1(n4037), .B2(n4281), .ZN(n3647)
         );
  XNOR2_X1 U4237 ( .A(n3648), .B(n3647), .ZN(n3838) );
  OR2_X1 U4238 ( .A1(n3835), .A2(n3838), .ZN(n3646) );
  NOR2_X1 U4239 ( .A1(n3648), .A2(n3647), .ZN(n3735) );
  NAND2_X1 U4240 ( .A1(n4277), .A2(n3719), .ZN(n3650) );
  NAND2_X1 U4241 ( .A1(n4259), .A2(n3718), .ZN(n3649) );
  NAND2_X1 U4242 ( .A1(n3650), .A2(n3649), .ZN(n3651) );
  XNOR2_X1 U4243 ( .A(n3651), .B(n3671), .ZN(n3653) );
  NOR2_X1 U4244 ( .A1(n4037), .A2(n4266), .ZN(n3652) );
  AOI21_X1 U4245 ( .B1(n4277), .B2(n3674), .A(n3652), .ZN(n3654) );
  XNOR2_X1 U4246 ( .A(n3653), .B(n3654), .ZN(n3734) );
  INV_X1 U4247 ( .A(n3653), .ZN(n3656) );
  INV_X1 U4248 ( .A(n3654), .ZN(n3655) );
  NAND2_X1 U4249 ( .A1(n3656), .A2(n3655), .ZN(n3660) );
  NAND2_X1 U4250 ( .A1(n4260), .A2(n3719), .ZN(n3658) );
  NAND2_X1 U4251 ( .A1(n4236), .A2(n3718), .ZN(n3657) );
  NAND2_X1 U4252 ( .A1(n3658), .A2(n3657), .ZN(n3659) );
  XNOR2_X1 U4253 ( .A(n3659), .B(n3671), .ZN(n3661) );
  OAI22_X1 U4254 ( .A1(n4222), .A2(n3664), .B1(n4037), .B2(n4241), .ZN(n3816)
         );
  NAND3_X1 U4255 ( .A1(n3736), .A2(n3661), .A3(n3660), .ZN(n3813) );
  OAI21_X2 U4256 ( .B1(n3814), .B2(n3816), .A(n3813), .ZN(n3783) );
  OAI22_X1 U4257 ( .A1(n3665), .A2(n4037), .B1(n3662), .B2(n4226), .ZN(n3663)
         );
  XOR2_X1 U4258 ( .A(n3720), .B(n3663), .Z(n3780) );
  NAND2_X1 U4259 ( .A1(n3783), .A2(n3780), .ZN(n3666) );
  OAI22_X1 U4260 ( .A1(n3665), .A2(n3664), .B1(n4037), .B2(n4226), .ZN(n3781)
         );
  INV_X1 U4261 ( .A(n3783), .ZN(n3668) );
  INV_X1 U4262 ( .A(n3780), .ZN(n3667) );
  NAND2_X1 U4263 ( .A1(n4219), .A2(n3719), .ZN(n3670) );
  NAND2_X1 U4264 ( .A1(n4207), .A2(n3718), .ZN(n3669) );
  NAND2_X1 U4265 ( .A1(n3670), .A2(n3669), .ZN(n3672) );
  XNOR2_X1 U4266 ( .A(n3672), .B(n3671), .ZN(n3676) );
  NOR2_X1 U4267 ( .A1(n4037), .A2(n4201), .ZN(n3673) );
  AOI21_X1 U4268 ( .B1(n4219), .B2(n3674), .A(n3673), .ZN(n3675) );
  NOR2_X1 U4269 ( .A1(n3676), .A2(n3675), .ZN(n3863) );
  NAND2_X1 U4270 ( .A1(n3676), .A2(n3675), .ZN(n3685) );
  NAND2_X1 U4271 ( .A1(n3687), .A2(n3685), .ZN(n3684) );
  NAND2_X1 U4272 ( .A1(n4198), .A2(n3719), .ZN(n3678) );
  NAND2_X1 U4273 ( .A1(n2744), .A2(n3718), .ZN(n3677) );
  NAND2_X1 U4274 ( .A1(n3678), .A2(n3677), .ZN(n3679) );
  XNOR2_X1 U4275 ( .A(n3679), .B(n3720), .ZN(n3683) );
  NAND2_X1 U4276 ( .A1(n4198), .A2(n2933), .ZN(n3681) );
  NAND2_X1 U4277 ( .A1(n2744), .A2(n3719), .ZN(n3680) );
  NAND2_X1 U4278 ( .A1(n3681), .A2(n3680), .ZN(n3682) );
  NAND2_X1 U4279 ( .A1(n3683), .A2(n3682), .ZN(n3712) );
  OAI21_X1 U4280 ( .B1(n3683), .B2(n3682), .A(n3712), .ZN(n3686) );
  AOI21_X1 U4281 ( .B1(n3684), .B2(n3686), .A(n3871), .ZN(n3693) );
  INV_X1 U4282 ( .A(n3685), .ZN(n3862) );
  NOR2_X1 U4283 ( .A1(n3686), .A2(n3862), .ZN(n3714) );
  NAND2_X1 U4284 ( .A1(n3687), .A2(n3714), .ZN(n3692) );
  INV_X1 U4285 ( .A(n4179), .ZN(n3690) );
  AOI22_X1 U4286 ( .A1(n4879), .A2(n2744), .B1(n3818), .B2(n4219), .ZN(n3689)
         );
  AOI22_X1 U4287 ( .A1(n3840), .A2(n4175), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3688) );
  OAI211_X1 U4288 ( .C1(n4891), .C2(n3690), .A(n3689), .B(n3688), .ZN(n3691)
         );
  AOI21_X1 U4289 ( .B1(n3693), .B2(n3692), .A(n3691), .ZN(n3694) );
  INV_X1 U4290 ( .A(n3694), .ZN(U3211) );
  INV_X1 U4291 ( .A(n4879), .ZN(n3761) );
  NAND2_X1 U4292 ( .A1(n3695), .A2(n4886), .ZN(n3697) );
  AOI22_X1 U4293 ( .A1(n3703), .A2(REG3_REG_0__SCAN_IN), .B1(n4877), .B2(n4057), .ZN(n3696) );
  OAI211_X1 U4294 ( .C1(n3761), .C2(n3698), .A(n3697), .B(n3696), .ZN(U3229)
         );
  AOI21_X1 U4295 ( .B1(n3701), .B2(n3700), .A(n3699), .ZN(n3706) );
  AOI22_X1 U4296 ( .A1(n3840), .A2(n4055), .B1(n4875), .B2(n4057), .ZN(n3705)
         );
  AOI22_X1 U4297 ( .A1(REG3_REG_2__SCAN_IN), .A2(n3703), .B1(n4879), .B2(n3702), .ZN(n3704) );
  OAI211_X1 U4298 ( .C1(n3706), .C2(n3871), .A(n3705), .B(n3704), .ZN(U3234)
         );
  INV_X1 U4299 ( .A(n3707), .ZN(n3711) );
  NAND3_X1 U4300 ( .A1(n3708), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3710) );
  OAI22_X1 U4301 ( .A1(n3711), .A2(n3710), .B1(STATE_REG_SCAN_IN), .B2(n3709), 
        .ZN(U3321) );
  INV_X1 U4302 ( .A(n3712), .ZN(n3715) );
  OR2_X1 U4303 ( .A1(n3863), .A2(n3715), .ZN(n3713) );
  NOR2_X1 U4304 ( .A1(n3865), .A2(n3713), .ZN(n3717) );
  NOR2_X1 U4305 ( .A1(n3715), .A2(n3714), .ZN(n3716) );
  NOR2_X1 U4306 ( .A1(n3717), .A2(n3716), .ZN(n3725) );
  AOI22_X1 U4307 ( .A1(n4175), .A2(n3719), .B1(n3718), .B2(n4162), .ZN(n3723)
         );
  AOI22_X1 U4308 ( .A1(n4175), .A2(n2933), .B1(n3719), .B2(n4162), .ZN(n3721)
         );
  XNOR2_X1 U4309 ( .A(n3721), .B(n3720), .ZN(n3722) );
  XOR2_X1 U4310 ( .A(n3723), .B(n3722), .Z(n3724) );
  XNOR2_X1 U4311 ( .A(n3725), .B(n3724), .ZN(n3733) );
  INV_X1 U4312 ( .A(n4154), .ZN(n3730) );
  AOI22_X1 U4313 ( .A1(n4879), .A2(n4162), .B1(n3818), .B2(n4198), .ZN(n3729)
         );
  NOR2_X1 U4314 ( .A1(n3726), .A2(STATE_REG_SCAN_IN), .ZN(n3727) );
  AOI21_X1 U4315 ( .B1(n4877), .B2(n4163), .A(n3727), .ZN(n3728) );
  OAI211_X1 U4316 ( .C1(n4891), .C2(n3730), .A(n3729), .B(n3728), .ZN(n3731)
         );
  INV_X1 U4317 ( .A(n3731), .ZN(n3732) );
  OAI21_X1 U4318 ( .B1(n3733), .B2(n3871), .A(n3732), .ZN(U3217) );
  OAI21_X1 U4319 ( .B1(n2266), .B2(n3735), .A(n3734), .ZN(n3737) );
  NAND3_X1 U4320 ( .A1(n3737), .A2(n4886), .A3(n3736), .ZN(n3742) );
  AOI22_X1 U4321 ( .A1(n4875), .A2(n4297), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3741) );
  AOI22_X1 U4322 ( .A1(n4879), .A2(n4259), .B1(n4877), .B2(n4260), .ZN(n3740)
         );
  INV_X1 U4323 ( .A(n4267), .ZN(n3738) );
  OR2_X1 U4324 ( .A1(n4891), .A2(n3738), .ZN(n3739) );
  NAND4_X1 U4325 ( .A1(n3742), .A2(n3741), .A3(n3740), .A4(n3739), .ZN(U3213)
         );
  AND2_X1 U4326 ( .A1(n3274), .A2(n3743), .ZN(n3746) );
  OAI211_X1 U4327 ( .C1(n3746), .C2(n3745), .A(n4886), .B(n3744), .ZN(n3752)
         );
  NOR2_X1 U4328 ( .A1(STATE_REG_SCAN_IN), .A2(n4582), .ZN(n4690) );
  AOI21_X1 U4329 ( .B1(n4877), .B2(n4048), .A(n4690), .ZN(n3751) );
  AOI22_X1 U4330 ( .A1(n4879), .A2(n3747), .B1(n3818), .B2(n4050), .ZN(n3750)
         );
  INV_X1 U4331 ( .A(n4848), .ZN(n3748) );
  OR2_X1 U4332 ( .A1(n4891), .A2(n3748), .ZN(n3749) );
  NAND4_X1 U4333 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(U3214)
         );
  NAND2_X1 U4334 ( .A1(n3847), .A2(n3753), .ZN(n3755) );
  AND2_X1 U4335 ( .A1(n3755), .A2(n3754), .ZN(n3759) );
  AOI21_X1 U4336 ( .B1(n3759), .B2(n3758), .A(n2276), .ZN(n3767) );
  AND2_X1 U4337 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4736) );
  OAI22_X1 U4338 ( .A1(n3761), .A2(n4327), .B1(n3760), .B2(n4325), .ZN(n3762)
         );
  AOI211_X1 U4339 ( .C1(n4877), .C2(n4321), .A(n4736), .B(n3762), .ZN(n3766)
         );
  INV_X1 U4340 ( .A(n4891), .ZN(n3764) );
  NAND2_X1 U4341 ( .A1(n3764), .A2(n3763), .ZN(n3765) );
  OAI211_X1 U4342 ( .C1(n3767), .C2(n3871), .A(n3766), .B(n3765), .ZN(U3216)
         );
  INV_X1 U4343 ( .A(n3825), .ZN(n3769) );
  OAI21_X1 U4344 ( .B1(n3768), .B2(n3769), .A(n3826), .ZN(n3773) );
  XNOR2_X1 U4345 ( .A(n3771), .B(n3770), .ZN(n3772) );
  XNOR2_X1 U4346 ( .A(n3773), .B(n3772), .ZN(n3778) );
  INV_X1 U4347 ( .A(n3774), .ZN(n4305) );
  AOI22_X1 U4348 ( .A1(n4879), .A2(n4296), .B1(n3818), .B2(n4321), .ZN(n3776)
         );
  AOI22_X1 U4349 ( .A1(n3840), .A2(n4297), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3775) );
  OAI211_X1 U4350 ( .C1(n4891), .C2(n4305), .A(n3776), .B(n3775), .ZN(n3777)
         );
  AOI21_X1 U4351 ( .B1(n3778), .B2(n4886), .A(n3777), .ZN(n3779) );
  INV_X1 U4352 ( .A(n3779), .ZN(U3220) );
  XOR2_X1 U4353 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR2_X1 U4354 ( .A(n3783), .B(n3782), .ZN(n3789) );
  INV_X1 U4355 ( .A(n3784), .ZN(n4223) );
  AOI22_X1 U4356 ( .A1(n4879), .A2(n4218), .B1(n3818), .B2(n4260), .ZN(n3786)
         );
  AOI22_X1 U4357 ( .A1(n4877), .A2(n4219), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3785) );
  OAI211_X1 U4358 ( .C1(n4891), .C2(n4223), .A(n3786), .B(n3785), .ZN(n3787)
         );
  INV_X1 U4359 ( .A(n3787), .ZN(n3788) );
  OAI21_X1 U4360 ( .B1(n3789), .B2(n3871), .A(n3788), .ZN(U3222) );
  NOR2_X1 U4361 ( .A1(n3791), .A2(n3790), .ZN(n3797) );
  INV_X1 U4362 ( .A(n3792), .ZN(n3795) );
  OAI21_X1 U4363 ( .B1(n3792), .B2(n4883), .A(n4884), .ZN(n3793) );
  OAI21_X1 U4364 ( .B1(n3795), .B2(n3794), .A(n3793), .ZN(n3796) );
  XOR2_X1 U4365 ( .A(n3797), .B(n3796), .Z(n3803) );
  AOI22_X1 U4366 ( .A1(n4879), .A2(n3798), .B1(n3840), .B2(n4044), .ZN(n3800)
         );
  NOR2_X1 U4367 ( .A1(STATE_REG_SCAN_IN), .A2(n4529), .ZN(n4730) );
  AOI21_X1 U4368 ( .B1(n3818), .B2(n4045), .A(n4730), .ZN(n3799) );
  OAI211_X1 U4369 ( .C1(n4891), .C2(n3801), .A(n3800), .B(n3799), .ZN(n3802)
         );
  AOI21_X1 U4370 ( .B1(n3803), .B2(n4886), .A(n3802), .ZN(n3804) );
  INV_X1 U4371 ( .A(n3804), .ZN(U3223) );
  NAND2_X1 U4372 ( .A1(n3846), .A2(n3848), .ZN(n3805) );
  XOR2_X1 U4373 ( .A(n3805), .B(n3847), .Z(n3811) );
  AOI22_X1 U4374 ( .A1(n4879), .A2(n3806), .B1(n3840), .B2(n4043), .ZN(n3808)
         );
  AND2_X1 U4375 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4124) );
  AOI21_X1 U4376 ( .B1(n4875), .B2(n4876), .A(n4124), .ZN(n3807) );
  OAI211_X1 U4377 ( .C1(n4891), .C2(n3809), .A(n3808), .B(n3807), .ZN(n3810)
         );
  AOI21_X1 U4378 ( .B1(n3811), .B2(n4886), .A(n3810), .ZN(n3812) );
  INV_X1 U4379 ( .A(n3812), .ZN(U3225) );
  INV_X1 U4380 ( .A(n3813), .ZN(n3815) );
  NOR2_X1 U4381 ( .A1(n3815), .A2(n3814), .ZN(n3817) );
  XNOR2_X1 U4382 ( .A(n3817), .B(n3816), .ZN(n3824) );
  INV_X1 U4383 ( .A(n4244), .ZN(n3821) );
  AOI22_X1 U4384 ( .A1(n4879), .A2(n4236), .B1(n3818), .B2(n4277), .ZN(n3820)
         );
  AOI22_X1 U4385 ( .A1(n4877), .A2(n4237), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3819) );
  OAI211_X1 U4386 ( .C1(n4891), .C2(n3821), .A(n3820), .B(n3819), .ZN(n3822)
         );
  INV_X1 U4387 ( .A(n3822), .ZN(n3823) );
  OAI21_X1 U4388 ( .B1(n3824), .B2(n3871), .A(n3823), .ZN(U3226) );
  NAND2_X1 U4389 ( .A1(n3826), .A2(n3825), .ZN(n3827) );
  XOR2_X1 U4390 ( .A(n3827), .B(n3768), .Z(n3833) );
  AOI22_X1 U4391 ( .A1(n4879), .A2(n3828), .B1(n4875), .B2(n4042), .ZN(n3830)
         );
  AOI22_X1 U4392 ( .A1(n3840), .A2(n4278), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3829) );
  OAI211_X1 U4393 ( .C1(n4891), .C2(n3831), .A(n3830), .B(n3829), .ZN(n3832)
         );
  AOI21_X1 U4394 ( .B1(n3833), .B2(n4886), .A(n3832), .ZN(n3834) );
  INV_X1 U4395 ( .A(n3834), .ZN(U3230) );
  OR2_X1 U4396 ( .A1(n3836), .A2(n3835), .ZN(n3837) );
  AOI21_X1 U4397 ( .B1(n3838), .B2(n3837), .A(n2266), .ZN(n3845) );
  INV_X1 U4398 ( .A(n3839), .ZN(n4285) );
  AOI22_X1 U4399 ( .A1(n4879), .A2(n4288), .B1(n3840), .B2(n4277), .ZN(n3842)
         );
  AOI22_X1 U4400 ( .A1(n4875), .A2(n4278), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3841) );
  OAI211_X1 U4401 ( .C1(n4891), .C2(n4285), .A(n3842), .B(n3841), .ZN(n3843)
         );
  INV_X1 U4402 ( .A(n3843), .ZN(n3844) );
  OAI21_X1 U4403 ( .B1(n3845), .B2(n3871), .A(n3844), .ZN(U3232) );
  NAND2_X1 U4404 ( .A1(n3847), .A2(n3846), .ZN(n3849) );
  NAND2_X1 U4405 ( .A1(n3849), .A2(n3848), .ZN(n3853) );
  XOR2_X1 U4406 ( .A(n3851), .B(n3850), .Z(n3852) );
  XNOR2_X1 U4407 ( .A(n3853), .B(n3852), .ZN(n3860) );
  AOI22_X1 U4408 ( .A1(n4879), .A2(n3854), .B1(n4875), .B2(n4044), .ZN(n3857)
         );
  NOR2_X1 U4409 ( .A1(STATE_REG_SCAN_IN), .A2(n3855), .ZN(n4135) );
  AOI21_X1 U4410 ( .B1(n4877), .B2(n4042), .A(n4135), .ZN(n3856) );
  OAI211_X1 U4411 ( .C1(n4891), .C2(n3858), .A(n3857), .B(n3856), .ZN(n3859)
         );
  AOI21_X1 U4412 ( .B1(n3860), .B2(n4886), .A(n3859), .ZN(n3861) );
  INV_X1 U4413 ( .A(n3861), .ZN(U3235) );
  NOR2_X1 U4414 ( .A1(n3863), .A2(n3862), .ZN(n3864) );
  XNOR2_X1 U4415 ( .A(n3865), .B(n3864), .ZN(n3872) );
  INV_X1 U4416 ( .A(n3866), .ZN(n4204) );
  AOI22_X1 U4417 ( .A1(n4879), .A2(n4207), .B1(n4875), .B2(n4237), .ZN(n3868)
         );
  AOI22_X1 U4418 ( .A1(n4877), .A2(n4198), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3867) );
  OAI211_X1 U4419 ( .C1(n4891), .C2(n4204), .A(n3868), .B(n3867), .ZN(n3869)
         );
  INV_X1 U4420 ( .A(n3869), .ZN(n3870) );
  OAI21_X1 U4421 ( .B1(n3872), .B2(n3871), .A(n3870), .ZN(U3237) );
  OR2_X1 U4422 ( .A1(n3935), .A2(n4339), .ZN(n3874) );
  NAND2_X1 U4423 ( .A1(n4019), .A2(n4022), .ZN(n3873) );
  AND2_X1 U4424 ( .A1(n3874), .A2(n3873), .ZN(n3991) );
  INV_X1 U4425 ( .A(n4003), .ZN(n3923) );
  NAND2_X1 U4426 ( .A1(n3876), .A2(n3875), .ZN(n3914) );
  AND2_X1 U4427 ( .A1(n3914), .A2(n3886), .ZN(n3997) );
  NAND3_X1 U4428 ( .A1(n3879), .A2(n3878), .A3(n3877), .ZN(n3908) );
  INV_X1 U4429 ( .A(n3905), .ZN(n3880) );
  OR3_X1 U4430 ( .A1(n3908), .A2(n3881), .A3(n3880), .ZN(n3884) );
  NAND2_X1 U4431 ( .A1(n3883), .A2(n3882), .ZN(n3918) );
  AOI21_X1 U4432 ( .B1(n3885), .B2(n3884), .A(n3918), .ZN(n3890) );
  NAND2_X1 U4433 ( .A1(n3887), .A2(n3886), .ZN(n4000) );
  INV_X1 U4434 ( .A(n3888), .ZN(n3889) );
  NOR3_X1 U4435 ( .A1(n3890), .A2(n4000), .A3(n3889), .ZN(n3920) );
  INV_X1 U4436 ( .A(n3891), .ZN(n3893) );
  OAI211_X1 U4437 ( .C1(n3894), .C2(n4023), .A(n3893), .B(n3892), .ZN(n3897)
         );
  NAND3_X1 U4438 ( .A1(n3897), .A2(n3896), .A3(n3895), .ZN(n3900) );
  NAND3_X1 U4439 ( .A1(n3900), .A2(n3899), .A3(n3898), .ZN(n3903) );
  NAND3_X1 U4440 ( .A1(n3903), .A2(n3902), .A3(n3901), .ZN(n3907) );
  NAND4_X1 U4441 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3910)
         );
  AOI21_X1 U4442 ( .B1(n3910), .B2(n3909), .A(n3908), .ZN(n3917) );
  AOI21_X1 U4443 ( .B1(n3913), .B2(n3912), .A(n3911), .ZN(n3916) );
  INV_X1 U4444 ( .A(n3914), .ZN(n3915) );
  OAI21_X1 U4445 ( .B1(n3917), .B2(n3916), .A(n3915), .ZN(n3919) );
  OAI22_X1 U4446 ( .A1(n3997), .A2(n3920), .B1(n3919), .B2(n3918), .ZN(n3922)
         );
  OAI211_X1 U4447 ( .C1(n3923), .C2(n3922), .A(n3999), .B(n3921), .ZN(n3925)
         );
  INV_X1 U4448 ( .A(n3924), .ZN(n4010) );
  OAI221_X1 U4449 ( .B1(n3946), .B2(n4005), .C1(n3946), .C2(n3925), .A(n4010), 
        .ZN(n3926) );
  AOI21_X1 U4450 ( .B1(n3927), .B2(n3926), .A(n4012), .ZN(n3930) );
  INV_X1 U4451 ( .A(n4011), .ZN(n3929) );
  INV_X1 U4452 ( .A(n3995), .ZN(n3928) );
  OAI21_X1 U4453 ( .B1(n3930), .B2(n3929), .A(n3928), .ZN(n3931) );
  NAND4_X1 U4454 ( .A1(n3991), .A2(n3932), .A3(n3992), .A4(n3931), .ZN(n3941)
         );
  NAND2_X1 U4455 ( .A1(n4163), .A2(n3938), .ZN(n3933) );
  AND2_X1 U4456 ( .A1(n3934), .A2(n3933), .ZN(n3993) );
  INV_X1 U4457 ( .A(n3993), .ZN(n3940) );
  NOR2_X1 U4458 ( .A1(n4019), .A2(n4022), .ZN(n3937) );
  NOR2_X1 U4459 ( .A1(n3991), .A2(n3937), .ZN(n3939) );
  AND2_X1 U4460 ( .A1(n3935), .A2(n4339), .ZN(n3936) );
  NOR2_X1 U4461 ( .A1(n3937), .A2(n3936), .ZN(n3957) );
  OAI21_X1 U4462 ( .B1(n4163), .B2(n3938), .A(n3957), .ZN(n3994) );
  AOI21_X1 U4463 ( .B1(n3993), .B2(n3996), .A(n3994), .ZN(n4017) );
  OAI22_X1 U4464 ( .A1(n3941), .A2(n3940), .B1(n3939), .B2(n4017), .ZN(n4031)
         );
  NAND2_X1 U4465 ( .A1(n4031), .A2(n4814), .ZN(n4029) );
  NAND2_X1 U4466 ( .A1(n3943), .A2(n3942), .ZN(n4316) );
  INV_X1 U4467 ( .A(n4316), .ZN(n3951) );
  NOR2_X1 U4468 ( .A1(n3945), .A2(n3944), .ZN(n3950) );
  INV_X1 U4469 ( .A(n3946), .ZN(n4255) );
  NAND2_X1 U4470 ( .A1(n4255), .A2(n4253), .ZN(n4294) );
  NOR4_X1 U4471 ( .A1(n4275), .A2(n3948), .A3(n4294), .A4(n3947), .ZN(n3949)
         );
  NAND4_X1 U4472 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3990)
         );
  INV_X1 U4473 ( .A(n4754), .ZN(n3956) );
  INV_X1 U4474 ( .A(n3953), .ZN(n3955) );
  NAND4_X1 U4475 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3963)
         );
  NAND4_X1 U4476 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3962)
         );
  NOR2_X1 U4477 ( .A1(n3963), .A2(n3962), .ZN(n3988) );
  NAND2_X1 U4478 ( .A1(n4193), .A2(n3964), .ZN(n4215) );
  INV_X1 U4479 ( .A(n4215), .ZN(n3969) );
  NAND2_X1 U4480 ( .A1(n3965), .A2(n4213), .ZN(n4234) );
  INV_X1 U4481 ( .A(n4234), .ZN(n3968) );
  NAND2_X1 U4482 ( .A1(n4232), .A2(n3966), .ZN(n4257) );
  INV_X1 U4483 ( .A(n4257), .ZN(n3967) );
  NAND4_X1 U4484 ( .A1(n3991), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(n3972)
         );
  NAND2_X1 U4485 ( .A1(n3970), .A2(n3992), .ZN(n4191) );
  INV_X1 U4486 ( .A(n4191), .ZN(n4196) );
  NAND2_X1 U4487 ( .A1(n4196), .A2(n4180), .ZN(n3971) );
  NOR2_X1 U4488 ( .A1(n3972), .A2(n3971), .ZN(n3987) );
  NOR2_X1 U4489 ( .A1(n3974), .A2(n3973), .ZN(n3976) );
  NAND3_X1 U4490 ( .A1(n3977), .A2(n3976), .A3(n3975), .ZN(n3982) );
  INV_X1 U4491 ( .A(n4160), .ZN(n3979) );
  NAND4_X1 U4492 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n4815), .ZN(n3981)
         );
  NOR2_X1 U4493 ( .A1(n3982), .A2(n3981), .ZN(n3986) );
  NOR2_X1 U4494 ( .A1(n3984), .A2(n3983), .ZN(n3985) );
  NAND4_X1 U4495 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3989)
         );
  NOR2_X1 U4496 ( .A1(n3990), .A2(n3989), .ZN(n4025) );
  INV_X1 U4497 ( .A(n3991), .ZN(n4021) );
  NAND3_X1 U4498 ( .A1(n4180), .A2(n3993), .A3(n3992), .ZN(n4016) );
  NOR3_X1 U4499 ( .A1(n3996), .A2(n3995), .A3(n3994), .ZN(n4015) );
  INV_X1 U4500 ( .A(n3997), .ZN(n3998) );
  OAI211_X1 U4501 ( .C1(n4001), .C2(n4000), .A(n3999), .B(n3998), .ZN(n4004)
         );
  AOI21_X1 U4502 ( .B1(n4004), .B2(n4003), .A(n4002), .ZN(n4007) );
  INV_X1 U4503 ( .A(n4005), .ZN(n4006) );
  NOR2_X1 U4504 ( .A1(n4007), .A2(n4006), .ZN(n4009) );
  AOI21_X1 U4505 ( .B1(n4010), .B2(n4009), .A(n4008), .ZN(n4013) );
  OAI21_X1 U4506 ( .B1(n4013), .B2(n4012), .A(n4011), .ZN(n4014) );
  AOI22_X1 U4507 ( .A1(n4017), .A2(n4016), .B1(n4015), .B2(n4014), .ZN(n4018)
         );
  AOI21_X1 U4508 ( .B1(n4019), .B2(n4339), .A(n4018), .ZN(n4020) );
  AOI21_X1 U4509 ( .B1(n4022), .B2(n4021), .A(n4020), .ZN(n4024) );
  MUX2_X1 U4510 ( .A(n4025), .B(n4024), .S(n4023), .Z(n4026) );
  XNOR2_X1 U4511 ( .A(n4026), .B(n4168), .ZN(n4028) );
  MUX2_X1 U4512 ( .A(n4029), .B(n4028), .S(n4027), .Z(n4030) );
  OAI21_X1 U4513 ( .B1(n4031), .B2(n4752), .A(n4030), .ZN(n4032) );
  INV_X1 U4514 ( .A(n4032), .ZN(n4041) );
  INV_X1 U4515 ( .A(n4033), .ZN(n4035) );
  NAND4_X1 U4516 ( .A1(n4060), .A2(STATE_REG_SCAN_IN), .A3(n4035), .A4(n4034), 
        .ZN(n4036) );
  NOR3_X1 U4517 ( .A1(n4037), .A2(n4895), .A3(n4036), .ZN(n4040) );
  OAI21_X1 U4518 ( .B1(n4433), .B2(n4038), .A(B_REG_SCAN_IN), .ZN(n4039) );
  OAI22_X1 U4519 ( .A1(n4041), .A2(n4433), .B1(n4040), .B2(n4039), .ZN(U3239)
         );
  MUX2_X1 U4520 ( .A(n4163), .B(DATAO_REG_29__SCAN_IN), .S(n4058), .Z(U3579)
         );
  MUX2_X1 U4521 ( .A(n4175), .B(DATAO_REG_28__SCAN_IN), .S(n4058), .Z(U3578)
         );
  MUX2_X1 U4522 ( .A(n4198), .B(DATAO_REG_27__SCAN_IN), .S(n4058), .Z(U3577)
         );
  MUX2_X1 U4523 ( .A(n4219), .B(DATAO_REG_26__SCAN_IN), .S(n4058), .Z(U3576)
         );
  MUX2_X1 U4524 ( .A(n4237), .B(DATAO_REG_25__SCAN_IN), .S(n4058), .Z(U3575)
         );
  MUX2_X1 U4525 ( .A(n4260), .B(DATAO_REG_24__SCAN_IN), .S(n4058), .Z(U3574)
         );
  MUX2_X1 U4526 ( .A(n4277), .B(DATAO_REG_23__SCAN_IN), .S(n4058), .Z(U3573)
         );
  MUX2_X1 U4527 ( .A(n4297), .B(DATAO_REG_22__SCAN_IN), .S(n4058), .Z(U3572)
         );
  MUX2_X1 U4528 ( .A(n4278), .B(DATAO_REG_21__SCAN_IN), .S(n4058), .Z(U3571)
         );
  MUX2_X1 U4529 ( .A(n4321), .B(DATAO_REG_20__SCAN_IN), .S(n4058), .Z(U3570)
         );
  MUX2_X1 U4530 ( .A(n4042), .B(DATAO_REG_19__SCAN_IN), .S(n4058), .Z(U3569)
         );
  MUX2_X1 U4531 ( .A(n4043), .B(DATAO_REG_18__SCAN_IN), .S(n4058), .Z(U3568)
         );
  MUX2_X1 U4532 ( .A(n4044), .B(DATAO_REG_17__SCAN_IN), .S(n4058), .Z(U3567)
         );
  MUX2_X1 U4533 ( .A(n4876), .B(DATAO_REG_16__SCAN_IN), .S(n4058), .Z(U3566)
         );
  MUX2_X1 U4534 ( .A(n4045), .B(DATAO_REG_15__SCAN_IN), .S(n4058), .Z(U3565)
         );
  MUX2_X1 U4535 ( .A(n4874), .B(DATAO_REG_14__SCAN_IN), .S(n4058), .Z(U3564)
         );
  MUX2_X1 U4536 ( .A(n4046), .B(DATAO_REG_13__SCAN_IN), .S(n4058), .Z(U3563)
         );
  MUX2_X1 U4537 ( .A(n4047), .B(DATAO_REG_12__SCAN_IN), .S(n4058), .Z(U3562)
         );
  MUX2_X1 U4538 ( .A(n4048), .B(DATAO_REG_11__SCAN_IN), .S(n4058), .Z(U3561)
         );
  MUX2_X1 U4539 ( .A(n4049), .B(DATAO_REG_10__SCAN_IN), .S(n4058), .Z(U3560)
         );
  MUX2_X1 U4540 ( .A(n4050), .B(DATAO_REG_9__SCAN_IN), .S(n4058), .Z(U3559) );
  MUX2_X1 U4541 ( .A(DATAO_REG_8__SCAN_IN), .B(n4051), .S(U4043), .Z(U3558) );
  MUX2_X1 U4542 ( .A(n4052), .B(DATAO_REG_7__SCAN_IN), .S(n4058), .Z(U3557) );
  MUX2_X1 U4543 ( .A(n4802), .B(DATAO_REG_6__SCAN_IN), .S(n4058), .Z(U3556) );
  MUX2_X1 U4544 ( .A(DATAO_REG_5__SCAN_IN), .B(n4053), .S(U4043), .Z(U3555) );
  MUX2_X1 U4545 ( .A(n4054), .B(DATAO_REG_4__SCAN_IN), .S(n4058), .Z(U3554) );
  MUX2_X1 U4546 ( .A(n4055), .B(DATAO_REG_3__SCAN_IN), .S(n4058), .Z(U3553) );
  MUX2_X1 U4547 ( .A(n4056), .B(DATAO_REG_2__SCAN_IN), .S(n4058), .Z(U3552) );
  MUX2_X1 U4548 ( .A(n4057), .B(DATAO_REG_1__SCAN_IN), .S(n4058), .Z(U3551) );
  MUX2_X1 U4549 ( .A(n2912), .B(DATAO_REG_0__SCAN_IN), .S(n4058), .Z(U3550) );
  AOI22_X1 U4550 ( .A1(n4737), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4067) );
  NAND3_X1 U4551 ( .A1(n4744), .A2(IR_REG_0__SCAN_IN), .A3(n4059), .ZN(n4066)
         );
  NOR2_X1 U4552 ( .A1(n4060), .A2(REG1_REG_0__SCAN_IN), .ZN(n4061) );
  OAI21_X1 U4553 ( .B1(IR_REG_0__SCAN_IN), .B2(n4061), .A(n4064), .ZN(n4063)
         );
  OAI211_X1 U4554 ( .C1(IR_REG_0__SCAN_IN), .C2(n4064), .A(n4063), .B(n4062), 
        .ZN(n4065) );
  NAND3_X1 U4555 ( .A1(n4067), .A2(n4066), .A3(n4065), .ZN(U3240) );
  INV_X1 U4556 ( .A(n4747), .ZN(n4125) );
  NAND2_X1 U4557 ( .A1(n4125), .A2(n4432), .ZN(n4079) );
  AOI22_X1 U4558 ( .A1(n4737), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4078) );
  MUX2_X1 U4559 ( .A(REG1_REG_1__SCAN_IN), .B(n4764), .S(n4068), .Z(n4070) );
  NAND2_X1 U4560 ( .A1(n4070), .A2(n4069), .ZN(n4071) );
  NAND3_X1 U4561 ( .A1(n4744), .A2(n4072), .A3(n4071), .ZN(n4077) );
  OAI211_X1 U4562 ( .C1(n4075), .C2(n4074), .A(n4710), .B(n4073), .ZN(n4076)
         );
  NAND4_X1 U4563 ( .A1(n4079), .A2(n4078), .A3(n4077), .A4(n4076), .ZN(U3241)
         );
  AOI22_X1 U4564 ( .A1(n4737), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4090) );
  OAI211_X1 U4565 ( .C1(n4082), .C2(n4081), .A(n4710), .B(n4080), .ZN(n4086)
         );
  NAND2_X1 U4566 ( .A1(n4744), .A2(n4084), .ZN(n4085) );
  AND2_X1 U4567 ( .A1(n4086), .A2(n4085), .ZN(n4089) );
  OR2_X1 U4568 ( .A1(n4747), .A2(n4087), .ZN(n4088) );
  NAND4_X1 U4569 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(U3242)
         );
  INV_X1 U4570 ( .A(n4744), .ZN(n4721) );
  XNOR2_X1 U4571 ( .A(n4107), .B(n4092), .ZN(n4109) );
  INV_X1 U4572 ( .A(n4093), .ZN(n4430) );
  NAND2_X1 U4573 ( .A1(n4430), .A2(n4094), .ZN(n4096) );
  NAND2_X1 U4574 ( .A1(n4096), .A2(n4095), .ZN(n4108) );
  XNOR2_X1 U4575 ( .A(n4109), .B(n4108), .ZN(n4106) );
  AND2_X1 U4576 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4873) );
  NOR2_X1 U4577 ( .A1(n4098), .A2(n4097), .ZN(n4102) );
  NAND2_X1 U4578 ( .A1(n4107), .A2(REG2_REG_15__SCAN_IN), .ZN(n4118) );
  OR2_X1 U4579 ( .A1(n4107), .A2(REG2_REG_15__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U4580 ( .A1(n4118), .A2(n4099), .ZN(n4101) );
  INV_X1 U4581 ( .A(n4119), .ZN(n4100) );
  AOI211_X1 U4582 ( .C1(n4102), .C2(n4101), .A(n4100), .B(n4748), .ZN(n4103)
         );
  AOI211_X1 U4583 ( .C1(n4737), .C2(ADDR_REG_15__SCAN_IN), .A(n4873), .B(n4103), .ZN(n4105) );
  NAND2_X1 U4584 ( .A1(n4125), .A2(n4107), .ZN(n4104) );
  OAI211_X1 U4585 ( .C1(n4721), .C2(n4106), .A(n4105), .B(n4104), .ZN(U3255)
         );
  AOI22_X1 U4586 ( .A1(n4109), .A2(n4108), .B1(REG1_REG_15__SCAN_IN), .B2(
        n4107), .ZN(n4110) );
  INV_X1 U4587 ( .A(n4110), .ZN(n4112) );
  NOR2_X1 U4588 ( .A1(n4111), .A2(n4112), .ZN(n4113) );
  INV_X1 U4589 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4115) );
  NOR2_X1 U4590 ( .A1(n4130), .A2(REG1_REG_17__SCAN_IN), .ZN(n4140) );
  INV_X1 U4591 ( .A(n4140), .ZN(n4114) );
  OAI21_X1 U4592 ( .B1(n4117), .B2(n4115), .A(n4114), .ZN(n4116) );
  AOI21_X1 U4593 ( .B1(n2274), .B2(n4116), .A(n4139), .ZN(n4128) );
  XNOR2_X1 U4594 ( .A(n4117), .B(REG2_REG_17__SCAN_IN), .ZN(n4122) );
  NAND2_X1 U4595 ( .A1(n2280), .A2(n4893), .ZN(n4120) );
  NAND2_X1 U4596 ( .A1(n4121), .A2(n4122), .ZN(n4129) );
  AOI221_X1 U4597 ( .B1(n4122), .B2(n4129), .C1(n4121), .C2(n4129), .A(n4748), 
        .ZN(n4123) );
  AOI211_X1 U4598 ( .C1(n4737), .C2(ADDR_REG_17__SCAN_IN), .A(n4124), .B(n4123), .ZN(n4127) );
  NAND2_X1 U4599 ( .A1(n4125), .A2(n4130), .ZN(n4126) );
  OAI211_X1 U4600 ( .C1(n4128), .C2(n4721), .A(n4127), .B(n4126), .ZN(U3257)
         );
  OAI21_X1 U4601 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4130), .A(n4129), .ZN(n4134) );
  INV_X1 U4602 ( .A(n4144), .ZN(n4738) );
  NOR2_X1 U4603 ( .A1(n4738), .A2(n4131), .ZN(n4132) );
  AOI21_X1 U4604 ( .B1(n4131), .B2(n4738), .A(n4132), .ZN(n4133) );
  INV_X1 U4605 ( .A(n4136), .ZN(n4137) );
  NOR2_X1 U4606 ( .A1(n4140), .A2(n4139), .ZN(n4739) );
  XNOR2_X1 U4607 ( .A(n4144), .B(REG1_REG_18__SCAN_IN), .ZN(n4740) );
  XOR2_X1 U4608 ( .A(n4739), .B(n4740), .Z(n4141) );
  NAND2_X1 U4609 ( .A1(n4744), .A2(n4141), .ZN(n4142) );
  OAI211_X1 U4610 ( .C1(n4144), .C2(n4747), .A(n4143), .B(n4142), .ZN(U3258)
         );
  INV_X1 U4611 ( .A(n4145), .ZN(n4152) );
  OAI22_X1 U4612 ( .A1(n4147), .A2(n4859), .B1(n4146), .B2(n4863), .ZN(n4148)
         );
  OAI21_X1 U4613 ( .B1(n4149), .B2(n4148), .A(n4333), .ZN(n4151) );
  NAND2_X1 U4614 ( .A1(n4900), .A2(REG2_REG_29__SCAN_IN), .ZN(n4150) );
  OAI211_X1 U4615 ( .C1(n4152), .C2(n4335), .A(n4151), .B(n4150), .ZN(U3354)
         );
  XNOR2_X1 U4616 ( .A(n4153), .B(n4160), .ZN(n4344) );
  AOI22_X1 U4617 ( .A1(n4900), .A2(REG2_REG_28__SCAN_IN), .B1(n4154), .B2(
        n4847), .ZN(n4171) );
  INV_X1 U4618 ( .A(n4155), .ZN(n4156) );
  OAI211_X1 U4619 ( .C1(n4183), .C2(n4157), .A(n4156), .B(n4811), .ZN(n4342)
         );
  INV_X1 U4620 ( .A(n4158), .ZN(n4159) );
  NOR2_X1 U4621 ( .A1(n4172), .A2(n4159), .ZN(n4161) );
  XNOR2_X1 U4622 ( .A(n4161), .B(n4160), .ZN(n4167) );
  AOI22_X1 U4623 ( .A1(n4163), .A2(n4320), .B1(n4162), .B2(n4800), .ZN(n4164)
         );
  OAI21_X1 U4624 ( .B1(n4165), .B2(n4324), .A(n4164), .ZN(n4166) );
  OAI21_X1 U4625 ( .B1(n4168), .B2(n4342), .A(n4343), .ZN(n4169) );
  NAND2_X1 U4626 ( .A1(n4169), .A2(n4333), .ZN(n4170) );
  OAI211_X1 U4627 ( .C1(n4344), .C2(n4335), .A(n4171), .B(n4170), .ZN(U3262)
         );
  AOI21_X1 U4628 ( .B1(n4174), .B2(n4173), .A(n4172), .ZN(n4178) );
  AOI22_X1 U4629 ( .A1(n4175), .A2(n4320), .B1(n2744), .B2(n4800), .ZN(n4177)
         );
  NAND2_X1 U4630 ( .A1(n4219), .A2(n4801), .ZN(n4176) );
  OAI211_X1 U4631 ( .C1(n4178), .C2(n4300), .A(n4177), .B(n4176), .ZN(n4345)
         );
  AOI21_X1 U4632 ( .B1(n4179), .B2(n4847), .A(n4345), .ZN(n4190) );
  XNOR2_X1 U4633 ( .A(n4181), .B(n4180), .ZN(n4346) );
  INV_X1 U4634 ( .A(n4335), .ZN(n4182) );
  NAND2_X1 U4635 ( .A1(n4346), .A2(n4182), .ZN(n4189) );
  INV_X1 U4636 ( .A(n4350), .ZN(n4186) );
  INV_X1 U4637 ( .A(n4183), .ZN(n4184) );
  OAI21_X1 U4638 ( .B1(n4186), .B2(n4185), .A(n4184), .ZN(n4400) );
  INV_X1 U4639 ( .A(n4400), .ZN(n4187) );
  AOI22_X1 U4640 ( .A1(n4187), .A2(n4896), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4900), .ZN(n4188) );
  OAI211_X1 U4641 ( .C1(n4900), .C2(n4190), .A(n4189), .B(n4188), .ZN(U3263)
         );
  XNOR2_X1 U4642 ( .A(n4192), .B(n4191), .ZN(n4353) );
  INV_X1 U4643 ( .A(n4193), .ZN(n4194) );
  OR2_X1 U4644 ( .A1(n4195), .A2(n4194), .ZN(n4197) );
  XNOR2_X1 U4645 ( .A(n4197), .B(n4196), .ZN(n4203) );
  NAND2_X1 U4646 ( .A1(n4237), .A2(n4801), .ZN(n4200) );
  NAND2_X1 U4647 ( .A1(n4198), .A2(n4320), .ZN(n4199) );
  OAI211_X1 U4648 ( .C1(n4282), .C2(n4201), .A(n4200), .B(n4199), .ZN(n4202)
         );
  AOI21_X1 U4649 ( .B1(n4203), .B2(n4807), .A(n4202), .ZN(n4352) );
  INV_X1 U4650 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4205) );
  OAI22_X1 U4651 ( .A1(n4333), .A2(n4205), .B1(n4204), .B2(n4863), .ZN(n4206)
         );
  INV_X1 U4652 ( .A(n4206), .ZN(n4209) );
  NAND2_X1 U4653 ( .A1(n4225), .A2(n4207), .ZN(n4349) );
  NAND3_X1 U4654 ( .A1(n4350), .A2(n4896), .A3(n4349), .ZN(n4208) );
  OAI211_X1 U4655 ( .C1(n4352), .C2(n4900), .A(n4209), .B(n4208), .ZN(n4210)
         );
  INV_X1 U4656 ( .A(n4210), .ZN(n4211) );
  OAI21_X1 U4657 ( .B1(n4353), .B2(n4335), .A(n4211), .ZN(U3264) );
  XOR2_X1 U4658 ( .A(n4215), .B(n4212), .Z(n4355) );
  INV_X1 U4659 ( .A(n4355), .ZN(n4230) );
  NAND2_X1 U4660 ( .A1(n4214), .A2(n4213), .ZN(n4216) );
  XNOR2_X1 U4661 ( .A(n4216), .B(n4215), .ZN(n4217) );
  NAND2_X1 U4662 ( .A1(n4217), .A2(n4807), .ZN(n4221) );
  AOI22_X1 U4663 ( .A1(n4219), .A2(n4320), .B1(n4800), .B2(n4218), .ZN(n4220)
         );
  OAI211_X1 U4664 ( .C1(n4222), .C2(n4324), .A(n4221), .B(n4220), .ZN(n4354)
         );
  INV_X1 U4665 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4224) );
  OAI22_X1 U4666 ( .A1(n4333), .A2(n4224), .B1(n4223), .B2(n4863), .ZN(n4228)
         );
  OAI21_X1 U4667 ( .B1(n4243), .B2(n4226), .A(n4225), .ZN(n4405) );
  NOR2_X1 U4668 ( .A1(n4405), .A2(n4859), .ZN(n4227) );
  AOI211_X1 U4669 ( .C1(n4354), .C2(n4333), .A(n4228), .B(n4227), .ZN(n4229)
         );
  OAI21_X1 U4670 ( .B1(n4230), .B2(n4335), .A(n4229), .ZN(U3265) );
  XOR2_X1 U4671 ( .A(n4234), .B(n4231), .Z(n4359) );
  INV_X1 U4672 ( .A(n4359), .ZN(n4248) );
  NAND2_X1 U4673 ( .A1(n4233), .A2(n4232), .ZN(n4235) );
  XNOR2_X1 U4674 ( .A(n4235), .B(n4234), .ZN(n4240) );
  AOI22_X1 U4675 ( .A1(n4237), .A2(n4320), .B1(n4800), .B2(n4236), .ZN(n4239)
         );
  NAND2_X1 U4676 ( .A1(n4277), .A2(n4801), .ZN(n4238) );
  OAI211_X1 U4677 ( .C1(n4240), .C2(n4300), .A(n4239), .B(n4238), .ZN(n4358)
         );
  NOR2_X1 U4678 ( .A1(n4264), .A2(n4241), .ZN(n4242) );
  OR2_X1 U4679 ( .A1(n4243), .A2(n4242), .ZN(n4409) );
  AOI22_X1 U4680 ( .A1(n4900), .A2(REG2_REG_24__SCAN_IN), .B1(n4244), .B2(
        n4847), .ZN(n4245) );
  OAI21_X1 U4681 ( .B1(n4409), .B2(n4859), .A(n4245), .ZN(n4246) );
  AOI21_X1 U4682 ( .B1(n4358), .B2(n4333), .A(n4246), .ZN(n4247) );
  OAI21_X1 U4683 ( .B1(n4248), .B2(n4335), .A(n4247), .ZN(U3266) );
  OAI21_X1 U4684 ( .B1(n4293), .B2(n4250), .A(n4249), .ZN(n4274) );
  AND2_X1 U4685 ( .A1(n4274), .A2(n4275), .ZN(n4272) );
  NOR2_X1 U4686 ( .A1(n4272), .A2(n4251), .ZN(n4252) );
  XNOR2_X1 U4687 ( .A(n4252), .B(n4257), .ZN(n4363) );
  INV_X1 U4688 ( .A(n4363), .ZN(n4271) );
  INV_X1 U4689 ( .A(n4253), .ZN(n4254) );
  AOI21_X1 U4690 ( .B1(n4295), .B2(n4255), .A(n4254), .ZN(n4276) );
  OAI21_X1 U4691 ( .B1(n4276), .B2(n4275), .A(n4256), .ZN(n4258) );
  XNOR2_X1 U4692 ( .A(n4258), .B(n4257), .ZN(n4263) );
  AOI22_X1 U4693 ( .A1(n4297), .A2(n4801), .B1(n4800), .B2(n4259), .ZN(n4262)
         );
  NAND2_X1 U4694 ( .A1(n4260), .A2(n4320), .ZN(n4261) );
  OAI211_X1 U4695 ( .C1(n4263), .C2(n4300), .A(n4262), .B(n4261), .ZN(n4362)
         );
  INV_X1 U4696 ( .A(n4264), .ZN(n4265) );
  OAI21_X1 U4697 ( .B1(n2304), .B2(n4266), .A(n4265), .ZN(n4413) );
  AOI22_X1 U4698 ( .A1(n4900), .A2(REG2_REG_23__SCAN_IN), .B1(n4267), .B2(
        n4847), .ZN(n4268) );
  OAI21_X1 U4699 ( .B1(n4413), .B2(n4859), .A(n4268), .ZN(n4269) );
  AOI21_X1 U4700 ( .B1(n4362), .B2(n4333), .A(n4269), .ZN(n4270) );
  OAI21_X1 U4701 ( .B1(n4271), .B2(n4335), .A(n4270), .ZN(U3267) );
  INV_X1 U4702 ( .A(n4272), .ZN(n4273) );
  OAI21_X1 U4703 ( .B1(n4274), .B2(n4275), .A(n4273), .ZN(n4370) );
  XNOR2_X1 U4704 ( .A(n4276), .B(n4275), .ZN(n4284) );
  NAND2_X1 U4705 ( .A1(n4277), .A2(n4320), .ZN(n4280) );
  NAND2_X1 U4706 ( .A1(n4278), .A2(n4801), .ZN(n4279) );
  OAI211_X1 U4707 ( .C1(n4282), .C2(n4281), .A(n4280), .B(n4279), .ZN(n4283)
         );
  AOI21_X1 U4708 ( .B1(n4284), .B2(n4807), .A(n4283), .ZN(n4369) );
  INV_X1 U4709 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4286) );
  OAI22_X1 U4710 ( .A1(n4333), .A2(n4286), .B1(n4285), .B2(n4863), .ZN(n4287)
         );
  INV_X1 U4711 ( .A(n4287), .ZN(n4290) );
  NAND2_X1 U4712 ( .A1(n4302), .A2(n4288), .ZN(n4366) );
  NAND3_X1 U4713 ( .A1(n4367), .A2(n4896), .A3(n4366), .ZN(n4289) );
  OAI211_X1 U4714 ( .C1(n4369), .C2(n4900), .A(n4290), .B(n4289), .ZN(n4291)
         );
  INV_X1 U4715 ( .A(n4291), .ZN(n4292) );
  OAI21_X1 U4716 ( .B1(n4370), .B2(n4335), .A(n4292), .ZN(U3268) );
  XNOR2_X1 U4717 ( .A(n4293), .B(n4294), .ZN(n4372) );
  INV_X1 U4718 ( .A(n4372), .ZN(n4310) );
  XNOR2_X1 U4719 ( .A(n4295), .B(n4294), .ZN(n4301) );
  AOI22_X1 U4720 ( .A1(n4297), .A2(n4320), .B1(n4800), .B2(n4296), .ZN(n4299)
         );
  NAND2_X1 U4721 ( .A1(n4321), .A2(n4801), .ZN(n4298) );
  OAI211_X1 U4722 ( .C1(n4301), .C2(n4300), .A(n4299), .B(n4298), .ZN(n4371)
         );
  OAI21_X1 U4723 ( .B1(n4304), .B2(n4303), .A(n4302), .ZN(n4418) );
  NOR2_X1 U4724 ( .A1(n4418), .A2(n4859), .ZN(n4308) );
  INV_X1 U4725 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4306) );
  OAI22_X1 U4726 ( .A1(n4333), .A2(n4306), .B1(n4305), .B2(n4863), .ZN(n4307)
         );
  AOI211_X1 U4727 ( .C1(n4371), .C2(n4333), .A(n4308), .B(n4307), .ZN(n4309)
         );
  OAI21_X1 U4728 ( .B1(n4310), .B2(n4335), .A(n4309), .ZN(U3269) );
  XNOR2_X1 U4729 ( .A(n4311), .B(n4316), .ZN(n4381) );
  INV_X1 U4730 ( .A(n4381), .ZN(n4336) );
  INV_X1 U4731 ( .A(n4312), .ZN(n4314) );
  OAI21_X1 U4732 ( .B1(n4315), .B2(n4314), .A(n4313), .ZN(n4317) );
  XNOR2_X1 U4733 ( .A(n4317), .B(n4316), .ZN(n4318) );
  NAND2_X1 U4734 ( .A1(n4318), .A2(n4807), .ZN(n4323) );
  AOI22_X1 U4735 ( .A1(n4321), .A2(n4320), .B1(n4800), .B2(n4319), .ZN(n4322)
         );
  OAI211_X1 U4736 ( .C1(n4325), .C2(n4324), .A(n4323), .B(n4322), .ZN(n4380)
         );
  OAI21_X1 U4737 ( .B1(n4328), .B2(n4327), .A(n4326), .ZN(n4424) );
  NOR2_X1 U4738 ( .A1(n4424), .A2(n4859), .ZN(n4332) );
  INV_X1 U4739 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4330) );
  OAI22_X1 U4740 ( .A1(n4333), .A2(n4330), .B1(n4329), .B2(n4863), .ZN(n4331)
         );
  AOI211_X1 U4741 ( .C1(n4380), .C2(n4333), .A(n4332), .B(n4331), .ZN(n4334)
         );
  OAI21_X1 U4742 ( .B1(n4336), .B2(n4335), .A(n4334), .ZN(U3271) );
  AOI21_X1 U4743 ( .B1(n4339), .B2(n2273), .A(n4337), .ZN(n4897) );
  INV_X1 U4744 ( .A(n4897), .ZN(n4395) );
  INV_X1 U4745 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4340) );
  AOI21_X1 U4746 ( .B1(n4339), .B2(n4800), .A(n4338), .ZN(n4899) );
  MUX2_X1 U4747 ( .A(n4340), .B(n4899), .S(n4831), .Z(n4341) );
  OAI21_X1 U4748 ( .B1(n4395), .B2(n4383), .A(n4341), .ZN(U3548) );
  INV_X1 U4749 ( .A(n4826), .ZN(n4391) );
  OAI211_X1 U4750 ( .C1(n4344), .C2(n4391), .A(n4343), .B(n4342), .ZN(n4396)
         );
  MUX2_X1 U4751 ( .A(REG1_REG_28__SCAN_IN), .B(n4396), .S(n4831), .Z(U3546) );
  INV_X1 U4752 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4347) );
  AOI21_X1 U4753 ( .B1(n4346), .B2(n4826), .A(n4345), .ZN(n4397) );
  MUX2_X1 U4754 ( .A(n4347), .B(n4397), .S(n4831), .Z(n4348) );
  OAI21_X1 U4755 ( .B1(n4383), .B2(n4400), .A(n4348), .ZN(U3545) );
  NAND3_X1 U4756 ( .A1(n4350), .A2(n4811), .A3(n4349), .ZN(n4351) );
  OAI211_X1 U4757 ( .C1(n4353), .C2(n4391), .A(n4352), .B(n4351), .ZN(n4401)
         );
  MUX2_X1 U4758 ( .A(REG1_REG_26__SCAN_IN), .B(n4401), .S(n4831), .Z(U3544) );
  INV_X1 U4759 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4356) );
  AOI21_X1 U4760 ( .B1(n4355), .B2(n4826), .A(n4354), .ZN(n4402) );
  MUX2_X1 U4761 ( .A(n4356), .B(n4402), .S(n4831), .Z(n4357) );
  OAI21_X1 U4762 ( .B1(n4383), .B2(n4405), .A(n4357), .ZN(U3543) );
  INV_X1 U4763 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4360) );
  AOI21_X1 U4764 ( .B1(n4359), .B2(n4826), .A(n4358), .ZN(n4406) );
  MUX2_X1 U4765 ( .A(n4360), .B(n4406), .S(n4831), .Z(n4361) );
  OAI21_X1 U4766 ( .B1(n4383), .B2(n4409), .A(n4361), .ZN(U3542) );
  INV_X1 U4767 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4364) );
  AOI21_X1 U4768 ( .B1(n4363), .B2(n4826), .A(n4362), .ZN(n4410) );
  MUX2_X1 U4769 ( .A(n4364), .B(n4410), .S(n4831), .Z(n4365) );
  OAI21_X1 U4770 ( .B1(n4383), .B2(n4413), .A(n4365), .ZN(U3541) );
  NAND3_X1 U4771 ( .A1(n4367), .A2(n4811), .A3(n4366), .ZN(n4368) );
  OAI211_X1 U4772 ( .C1(n4370), .C2(n4391), .A(n4369), .B(n4368), .ZN(n4414)
         );
  MUX2_X1 U4773 ( .A(REG1_REG_22__SCAN_IN), .B(n4414), .S(n4831), .Z(U3540) );
  INV_X1 U4774 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4373) );
  AOI21_X1 U4775 ( .B1(n4372), .B2(n4826), .A(n4371), .ZN(n4415) );
  MUX2_X1 U4776 ( .A(n4373), .B(n4415), .S(n4831), .Z(n4374) );
  OAI21_X1 U4777 ( .B1(n4383), .B2(n4418), .A(n4374), .ZN(U3539) );
  NAND3_X1 U4778 ( .A1(n4376), .A2(n4811), .A3(n4375), .ZN(n4377) );
  OAI211_X1 U4779 ( .C1(n4379), .C2(n4760), .A(n4378), .B(n4377), .ZN(n4419)
         );
  MUX2_X1 U4780 ( .A(REG1_REG_20__SCAN_IN), .B(n4419), .S(n4831), .Z(U3538) );
  INV_X1 U4781 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4741) );
  AOI21_X1 U4782 ( .B1(n4381), .B2(n4826), .A(n4380), .ZN(n4420) );
  MUX2_X1 U4783 ( .A(n4741), .B(n4420), .S(n4831), .Z(n4382) );
  OAI21_X1 U4784 ( .B1(n4383), .B2(n4424), .A(n4382), .ZN(U3537) );
  OAI211_X1 U4785 ( .C1(n4386), .C2(n4391), .A(n4385), .B(n4384), .ZN(n4425)
         );
  MUX2_X1 U4786 ( .A(REG1_REG_18__SCAN_IN), .B(n4425), .S(n4831), .Z(U3536) );
  NAND3_X1 U4787 ( .A1(n4388), .A2(n4811), .A3(n4387), .ZN(n4389) );
  OAI211_X1 U4788 ( .C1(n4392), .C2(n4391), .A(n4390), .B(n4389), .ZN(n4426)
         );
  MUX2_X1 U4789 ( .A(REG1_REG_16__SCAN_IN), .B(n4426), .S(n4831), .Z(U3534) );
  INV_X1 U4790 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4393) );
  MUX2_X1 U4791 ( .A(n4393), .B(n4899), .S(n4835), .Z(n4394) );
  OAI21_X1 U4792 ( .B1(n4395), .B2(n4423), .A(n4394), .ZN(U3516) );
  MUX2_X1 U4793 ( .A(REG0_REG_28__SCAN_IN), .B(n4396), .S(n4835), .Z(U3514) );
  INV_X1 U4794 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4398) );
  MUX2_X1 U4795 ( .A(n4398), .B(n4397), .S(n4835), .Z(n4399) );
  OAI21_X1 U4796 ( .B1(n4400), .B2(n4423), .A(n4399), .ZN(U3513) );
  MUX2_X1 U4797 ( .A(REG0_REG_26__SCAN_IN), .B(n4401), .S(n4835), .Z(U3512) );
  INV_X1 U4798 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4403) );
  MUX2_X1 U4799 ( .A(n4403), .B(n4402), .S(n4835), .Z(n4404) );
  OAI21_X1 U4800 ( .B1(n4405), .B2(n4423), .A(n4404), .ZN(U3511) );
  INV_X1 U4801 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4407) );
  MUX2_X1 U4802 ( .A(n4407), .B(n4406), .S(n4835), .Z(n4408) );
  OAI21_X1 U4803 ( .B1(n4409), .B2(n4423), .A(n4408), .ZN(U3510) );
  INV_X1 U4804 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4411) );
  MUX2_X1 U4805 ( .A(n4411), .B(n4410), .S(n4835), .Z(n4412) );
  OAI21_X1 U4806 ( .B1(n4413), .B2(n4423), .A(n4412), .ZN(U3509) );
  MUX2_X1 U4807 ( .A(REG0_REG_22__SCAN_IN), .B(n4414), .S(n4835), .Z(U3508) );
  INV_X1 U4808 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4416) );
  MUX2_X1 U4809 ( .A(n4416), .B(n4415), .S(n4835), .Z(n4417) );
  OAI21_X1 U4810 ( .B1(n4418), .B2(n4423), .A(n4417), .ZN(U3507) );
  MUX2_X1 U4811 ( .A(REG0_REG_20__SCAN_IN), .B(n4419), .S(n4835), .Z(U3506) );
  INV_X1 U4812 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4421) );
  MUX2_X1 U4813 ( .A(n4421), .B(n4420), .S(n4835), .Z(n4422) );
  OAI21_X1 U4814 ( .B1(n4424), .B2(n4423), .A(n4422), .ZN(U3505) );
  MUX2_X1 U4815 ( .A(REG0_REG_18__SCAN_IN), .B(n4425), .S(n4835), .Z(U3503) );
  MUX2_X1 U4816 ( .A(REG0_REG_16__SCAN_IN), .B(n4426), .S(n4835), .Z(U3499) );
  MUX2_X1 U4817 ( .A(n4427), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4818 ( .A(n4428), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4819 ( .A(DATAI_25_), .B(n4429), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4820 ( .A(DATAI_24_), .B(n2838), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4821 ( .A(n4738), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U4822 ( .A(DATAI_14_), .B(n4430), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U4823 ( .A(n4682), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U4824 ( .A(DATAI_3_), .B(n4431), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4825 ( .A(n2349), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4826 ( .A(n4432), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U4827 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U4828 ( .A(DATAI_23_), .ZN(n4552) );
  OAI21_X1 U4829 ( .B1(STATE_REG_SCAN_IN), .B2(n4552), .A(n4433), .ZN(U3329)
         );
  AND2_X1 U4830 ( .A1(D_REG_2__SCAN_IN), .A2(n4434), .ZN(U3320) );
  AND2_X1 U4831 ( .A1(D_REG_3__SCAN_IN), .A2(n4434), .ZN(U3319) );
  AND2_X1 U4832 ( .A1(D_REG_4__SCAN_IN), .A2(n4434), .ZN(U3318) );
  AND2_X1 U4833 ( .A1(D_REG_5__SCAN_IN), .A2(n4434), .ZN(U3317) );
  AND2_X1 U4834 ( .A1(D_REG_6__SCAN_IN), .A2(n4434), .ZN(U3316) );
  AND2_X1 U4835 ( .A1(D_REG_7__SCAN_IN), .A2(n4434), .ZN(U3315) );
  AND2_X1 U4836 ( .A1(D_REG_8__SCAN_IN), .A2(n4434), .ZN(U3314) );
  AND2_X1 U4837 ( .A1(D_REG_9__SCAN_IN), .A2(n4434), .ZN(U3313) );
  AND2_X1 U4838 ( .A1(D_REG_10__SCAN_IN), .A2(n4434), .ZN(U3312) );
  AND2_X1 U4839 ( .A1(D_REG_11__SCAN_IN), .A2(n4434), .ZN(U3311) );
  AND2_X1 U4840 ( .A1(D_REG_12__SCAN_IN), .A2(n4434), .ZN(U3310) );
  AND2_X1 U4841 ( .A1(D_REG_13__SCAN_IN), .A2(n4434), .ZN(U3309) );
  AND2_X1 U4842 ( .A1(D_REG_14__SCAN_IN), .A2(n4434), .ZN(U3308) );
  AND2_X1 U4843 ( .A1(D_REG_15__SCAN_IN), .A2(n4434), .ZN(U3307) );
  AND2_X1 U4844 ( .A1(D_REG_16__SCAN_IN), .A2(n4434), .ZN(U3306) );
  AND2_X1 U4845 ( .A1(D_REG_17__SCAN_IN), .A2(n4434), .ZN(U3305) );
  AND2_X1 U4846 ( .A1(D_REG_18__SCAN_IN), .A2(n4434), .ZN(U3304) );
  AND2_X1 U4847 ( .A1(D_REG_19__SCAN_IN), .A2(n4434), .ZN(U3303) );
  AND2_X1 U4848 ( .A1(D_REG_20__SCAN_IN), .A2(n4434), .ZN(U3302) );
  AND2_X1 U4849 ( .A1(D_REG_21__SCAN_IN), .A2(n4434), .ZN(U3301) );
  AND2_X1 U4850 ( .A1(D_REG_22__SCAN_IN), .A2(n4434), .ZN(U3300) );
  AND2_X1 U4851 ( .A1(D_REG_23__SCAN_IN), .A2(n4434), .ZN(U3299) );
  AND2_X1 U4852 ( .A1(D_REG_24__SCAN_IN), .A2(n4434), .ZN(U3298) );
  AND2_X1 U4853 ( .A1(D_REG_26__SCAN_IN), .A2(n4434), .ZN(U3296) );
  AND2_X1 U4854 ( .A1(D_REG_27__SCAN_IN), .A2(n4434), .ZN(U3295) );
  AND2_X1 U4855 ( .A1(D_REG_28__SCAN_IN), .A2(n4434), .ZN(U3294) );
  AND2_X1 U4856 ( .A1(D_REG_29__SCAN_IN), .A2(n4434), .ZN(U3293) );
  AND2_X1 U4857 ( .A1(D_REG_30__SCAN_IN), .A2(n4434), .ZN(U3292) );
  AND2_X1 U4858 ( .A1(D_REG_31__SCAN_IN), .A2(n4434), .ZN(U3291) );
  NAND2_X1 U4859 ( .A1(n4434), .A2(D_REG_25__SCAN_IN), .ZN(n4630) );
  INV_X1 U4860 ( .A(keyinput_54), .ZN(n4508) );
  OAI22_X1 U4861 ( .A1(n4436), .A2(keyinput_49), .B1(keyinput_48), .B2(
        REG3_REG_17__SCAN_IN), .ZN(n4435) );
  AOI221_X1 U4862 ( .B1(n4436), .B2(keyinput_49), .C1(REG3_REG_17__SCAN_IN), 
        .C2(keyinput_48), .A(n4435), .ZN(n4506) );
  XOR2_X1 U4863 ( .A(n4598), .B(keyinput_45), .Z(n4500) );
  INV_X1 U4864 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4531) );
  AOI22_X1 U4865 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_34), .B1(n4531), 
        .B2(keyinput_35), .ZN(n4437) );
  OAI221_X1 U4866 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_34), .C1(n4531), 
        .C2(keyinput_35), .A(n4437), .ZN(n4487) );
  INV_X1 U4867 ( .A(DATAI_0_), .ZN(n4439) );
  AOI22_X1 U4868 ( .A1(U3149), .A2(keyinput_32), .B1(keyinput_31), .B2(n4439), 
        .ZN(n4438) );
  OAI221_X1 U4869 ( .B1(U3149), .B2(keyinput_32), .C1(n4439), .C2(keyinput_31), 
        .A(n4438), .ZN(n4481) );
  OAI22_X1 U4870 ( .A1(n2603), .A2(keyinput_20), .B1(keyinput_19), .B2(
        DATAI_12_), .ZN(n4440) );
  AOI221_X1 U4871 ( .B1(n2603), .B2(keyinput_20), .C1(DATAI_12_), .C2(
        keyinput_19), .A(n4440), .ZN(n4471) );
  OAI22_X1 U4872 ( .A1(DATAI_25_), .A2(keyinput_6), .B1(DATAI_24_), .B2(
        keyinput_7), .ZN(n4441) );
  AOI221_X1 U4873 ( .B1(DATAI_25_), .B2(keyinput_6), .C1(keyinput_7), .C2(
        DATAI_24_), .A(n4441), .ZN(n4451) );
  INV_X1 U4874 ( .A(DATAI_26_), .ZN(n4546) );
  INV_X1 U4875 ( .A(keyinput_5), .ZN(n4449) );
  OAI22_X1 U4876 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        DATAI_31_), .ZN(n4442) );
  AOI221_X1 U4877 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n4442), .ZN(n4446) );
  INV_X1 U4878 ( .A(DATAI_28_), .ZN(n4894) );
  AOI22_X1 U4879 ( .A1(n4894), .A2(keyinput_3), .B1(n4444), .B2(keyinput_2), 
        .ZN(n4443) );
  OAI221_X1 U4880 ( .B1(n4894), .B2(keyinput_3), .C1(n4444), .C2(keyinput_2), 
        .A(n4443), .ZN(n4445) );
  AOI211_X1 U4881 ( .C1(DATAI_27_), .C2(keyinput_4), .A(n4446), .B(n4445), 
        .ZN(n4447) );
  OAI21_X1 U4882 ( .B1(DATAI_27_), .B2(keyinput_4), .A(n4447), .ZN(n4448) );
  OAI221_X1 U4883 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(n4546), .C2(n4449), 
        .A(n4448), .ZN(n4450) );
  AOI22_X1 U4884 ( .A1(n4451), .A2(n4450), .B1(keyinput_10), .B2(n4553), .ZN(
        n4452) );
  OAI21_X1 U4885 ( .B1(keyinput_10), .B2(n4553), .A(n4452), .ZN(n4465) );
  AOI22_X1 U4886 ( .A1(DATAI_22_), .A2(keyinput_9), .B1(DATAI_23_), .B2(
        keyinput_8), .ZN(n4453) );
  OAI221_X1 U4887 ( .B1(DATAI_22_), .B2(keyinput_9), .C1(DATAI_23_), .C2(
        keyinput_8), .A(n4453), .ZN(n4464) );
  AOI22_X1 U4888 ( .A1(n4892), .A2(keyinput_15), .B1(n2692), .B2(keyinput_12), 
        .ZN(n4454) );
  OAI221_X1 U4889 ( .B1(n4892), .B2(keyinput_15), .C1(n2692), .C2(keyinput_12), 
        .A(n4454), .ZN(n4462) );
  AOI22_X1 U4890 ( .A1(n2676), .A2(keyinput_14), .B1(n4456), .B2(keyinput_13), 
        .ZN(n4455) );
  OAI221_X1 U4891 ( .B1(n2676), .B2(keyinput_14), .C1(n4456), .C2(keyinput_13), 
        .A(n4455), .ZN(n4461) );
  AOI22_X1 U4892 ( .A1(DATAI_15_), .A2(keyinput_16), .B1(DATAI_20_), .B2(
        keyinput_11), .ZN(n4457) );
  OAI221_X1 U4893 ( .B1(DATAI_15_), .B2(keyinput_16), .C1(DATAI_20_), .C2(
        keyinput_11), .A(n4457), .ZN(n4460) );
  AOI22_X1 U4894 ( .A1(DATAI_13_), .A2(keyinput_18), .B1(DATAI_14_), .B2(
        keyinput_17), .ZN(n4458) );
  OAI221_X1 U4895 ( .B1(DATAI_13_), .B2(keyinput_18), .C1(DATAI_14_), .C2(
        keyinput_17), .A(n4458), .ZN(n4459) );
  NOR4_X1 U4896 ( .A1(n4462), .A2(n4461), .A3(n4460), .A4(n4459), .ZN(n4463)
         );
  OAI21_X1 U4897 ( .B1(n4465), .B2(n4464), .A(n4463), .ZN(n4470) );
  INV_X1 U4898 ( .A(DATAI_10_), .ZN(n4566) );
  AOI22_X1 U4899 ( .A1(DATAI_7_), .A2(keyinput_24), .B1(n4566), .B2(
        keyinput_21), .ZN(n4466) );
  OAI221_X1 U4900 ( .B1(DATAI_7_), .B2(keyinput_24), .C1(n4566), .C2(
        keyinput_21), .A(n4466), .ZN(n4469) );
  INV_X1 U4901 ( .A(DATAI_6_), .ZN(n4786) );
  INV_X1 U4902 ( .A(DATAI_9_), .ZN(n4845) );
  AOI22_X1 U4903 ( .A1(n4786), .A2(keyinput_25), .B1(n4845), .B2(keyinput_22), 
        .ZN(n4467) );
  OAI221_X1 U4904 ( .B1(n4786), .B2(keyinput_25), .C1(n4845), .C2(keyinput_22), 
        .A(n4467), .ZN(n4468) );
  AOI211_X1 U4905 ( .C1(n4471), .C2(n4470), .A(n4469), .B(n4468), .ZN(n4479)
         );
  OAI22_X1 U4906 ( .A1(n4836), .A2(keyinput_23), .B1(keyinput_26), .B2(
        DATAI_5_), .ZN(n4472) );
  AOI221_X1 U4907 ( .B1(n4836), .B2(keyinput_23), .C1(DATAI_5_), .C2(
        keyinput_26), .A(n4472), .ZN(n4478) );
  INV_X1 U4908 ( .A(DATAI_3_), .ZN(n4572) );
  AOI22_X1 U4909 ( .A1(DATAI_4_), .A2(keyinput_27), .B1(n4572), .B2(
        keyinput_28), .ZN(n4473) );
  OAI221_X1 U4910 ( .B1(DATAI_4_), .B2(keyinput_27), .C1(n4572), .C2(
        keyinput_28), .A(n4473), .ZN(n4477) );
  XOR2_X1 U4911 ( .A(n2489), .B(keyinput_30), .Z(n4475) );
  XNOR2_X1 U4912 ( .A(DATAI_2_), .B(keyinput_29), .ZN(n4474) );
  NAND2_X1 U4913 ( .A1(n4475), .A2(n4474), .ZN(n4476) );
  AOI211_X1 U4914 ( .C1(n4479), .C2(n4478), .A(n4477), .B(n4476), .ZN(n4480)
         );
  OAI22_X1 U4915 ( .A1(keyinput_33), .A2(n2549), .B1(n4481), .B2(n4480), .ZN(
        n4482) );
  AOI21_X1 U4916 ( .B1(keyinput_33), .B2(n2549), .A(n4482), .ZN(n4486) );
  XNOR2_X1 U4917 ( .A(keyinput_37), .B(n4582), .ZN(n4485) );
  OAI22_X1 U4918 ( .A1(n4772), .A2(keyinput_38), .B1(keyinput_36), .B2(
        REG3_REG_23__SCAN_IN), .ZN(n4483) );
  AOI221_X1 U4919 ( .B1(n4772), .B2(keyinput_38), .C1(REG3_REG_23__SCAN_IN), 
        .C2(keyinput_36), .A(n4483), .ZN(n4484) );
  OAI211_X1 U4920 ( .C1(n4487), .C2(n4486), .A(n4485), .B(n4484), .ZN(n4496)
         );
  OAI22_X1 U4921 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_39), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_40), .ZN(n4488) );
  AOI221_X1 U4922 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_39), .C1(
        keyinput_40), .C2(REG3_REG_28__SCAN_IN), .A(n4488), .ZN(n4495) );
  AOI22_X1 U4923 ( .A1(n4490), .A2(keyinput_44), .B1(keyinput_43), .B2(n2705), 
        .ZN(n4489) );
  OAI221_X1 U4924 ( .B1(n4490), .B2(keyinput_44), .C1(n2705), .C2(keyinput_43), 
        .A(n4489), .ZN(n4494) );
  XNOR2_X1 U4925 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_41), .ZN(n4492) );
  XNOR2_X1 U4926 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .ZN(n4491) );
  NAND2_X1 U4927 ( .A1(n4492), .A2(n4491), .ZN(n4493) );
  AOI211_X1 U4928 ( .C1(n4496), .C2(n4495), .A(n4494), .B(n4493), .ZN(n4499)
         );
  OAI22_X1 U4929 ( .A1(n2527), .A2(keyinput_47), .B1(keyinput_46), .B2(
        REG3_REG_16__SCAN_IN), .ZN(n4497) );
  AOI221_X1 U4930 ( .B1(n2527), .B2(keyinput_47), .C1(REG3_REG_16__SCAN_IN), 
        .C2(keyinput_46), .A(n4497), .ZN(n4498) );
  OAI21_X1 U4931 ( .B1(n4500), .B2(n4499), .A(n4498), .ZN(n4505) );
  AOI22_X1 U4932 ( .A1(n2570), .A2(keyinput_51), .B1(keyinput_53), .B2(n4605), 
        .ZN(n4501) );
  OAI221_X1 U4933 ( .B1(n2570), .B2(keyinput_51), .C1(n4605), .C2(keyinput_53), 
        .A(n4501), .ZN(n4504) );
  AOI22_X1 U4934 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_52), .B1(
        REG3_REG_4__SCAN_IN), .B2(keyinput_50), .ZN(n4502) );
  OAI221_X1 U4935 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_52), .C1(
        REG3_REG_4__SCAN_IN), .C2(keyinput_50), .A(n4502), .ZN(n4503) );
  AOI211_X1 U4936 ( .C1(n4506), .C2(n4505), .A(n4504), .B(n4503), .ZN(n4507)
         );
  AOI221_X1 U4937 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_54), .C1(n4609), 
        .C2(n4508), .A(n4507), .ZN(n4511) );
  INV_X1 U4938 ( .A(keyinput_55), .ZN(n4509) );
  MUX2_X1 U4939 ( .A(n4509), .B(keyinput_55), .S(IR_REG_0__SCAN_IN), .Z(n4510)
         );
  NOR2_X1 U4940 ( .A1(n4511), .A2(n4510), .ZN(n4514) );
  INV_X1 U4941 ( .A(keyinput_56), .ZN(n4512) );
  MUX2_X1 U4942 ( .A(keyinput_56), .B(n4512), .S(IR_REG_1__SCAN_IN), .Z(n4513)
         );
  NOR2_X1 U4943 ( .A1(n4514), .A2(n4513), .ZN(n4520) );
  AOI22_X1 U4944 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_58), .B1(n4617), .B2(
        keyinput_57), .ZN(n4515) );
  OAI221_X1 U4945 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_58), .C1(n4617), .C2(
        keyinput_57), .A(n4515), .ZN(n4519) );
  OAI22_X1 U4946 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_61), .B1(keyinput_59), 
        .B2(IR_REG_4__SCAN_IN), .ZN(n4516) );
  AOI221_X1 U4947 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_61), .C1(
        IR_REG_4__SCAN_IN), .C2(keyinput_59), .A(n4516), .ZN(n4518) );
  XNOR2_X1 U4948 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n4517) );
  OAI211_X1 U4949 ( .C1(n4520), .C2(n4519), .A(n4518), .B(n4517), .ZN(n4523)
         );
  XNOR2_X1 U4950 ( .A(n4521), .B(keyinput_62), .ZN(n4522) );
  NAND2_X1 U4951 ( .A1(n4523), .A2(n4522), .ZN(n4526) );
  INV_X1 U4952 ( .A(keyinput_63), .ZN(n4524) );
  MUX2_X1 U4953 ( .A(keyinput_63), .B(n4524), .S(IR_REG_8__SCAN_IN), .Z(n4525)
         );
  NAND2_X1 U4954 ( .A1(n4526), .A2(n4525), .ZN(n4627) );
  AOI22_X1 U4955 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_113), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput_112), .ZN(n4527) );
  OAI221_X1 U4956 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_113), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput_112), .A(n4527), .ZN(n4603) );
  OAI22_X1 U4957 ( .A1(n4529), .A2(keyinput_110), .B1(keyinput_111), .B2(
        REG3_REG_5__SCAN_IN), .ZN(n4528) );
  AOI221_X1 U4958 ( .B1(n4529), .B2(keyinput_110), .C1(REG3_REG_5__SCAN_IN), 
        .C2(keyinput_111), .A(n4528), .ZN(n4602) );
  INV_X1 U4959 ( .A(keyinput_109), .ZN(n4597) );
  OAI22_X1 U4960 ( .A1(n4531), .A2(keyinput_99), .B1(REG3_REG_27__SCAN_IN), 
        .B2(keyinput_98), .ZN(n4530) );
  AOI221_X1 U4961 ( .B1(n4531), .B2(keyinput_99), .C1(keyinput_98), .C2(
        REG3_REG_27__SCAN_IN), .A(n4530), .ZN(n4586) );
  OAI22_X1 U4962 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_96), .B1(keyinput_95), 
        .B2(DATAI_0_), .ZN(n4532) );
  AOI221_X1 U4963 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_96), .C1(DATAI_0_), 
        .C2(keyinput_95), .A(n4532), .ZN(n4579) );
  INV_X1 U4964 ( .A(DATAI_7_), .ZN(n4794) );
  AOI22_X1 U4965 ( .A1(n2537), .A2(keyinput_90), .B1(n4794), .B2(keyinput_88), 
        .ZN(n4533) );
  OAI221_X1 U4966 ( .B1(n2537), .B2(keyinput_90), .C1(n4794), .C2(keyinput_88), 
        .A(n4533), .ZN(n4577) );
  AOI22_X1 U4967 ( .A1(DATAI_13_), .A2(keyinput_82), .B1(n4535), .B2(
        keyinput_81), .ZN(n4534) );
  OAI221_X1 U4968 ( .B1(DATAI_13_), .B2(keyinput_82), .C1(n4535), .C2(
        keyinput_81), .A(n4534), .ZN(n4562) );
  AOI22_X1 U4969 ( .A1(n4537), .A2(keyinput_80), .B1(n2692), .B2(keyinput_76), 
        .ZN(n4536) );
  OAI221_X1 U4970 ( .B1(n4537), .B2(keyinput_80), .C1(n2692), .C2(keyinput_76), 
        .A(n4536), .ZN(n4561) );
  AOI22_X1 U4971 ( .A1(DATAI_24_), .A2(keyinput_71), .B1(DATAI_25_), .B2(
        keyinput_70), .ZN(n4538) );
  OAI221_X1 U4972 ( .B1(DATAI_24_), .B2(keyinput_71), .C1(DATAI_25_), .C2(
        keyinput_70), .A(n4538), .ZN(n4550) );
  INV_X1 U4973 ( .A(keyinput_69), .ZN(n4547) );
  XOR2_X1 U4974 ( .A(DATAI_29_), .B(keyinput_66), .Z(n4544) );
  OAI22_X1 U4975 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        DATAI_31_), .ZN(n4539) );
  AOI221_X1 U4976 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n4539), .ZN(n4543) );
  AOI22_X1 U4977 ( .A1(n4541), .A2(keyinput_68), .B1(n4894), .B2(keyinput_67), 
        .ZN(n4540) );
  OAI221_X1 U4978 ( .B1(n4541), .B2(keyinput_68), .C1(n4894), .C2(keyinput_67), 
        .A(n4540), .ZN(n4542) );
  NOR3_X1 U4979 ( .A1(n4544), .A2(n4543), .A3(n4542), .ZN(n4545) );
  AOI221_X1 U4980 ( .B1(DATAI_26_), .B2(n4547), .C1(n4546), .C2(keyinput_69), 
        .A(n4545), .ZN(n4549) );
  NAND2_X1 U4981 ( .A1(keyinput_73), .A2(DATAI_22_), .ZN(n4548) );
  OAI221_X1 U4982 ( .B1(n4550), .B2(n4549), .C1(keyinput_73), .C2(DATAI_22_), 
        .A(n4548), .ZN(n4559) );
  AOI22_X1 U4983 ( .A1(n4553), .A2(keyinput_74), .B1(n4552), .B2(keyinput_72), 
        .ZN(n4551) );
  OAI221_X1 U4984 ( .B1(n4553), .B2(keyinput_74), .C1(n4552), .C2(keyinput_72), 
        .A(n4551), .ZN(n4558) );
  OAI22_X1 U4985 ( .A1(DATAI_17_), .A2(keyinput_78), .B1(DATAI_16_), .B2(
        keyinput_79), .ZN(n4554) );
  AOI221_X1 U4986 ( .B1(DATAI_17_), .B2(keyinput_78), .C1(keyinput_79), .C2(
        DATAI_16_), .A(n4554), .ZN(n4557) );
  OAI22_X1 U4987 ( .A1(DATAI_20_), .A2(keyinput_75), .B1(DATAI_18_), .B2(
        keyinput_77), .ZN(n4555) );
  AOI221_X1 U4988 ( .B1(DATAI_20_), .B2(keyinput_75), .C1(keyinput_77), .C2(
        DATAI_18_), .A(n4555), .ZN(n4556) );
  OAI211_X1 U4989 ( .C1(n4559), .C2(n4558), .A(n4557), .B(n4556), .ZN(n4560)
         );
  NOR3_X1 U4990 ( .A1(n4562), .A2(n4561), .A3(n4560), .ZN(n4570) );
  INV_X1 U4991 ( .A(DATAI_12_), .ZN(n4869) );
  AOI22_X1 U4992 ( .A1(n2603), .A2(keyinput_84), .B1(n4869), .B2(keyinput_83), 
        .ZN(n4563) );
  OAI221_X1 U4993 ( .B1(n2603), .B2(keyinput_84), .C1(n4869), .C2(keyinput_83), 
        .A(n4563), .ZN(n4569) );
  OAI22_X1 U4994 ( .A1(DATAI_8_), .A2(keyinput_87), .B1(keyinput_89), .B2(
        DATAI_6_), .ZN(n4564) );
  AOI221_X1 U4995 ( .B1(DATAI_8_), .B2(keyinput_87), .C1(DATAI_6_), .C2(
        keyinput_89), .A(n4564), .ZN(n4568) );
  OAI22_X1 U4996 ( .A1(n4566), .A2(keyinput_85), .B1(n4845), .B2(keyinput_86), 
        .ZN(n4565) );
  AOI221_X1 U4997 ( .B1(n4566), .B2(keyinput_85), .C1(keyinput_86), .C2(n4845), 
        .A(n4565), .ZN(n4567) );
  OAI211_X1 U4998 ( .C1(n4570), .C2(n4569), .A(n4568), .B(n4567), .ZN(n4576)
         );
  OAI22_X1 U4999 ( .A1(n4572), .A2(keyinput_92), .B1(keyinput_91), .B2(
        DATAI_4_), .ZN(n4571) );
  AOI221_X1 U5000 ( .B1(n4572), .B2(keyinput_92), .C1(DATAI_4_), .C2(
        keyinput_91), .A(n4571), .ZN(n4575) );
  OAI22_X1 U5001 ( .A1(DATAI_2_), .A2(keyinput_93), .B1(DATAI_1_), .B2(
        keyinput_94), .ZN(n4573) );
  AOI221_X1 U5002 ( .B1(DATAI_2_), .B2(keyinput_93), .C1(keyinput_94), .C2(
        DATAI_1_), .A(n4573), .ZN(n4574) );
  OAI211_X1 U5003 ( .C1(n4577), .C2(n4576), .A(n4575), .B(n4574), .ZN(n4578)
         );
  AOI22_X1 U5004 ( .A1(n4579), .A2(n4578), .B1(keyinput_97), .B2(
        REG3_REG_7__SCAN_IN), .ZN(n4580) );
  OAI21_X1 U5005 ( .B1(keyinput_97), .B2(REG3_REG_7__SCAN_IN), .A(n4580), .ZN(
        n4585) );
  XOR2_X1 U5006 ( .A(keyinput_100), .B(REG3_REG_23__SCAN_IN), .Z(n4584) );
  AOI22_X1 U5007 ( .A1(n4582), .A2(keyinput_101), .B1(n4772), .B2(keyinput_102), .ZN(n4581) );
  OAI221_X1 U5008 ( .B1(n4582), .B2(keyinput_101), .C1(n4772), .C2(
        keyinput_102), .A(n4581), .ZN(n4583) );
  AOI211_X1 U5009 ( .C1(n4586), .C2(n4585), .A(n4584), .B(n4583), .ZN(n4589)
         );
  AOI22_X1 U5010 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput_104), .B1(
        REG3_REG_19__SCAN_IN), .B2(keyinput_103), .ZN(n4587) );
  OAI221_X1 U5011 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_104), .C1(
        REG3_REG_19__SCAN_IN), .C2(keyinput_103), .A(n4587), .ZN(n4588) );
  OR2_X1 U5012 ( .A1(n4589), .A2(n4588), .ZN(n4595) );
  OAI22_X1 U5013 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_105), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_108), .ZN(n4590) );
  AOI221_X1 U5014 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_105), .C1(
        keyinput_108), .C2(REG3_REG_12__SCAN_IN), .A(n4590), .ZN(n4594) );
  INV_X1 U5015 ( .A(keyinput_107), .ZN(n4591) );
  XNOR2_X1 U5016 ( .A(n4591), .B(REG3_REG_21__SCAN_IN), .ZN(n4593) );
  XNOR2_X1 U5017 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_106), .ZN(n4592) );
  NAND4_X1 U5018 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(n4596)
         );
  OAI221_X1 U5019 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_109), .C1(n4598), 
        .C2(n4597), .A(n4596), .ZN(n4601) );
  OAI22_X1 U5020 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_114), .B1(
        REG3_REG_0__SCAN_IN), .B2(keyinput_116), .ZN(n4599) );
  AOI221_X1 U5021 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_114), .C1(
        keyinput_116), .C2(REG3_REG_0__SCAN_IN), .A(n4599), .ZN(n4600) );
  OAI221_X1 U5022 ( .B1(n4603), .B2(n4602), .C1(n4603), .C2(n4601), .A(n4600), 
        .ZN(n4607) );
  AOI22_X1 U5023 ( .A1(n2570), .A2(keyinput_115), .B1(keyinput_117), .B2(n4605), .ZN(n4604) );
  OAI221_X1 U5024 ( .B1(n2570), .B2(keyinput_115), .C1(n4605), .C2(
        keyinput_117), .A(n4604), .ZN(n4606) );
  OAI22_X1 U5025 ( .A1(keyinput_118), .A2(n4609), .B1(n4607), .B2(n4606), .ZN(
        n4608) );
  AOI21_X1 U5026 ( .B1(keyinput_118), .B2(n4609), .A(n4608), .ZN(n4612) );
  INV_X1 U5027 ( .A(keyinput_119), .ZN(n4610) );
  MUX2_X1 U5028 ( .A(keyinput_119), .B(n4610), .S(IR_REG_0__SCAN_IN), .Z(n4611) );
  NOR2_X1 U5029 ( .A1(n4612), .A2(n4611), .ZN(n4615) );
  INV_X1 U5030 ( .A(keyinput_120), .ZN(n4613) );
  MUX2_X1 U5031 ( .A(n4613), .B(keyinput_120), .S(IR_REG_1__SCAN_IN), .Z(n4614) );
  NOR2_X1 U5032 ( .A1(n4615), .A2(n4614), .ZN(n4622) );
  AOI22_X1 U5033 ( .A1(n2519), .A2(keyinput_122), .B1(n4617), .B2(keyinput_121), .ZN(n4616) );
  OAI221_X1 U5034 ( .B1(n2519), .B2(keyinput_122), .C1(n4617), .C2(
        keyinput_121), .A(n4616), .ZN(n4621) );
  XNOR2_X1 U5035 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_123), .ZN(n4620) );
  OAI22_X1 U5036 ( .A1(n2557), .A2(keyinput_125), .B1(IR_REG_5__SCAN_IN), .B2(
        keyinput_124), .ZN(n4618) );
  AOI221_X1 U5037 ( .B1(n2557), .B2(keyinput_125), .C1(keyinput_124), .C2(
        IR_REG_5__SCAN_IN), .A(n4618), .ZN(n4619) );
  OAI211_X1 U5038 ( .C1(n4622), .C2(n4621), .A(n4620), .B(n4619), .ZN(n4625)
         );
  INV_X1 U5039 ( .A(keyinput_126), .ZN(n4623) );
  MUX2_X1 U5040 ( .A(keyinput_126), .B(n4623), .S(IR_REG_7__SCAN_IN), .Z(n4624) );
  NAND2_X1 U5041 ( .A1(n4625), .A2(n4624), .ZN(n4626) );
  OAI211_X1 U5042 ( .C1(IR_REG_8__SCAN_IN), .C2(keyinput_127), .A(n4627), .B(
        n4626), .ZN(n4628) );
  AOI21_X1 U5043 ( .B1(keyinput_127), .B2(IR_REG_8__SCAN_IN), .A(n4628), .ZN(
        n4629) );
  XNOR2_X1 U5044 ( .A(n4630), .B(n4629), .ZN(U3297) );
  AOI211_X1 U5045 ( .C1(n4632), .C2(n4631), .A(n2289), .B(n4748), .ZN(n4634)
         );
  AOI211_X1 U5046 ( .C1(n4737), .C2(ADDR_REG_5__SCAN_IN), .A(n4634), .B(n4633), 
        .ZN(n4639) );
  OAI211_X1 U5047 ( .C1(n4637), .C2(n4636), .A(n4744), .B(n4635), .ZN(n4638)
         );
  OAI211_X1 U5048 ( .C1(n4747), .C2(n4785), .A(n4639), .B(n4638), .ZN(U3245)
         );
  AOI211_X1 U5049 ( .C1(n4642), .C2(n4641), .A(n4640), .B(n4748), .ZN(n4644)
         );
  AOI211_X1 U5050 ( .C1(n4737), .C2(ADDR_REG_6__SCAN_IN), .A(n4644), .B(n4643), 
        .ZN(n4648) );
  OAI211_X1 U5051 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4646), .A(n4744), .B(n4645), 
        .ZN(n4647) );
  OAI211_X1 U5052 ( .C1(n4747), .C2(n4787), .A(n4648), .B(n4647), .ZN(U3246)
         );
  AOI22_X1 U5053 ( .A1(n4650), .A2(n4649), .B1(REG2_REG_7__SCAN_IN), .B2(n4795), .ZN(n4652) );
  OAI21_X1 U5054 ( .B1(n4653), .B2(n4652), .A(n4710), .ZN(n4651) );
  AOI21_X1 U5055 ( .B1(n4653), .B2(n4652), .A(n4651), .ZN(n4655) );
  AOI211_X1 U5056 ( .C1(n4737), .C2(ADDR_REG_7__SCAN_IN), .A(n4655), .B(n4654), 
        .ZN(n4661) );
  AOI21_X1 U5057 ( .B1(n4795), .B2(n4830), .A(n4656), .ZN(n4659) );
  AOI21_X1 U5058 ( .B1(n4659), .B2(n4658), .A(n4721), .ZN(n4657) );
  OAI21_X1 U5059 ( .B1(n4659), .B2(n4658), .A(n4657), .ZN(n4660) );
  OAI211_X1 U5060 ( .C1(n4747), .C2(n4795), .A(n4661), .B(n4660), .ZN(U3247)
         );
  AOI211_X1 U5061 ( .C1(n4664), .C2(n4663), .A(n4662), .B(n4721), .ZN(n4666)
         );
  AOI211_X1 U5062 ( .C1(n4737), .C2(ADDR_REG_8__SCAN_IN), .A(n4666), .B(n4665), 
        .ZN(n4670) );
  OAI211_X1 U5063 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4668), .A(n4710), .B(n4667), 
        .ZN(n4669) );
  OAI211_X1 U5064 ( .C1(n4747), .C2(n4837), .A(n4670), .B(n4669), .ZN(U3248)
         );
  AOI22_X1 U5065 ( .A1(n4671), .A2(n2316), .B1(REG1_REG_9__SCAN_IN), .B2(n4846), .ZN(n4673) );
  OAI21_X1 U5066 ( .B1(n4674), .B2(n4673), .A(n4744), .ZN(n4672) );
  AOI21_X1 U5067 ( .B1(n4674), .B2(n4673), .A(n4672), .ZN(n4676) );
  AOI211_X1 U5068 ( .C1(n4737), .C2(ADDR_REG_9__SCAN_IN), .A(n4676), .B(n4675), 
        .ZN(n4681) );
  OAI211_X1 U5069 ( .C1(n4679), .C2(n4678), .A(n4710), .B(n4677), .ZN(n4680)
         );
  OAI211_X1 U5070 ( .C1(n4747), .C2(n4846), .A(n4681), .B(n4680), .ZN(U3249)
         );
  OAI211_X1 U5071 ( .C1(n4684), .C2(REG2_REG_10__SCAN_IN), .A(n4683), .B(n4710), .ZN(n4688) );
  OAI211_X1 U5072 ( .C1(n4686), .C2(REG1_REG_10__SCAN_IN), .A(n4744), .B(n4685), .ZN(n4687) );
  OAI211_X1 U5073 ( .C1(n4747), .C2(n3436), .A(n4688), .B(n4687), .ZN(n4689)
         );
  AOI211_X1 U5074 ( .C1(n4737), .C2(ADDR_REG_10__SCAN_IN), .A(n4690), .B(n4689), .ZN(n4691) );
  INV_X1 U5075 ( .A(n4691), .ZN(U3250) );
  INV_X1 U5076 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4692) );
  AOI22_X1 U5077 ( .A1(n4693), .A2(REG1_REG_11__SCAN_IN), .B1(n4692), .B2(
        n4856), .ZN(n4696) );
  OAI21_X1 U5078 ( .B1(n4696), .B2(n4695), .A(n4744), .ZN(n4694) );
  AOI21_X1 U5079 ( .B1(n4696), .B2(n4695), .A(n4694), .ZN(n4698) );
  AOI211_X1 U5080 ( .C1(n4737), .C2(ADDR_REG_11__SCAN_IN), .A(n4698), .B(n4697), .ZN(n4703) );
  OAI211_X1 U5081 ( .C1(n4701), .C2(n4700), .A(n4710), .B(n4699), .ZN(n4702)
         );
  OAI211_X1 U5082 ( .C1(n4747), .C2(n4856), .A(n4703), .B(n4702), .ZN(U3251)
         );
  AOI211_X1 U5083 ( .C1(n4706), .C2(n4705), .A(n4704), .B(n4721), .ZN(n4708)
         );
  AOI211_X1 U5084 ( .C1(n4737), .C2(ADDR_REG_12__SCAN_IN), .A(n4708), .B(n4707), .ZN(n4713) );
  OAI211_X1 U5085 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4711), .A(n4710), .B(n4709), .ZN(n4712) );
  OAI211_X1 U5086 ( .C1(n4747), .C2(n4870), .A(n4713), .B(n4712), .ZN(U3252)
         );
  AOI21_X1 U5087 ( .B1(n4722), .B2(n3360), .A(n4714), .ZN(n4715) );
  XNOR2_X1 U5088 ( .A(n4716), .B(n4715), .ZN(n4726) );
  NAND2_X1 U5089 ( .A1(n4717), .A2(n2264), .ZN(n4718) );
  XNOR2_X1 U5090 ( .A(n4719), .B(n4718), .ZN(n4720) );
  OAI22_X1 U5091 ( .A1(n4722), .A2(n4747), .B1(n4721), .B2(n4720), .ZN(n4723)
         );
  AOI211_X1 U5092 ( .C1(n4737), .C2(ADDR_REG_13__SCAN_IN), .A(n4724), .B(n4723), .ZN(n4725) );
  OAI21_X1 U5093 ( .B1(n4726), .B2(n4748), .A(n4725), .ZN(U3253) );
  AOI221_X1 U5094 ( .B1(n4728), .B2(n4727), .C1(n3373), .C2(n4727), .A(n4748), 
        .ZN(n4729) );
  AOI211_X1 U5095 ( .C1(n4737), .C2(ADDR_REG_16__SCAN_IN), .A(n4730), .B(n4729), .ZN(n4734) );
  OAI221_X1 U5096 ( .B1(n4732), .B2(REG1_REG_16__SCAN_IN), .C1(n4732), .C2(
        n4731), .A(n4744), .ZN(n4733) );
  OAI211_X1 U5097 ( .C1(n4747), .C2(n4893), .A(n4734), .B(n4733), .ZN(U3256)
         );
  MUX2_X1 U5098 ( .A(REG2_REG_19__SCAN_IN), .B(n4330), .S(n4814), .Z(n4735) );
  AOI21_X1 U5099 ( .B1(n4737), .B2(ADDR_REG_19__SCAN_IN), .A(n4736), .ZN(n4746) );
  AOI22_X1 U5100 ( .A1(n4740), .A2(n4739), .B1(REG1_REG_18__SCAN_IN), .B2(
        n4738), .ZN(n4743) );
  MUX2_X1 U5101 ( .A(n4741), .B(REG1_REG_19__SCAN_IN), .S(n4814), .Z(n4742) );
  XNOR2_X1 U5102 ( .A(n4743), .B(n4742), .ZN(n4745) );
  INV_X1 U5103 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4749) );
  AOI22_X1 U5104 ( .A1(n4835), .A2(n4750), .B1(n4749), .B2(n4832), .ZN(U3467)
         );
  AOI21_X1 U5105 ( .B1(n4753), .B2(n4752), .A(n4751), .ZN(n4757) );
  AOI22_X1 U5106 ( .A1(n4754), .A2(n4851), .B1(REG3_REG_0__SCAN_IN), .B2(n4847), .ZN(n4755) );
  OAI221_X1 U5107 ( .B1(n4900), .B2(n4757), .C1(n4333), .C2(n4756), .A(n4755), 
        .ZN(U3290) );
  OAI22_X1 U5108 ( .A1(n4761), .A2(n4760), .B1(n4759), .B2(n4758), .ZN(n4762)
         );
  NOR2_X1 U5109 ( .A1(n4763), .A2(n4762), .ZN(n4766) );
  AOI22_X1 U5110 ( .A1(n4831), .A2(n4766), .B1(n4764), .B2(n2856), .ZN(U3519)
         );
  INV_X1 U5111 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5112 ( .A1(n4835), .A2(n4766), .B1(n4765), .B2(n4832), .ZN(U3469)
         );
  AOI22_X1 U5113 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4900), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4847), .ZN(n4770) );
  AOI22_X1 U5114 ( .A1(n4768), .A2(n4851), .B1(n4896), .B2(n4767), .ZN(n4769)
         );
  OAI211_X1 U5115 ( .C1(n4900), .C2(n4771), .A(n4770), .B(n4769), .ZN(U3288)
         );
  AOI22_X1 U5116 ( .A1(n4900), .A2(REG2_REG_3__SCAN_IN), .B1(n4847), .B2(n4772), .ZN(n4776) );
  AOI22_X1 U5117 ( .A1(n4774), .A2(n4851), .B1(n4896), .B2(n4773), .ZN(n4775)
         );
  OAI211_X1 U5118 ( .C1(n4900), .C2(n4777), .A(n4776), .B(n4775), .ZN(U3287)
         );
  INV_X1 U5119 ( .A(n4778), .ZN(n4780) );
  AOI211_X1 U5120 ( .C1(n4782), .C2(n4781), .A(n4780), .B(n4779), .ZN(n4784)
         );
  AOI22_X1 U5121 ( .A1(n4831), .A2(n4784), .B1(n3449), .B2(n2856), .ZN(U3522)
         );
  INV_X1 U5122 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4783) );
  AOI22_X1 U5123 ( .A1(n4835), .A2(n4784), .B1(n4783), .B2(n4832), .ZN(U3475)
         );
  AOI22_X1 U5124 ( .A1(STATE_REG_SCAN_IN), .A2(n4785), .B1(n2537), .B2(U3149), 
        .ZN(U3347) );
  AOI22_X1 U5125 ( .A1(STATE_REG_SCAN_IN), .A2(n4787), .B1(n4786), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5126 ( .A1(n4788), .A2(n4847), .B1(REG2_REG_6__SCAN_IN), .B2(n4900), .ZN(n4792) );
  AOI22_X1 U5127 ( .A1(n4790), .A2(n4851), .B1(n4896), .B2(n4789), .ZN(n4791)
         );
  OAI211_X1 U5128 ( .C1(n4900), .C2(n4793), .A(n4792), .B(n4791), .ZN(U3284)
         );
  AOI22_X1 U5129 ( .A1(STATE_REG_SCAN_IN), .A2(n4795), .B1(n4794), .B2(U3149), 
        .ZN(U3345) );
  NAND2_X1 U5130 ( .A1(n4797), .A2(n4796), .ZN(n4798) );
  XNOR2_X1 U5131 ( .A(n4798), .B(n4815), .ZN(n4808) );
  AOI22_X1 U5132 ( .A1(n4802), .A2(n4801), .B1(n4800), .B2(n4799), .ZN(n4803)
         );
  OAI21_X1 U5133 ( .B1(n4805), .B2(n4804), .A(n4803), .ZN(n4806) );
  AOI21_X1 U5134 ( .B1(n4808), .B2(n4807), .A(n4806), .ZN(n4828) );
  OR2_X1 U5135 ( .A1(n4810), .A2(n4809), .ZN(n4812) );
  AND3_X1 U5136 ( .A1(n4813), .A2(n4812), .A3(n4811), .ZN(n4825) );
  AOI21_X1 U5137 ( .B1(n4825), .B2(n4814), .A(n4900), .ZN(n4821) );
  NAND2_X1 U5138 ( .A1(n4816), .A2(n4815), .ZN(n4817) );
  AND2_X1 U5139 ( .A1(n4818), .A2(n4817), .ZN(n4827) );
  NAND2_X1 U5140 ( .A1(n4827), .A2(n4819), .ZN(n4820) );
  NAND3_X1 U5141 ( .A1(n4828), .A2(n4821), .A3(n4820), .ZN(n4822) );
  OAI21_X1 U5142 ( .B1(REG2_REG_7__SCAN_IN), .B2(n4333), .A(n4822), .ZN(n4823)
         );
  OAI21_X1 U5143 ( .B1(n4824), .B2(n4863), .A(n4823), .ZN(U3283) );
  AOI21_X1 U5144 ( .B1(n4827), .B2(n4826), .A(n4825), .ZN(n4829) );
  AND2_X1 U5145 ( .A1(n4829), .A2(n4828), .ZN(n4834) );
  AOI22_X1 U5146 ( .A1(n4831), .A2(n4834), .B1(n4830), .B2(n2856), .ZN(U3525)
         );
  INV_X1 U5147 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U5148 ( .A1(n4835), .A2(n4834), .B1(n4833), .B2(n4832), .ZN(U3481)
         );
  AOI22_X1 U5149 ( .A1(STATE_REG_SCAN_IN), .A2(n4837), .B1(n4836), .B2(U3149), 
        .ZN(U3344) );
  AOI22_X1 U5150 ( .A1(n4838), .A2(n4847), .B1(REG2_REG_8__SCAN_IN), .B2(n4900), .ZN(n4843) );
  INV_X1 U5151 ( .A(n4839), .ZN(n4840) );
  AOI22_X1 U5152 ( .A1(n4841), .A2(n4851), .B1(n4896), .B2(n4840), .ZN(n4842)
         );
  OAI211_X1 U5153 ( .C1(n4900), .C2(n4844), .A(n4843), .B(n4842), .ZN(U3282)
         );
  AOI22_X1 U5154 ( .A1(STATE_REG_SCAN_IN), .A2(n4846), .B1(n4845), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5155 ( .A1(n4848), .A2(n4847), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4900), .ZN(n4854) );
  INV_X1 U5156 ( .A(n4849), .ZN(n4850) );
  AOI22_X1 U5157 ( .A1(n4852), .A2(n4851), .B1(n4896), .B2(n4850), .ZN(n4853)
         );
  OAI211_X1 U5158 ( .C1(n4900), .C2(n4855), .A(n4854), .B(n4853), .ZN(U3280)
         );
  AOI22_X1 U5159 ( .A1(STATE_REG_SCAN_IN), .A2(n4856), .B1(n2603), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5160 ( .A(n4857), .ZN(n4861) );
  OAI22_X1 U5161 ( .A1(n4861), .A2(n4860), .B1(n4859), .B2(n4858), .ZN(n4866)
         );
  OAI22_X1 U5162 ( .A1(n4864), .A2(n4863), .B1(n4862), .B2(n4333), .ZN(n4865)
         );
  NOR2_X1 U5163 ( .A1(n4866), .A2(n4865), .ZN(n4867) );
  OAI21_X1 U5164 ( .B1(n4868), .B2(n4900), .A(n4867), .ZN(U3279) );
  AOI22_X1 U5165 ( .A1(STATE_REG_SCAN_IN), .A2(n4870), .B1(n4869), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5166 ( .A1(U3149), .A2(n4871), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4872) );
  INV_X1 U5167 ( .A(n4872), .ZN(U3339) );
  AOI21_X1 U5168 ( .B1(n4875), .B2(n4874), .A(n4873), .ZN(n4882) );
  NAND2_X1 U5169 ( .A1(n4877), .A2(n4876), .ZN(n4881) );
  NAND2_X1 U5170 ( .A1(n4879), .A2(n4878), .ZN(n4880) );
  AND3_X1 U5171 ( .A1(n4882), .A2(n4881), .A3(n4880), .ZN(n4889) );
  XNOR2_X1 U5172 ( .A(n4884), .B(n4883), .ZN(n4885) );
  XNOR2_X1 U5173 ( .A(n3792), .B(n4885), .ZN(n4887) );
  NAND2_X1 U5174 ( .A1(n4887), .A2(n4886), .ZN(n4888) );
  OAI211_X1 U5175 ( .C1(n4891), .C2(n4890), .A(n4889), .B(n4888), .ZN(U3238)
         );
  AOI22_X1 U5176 ( .A1(STATE_REG_SCAN_IN), .A2(n4893), .B1(n4892), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5177 ( .A1(STATE_REG_SCAN_IN), .A2(n4895), .B1(n4894), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U5178 ( .A1(n4897), .A2(n4896), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4900), .ZN(n4898) );
  OAI21_X1 U5179 ( .B1(n4900), .B2(n4899), .A(n4898), .ZN(U3261) );
  CLKBUF_X1 U2293 ( .A(n2495), .Z(n2753) );
  CLKBUF_X3 U2396 ( .A(n2496), .Z(n2513) );
endmodule

