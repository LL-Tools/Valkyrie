

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698;

  OAI211_X1 U10990 ( .C1(n20371), .C2(n20368), .A(n20419), .B(n20367), .ZN(
        n20404) );
  NOR2_X1 U10991 ( .A1(n10190), .A2(n10087), .ZN(n21375) );
  NOR2_X1 U10992 ( .A1(n14508), .A2(n18522), .ZN(n18531) );
  INV_X1 U10993 ( .A(n18015), .ZN(n18032) );
  AOI211_X1 U10994 ( .C1(n20016), .C2(n20607), .A(n20035), .B(n20606), .ZN(
        n20017) );
  AND2_X1 U10995 ( .A1(n11145), .A2(n13189), .ZN(n20419) );
  AOI21_X1 U10996 ( .B1(n16607), .B2(n16608), .A(n10006), .ZN(n11035) );
  OR2_X1 U10997 ( .A1(n15816), .A2(n20811), .ZN(n20826) );
  NOR2_X1 U10998 ( .A1(n10649), .A2(n10646), .ZN(n20209) );
  NAND2_X1 U10999 ( .A1(n10236), .A2(n10234), .ZN(n12146) );
  AND2_X1 U11000 ( .A1(n9574), .A2(n13350), .ZN(n10657) );
  CLKBUF_X3 U11001 ( .A(n13299), .Z(n9548) );
  INV_X2 U11002 ( .A(n13350), .ZN(n16366) );
  INV_X1 U11003 ( .A(n19166), .ZN(n18396) );
  NOR2_X1 U11004 ( .A1(n11805), .A2(n11804), .ZN(n19153) );
  CLKBUF_X1 U11005 ( .A(n12050), .Z(n12592) );
  CLKBUF_X2 U11006 ( .A(n12244), .Z(n12746) );
  CLKBUF_X2 U11007 ( .A(n12160), .Z(n12743) );
  CLKBUF_X2 U11008 ( .A(n12149), .Z(n12744) );
  INV_X1 U11009 ( .A(n13534), .ZN(n10733) );
  AND2_X1 U11010 ( .A1(n14202), .A2(n14550), .ZN(n13542) );
  AND2_X1 U11011 ( .A1(n14202), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13527) );
  INV_X1 U11012 ( .A(n10496), .ZN(n9595) );
  INV_X4 U11013 ( .A(n11727), .ZN(n18334) );
  AND2_X2 U11014 ( .A1(n11559), .A2(n17351), .ZN(n11684) );
  CLKBUF_X2 U11015 ( .A(n10575), .Z(n11287) );
  AND2_X2 U11016 ( .A1(n14033), .A2(n11561), .ZN(n11606) );
  INV_X1 U11017 ( .A(n18256), .ZN(n17449) );
  INV_X2 U11018 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17345) );
  BUF_X4 U11019 ( .A(n12263), .Z(n9551) );
  AND2_X2 U11020 ( .A1(n11963), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14355) );
  NAND2_X2 U11021 ( .A1(n15010), .A2(n15012), .ZN(n14988) );
  NOR2_X2 U11022 ( .A1(n20768), .A2(n12094), .ZN(n20756) );
  AND2_X2 U11023 ( .A1(n14498), .A2(n12094), .ZN(n14493) );
  AND2_X1 U11024 ( .A1(n14556), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9592) );
  AND2_X1 U11025 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11979) );
  AND2_X2 U11026 ( .A1(n10107), .A2(n14341), .ZN(n12068) );
  AND2_X1 U11027 ( .A1(n9850), .A2(n9849), .ZN(n10134) );
  INV_X1 U11028 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10490) );
  AOI21_X1 U11029 ( .B1(n10624), .B2(P2_EBX_REG_2__SCAN_IN), .A(n10483), .ZN(
        n10617) );
  INV_X1 U11030 ( .A(n10649), .ZN(n10647) );
  NAND2_X2 U11031 ( .A1(n12239), .A2(n12238), .ZN(n12834) );
  AND2_X1 U11032 ( .A1(n9881), .A2(n9765), .ZN(n9945) );
  INV_X1 U11033 ( .A(n13297), .ZN(n11223) );
  AND2_X1 U11034 ( .A1(n13507), .A2(n14556), .ZN(n13540) );
  AND2_X1 U11035 ( .A1(n16405), .A2(n14580), .ZN(n13701) );
  AND2_X1 U11036 ( .A1(n10052), .A2(n9601), .ZN(n10659) );
  NOR2_X2 U11037 ( .A1(n14074), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11559) );
  AND2_X1 U11038 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11561) );
  CLKBUF_X2 U11039 ( .A(n9565), .Z(n9577) );
  NAND2_X1 U11040 ( .A1(n12252), .A2(n12251), .ZN(n10178) );
  CLKBUF_X2 U11042 ( .A(n13719), .Z(n9591) );
  INV_X1 U11043 ( .A(n16362), .ZN(n16305) );
  INV_X1 U11044 ( .A(n13243), .ZN(n16249) );
  NAND2_X1 U11045 ( .A1(n13365), .A2(n13364), .ZN(n13368) );
  NOR2_X2 U11047 ( .A1(n14679), .A2(n10012), .ZN(n15220) );
  NAND2_X1 U11048 ( .A1(n15703), .A2(n15802), .ZN(n15816) );
  NAND2_X1 U11049 ( .A1(n12253), .A2(n12901), .ZN(n15870) );
  OR2_X1 U11050 ( .A1(n16400), .A2(n16399), .ZN(n16397) );
  OAI21_X1 U11051 ( .B1(n11020), .B2(n11513), .A(n16974), .ZN(n16688) );
  NAND2_X1 U11052 ( .A1(n13370), .A2(n13369), .ZN(n14197) );
  XNOR2_X1 U11053 ( .A(n11918), .B(n11917), .ZN(n13808) );
  NOR2_X1 U11054 ( .A1(n11776), .A2(n11775), .ZN(n9695) );
  INV_X1 U11055 ( .A(n15255), .ZN(n20668) );
  AND2_X1 U11056 ( .A1(n15184), .A2(n13031), .ZN(n15139) );
  INV_X1 U11057 ( .A(n9593), .ZN(n17491) );
  AND2_X1 U11058 ( .A1(n9789), .A2(n11503), .ZN(n16874) );
  AND2_X1 U11059 ( .A1(n16691), .A2(n10216), .ZN(n16971) );
  OAI21_X1 U11060 ( .B1(n16741), .B2(n16717), .A(n16716), .ZN(n16728) );
  INV_X1 U11061 ( .A(n20014), .ZN(n20037) );
  INV_X1 U11062 ( .A(n20272), .ZN(n20286) );
  OAI21_X1 U11063 ( .B1(n20371), .B2(n20370), .A(n20369), .ZN(n20403) );
  OR2_X1 U11064 ( .A1(n17683), .A2(n17682), .ZN(n17684) );
  INV_X1 U11065 ( .A(n18533), .ZN(n18522) );
  INV_X1 U11066 ( .A(n18712), .ZN(n10316) );
  INV_X1 U11067 ( .A(n17314), .ZN(n19122) );
  INV_X1 U11068 ( .A(n20693), .ZN(n20678) );
  AOI211_X1 U11069 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17724), .A(n17698), 
        .B(n17697), .ZN(n17701) );
  INV_X1 U11070 ( .A(n18904), .ZN(n18811) );
  INV_X4 U11071 ( .A(n15595), .ZN(n15583) );
  INV_X1 U11072 ( .A(n18214), .ZN(n9556) );
  AND2_X2 U11073 ( .A1(n14355), .A2(n14341), .ZN(n12263) );
  BUF_X4 U11074 ( .A(n10624), .Z(n11523) );
  AND3_X1 U11075 ( .A1(n10660), .A2(n10272), .A3(n10271), .ZN(n9546) );
  NAND2_X2 U11076 ( .A1(n10274), .A2(n10273), .ZN(n11279) );
  AND2_X2 U11077 ( .A1(n9986), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10670) );
  NOR3_X4 U11078 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n18017) );
  AND2_X1 U11079 ( .A1(n11253), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9547) );
  AND2_X4 U11080 ( .A1(n11253), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10624) );
  NAND2_X2 U11081 ( .A1(n10182), .A2(n10669), .ZN(n10181) );
  AND2_X2 U11082 ( .A1(n10910), .A2(n10926), .ZN(n10907) );
  NAND4_X4 U11083 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12111) );
  NAND2_X4 U11084 ( .A1(n10181), .A2(n10172), .ZN(n19875) );
  NAND2_X2 U11085 ( .A1(n10180), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10172) );
  INV_X2 U11086 ( .A(n9594), .ZN(n13719) );
  AOI21_X2 U11087 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15451), .A(
        n15443), .ZN(n15444) );
  AND3_X2 U11088 ( .A1(n10238), .A2(n10239), .A3(n9710), .ZN(n11922) );
  OAI21_X2 U11089 ( .B1(n12220), .B2(n10438), .A(n10436), .ZN(n14107) );
  XNOR2_X2 U11090 ( .A(n16578), .B(n16576), .ZN(n16588) );
  AND4_X2 U11091 ( .A1(n10713), .A2(n10712), .A3(n9705), .A4(n10711), .ZN(
        n10722) );
  AND2_X1 U11092 ( .A1(n10659), .A2(n13361), .ZN(n20324) );
  AND2_X2 U11093 ( .A1(n9825), .A2(n10658), .ZN(n19978) );
  XNOR2_X2 U11094 ( .A(n12146), .B(n12145), .ZN(n12203) );
  OR2_X2 U11095 ( .A1(n13808), .A2(n10241), .ZN(n10238) );
  NAND3_X2 U11096 ( .A1(n10016), .A2(n10300), .A3(n10661), .ZN(n10051) );
  AND2_X2 U11097 ( .A1(n9670), .A2(n9546), .ZN(n10016) );
  AND2_X1 U11098 ( .A1(n10107), .A2(n14341), .ZN(n9549) );
  AND2_X2 U11099 ( .A1(n10107), .A2(n14341), .ZN(n9550) );
  XNOR2_X2 U11100 ( .A(n12199), .B(n12197), .ZN(n12210) );
  NAND2_X2 U11101 ( .A1(n12216), .A2(n12177), .ZN(n12199) );
  INV_X1 U11102 ( .A(n11493), .ZN(n9805) );
  NAND2_X2 U11103 ( .A1(n9605), .A2(n9851), .ZN(n17493) );
  AND2_X2 U11104 ( .A1(n13708), .A2(n10558), .ZN(n9851) );
  NOR2_X4 U11106 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14365) );
  NAND2_X2 U11107 ( .A1(n9621), .A2(n11495), .ZN(n10600) );
  OAI21_X2 U11108 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16739), .A(
        n16738), .ZN(n17040) );
  AND2_X4 U11109 ( .A1(n10077), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11974) );
  NAND2_X2 U11110 ( .A1(n10578), .A2(n11279), .ZN(n13271) );
  NAND2_X4 U11111 ( .A1(n10275), .A2(n10551), .ZN(n10578) );
  NOR2_X2 U11112 ( .A1(n14686), .A2(n16434), .ZN(n16428) );
  AND2_X1 U11113 ( .A1(n10111), .A2(n14341), .ZN(n9554) );
  INV_X1 U11114 ( .A(n18214), .ZN(n9555) );
  INV_X1 U11115 ( .A(n9555), .ZN(n9557) );
  AND2_X1 U11116 ( .A1(n11559), .A2(n14033), .ZN(n18294) );
  AND2_X4 U11117 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14341) );
  OAI21_X1 U11118 ( .B1(n16664), .B2(n10429), .A(n10424), .ZN(n14840) );
  OAI21_X1 U11119 ( .B1(n9975), .B2(n9977), .A(n14810), .ZN(n16664) );
  AND2_X1 U11120 ( .A1(n10268), .A2(n10352), .ZN(n16575) );
  OAI21_X1 U11121 ( .B1(n15437), .B2(n20837), .A(n10380), .ZN(n10309) );
  OR2_X1 U11122 ( .A1(n17189), .A2(n18712), .ZN(n10314) );
  XNOR2_X1 U11123 ( .A(n13088), .B(n14933), .ZN(n14960) );
  AND2_X1 U11124 ( .A1(n10353), .A2(n9624), .ZN(n10268) );
  AND2_X1 U11125 ( .A1(n18677), .A2(n9664), .ZN(n17332) );
  NAND2_X1 U11126 ( .A1(n20362), .A2(n20332), .ZN(n20360) );
  XNOR2_X1 U11127 ( .A(n10936), .B(n10939), .ZN(n9790) );
  NAND2_X1 U11128 ( .A1(n20362), .A2(n20250), .ZN(n20272) );
  AOI21_X1 U11129 ( .B1(n10355), .B2(n10358), .A(n10354), .ZN(n10353) );
  XNOR2_X1 U11130 ( .A(n14197), .B(n14199), .ZN(n20567) );
  INV_X4 U11131 ( .A(n15294), .ZN(n9558) );
  NOR2_X1 U11132 ( .A1(n10254), .A2(n17315), .ZN(n17267) );
  AND2_X1 U11133 ( .A1(n10048), .A2(n10651), .ZN(n20016) );
  INV_X1 U11134 ( .A(n17139), .ZN(n9563) );
  AND2_X1 U11135 ( .A1(n12967), .A2(n13767), .ZN(n13115) );
  NAND2_X1 U11136 ( .A1(n11505), .A2(n20602), .ZN(n17139) );
  AND2_X1 U11137 ( .A1(n18366), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n18364) );
  NAND2_X1 U11138 ( .A1(n19029), .A2(n17314), .ZN(n18995) );
  NAND2_X1 U11139 ( .A1(n10610), .A2(n10611), .ZN(n10189) );
  OAI22_X1 U11140 ( .A1(n12832), .A2(n12831), .B1(n12847), .B2(n12830), .ZN(
        n12836) );
  NAND2_X1 U11141 ( .A1(n18383), .A2(P3_EBX_REG_2__SCAN_IN), .ZN(n18381) );
  AND2_X1 U11142 ( .A1(n10591), .A2(n10590), .ZN(n11253) );
  OR2_X1 U11143 ( .A1(n11843), .A2(n11888), .ZN(n11940) );
  NAND2_X1 U11144 ( .A1(n10055), .A2(n18396), .ZN(n14070) );
  NOR2_X1 U11145 ( .A1(n10596), .A2(n13271), .ZN(n10590) );
  NAND2_X1 U11146 ( .A1(n9609), .A2(n9647), .ZN(n14335) );
  BUF_X1 U11148 ( .A(n12093), .Z(n9580) );
  INV_X1 U11149 ( .A(n9801), .ZN(n10584) );
  OR2_X1 U11150 ( .A1(n11634), .A2(n11633), .ZN(n18529) );
  BUF_X1 U11151 ( .A(n13080), .Z(n9573) );
  CLKBUF_X2 U11152 ( .A(n12111), .Z(n20854) );
  CLKBUF_X2 U11153 ( .A(n12086), .Z(n20869) );
  INV_X8 U11154 ( .A(n11799), .ZN(n18349) );
  INV_X2 U11155 ( .A(n13533), .ZN(n13465) );
  INV_X1 U11156 ( .A(n11684), .ZN(n9567) );
  INV_X1 U11157 ( .A(n11649), .ZN(n18325) );
  INV_X2 U11158 ( .A(n17376), .ZN(n11799) );
  CLKBUF_X2 U11159 ( .A(n12045), .Z(n12603) );
  INV_X4 U11160 ( .A(n18323), .ZN(n9559) );
  INV_X1 U11161 ( .A(n10379), .ZN(n12149) );
  BUF_X2 U11162 ( .A(n12719), .Z(n12756) );
  BUF_X2 U11163 ( .A(n12747), .Z(n12591) );
  CLKBUF_X2 U11164 ( .A(n12063), .Z(n12720) );
  INV_X4 U11165 ( .A(n11623), .ZN(n9560) );
  INV_X4 U11166 ( .A(n17408), .ZN(n9561) );
  INV_X1 U11167 ( .A(n13511), .ZN(n9562) );
  CLKBUF_X2 U11168 ( .A(n12754), .Z(n12664) );
  NAND2_X2 U11169 ( .A1(n9576), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10727) );
  AND2_X4 U11170 ( .A1(n14365), .A2(n11979), .ZN(n12753) );
  INV_X2 U11171 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14074) );
  INV_X2 U11172 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10077) );
  NOR2_X4 U11173 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10150) );
  AND2_X1 U11174 ( .A1(n10142), .A2(n10141), .ZN(n16623) );
  AND2_X1 U11175 ( .A1(n10100), .A2(n10099), .ZN(n16677) );
  AOI21_X1 U11176 ( .B1(n9653), .B2(n9823), .A(n16944), .ZN(n16945) );
  AOI21_X1 U11177 ( .B1(n9653), .B2(n9824), .A(n16659), .ZN(n16660) );
  NAND2_X1 U11178 ( .A1(n16738), .A2(n16730), .ZN(n17013) );
  AND2_X1 U11179 ( .A1(n13171), .A2(n10336), .ZN(n10335) );
  AND2_X1 U11180 ( .A1(n9993), .A2(n10054), .ZN(n16932) );
  AND2_X1 U11181 ( .A1(n9965), .A2(n9964), .ZN(n16629) );
  AOI21_X1 U11182 ( .B1(n17008), .B2(n16836), .A(n16723), .ZN(n16724) );
  AND2_X1 U11183 ( .A1(n9788), .A2(n9787), .ZN(n9786) );
  NAND2_X1 U11184 ( .A1(n10329), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9857) );
  OAI21_X1 U11185 ( .B1(n16594), .B2(n10153), .A(n10325), .ZN(n10152) );
  AND2_X1 U11186 ( .A1(n10031), .A2(n10030), .ZN(n16573) );
  AOI21_X1 U11187 ( .B1(n10306), .B2(n10305), .A(n10302), .ZN(n10301) );
  OR2_X1 U11188 ( .A1(n9966), .A2(n16911), .ZN(n9965) );
  XNOR2_X1 U11189 ( .A(n16664), .B(n9719), .ZN(n16947) );
  AOI21_X1 U11190 ( .B1(n14815), .B2(n13168), .A(n13167), .ZN(n16970) );
  XNOR2_X1 U11191 ( .A(n9903), .B(n9720), .ZN(n17008) );
  AND2_X1 U11192 ( .A1(n16794), .A2(n16793), .ZN(n16796) );
  OR2_X1 U11193 ( .A1(n11040), .A2(n9862), .ZN(n9856) );
  NAND2_X1 U11194 ( .A1(n16617), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16594) );
  AND2_X1 U11195 ( .A1(n9807), .A2(n9806), .ZN(n16617) );
  INV_X1 U11196 ( .A(n13160), .ZN(n9975) );
  NAND2_X1 U11197 ( .A1(n9961), .A2(n9959), .ZN(n16912) );
  AND2_X1 U11198 ( .A1(n9822), .A2(n13175), .ZN(n9877) );
  OAI21_X1 U11199 ( .B1(n9771), .B2(n14858), .A(n14974), .ZN(n15437) );
  NAND2_X1 U11200 ( .A1(n15435), .A2(n13126), .ZN(n13173) );
  OAI22_X1 U11201 ( .A1(n10330), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n13307), .B2(n16592), .ZN(n10328) );
  AOI21_X1 U11202 ( .B1(n14975), .B2(n14974), .A(n14973), .ZN(n15430) );
  OAI21_X1 U11203 ( .B1(n15148), .B2(n15136), .A(n15135), .ZN(n15543) );
  NOR2_X1 U11204 ( .A1(n14962), .A2(n13140), .ZN(n12774) );
  OAI21_X1 U11205 ( .B1(n14992), .B2(n14991), .A(n14990), .ZN(n15353) );
  NAND2_X1 U11206 ( .A1(n15540), .A2(n9815), .ZN(n15525) );
  NAND2_X1 U11207 ( .A1(n13750), .A2(n12740), .ZN(n14962) );
  INV_X1 U11208 ( .A(n16592), .ZN(n10331) );
  OR2_X1 U11209 ( .A1(n16883), .A2(n16884), .ZN(n10151) );
  OAI21_X1 U11210 ( .B1(n15054), .B2(n9645), .A(n15040), .ZN(n15491) );
  NAND2_X1 U11211 ( .A1(n10314), .A2(n10313), .ZN(n17286) );
  OAI21_X1 U11212 ( .B1(n15025), .B2(n15024), .A(n15023), .ZN(n15461) );
  AND2_X1 U11213 ( .A1(n15166), .A2(n15147), .ZN(n15148) );
  OAI211_X1 U11214 ( .C1(n20102), .C2(n20086), .A(n20085), .B(n20419), .ZN(
        n20105) );
  XNOR2_X1 U11215 ( .A(n13301), .B(n13300), .ZN(n16369) );
  XNOR2_X1 U11216 ( .A(n10403), .B(n10402), .ZN(n14806) );
  AND3_X1 U11217 ( .A1(n15134), .A2(n15179), .A3(n15165), .ZN(n15166) );
  OR2_X1 U11218 ( .A1(n15098), .A2(n15039), .ZN(n15040) );
  CLKBUF_X1 U11219 ( .A(n15010), .Z(n15011) );
  NAND2_X1 U11220 ( .A1(n10073), .A2(n10072), .ZN(n13752) );
  INV_X1 U11221 ( .A(n10299), .ZN(n10935) );
  OAI211_X1 U11222 ( .C1(n20185), .C2(n20181), .A(n20419), .B(n20180), .ZN(
        n20205) );
  NAND2_X1 U11223 ( .A1(n9846), .A2(n9845), .ZN(n16835) );
  OR2_X1 U11224 ( .A1(n10231), .A2(n9820), .ZN(n15594) );
  NOR2_X1 U11225 ( .A1(n20213), .A2(n10165), .ZN(n20214) );
  NAND2_X1 U11226 ( .A1(n13762), .A2(n12587), .ZN(n13764) );
  NAND2_X1 U11227 ( .A1(n10850), .A2(n13293), .ZN(n16795) );
  NAND2_X1 U11228 ( .A1(n10825), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10827) );
  OAI211_X1 U11229 ( .C1(n19949), .C2(n20570), .A(n20419), .B(n19948), .ZN(
        n19967) );
  AOI21_X1 U11230 ( .B1(n10362), .B2(n10364), .A(n9837), .ZN(n10360) );
  INV_X1 U11231 ( .A(n10828), .ZN(n16832) );
  AND2_X1 U11232 ( .A1(n10363), .A2(n11171), .ZN(n10362) );
  NOR2_X1 U11233 ( .A1(n9911), .A2(n9910), .ZN(n9909) );
  NAND2_X1 U11234 ( .A1(n9945), .A2(n9912), .ZN(n10070) );
  NAND2_X1 U11235 ( .A1(n10063), .A2(n16284), .ZN(n10299) );
  NOR2_X1 U11236 ( .A1(n9790), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16830) );
  NAND3_X1 U11237 ( .A1(n12928), .A2(n9764), .A3(n9880), .ZN(n9912) );
  NAND2_X1 U11238 ( .A1(n15973), .A2(n10341), .ZN(n15966) );
  INV_X1 U11239 ( .A(n20455), .ZN(n20468) );
  AND2_X1 U11240 ( .A1(n10018), .A2(n10017), .ZN(n9830) );
  NAND2_X1 U11241 ( .A1(n13087), .A2(n13086), .ZN(n13088) );
  OR2_X1 U11242 ( .A1(n17332), .A2(n10316), .ZN(n9927) );
  NOR2_X2 U11243 ( .A1(n20335), .A2(n20178), .ZN(n20231) );
  XNOR2_X1 U11244 ( .A(n14937), .B(n14936), .ZN(n15627) );
  NAND2_X1 U11245 ( .A1(n20251), .A2(n20361), .ZN(n20472) );
  OR2_X1 U11246 ( .A1(n20115), .A2(n20562), .ZN(n20014) );
  OR2_X1 U11247 ( .A1(n15962), .A2(n11513), .ZN(n16579) );
  NAND2_X1 U11248 ( .A1(n10183), .A2(n10822), .ZN(n10937) );
  OR2_X1 U11249 ( .A1(n20567), .A2(n19840), .ZN(n20010) );
  AND2_X1 U11250 ( .A1(n20567), .A2(n21692), .ZN(n20362) );
  AND2_X1 U11251 ( .A1(n20567), .A2(n19840), .ZN(n20251) );
  AND2_X1 U11252 ( .A1(n9701), .A2(n15527), .ZN(n9880) );
  NOR2_X1 U11253 ( .A1(n9883), .A2(n9882), .ZN(n9881) );
  OR2_X1 U11254 ( .A1(n15654), .A2(n15646), .ZN(n15631) );
  AOI21_X1 U11255 ( .B1(n11035), .B2(n10357), .A(n10356), .ZN(n10355) );
  OAI21_X2 U11256 ( .B1(n15675), .B2(n13125), .A(n15622), .ZN(n15653) );
  AND2_X1 U11257 ( .A1(n9602), .A2(n9757), .ZN(n10074) );
  INV_X1 U11258 ( .A(n14678), .ZN(n10014) );
  NOR2_X1 U11259 ( .A1(n9600), .A2(n10434), .ZN(n10432) );
  NAND2_X1 U11260 ( .A1(n9766), .A2(n12284), .ZN(n14424) );
  OR2_X1 U11261 ( .A1(n20578), .A2(n20009), .ZN(n20562) );
  NOR2_X1 U11262 ( .A1(n9955), .A2(n9871), .ZN(n9870) );
  AND2_X1 U11263 ( .A1(n9676), .A2(n10465), .ZN(n9915) );
  NAND2_X1 U11264 ( .A1(n12923), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12924) );
  OR2_X1 U11265 ( .A1(n20578), .A2(n20585), .ZN(n20178) );
  AND2_X1 U11266 ( .A1(n15537), .A2(n15524), .ZN(n15527) );
  NAND2_X1 U11267 ( .A1(n11706), .A2(n10462), .ZN(n18770) );
  AND4_X1 U11268 ( .A1(n10187), .A2(n10802), .A3(n10799), .A4(n10186), .ZN(
        n10185) );
  NAND2_X1 U11269 ( .A1(n9818), .A2(n12908), .ZN(n12923) );
  OR2_X1 U11270 ( .A1(n9664), .A2(n11717), .ZN(n10322) );
  NAND2_X1 U11271 ( .A1(n11157), .A2(n11158), .ZN(n11165) );
  NAND2_X1 U11272 ( .A1(n18147), .A2(n11836), .ZN(n18149) );
  AND2_X1 U11273 ( .A1(n15563), .A2(n15560), .ZN(n15514) );
  AND3_X1 U11274 ( .A1(n10776), .A2(n10772), .A3(n10161), .ZN(n9868) );
  NAND2_X1 U11275 ( .A1(n13326), .A2(n13330), .ZN(n17704) );
  AND3_X1 U11276 ( .A1(n10261), .A2(n10260), .A3(n10259), .ZN(n10300) );
  AND2_X1 U11277 ( .A1(n9918), .A2(n12278), .ZN(n9622) );
  AOI21_X1 U11278 ( .B1(n20016), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A(n9833), .ZN(n10802) );
  INV_X1 U11279 ( .A(n15326), .ZN(n10013) );
  NAND2_X1 U11280 ( .A1(n9581), .A2(n12934), .ZN(n14615) );
  OR2_X1 U11281 ( .A1(n18713), .A2(n18973), .ZN(n11717) );
  NOR2_X1 U11282 ( .A1(n14078), .A2(n14165), .ZN(n14163) );
  AND2_X1 U11283 ( .A1(n14006), .A2(n13358), .ZN(n14099) );
  OR2_X1 U11284 ( .A1(n19904), .A2(n13436), .ZN(n9678) );
  OAI21_X1 U11285 ( .B1(n18713), .B2(n18669), .A(n11715), .ZN(n11716) );
  OR2_X1 U11286 ( .A1(n14385), .A2(n10323), .ZN(n18788) );
  NAND2_X1 U11287 ( .A1(n15009), .A2(n14993), .ZN(n14995) );
  OAI21_X2 U11288 ( .B1(n16004), .B2(n16602), .A(n16249), .ZN(n15992) );
  OAI21_X1 U11289 ( .B1(n15867), .B2(n12897), .A(n12887), .ZN(n14255) );
  NAND2_X2 U11290 ( .A1(n9772), .A2(n10178), .ZN(n12901) );
  AOI21_X1 U11291 ( .B1(n10382), .B2(n12209), .A(n10383), .ZN(n10381) );
  OR2_X1 U11292 ( .A1(n18824), .A2(n18730), .ZN(n18884) );
  NAND2_X1 U11293 ( .A1(n10647), .A2(n10646), .ZN(n20140) );
  AND2_X1 U11294 ( .A1(n15036), .A2(n15007), .ZN(n15009) );
  AND2_X1 U11295 ( .A1(n10048), .A2(n10657), .ZN(n10798) );
  AND2_X1 U11296 ( .A1(n16083), .A2(n13293), .ZN(n11027) );
  AND3_X1 U11297 ( .A1(n10032), .A2(n10178), .A3(n10033), .ZN(n12322) );
  OR2_X1 U11298 ( .A1(n20826), .A2(n15817), .ZN(n17528) );
  NOR2_X1 U11299 ( .A1(n10646), .A2(n14784), .ZN(n10116) );
  AND2_X1 U11300 ( .A1(n9825), .A2(n10657), .ZN(n10796) );
  AND2_X1 U11301 ( .A1(n13358), .A2(n13355), .ZN(n14005) );
  NAND2_X1 U11302 ( .A1(n12214), .A2(n12213), .ZN(n14133) );
  NAND2_X1 U11303 ( .A1(n18906), .A2(n18799), .ZN(n18860) );
  NAND2_X1 U11304 ( .A1(n14728), .A2(n18515), .ZN(n18810) );
  AND2_X1 U11305 ( .A1(n15816), .A2(n20825), .ZN(n15823) );
  AND2_X1 U11306 ( .A1(n11011), .A2(n9656), .ZN(n16083) );
  NAND2_X1 U11307 ( .A1(n16249), .A2(n16292), .ZN(n16362) );
  NOR2_X1 U11308 ( .A1(n16069), .A2(n11513), .ZN(n11013) );
  AND2_X1 U11309 ( .A1(n10650), .A2(n16366), .ZN(n9601) );
  NOR2_X1 U11310 ( .A1(n9644), .A2(n18578), .ZN(n14728) );
  NAND2_X1 U11311 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18851), .ZN(
        n11930) );
  BUF_X2 U11312 ( .A(n16347), .Z(n9574) );
  CLKBUF_X1 U11313 ( .A(n15864), .Z(n9599) );
  INV_X1 U11314 ( .A(n11325), .ZN(n14002) );
  OR3_X1 U11315 ( .A1(n19596), .A2(n19595), .A3(n19734), .ZN(n19608) );
  AND2_X1 U11316 ( .A1(n14786), .A2(n14791), .ZN(n17098) );
  NAND2_X2 U11317 ( .A1(n20712), .A2(n12036), .ZN(n15328) );
  AOI21_X1 U11318 ( .B1(n10112), .B2(n14376), .A(n9604), .ZN(n10307) );
  AND2_X1 U11319 ( .A1(n17763), .A2(n13330), .ZN(n17753) );
  NAND2_X1 U11320 ( .A1(n15139), .A2(n13038), .ZN(n15121) );
  NOR2_X1 U11321 ( .A1(n18368), .A2(n14712), .ZN(n18366) );
  NAND2_X1 U11322 ( .A1(n10990), .A2(n10999), .ZN(n11005) );
  OR2_X1 U11323 ( .A1(n14657), .A2(n14608), .ZN(n14653) );
  NAND2_X1 U11324 ( .A1(n10177), .A2(n12132), .ZN(n12129) );
  NAND2_X2 U11325 ( .A1(n12836), .A2(n12835), .ZN(n14013) );
  XNOR2_X1 U11326 ( .A(n11658), .B(n11656), .ZN(n14159) );
  NAND2_X1 U11327 ( .A1(n12195), .A2(n12194), .ZN(n20893) );
  AND2_X2 U11328 ( .A1(n10984), .A2(n10965), .ZN(n10990) );
  NAND2_X1 U11329 ( .A1(n14798), .A2(n14797), .ZN(n14800) );
  NAND2_X1 U11330 ( .A1(n10582), .A2(n10044), .ZN(n10636) );
  NAND2_X1 U11331 ( .A1(n11639), .A2(n11638), .ZN(n11658) );
  NAND2_X1 U11332 ( .A1(n20959), .A2(n12193), .ZN(n10177) );
  NOR2_X2 U11333 ( .A1(n14531), .A2(n12998), .ZN(n14617) );
  INV_X2 U11334 ( .A(n18385), .ZN(n9564) );
  AND2_X1 U11335 ( .A1(n11069), .A2(n11068), .ZN(n14401) );
  AND2_X1 U11336 ( .A1(n17348), .A2(n11945), .ZN(n17314) );
  AND2_X1 U11337 ( .A1(n11052), .A2(n11051), .ZN(n14190) );
  NAND2_X1 U11338 ( .A1(n10628), .A2(n10627), .ZN(n11048) );
  AOI21_X1 U11339 ( .B1(n12818), .B2(n12817), .A(n12816), .ZN(n12832) );
  AND2_X1 U11340 ( .A1(n10626), .A2(n10625), .ZN(n10627) );
  NAND2_X1 U11341 ( .A1(n10595), .A2(n10594), .ZN(n10635) );
  OR2_X1 U11342 ( .A1(n12810), .A2(n12809), .ZN(n12818) );
  AND2_X1 U11343 ( .A1(n9933), .A2(n13810), .ZN(n9932) );
  NAND2_X1 U11344 ( .A1(n12988), .A2(n10453), .ZN(n14531) );
  OR2_X1 U11345 ( .A1(n17350), .A2(n14069), .ZN(n9902) );
  OR2_X1 U11346 ( .A1(n10373), .A2(n9606), .ZN(n10961) );
  INV_X1 U11347 ( .A(n12147), .ZN(n9770) );
  NAND2_X1 U11348 ( .A1(n12120), .A2(n12119), .ZN(n12147) );
  NAND2_X1 U11349 ( .A1(n14504), .A2(n14503), .ZN(n10222) );
  NAND2_X1 U11350 ( .A1(n19587), .A2(n11938), .ZN(n17350) );
  INV_X1 U11351 ( .A(n11084), .ZN(n13297) );
  AND2_X1 U11352 ( .A1(n10217), .A2(n9901), .ZN(n19587) );
  INV_X2 U11353 ( .A(n10614), .ZN(n11084) );
  XNOR2_X1 U11354 ( .A(n11679), .B(n11897), .ZN(n11675) );
  OAI21_X1 U11355 ( .B1(n12110), .B2(n15253), .A(n9767), .ZN(n12120) );
  INV_X1 U11356 ( .A(n9804), .ZN(n9803) );
  NOR2_X1 U11357 ( .A1(n11946), .A2(n14070), .ZN(n14024) );
  NOR2_X1 U11358 ( .A1(n10918), .A2(n10911), .ZN(n10910) );
  OR2_X1 U11359 ( .A1(n14152), .A2(n14157), .ZN(n10241) );
  NAND2_X1 U11360 ( .A1(n11598), .A2(n11597), .ZN(n11615) );
  AND2_X1 U11361 ( .A1(n11212), .A2(n13930), .ZN(n10110) );
  XNOR2_X1 U11362 ( .A(n13319), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13331) );
  OAI21_X1 U11363 ( .B1(n10589), .B2(n13189), .A(n10464), .ZN(n9804) );
  NAND2_X1 U11364 ( .A1(n9852), .A2(n9673), .ZN(n10589) );
  NAND2_X1 U11365 ( .A1(n11940), .A2(n11949), .ZN(n11946) );
  NOR2_X1 U11366 ( .A1(n17657), .A2(n11935), .ZN(n14023) );
  OR2_X1 U11367 ( .A1(n12218), .A2(n12219), .ZN(n12215) );
  AND2_X1 U11368 ( .A1(n11912), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11913) );
  AND2_X1 U11369 ( .A1(n9708), .A2(n9907), .ZN(n13096) );
  AND2_X1 U11370 ( .A1(n14333), .A2(n12088), .ZN(n12117) );
  NOR2_X1 U11371 ( .A1(n10137), .A2(n11279), .ZN(n10136) );
  OR2_X1 U11372 ( .A1(n14334), .A2(n12950), .ZN(n13089) );
  INV_X1 U11373 ( .A(n10571), .ZN(n13708) );
  AND3_X1 U11374 ( .A1(n14070), .A2(n11936), .A3(n9695), .ZN(n11843) );
  AND2_X1 U11375 ( .A1(n10587), .A2(n14046), .ZN(n10269) );
  INV_X1 U11376 ( .A(n10095), .ZN(n14114) );
  NOR2_X1 U11377 ( .A1(n18396), .A2(n19162), .ZN(n11846) );
  NOR2_X1 U11378 ( .A1(n11836), .A2(n18538), .ZN(n11847) );
  NOR2_X1 U11379 ( .A1(n11836), .A2(n19153), .ZN(n11949) );
  INV_X1 U11380 ( .A(n10586), .ZN(n19869) );
  AND2_X1 U11381 ( .A1(n10586), .A2(n19862), .ZN(n10558) );
  NAND2_X1 U11382 ( .A1(n18687), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18644) );
  INV_X1 U11383 ( .A(n10584), .ZN(n13347) );
  NOR2_X1 U11384 ( .A1(n12174), .A2(n14376), .ZN(n12929) );
  INV_X1 U11385 ( .A(n13177), .ZN(n10192) );
  AND2_X1 U11386 ( .A1(n10114), .A2(n20885), .ZN(n12113) );
  INV_X2 U11387 ( .A(n12815), .ZN(n12820) );
  AND2_X1 U11388 ( .A1(n10114), .A2(n9702), .ZN(n10115) );
  NAND2_X1 U11389 ( .A1(n10191), .A2(n13177), .ZN(n14333) );
  NAND2_X1 U11390 ( .A1(n12087), .A2(n12106), .ZN(n9761) );
  NAND2_X1 U11391 ( .A1(n10586), .A2(n11205), .ZN(n10596) );
  CLKBUF_X3 U11392 ( .A(n13719), .Z(n9590) );
  NAND2_X1 U11393 ( .A1(n14666), .A2(n14512), .ZN(n11904) );
  CLKBUF_X1 U11394 ( .A(n10584), .Z(n14046) );
  OR2_X1 U11395 ( .A1(n10681), .A2(n10680), .ZN(n11277) );
  CLKBUF_X1 U11396 ( .A(n12109), .Z(n15253) );
  NAND2_X1 U11397 ( .A1(n12091), .A2(n9584), .ZN(n12971) );
  OR2_X1 U11398 ( .A1(n11581), .A2(n11580), .ZN(n14512) );
  NAND4_X2 U11399 ( .A1(n10849), .A2(n10848), .A3(n10847), .A4(n10846), .ZN(
        n13293) );
  NAND2_X1 U11400 ( .A1(n12171), .A2(n20869), .ZN(n12815) );
  AND2_X1 U11401 ( .A1(n20869), .A2(n20885), .ZN(n12087) );
  INV_X2 U11402 ( .A(n10191), .ZN(n9565) );
  OR2_X1 U11403 ( .A1(n11612), .A2(n11611), .ZN(n14509) );
  NAND4_X2 U11404 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n19736) );
  NAND2_X1 U11405 ( .A1(n10319), .A2(n10318), .ZN(n14516) );
  AND2_X1 U11406 ( .A1(n9618), .A2(n9679), .ZN(n19162) );
  NAND2_X1 U11407 ( .A1(n9899), .A2(n9661), .ZN(n18538) );
  AND2_X1 U11408 ( .A1(n9972), .A2(n9970), .ZN(n10586) );
  OR2_X2 U11409 ( .A1(n11790), .A2(n11789), .ZN(n19171) );
  CLKBUF_X2 U11410 ( .A(n12081), .Z(n20878) );
  OR2_X1 U11411 ( .A1(n12170), .A2(n12169), .ZN(n12877) );
  OR2_X1 U11412 ( .A1(n12159), .A2(n12158), .ZN(n12932) );
  AND4_X1 U11413 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(
        n9610) );
  NAND2_X2 U11414 ( .A1(n10555), .A2(n10554), .ZN(n19895) );
  BUF_X2 U11415 ( .A(n12082), .Z(n20859) );
  AND3_X1 U11416 ( .A1(n10056), .A2(n9612), .A3(n9693), .ZN(n19157) );
  INV_X1 U11417 ( .A(n12086), .ZN(n12969) );
  NAND2_X1 U11418 ( .A1(n10544), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10275) );
  INV_X1 U11419 ( .A(n12359), .ZN(n12367) );
  OR2_X2 U11420 ( .A1(n12035), .A2(n12034), .ZN(n20885) );
  OR2_X2 U11421 ( .A1(n12025), .A2(n12024), .ZN(n12107) );
  NAND2_X1 U11422 ( .A1(n12007), .A2(n12006), .ZN(n12082) );
  NAND4_X2 U11423 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n12083) );
  NAND2_X1 U11424 ( .A1(n9971), .A2(n9669), .ZN(n10557) );
  NAND4_X1 U11425 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n11984), .ZN(
        n12086) );
  NAND2_X1 U11426 ( .A1(n10488), .A2(n10487), .ZN(n12081) );
  NAND2_X1 U11427 ( .A1(n10495), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10065) );
  NAND2_X1 U11428 ( .A1(n9969), .A2(n9968), .ZN(n11205) );
  NAND2_X1 U11429 ( .A1(n10501), .A2(n10669), .ZN(n10064) );
  AND4_X1 U11430 ( .A1(n11973), .A2(n11972), .A3(n11971), .A4(n11970), .ZN(
        n11986) );
  AND4_X1 U11431 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n11997) );
  AND2_X1 U11432 ( .A1(n10522), .A2(n10519), .ZN(n9971) );
  AND4_X1 U11433 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .ZN(
        n12057) );
  AND4_X1 U11434 ( .A1(n12067), .A2(n12066), .A3(n12065), .A4(n12064), .ZN(
        n12079) );
  AND3_X1 U11435 ( .A1(n12001), .A2(n12000), .A3(n10486), .ZN(n12007) );
  NAND2_X1 U11436 ( .A1(n17232), .A2(n10457), .ZN(n17212) );
  AND4_X1 U11437 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n12006) );
  AND3_X1 U11438 ( .A1(n10531), .A2(n10669), .A3(n10530), .ZN(n10532) );
  INV_X2 U11439 ( .A(n18325), .ZN(n17450) );
  AND4_X1 U11440 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n11996) );
  AND4_X1 U11441 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n10488) );
  AND4_X1 U11442 ( .A1(n12072), .A2(n12071), .A3(n12070), .A4(n12069), .ZN(
        n12078) );
  AND4_X1 U11443 ( .A1(n12040), .A2(n12039), .A3(n12038), .A4(n12037), .ZN(
        n12058) );
  AND4_X1 U11444 ( .A1(n11983), .A2(n11982), .A3(n11981), .A4(n11980), .ZN(
        n11984) );
  NOR2_X2 U11445 ( .A1(n20838), .A2(n20837), .ZN(n20839) );
  AND4_X1 U11446 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11985) );
  AND4_X1 U11447 ( .A1(n12076), .A2(n12075), .A3(n12074), .A4(n12073), .ZN(
        n12077) );
  AND4_X1 U11448 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12080) );
  AND4_X1 U11449 ( .A1(n12054), .A2(n12053), .A3(n12052), .A4(n12051), .ZN(
        n12055) );
  AND4_X1 U11450 ( .A1(n12049), .A2(n12048), .A3(n12047), .A4(n12046), .ZN(
        n12056) );
  AND4_X1 U11451 ( .A1(n11968), .A2(n11967), .A3(n11966), .A4(n11965), .ZN(
        n11987) );
  INV_X2 U11452 ( .A(n17638), .ZN(U215) );
  NAND2_X2 U11453 ( .A1(n19749), .A2(n19650), .ZN(n19706) );
  CLKBUF_X1 U11454 ( .A(n13506), .Z(n13636) );
  AND2_X2 U11455 ( .A1(n9595), .A2(n10669), .ZN(n13526) );
  BUF_X2 U11456 ( .A(n12264), .Z(n12752) );
  AND2_X1 U11457 ( .A1(n11560), .A2(n11559), .ZN(n11649) );
  AND2_X2 U11458 ( .A1(n11557), .A2(n11560), .ZN(n17465) );
  NAND2_X2 U11459 ( .A1(n11562), .A2(n11560), .ZN(n11727) );
  AND2_X2 U11460 ( .A1(n11557), .A2(n14033), .ZN(n18054) );
  AND2_X2 U11461 ( .A1(n14355), .A2(n10078), .ZN(n12747) );
  CLKBUF_X1 U11462 ( .A(n10668), .Z(n13511) );
  NOR2_X1 U11463 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18010), .ZN(n17984) );
  INV_X2 U11464 ( .A(n17641), .ZN(n17643) );
  AND2_X2 U11465 ( .A1(n10107), .A2(n14365), .ZN(n12754) );
  AND2_X2 U11466 ( .A1(n14556), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10668) );
  NOR2_X1 U11467 ( .A1(n18820), .A2(n18803), .ZN(n18805) );
  NAND2_X1 U11468 ( .A1(n14556), .A2(n14541), .ZN(n13549) );
  AND2_X2 U11469 ( .A1(n11964), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10111) );
  NOR2_X1 U11470 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n17345), .ZN(
        n11558) );
  AND2_X1 U11471 ( .A1(n14074), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11557) );
  AND2_X2 U11472 ( .A1(n11979), .A2(n14341), .ZN(n12244) );
  AND2_X1 U11473 ( .A1(n11969), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10078) );
  NOR2_X2 U11474 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10107) );
  INV_X1 U11475 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10489) );
  INV_X1 U11476 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9986) );
  CLKBUF_X1 U11477 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n17154) );
  AND2_X1 U11478 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17351) );
  NOR2_X2 U11479 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14033) );
  NAND2_X1 U11480 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14065) );
  NAND2_X1 U11481 ( .A1(n9763), .A2(n9600), .ZN(n10026) );
  AND4_X1 U11482 ( .A1(n12091), .A2(n20859), .A3(n10083), .A4(n20878), .ZN(
        n9609) );
  CLKBUF_X1 U11483 ( .A(n10109), .Z(n9568) );
  AND2_X1 U11484 ( .A1(n10070), .A2(n15506), .ZN(n15496) );
  AND2_X1 U11485 ( .A1(n16637), .A2(n10446), .ZN(n10445) );
  INV_X1 U11486 ( .A(n16700), .ZN(n9874) );
  NAND2_X1 U11487 ( .A1(n12220), .A2(n10467), .ZN(n12880) );
  NAND2_X1 U11488 ( .A1(n16823), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9569) );
  NAND2_X1 U11489 ( .A1(n16823), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16824) );
  AND2_X1 U11490 ( .A1(n10460), .A2(n10578), .ZN(n10098) );
  AND2_X1 U11491 ( .A1(n9578), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13533) );
  NAND2_X2 U11492 ( .A1(n9831), .A2(n16269), .ZN(n10942) );
  NOR2_X2 U11493 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17854), .ZN(n17835) );
  NAND2_X2 U11494 ( .A1(n14254), .A2(n12889), .ZN(n14520) );
  OAI21_X1 U11495 ( .B1(n9805), .B2(n13189), .A(n9803), .ZN(n10045) );
  AOI21_X1 U11496 ( .B1(n10152), .B2(n17136), .A(n10151), .ZN(n16885) );
  NAND2_X2 U11497 ( .A1(n12277), .A2(n12204), .ZN(n15867) );
  AOI211_X1 U11498 ( .C1(n13682), .C2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n13638), .B(n13637), .ZN(n13641) );
  OAI211_X1 U11499 ( .C1(n14841), .C2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10149), .B(n10148), .ZN(n14764) );
  NAND2_X1 U11500 ( .A1(n14841), .A2(n9634), .ZN(n10030) );
  NAND2_X1 U11501 ( .A1(n14841), .A2(n9637), .ZN(n10326) );
  INV_X1 U11502 ( .A(n12587), .ZN(n9570) );
  AND2_X1 U11503 ( .A1(n9571), .A2(n13762), .ZN(n15010) );
  NOR2_X1 U11504 ( .A1(n12619), .A2(n9570), .ZN(n9571) );
  AND2_X2 U11505 ( .A1(n14296), .A2(n14424), .ZN(n9572) );
  AND2_X2 U11506 ( .A1(n15220), .A2(n10387), .ZN(n13762) );
  AND2_X4 U11507 ( .A1(n10150), .A2(n14541), .ZN(n9589) );
  AND2_X1 U11508 ( .A1(n12084), .A2(n12969), .ZN(n13177) );
  INV_X1 U11509 ( .A(n12084), .ZN(n14861) );
  NAND4_X1 U11510 ( .A1(n10081), .A2(n13111), .A3(n12107), .A4(n12221), .ZN(
        n13941) );
  AND2_X1 U11511 ( .A1(n12111), .A2(n9585), .ZN(n13080) );
  OAI21_X1 U11512 ( .B1(n10644), .B2(n9838), .A(n10645), .ZN(n16347) );
  AND2_X2 U11513 ( .A1(n10662), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11346) );
  NAND2_X1 U11514 ( .A1(n10173), .A2(n9801), .ZN(n9791) );
  AND2_X2 U11515 ( .A1(n10670), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9575) );
  NAND3_X1 U11516 ( .A1(n13089), .A2(n10106), .A3(n10103), .ZN(n12101) );
  INV_X4 U11517 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14541) );
  OAI21_X1 U11518 ( .B1(n9917), .B2(n12901), .A(n9916), .ZN(n12892) );
  AND3_X4 U11519 ( .A1(n10490), .A2(n10489), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9576) );
  OR2_X1 U11520 ( .A1(n11944), .A2(n9695), .ZN(n17657) );
  INV_X2 U11521 ( .A(n18884), .ZN(n18900) );
  AND2_X4 U11522 ( .A1(n14556), .A2(n14541), .ZN(n9578) );
  AND2_X1 U11523 ( .A1(n14556), .A2(n14541), .ZN(n9579) );
  INV_X2 U11524 ( .A(n13549), .ZN(n13682) );
  AND2_X1 U11525 ( .A1(n12148), .A2(n12147), .ZN(n12193) );
  NAND2_X1 U11526 ( .A1(n12105), .A2(n12104), .ZN(n12148) );
  NOR2_X2 U11527 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17779), .ZN(n17762) );
  AND2_X1 U11528 ( .A1(n12216), .A2(n12215), .ZN(n12220) );
  NOR2_X1 U11529 ( .A1(n12107), .A2(n20859), .ZN(n12093) );
  NAND2_X1 U11530 ( .A1(n10233), .A2(n10232), .ZN(n13868) );
  OAI21_X1 U11531 ( .B1(n15041), .B2(n13765), .A(n13764), .ZN(n15472) );
  OAI211_X2 U11532 ( .C1(n17503), .C2(n17508), .A(n12927), .B(n12926), .ZN(
        n12928) );
  AND2_X2 U11533 ( .A1(n11562), .A2(n17351), .ZN(n11628) );
  INV_X2 U11534 ( .A(n15595), .ZN(n9581) );
  AND2_X4 U11535 ( .A1(n9906), .A2(n12930), .ZN(n15595) );
  OR2_X1 U11536 ( .A1(n15870), .A2(n15871), .ZN(n21211) );
  NOR2_X4 U11537 ( .A1(n18644), .A2(n18647), .ZN(n13313) );
  INV_X4 U11538 ( .A(n9590), .ZN(n10902) );
  OAI21_X1 U11539 ( .B1(n14973), .B2(n14963), .A(n14962), .ZN(n15343) );
  XNOR2_X1 U11540 ( .A(n14962), .B(n10015), .ZN(n14950) );
  NAND2_X4 U11541 ( .A1(n10065), .A2(n10064), .ZN(n9594) );
  NAND2_X2 U11542 ( .A1(n12129), .A2(n12130), .ZN(n12232) );
  INV_X2 U11543 ( .A(n18325), .ZN(n9582) );
  NOR2_X2 U11544 ( .A1(n13941), .A2(n12036), .ZN(n12949) );
  AND2_X2 U11545 ( .A1(n14297), .A2(n14298), .ZN(n14296) );
  NAND4_X1 U11546 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n9584) );
  NAND4_X1 U11547 ( .A1(n12058), .A2(n12057), .A3(n12056), .A4(n12055), .ZN(
        n9585) );
  AND2_X4 U11548 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14556) );
  NOR2_X2 U11549 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17718), .ZN(n17717) );
  AND2_X1 U11550 ( .A1(n10670), .A2(n14541), .ZN(n9586) );
  AND2_X1 U11551 ( .A1(n10670), .A2(n14541), .ZN(n9587) );
  INV_X1 U11552 ( .A(n9586), .ZN(n9588) );
  AND2_X1 U11553 ( .A1(n13750), .A2(n14961), .ZN(n14973) );
  INV_X1 U11554 ( .A(n18824), .ZN(n18749) );
  NAND2_X2 U11555 ( .A1(n12201), .A2(n12200), .ZN(n12202) );
  BUF_X4 U11556 ( .A(n16405), .Z(n9593) );
  INV_X1 U11557 ( .A(n11279), .ZN(n16405) );
  AOI211_X2 U11558 ( .C1(n19610), .C2(n19609), .A(n19608), .B(n19607), .ZN(
        n19624) );
  XNOR2_X2 U11559 ( .A(n10942), .B(n17100), .ZN(n16819) );
  XNOR2_X1 U11560 ( .A(n14098), .B(n14100), .ZN(n20578) );
  INV_X1 U11561 ( .A(n10496), .ZN(n9596) );
  AND2_X1 U11562 ( .A1(n10047), .A2(n10648), .ZN(n20046) );
  AND3_X1 U11563 ( .A1(n10648), .A2(n10658), .A3(n13361), .ZN(n10806) );
  XNOR2_X2 U11564 ( .A(n13609), .B(n13593), .ZN(n16400) );
  OAI21_X2 U11565 ( .B1(n16423), .B2(n9632), .A(n13575), .ZN(n13609) );
  AND2_X1 U11566 ( .A1(n10111), .A2(n14341), .ZN(n9597) );
  AND2_X1 U11567 ( .A1(n10111), .A2(n14341), .ZN(n9598) );
  NOR2_X4 U11568 ( .A1(n13320), .A2(n13321), .ZN(n17232) );
  AND2_X1 U11569 ( .A1(n19895), .A2(n20607), .ZN(n11288) );
  NAND2_X1 U11570 ( .A1(n11034), .A2(n16630), .ZN(n10006) );
  NAND2_X1 U11571 ( .A1(n12092), .A2(n9761), .ZN(n12957) );
  NAND2_X1 U11572 ( .A1(n10014), .A2(n9672), .ZN(n10012) );
  AND3_X1 U11573 ( .A1(n9671), .A2(n12838), .A3(n12837), .ZN(n13178) );
  AND4_X1 U11574 ( .A1(n10837), .A2(n10836), .A3(n10835), .A4(n10834), .ZN(
        n10848) );
  NAND2_X1 U11575 ( .A1(n10829), .A2(n10824), .ZN(n10179) );
  INV_X1 U11576 ( .A(n11307), .ZN(n11462) );
  NOR2_X1 U11577 ( .A1(n11279), .A2(n9594), .ZN(n11273) );
  NOR2_X1 U11578 ( .A1(n10648), .A2(n16366), .ZN(n10334) );
  AOI21_X1 U11579 ( .B1(n20016), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A(n9687), .ZN(n10778) );
  AOI22_X1 U11580 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9675), .B2(n10657), .ZN(n10272) );
  NAND2_X1 U11581 ( .A1(n20324), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10128) );
  INV_X1 U11582 ( .A(n15203), .ZN(n10389) );
  NAND2_X1 U11583 ( .A1(n12296), .A2(n12295), .ZN(n12899) );
  AND2_X1 U11584 ( .A1(n15551), .A2(n9915), .ZN(n9764) );
  INV_X1 U11585 ( .A(n12203), .ZN(n10033) );
  INV_X1 U11586 ( .A(n12082), .ZN(n13111) );
  OAI21_X1 U11587 ( .B1(n10575), .B2(n19875), .A(n10529), .ZN(n9839) );
  INV_X1 U11588 ( .A(n11038), .ZN(n10356) );
  INV_X1 U11589 ( .A(n16607), .ZN(n10357) );
  NOR2_X1 U11590 ( .A1(n10267), .A2(n10266), .ZN(n10265) );
  INV_X1 U11591 ( .A(n10744), .ZN(n10267) );
  AND3_X1 U11592 ( .A1(n11246), .A2(n11208), .A3(n11207), .ZN(n11241) );
  NAND2_X1 U11593 ( .A1(n10584), .A2(n9594), .ZN(n10575) );
  NAND2_X1 U11594 ( .A1(n9836), .A2(n9835), .ZN(n10574) );
  OR2_X1 U11595 ( .A1(n11660), .A2(n18524), .ZN(n11679) );
  INV_X1 U11596 ( .A(n19157), .ZN(n10055) );
  INV_X1 U11597 ( .A(n10084), .ZN(n12112) );
  NAND2_X1 U11598 ( .A1(n9889), .A2(n9887), .ZN(n9943) );
  NAND2_X1 U11599 ( .A1(n15477), .A2(n10024), .ZN(n9889) );
  NOR2_X1 U11600 ( .A1(n9888), .A2(n9686), .ZN(n9887) );
  OR2_X1 U11601 ( .A1(n15583), .A2(n15716), .ZN(n12946) );
  AND2_X1 U11602 ( .A1(n12946), .A2(n10431), .ZN(n9602) );
  NAND2_X1 U11603 ( .A1(n10434), .A2(n9750), .ZN(n10431) );
  OR2_X1 U11604 ( .A1(n13178), .A2(n12958), .ZN(n12960) );
  NAND2_X1 U11605 ( .A1(n13347), .A2(n9594), .ZN(n10580) );
  NOR2_X1 U11606 ( .A1(n11165), .A2(n11166), .ZN(n11511) );
  NOR2_X1 U11607 ( .A1(n10944), .A2(n10369), .ZN(n10368) );
  NAND2_X1 U11608 ( .A1(n10908), .A2(n10370), .ZN(n10369) );
  AND2_X1 U11609 ( .A1(n10947), .A2(n14272), .ZN(n10370) );
  AND2_X1 U11610 ( .A1(n13225), .A2(n9742), .ZN(n13232) );
  NAND2_X1 U11611 ( .A1(n10110), .A2(n10109), .ZN(n9841) );
  NAND2_X1 U11612 ( .A1(n9685), .A2(n9605), .ZN(n9850) );
  OAI21_X1 U11613 ( .B1(n16577), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16595), .ZN(n11162) );
  INV_X1 U11614 ( .A(n16090), .ZN(n10409) );
  NOR2_X1 U11615 ( .A1(n13158), .A2(n10420), .ZN(n10419) );
  INV_X1 U11616 ( .A(n10959), .ZN(n10420) );
  INV_X1 U11617 ( .A(n14383), .ZN(n10347) );
  INV_X1 U11618 ( .A(n14406), .ZN(n10392) );
  NAND2_X1 U11619 ( .A1(n16766), .A2(n10955), .ZN(n10960) );
  AND2_X1 U11620 ( .A1(n16767), .A2(n16768), .ZN(n10955) );
  NAND2_X1 U11621 ( .A1(n9992), .A2(n10827), .ZN(n9954) );
  NAND2_X1 U11622 ( .A1(n14186), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13377) );
  NAND2_X1 U11623 ( .A1(n13376), .A2(n13375), .ZN(n13379) );
  OR2_X1 U11624 ( .A1(n10648), .A2(n13371), .ZN(n13376) );
  NAND2_X1 U11625 ( .A1(n10569), .A2(n10669), .ZN(n10274) );
  NAND2_X1 U11626 ( .A1(n10563), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10273) );
  NAND2_X1 U11627 ( .A1(n9825), .A2(n9601), .ZN(n19904) );
  AND2_X1 U11628 ( .A1(n10648), .A2(n14784), .ZN(n9825) );
  AND2_X1 U11629 ( .A1(n10648), .A2(n13361), .ZN(n10048) );
  NOR2_X1 U11630 ( .A1(n10156), .A2(n13361), .ZN(n20237) );
  NAND2_X1 U11631 ( .A1(n10556), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9972) );
  NAND2_X1 U11632 ( .A1(n10557), .A2(n10669), .ZN(n9970) );
  NAND3_X1 U11633 ( .A1(n11846), .A2(n9681), .A3(n11847), .ZN(n11944) );
  INV_X1 U11634 ( .A(n19587), .ZN(n11948) );
  OR2_X1 U11635 ( .A1(n11916), .A2(n11915), .ZN(n11917) );
  INV_X1 U11636 ( .A(n14344), .ZN(n13944) );
  NAND2_X1 U11637 ( .A1(n12834), .A2(n12833), .ZN(n12835) );
  INV_X1 U11638 ( .A(n12847), .ZN(n12833) );
  NAND2_X1 U11639 ( .A1(n13750), .A2(n13749), .ZN(n14855) );
  AOI21_X1 U11640 ( .B1(n12915), .B2(n12464), .A(n12334), .ZN(n15326) );
  NAND2_X1 U11641 ( .A1(n12279), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12299) );
  NAND2_X1 U11642 ( .A1(n12971), .A2(n12108), .ZN(n10095) );
  NAND2_X1 U11643 ( .A1(n9943), .A2(n13752), .ZN(n15435) );
  NOR2_X1 U11644 ( .A1(n9817), .A2(n9816), .ZN(n9815) );
  INV_X1 U11645 ( .A(n15538), .ZN(n9816) );
  INV_X1 U11646 ( .A(n15539), .ZN(n9817) );
  NAND2_X1 U11647 ( .A1(n13101), .A2(n10192), .ZN(n12968) );
  NAND2_X1 U11648 ( .A1(n11511), .A2(n11510), .ZN(n13290) );
  NOR2_X1 U11649 ( .A1(n15959), .A2(n16583), .ZN(n15949) );
  NAND2_X1 U11650 ( .A1(n10946), .A2(n10902), .ZN(n11043) );
  NAND2_X1 U11651 ( .A1(n10992), .A2(n11043), .ZN(n10984) );
  INV_X1 U11652 ( .A(n16617), .ZN(n10146) );
  AND4_X1 U11653 ( .A1(n10833), .A2(n10832), .A3(n10831), .A4(n10830), .ZN(
        n10849) );
  OR2_X1 U11654 ( .A1(n9624), .A2(n16597), .ZN(n9862) );
  AND2_X1 U11655 ( .A1(n9624), .A2(n16595), .ZN(n9858) );
  NAND2_X1 U11656 ( .A1(n10146), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10144) );
  AND2_X1 U11657 ( .A1(n14842), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10053) );
  NAND2_X1 U11658 ( .A1(n14841), .A2(n14842), .ZN(n16637) );
  NAND2_X1 U11659 ( .A1(n14841), .A2(n10158), .ZN(n16661) );
  AND2_X1 U11660 ( .A1(n11505), .A2(n11254), .ZN(n13164) );
  AND3_X1 U11661 ( .A1(n11362), .A2(n11361), .A3(n11360), .ZN(n14079) );
  AND2_X1 U11662 ( .A1(n13361), .A2(n9601), .ZN(n10047) );
  NOR2_X1 U11663 ( .A1(n14784), .A2(n9574), .ZN(n10653) );
  INV_X1 U11664 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17141) );
  NAND2_X1 U11665 ( .A1(n18818), .A2(n14733), .ZN(n9811) );
  OAI211_X1 U11666 ( .C1(n16571), .C2(n16304), .A(n15956), .B(n10287), .ZN(
        n10286) );
  AOI21_X1 U11667 ( .B1(n16359), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15948), .ZN(n10287) );
  NAND2_X1 U11668 ( .A1(n10331), .A2(n16864), .ZN(n10330) );
  AND2_X1 U11669 ( .A1(n10443), .A2(n9895), .ZN(n9891) );
  INV_X1 U11670 ( .A(n14900), .ZN(n9895) );
  OAI211_X1 U11671 ( .C1(n12781), .C2(n10192), .A(n12799), .B(n12780), .ZN(
        n12782) );
  NAND2_X1 U11672 ( .A1(n20878), .A2(n14861), .ZN(n10114) );
  NAND2_X1 U11673 ( .A1(n10779), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10131) );
  AOI22_X1 U11674 ( .A1(n20182), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n20237), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10777) );
  NAND2_X1 U11675 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10132) );
  OR2_X1 U11676 ( .A1(n9627), .A2(n9711), .ZN(n10097) );
  NAND2_X1 U11677 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10203) );
  NAND2_X1 U11678 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10195) );
  NAND2_X1 U11679 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10214) );
  INV_X1 U11680 ( .A(n15514), .ZN(n9882) );
  NAND2_X1 U11681 ( .A1(n15539), .A2(n9884), .ZN(n9883) );
  AND2_X1 U11682 ( .A1(n15512), .A2(n12945), .ZN(n9884) );
  AND2_X1 U11683 ( .A1(n9584), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12171) );
  XNOR2_X1 U11684 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12813) );
  INV_X1 U11685 ( .A(n10074), .ZN(n9910) );
  OAI21_X1 U11686 ( .B1(n12901), .B2(n12900), .A(n10471), .ZN(n9819) );
  INV_X1 U11687 ( .A(n12884), .ZN(n10235) );
  INV_X1 U11688 ( .A(n12189), .ZN(n12239) );
  NAND2_X1 U11689 ( .A1(n9768), .A2(n15253), .ZN(n9767) );
  AOI22_X1 U11690 ( .A1(n13094), .A2(n20854), .B1(n13093), .B2(n10192), .ZN(
        n13095) );
  NOR2_X1 U11691 ( .A1(n12083), .A2(n14376), .ZN(n12189) );
  NAND2_X1 U11692 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12054) );
  NAND2_X1 U11693 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12072) );
  AOI22_X1 U11694 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12063), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U11695 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U11696 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12747), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12009) );
  NAND3_X1 U11697 ( .A1(n10721), .A2(n10722), .A3(n10456), .ZN(n9802) );
  INV_X1 U11698 ( .A(n18518), .ZN(n11897) );
  INV_X1 U11699 ( .A(n14516), .ZN(n11898) );
  NAND2_X1 U11700 ( .A1(n14516), .A2(n14666), .ZN(n11617) );
  NOR2_X1 U11701 ( .A1(n12086), .A2(n12084), .ZN(n10081) );
  NAND2_X1 U11702 ( .A1(n12829), .A2(n12828), .ZN(n12847) );
  OR2_X1 U11703 ( .A1(n12826), .A2(n12825), .ZN(n12829) );
  AND2_X1 U11704 ( .A1(n10452), .A2(n9728), .ZN(n10388) );
  NAND2_X1 U11705 ( .A1(n10113), .A2(n10439), .ZN(n12881) );
  AND2_X1 U11706 ( .A1(n12876), .A2(n10440), .ZN(n10439) );
  OR2_X1 U11707 ( .A1(n20885), .A2(n21373), .ZN(n12765) );
  AOI21_X1 U11708 ( .B1(n9941), .B2(n13126), .A(n15637), .ZN(n9942) );
  INV_X1 U11709 ( .A(n13752), .ZN(n9941) );
  INV_X1 U11710 ( .A(n15661), .ZN(n10075) );
  NOR2_X1 U11711 ( .A1(n13055), .A2(n10126), .ZN(n10125) );
  INV_X1 U11712 ( .A(n15043), .ZN(n10126) );
  NAND2_X1 U11713 ( .A1(n12321), .A2(n9920), .ZN(n10035) );
  NOR2_X1 U11714 ( .A1(n12320), .A2(n12319), .ZN(n12321) );
  NAND2_X1 U11715 ( .A1(n20878), .A2(n20885), .ZN(n12950) );
  NAND2_X1 U11716 ( .A1(n10086), .A2(n10190), .ZN(n10085) );
  INV_X1 U11717 ( .A(n14333), .ZN(n10086) );
  INV_X1 U11718 ( .A(n12081), .ZN(n12221) );
  NAND2_X1 U11719 ( .A1(n12223), .A2(n14376), .ZN(n12216) );
  NAND2_X1 U11720 ( .A1(n12128), .A2(n12127), .ZN(n12130) );
  NOR2_X1 U11721 ( .A1(n12036), .A2(n10083), .ZN(n10233) );
  OR2_X1 U11722 ( .A1(n10709), .A2(n10708), .ZN(n10873) );
  NAND2_X1 U11723 ( .A1(n11160), .A2(n11043), .ZN(n11157) );
  NAND2_X1 U11724 ( .A1(n11030), .A2(n11043), .ZN(n11029) );
  NOR2_X1 U11725 ( .A1(n10377), .A2(n10973), .ZN(n10376) );
  NAND2_X1 U11726 ( .A1(n10470), .A2(n16431), .ZN(n10377) );
  AND2_X1 U11727 ( .A1(n10962), .A2(n10964), .ZN(n10365) );
  AND2_X1 U11728 ( .A1(n11477), .A2(n14824), .ZN(n14825) );
  NOR2_X1 U11729 ( .A1(n10399), .A2(n14675), .ZN(n10398) );
  INV_X1 U11730 ( .A(n14659), .ZN(n10399) );
  AND2_X1 U11731 ( .A1(n11241), .A2(n11240), .ZN(n14206) );
  AND2_X1 U11732 ( .A1(n14844), .A2(n14817), .ZN(n14843) );
  OR2_X1 U11733 ( .A1(n16126), .A2(n11513), .ZN(n11019) );
  NAND2_X1 U11734 ( .A1(n16575), .A2(n11163), .ZN(n13285) );
  AOI21_X1 U11735 ( .B1(n16579), .B2(n16582), .A(n13280), .ZN(n13283) );
  INV_X1 U11736 ( .A(n16613), .ZN(n10354) );
  INV_X1 U11737 ( .A(n11035), .ZN(n10358) );
  INV_X1 U11738 ( .A(n14689), .ZN(n10410) );
  INV_X1 U11739 ( .A(n16702), .ZN(n10418) );
  INV_X1 U11740 ( .A(n14400), .ZN(n10393) );
  INV_X1 U11741 ( .A(n13293), .ZN(n11513) );
  NAND2_X1 U11742 ( .A1(n10935), .A2(n17110), .ZN(n10940) );
  NAND4_X1 U11743 ( .A1(n10185), .A2(n9654), .A3(n10188), .A4(n10184), .ZN(
        n10183) );
  AND2_X1 U11744 ( .A1(n9951), .A2(n10828), .ZN(n9950) );
  NOR2_X1 U11745 ( .A1(n10933), .A2(n9848), .ZN(n9847) );
  INV_X1 U11746 ( .A(n16313), .ZN(n9848) );
  NAND2_X1 U11747 ( .A1(n9829), .A2(n10756), .ZN(n9844) );
  OR2_X1 U11748 ( .A1(n10740), .A2(n10739), .ZN(n10741) );
  NAND2_X1 U11749 ( .A1(n9692), .A2(n10858), .ZN(n10109) );
  INV_X1 U11750 ( .A(n10619), .ZN(n10639) );
  AND2_X1 U11751 ( .A1(n10897), .A2(n10896), .ZN(n11220) );
  AND2_X1 U11752 ( .A1(n11505), .A2(n14206), .ZN(n11258) );
  NAND2_X1 U11753 ( .A1(n13348), .A2(n20607), .ZN(n13374) );
  NAND2_X1 U11754 ( .A1(n14186), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13366) );
  INV_X1 U11755 ( .A(n10644), .ZN(n10650) );
  AND2_X1 U11756 ( .A1(n16366), .A2(n10644), .ZN(n10658) );
  AOI22_X1 U11757 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10510) );
  INV_X1 U11758 ( .A(n14582), .ZN(n14565) );
  AOI21_X1 U11759 ( .B1(n9561), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(n9946), 
        .ZN(n11592) );
  AND2_X1 U11760 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n9946) );
  NAND2_X1 U11761 ( .A1(n11680), .A2(n18518), .ZN(n11695) );
  NAND2_X1 U11762 ( .A1(n11900), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11899) );
  AND2_X1 U11763 ( .A1(n11845), .A2(n11844), .ZN(n11943) );
  AND2_X1 U11764 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11552) );
  NAND2_X1 U11765 ( .A1(n12107), .A2(n12111), .ZN(n12108) );
  AND2_X1 U11766 ( .A1(n13177), .A2(n10190), .ZN(n12956) );
  OR2_X1 U11767 ( .A1(n21521), .A2(n13770), .ZN(n15270) );
  INV_X1 U11768 ( .A(n21521), .ZN(n15261) );
  OR2_X1 U11769 ( .A1(n15400), .A2(n12950), .ZN(n12861) );
  OR3_X1 U11770 ( .A1(n14013), .A2(n15940), .A3(n13868), .ZN(n14448) );
  AND2_X1 U11771 ( .A1(n21373), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12771) );
  AND2_X1 U11772 ( .A1(n12586), .A2(n15099), .ZN(n12587) );
  NAND2_X1 U11773 ( .A1(n13762), .A2(n15099), .ZN(n15098) );
  AND2_X1 U11774 ( .A1(n12485), .A2(n12484), .ZN(n15112) );
  NAND2_X1 U11775 ( .A1(n10014), .A2(n10013), .ZN(n10011) );
  NAND2_X1 U11776 ( .A1(n12324), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12330) );
  NAND2_X1 U11777 ( .A1(n9622), .A2(n12464), .ZN(n9766) );
  NAND2_X1 U11778 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12255) );
  NAND2_X1 U11779 ( .A1(n14257), .A2(n12231), .ZN(n14298) );
  OAI21_X1 U11780 ( .B1(n12277), .B2(n10386), .A(n10381), .ZN(n14259) );
  INV_X1 U11781 ( .A(n10384), .ZN(n10383) );
  NAND2_X1 U11782 ( .A1(n14976), .A2(n14964), .ZN(n14932) );
  AOI22_X1 U11783 ( .A1(n14934), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n10095), .ZN(n14933) );
  NAND2_X1 U11784 ( .A1(n9943), .A2(n9885), .ZN(n13172) );
  AND2_X1 U11785 ( .A1(n13752), .A2(n9886), .ZN(n9885) );
  INV_X1 U11786 ( .A(n15645), .ZN(n9886) );
  AND2_X1 U11787 ( .A1(n9581), .A2(n15642), .ZN(n10039) );
  AOI21_X1 U11788 ( .B1(n10043), .B2(n15583), .A(n15642), .ZN(n10041) );
  NAND2_X1 U11789 ( .A1(n15426), .A2(n9631), .ZN(n10040) );
  NAND2_X1 U11790 ( .A1(n10026), .A2(n10024), .ZN(n15441) );
  INV_X1 U11791 ( .A(n10432), .ZN(n9914) );
  NAND2_X1 U11792 ( .A1(n13060), .A2(n10094), .ZN(n13772) );
  NAND2_X1 U11793 ( .A1(n14114), .A2(n15716), .ZN(n10094) );
  NOR2_X1 U11794 ( .A1(n15104), .A2(n15084), .ZN(n13044) );
  INV_X1 U11795 ( .A(n15121), .ZN(n13045) );
  NAND2_X1 U11796 ( .A1(n15595), .A2(n10088), .ZN(n15516) );
  NAND2_X1 U11797 ( .A1(n15552), .A2(n9648), .ZN(n15540) );
  NAND2_X1 U11798 ( .A1(n15595), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15549) );
  INV_X1 U11799 ( .A(n10437), .ZN(n10436) );
  OAI21_X1 U11800 ( .B1(n9650), .B2(n10438), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10437) );
  INV_X1 U11801 ( .A(n12879), .ZN(n10438) );
  INV_X1 U11802 ( .A(n15284), .ZN(n21329) );
  INV_X1 U11803 ( .A(n21211), .ZN(n21204) );
  OAI21_X1 U11804 ( .B1(n21526), .B2(n14378), .A(n15931), .ZN(n14375) );
  NOR2_X1 U11805 ( .A1(n21174), .A2(n21000), .ZN(n21336) );
  OR2_X1 U11806 ( .A1(n9599), .A2(n12880), .ZN(n21301) );
  INV_X1 U11807 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21372) );
  INV_X1 U11808 ( .A(n12083), .ZN(n10190) );
  NOR2_X1 U11809 ( .A1(n21000), .A2(n21248), .ZN(n20884) );
  OR2_X1 U11810 ( .A1(n15867), .A2(n15873), .ZN(n21379) );
  XNOR2_X1 U11811 ( .A(n13290), .B(n11512), .ZN(n13273) );
  AOI21_X1 U11812 ( .B1(n15949), .B2(n16567), .A(n13243), .ZN(n14756) );
  XNOR2_X1 U11813 ( .A(n11511), .B(n11172), .ZN(n15950) );
  AND2_X1 U11814 ( .A1(n16589), .A2(n15993), .ZN(n10295) );
  NAND2_X1 U11815 ( .A1(n10367), .A2(n9723), .ZN(n16008) );
  NAND2_X1 U11816 ( .A1(n16249), .A2(n9617), .ZN(n16025) );
  OR2_X1 U11817 ( .A1(n13231), .A2(n10284), .ZN(n9617) );
  INV_X1 U11818 ( .A(n11041), .ZN(n10367) );
  INV_X1 U11819 ( .A(n16008), .ZN(n16028) );
  INV_X1 U11820 ( .A(n10985), .ZN(n10963) );
  NAND2_X1 U11821 ( .A1(n10908), .A2(n10947), .ZN(n10372) );
  NOR2_X1 U11822 ( .A1(n10944), .A2(n10371), .ZN(n10008) );
  AND2_X1 U11823 ( .A1(n13243), .A2(n16292), .ZN(n16358) );
  AND2_X1 U11824 ( .A1(n11227), .A2(n11226), .ZN(n15974) );
  NOR2_X1 U11825 ( .A1(n15966), .A2(n11517), .ZN(n11520) );
  AND2_X1 U11826 ( .A1(n16103), .A2(n10349), .ZN(n16015) );
  AND2_X1 U11827 ( .A1(n9718), .A2(n10350), .ZN(n10349) );
  INV_X1 U11828 ( .A(n16013), .ZN(n10350) );
  NOR2_X1 U11829 ( .A1(n10346), .A2(n10344), .ZN(n10343) );
  INV_X1 U11830 ( .A(n16154), .ZN(n10344) );
  AND2_X1 U11831 ( .A1(n11466), .A2(n11465), .ZN(n16132) );
  NAND2_X1 U11832 ( .A1(n14197), .A2(n14198), .ZN(n9779) );
  XNOR2_X1 U11833 ( .A(n10282), .B(n14758), .ZN(n13303) );
  NAND2_X1 U11834 ( .A1(n13246), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10282) );
  AND2_X1 U11835 ( .A1(n11115), .A2(n11114), .ZN(n16053) );
  AND2_X1 U11836 ( .A1(n11063), .A2(n11062), .ZN(n14417) );
  AND2_X1 U11837 ( .A1(n11053), .A2(n11048), .ZN(n10406) );
  INV_X1 U11838 ( .A(n11297), .ZN(n13734) );
  NAND2_X1 U11839 ( .A1(n11520), .A2(n11519), .ZN(n13736) );
  OR2_X1 U11840 ( .A1(n10362), .A2(n9625), .ZN(n10361) );
  INV_X1 U11841 ( .A(n10360), .ZN(n10359) );
  AOI21_X1 U11842 ( .B1(n9828), .B2(n10853), .A(n10332), .ZN(n9806) );
  INV_X1 U11843 ( .A(n10856), .ZN(n10332) );
  NAND2_X1 U11844 ( .A1(n9960), .A2(n16609), .ZN(n9959) );
  NAND2_X1 U11845 ( .A1(n16632), .A2(n9962), .ZN(n9961) );
  NOR2_X1 U11846 ( .A1(n16627), .A2(n9963), .ZN(n9962) );
  NAND2_X1 U11847 ( .A1(n16637), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10443) );
  NAND2_X1 U11848 ( .A1(n14841), .A2(n9754), .ZN(n16654) );
  OR2_X1 U11849 ( .A1(n11015), .A2(n16939), .ZN(n16651) );
  OAI21_X1 U11850 ( .B1(n9975), .B2(n9737), .A(n9974), .ZN(n16648) );
  NAND2_X1 U11851 ( .A1(n16663), .A2(n13161), .ZN(n9974) );
  INV_X1 U11852 ( .A(n16663), .ZN(n9976) );
  NAND2_X1 U11853 ( .A1(n10423), .A2(n13157), .ZN(n16705) );
  AND3_X1 U11854 ( .A1(n11431), .A2(n11430), .A3(n11429), .ZN(n14383) );
  NAND2_X1 U11855 ( .A1(n9608), .A2(n10391), .ZN(n10390) );
  INV_X1 U11856 ( .A(n14326), .ZN(n10391) );
  INV_X1 U11857 ( .A(n16606), .ZN(n16714) );
  AND3_X1 U11858 ( .A1(n11344), .A2(n11343), .A3(n11342), .ZN(n14041) );
  AND3_X1 U11859 ( .A1(n9734), .A2(n11252), .A3(n11251), .ZN(n14535) );
  AND2_X1 U11860 ( .A1(n13508), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14202) );
  INV_X1 U11861 ( .A(n20010), .ZN(n20077) );
  INV_X1 U11862 ( .A(n20178), .ZN(n20136) );
  NOR2_X1 U11863 ( .A1(n20237), .A2(n20236), .ZN(n20245) );
  NOR2_X2 U11864 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20606) );
  AND2_X1 U11865 ( .A1(n20578), .A2(n20009), .ZN(n20332) );
  INV_X1 U11866 ( .A(n20419), .ZN(n20328) );
  NOR3_X1 U11867 ( .A1(n20324), .A2(n20365), .A3(n20326), .ZN(n20327) );
  INV_X1 U11868 ( .A(n20332), .ZN(n20334) );
  INV_X1 U11869 ( .A(n20251), .ZN(n20335) );
  AND2_X1 U11870 ( .A1(n20578), .A2(n20585), .ZN(n20361) );
  NAND2_X1 U11871 ( .A1(n10442), .A2(n13361), .ZN(n20417) );
  INV_X1 U11872 ( .A(n20417), .ZN(n10779) );
  INV_X1 U11873 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n10224) );
  AND2_X1 U11874 ( .A1(n18164), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n18147) );
  AND2_X1 U11875 ( .A1(n14710), .A2(n19743), .ZN(n10221) );
  INV_X1 U11876 ( .A(n19162), .ZN(n10218) );
  NAND2_X1 U11877 ( .A1(n14507), .A2(n14506), .ZN(n18395) );
  AND2_X1 U11878 ( .A1(n10222), .A2(n19743), .ZN(n14711) );
  NOR2_X1 U11879 ( .A1(n11808), .A2(n9900), .ZN(n9899) );
  XNOR2_X1 U11880 ( .A(n11722), .B(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17189) );
  AOI21_X1 U11881 ( .B1(n10322), .B2(n9616), .A(n9929), .ZN(n9928) );
  NAND2_X1 U11882 ( .A1(n10469), .A2(n9930), .ZN(n9929) );
  NAND2_X1 U11883 ( .A1(n9636), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9930) );
  NAND2_X1 U11884 ( .A1(n10252), .A2(n10250), .ZN(n18947) );
  AOI21_X1 U11885 ( .B1(n10253), .B2(n9743), .A(n10251), .ZN(n10250) );
  INV_X1 U11886 ( .A(n19077), .ZN(n10253) );
  OR2_X1 U11887 ( .A1(n10316), .A2(n11704), .ZN(n10324) );
  NAND2_X1 U11888 ( .A1(n11702), .A2(n21579), .ZN(n14385) );
  NAND2_X1 U11889 ( .A1(n11919), .A2(n10240), .ZN(n10239) );
  INV_X1 U11890 ( .A(n14152), .ZN(n10240) );
  OR2_X1 U11891 ( .A1(n13808), .A2(n14157), .ZN(n10243) );
  AND2_X1 U11892 ( .A1(n9695), .A2(n10218), .ZN(n11888) );
  AND2_X1 U11893 ( .A1(n11887), .A2(n11886), .ZN(n19592) );
  INV_X1 U11894 ( .A(n19585), .ZN(n19077) );
  AND4_X1 U11895 ( .A1(n11823), .A2(n11822), .A3(n11821), .A4(n11820), .ZN(
        n11833) );
  AND4_X1 U11896 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(
        n11834) );
  OR2_X1 U11897 ( .A1(n13141), .A2(n14934), .ZN(n13142) );
  NOR2_X2 U11898 ( .A1(n12861), .A2(n20838), .ZN(n15393) );
  INV_X1 U11899 ( .A(n15387), .ZN(n15392) );
  NAND2_X1 U11900 ( .A1(n20721), .A2(n9585), .ZN(n20713) );
  INV_X1 U11901 ( .A(n13140), .ZN(n10015) );
  NOR2_X1 U11902 ( .A1(n20633), .A2(n9924), .ZN(n9922) );
  NAND2_X1 U11903 ( .A1(n14855), .A2(n13751), .ZN(n14922) );
  NAND2_X1 U11904 ( .A1(n15530), .A2(n14109), .ZN(n20783) );
  INV_X1 U11905 ( .A(n20783), .ZN(n15533) );
  XNOR2_X1 U11906 ( .A(n15436), .B(n15652), .ZN(n15659) );
  AND2_X1 U11907 ( .A1(n10021), .A2(n10022), .ZN(n15433) );
  OR2_X1 U11908 ( .A1(n13753), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9921) );
  AND2_X1 U11909 ( .A1(n15739), .A2(n20823), .ZN(n10067) );
  XNOR2_X1 U11910 ( .A(n15489), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15737) );
  INV_X1 U11911 ( .A(n20808), .ZN(n20823) );
  OR2_X1 U11912 ( .A1(n12970), .A2(n9744), .ZN(n15862) );
  INV_X1 U11913 ( .A(n10105), .ZN(n10104) );
  CLKBUF_X1 U11914 ( .A(n15283), .Z(n15284) );
  INV_X1 U11915 ( .A(n21375), .ZN(n21241) );
  NAND2_X1 U11916 ( .A1(n13273), .A2(n16357), .ZN(n13274) );
  NAND2_X1 U11917 ( .A1(n15950), .A2(n16357), .ZN(n15951) );
  INV_X1 U11918 ( .A(n15949), .ZN(n10289) );
  NOR2_X1 U11919 ( .A1(n16362), .A2(n15947), .ZN(n10288) );
  OR2_X1 U11920 ( .A1(n13823), .A2(n13255), .ZN(n16351) );
  AND2_X1 U11921 ( .A1(n13823), .A2(n14587), .ZN(n16342) );
  AND2_X1 U11922 ( .A1(n14442), .A2(n14436), .ZN(n10411) );
  NAND2_X1 U11923 ( .A1(n13736), .A2(n11521), .ZN(n13707) );
  OR2_X1 U11924 ( .A1(n11520), .A2(n11519), .ZN(n11521) );
  XNOR2_X1 U11925 ( .A(n15966), .B(n11492), .ZN(n15955) );
  INV_X1 U11926 ( .A(n19797), .ZN(n16459) );
  AND2_X1 U11927 ( .A1(n13985), .A2(n19837), .ZN(n16541) );
  AND2_X1 U11928 ( .A1(n13704), .A2(n14601), .ZN(n19795) );
  OR2_X1 U11929 ( .A1(n14215), .A2(n13703), .ZN(n13704) );
  AND2_X1 U11930 ( .A1(n19795), .A2(n13706), .ZN(n19797) );
  NAND2_X1 U11931 ( .A1(n10030), .A2(n9643), .ZN(n9982) );
  INV_X1 U11932 ( .A(n13295), .ZN(n10402) );
  OR2_X1 U11933 ( .A1(n9634), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10149) );
  INV_X1 U11934 ( .A(n10328), .ZN(n10010) );
  INV_X1 U11935 ( .A(n16594), .ZN(n10329) );
  NOR2_X1 U11936 ( .A1(n16637), .A2(n10139), .ZN(n10138) );
  NAND2_X1 U11937 ( .A1(n13307), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10139) );
  OAI21_X1 U11938 ( .B1(n10144), .B2(n16846), .A(n9690), .ZN(n10143) );
  INV_X1 U11939 ( .A(n16622), .ZN(n10145) );
  NAND2_X1 U11940 ( .A1(n9967), .A2(n16836), .ZN(n9966) );
  NAND2_X1 U11941 ( .A1(n9958), .A2(n9680), .ZN(n9967) );
  OR2_X1 U11942 ( .A1(n16632), .A2(n16609), .ZN(n9958) );
  OR2_X1 U11943 ( .A1(n16935), .A2(n16863), .ZN(n9799) );
  NAND2_X1 U11944 ( .A1(n16691), .A2(n16969), .ZN(n10258) );
  NOR2_X1 U11945 ( .A1(n16684), .A2(n16846), .ZN(n10257) );
  INV_X1 U11946 ( .A(n14815), .ZN(n16684) );
  NAND2_X1 U11947 ( .A1(n16839), .A2(n13874), .ZN(n16856) );
  XNOR2_X1 U11948 ( .A(n11048), .B(n10632), .ZN(n10633) );
  NAND2_X1 U11949 ( .A1(n20587), .A2(n20419), .ZN(n19838) );
  INV_X1 U11950 ( .A(n16856), .ZN(n16842) );
  INV_X1 U11951 ( .A(n16839), .ZN(n16858) );
  OAI211_X1 U11952 ( .C1(n10030), .C2(n9985), .A(n9984), .B(n9981), .ZN(n13308) );
  NAND2_X1 U11953 ( .A1(n10030), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9981) );
  XNOR2_X1 U11954 ( .A(n10119), .B(n10480), .ZN(n13731) );
  NAND2_X1 U11955 ( .A1(n13289), .A2(n9649), .ZN(n10119) );
  NAND2_X1 U11956 ( .A1(n11234), .A2(n10403), .ZN(n16571) );
  OR2_X1 U11957 ( .A1(n11233), .A2(n11232), .ZN(n11234) );
  NAND2_X1 U11958 ( .A1(n11503), .A2(n11504), .ZN(n10031) );
  NAND2_X1 U11959 ( .A1(n10326), .A2(n16582), .ZN(n9789) );
  AND2_X1 U11960 ( .A1(n9859), .A2(n9563), .ZN(n9855) );
  AOI21_X1 U11961 ( .B1(n16632), .B2(n16630), .A(n9956), .ZN(n16911) );
  NAND2_X1 U11962 ( .A1(n16631), .A2(n16627), .ZN(n9956) );
  NAND2_X1 U11963 ( .A1(n16921), .A2(n17121), .ZN(n10304) );
  INV_X1 U11964 ( .A(n16920), .ZN(n10303) );
  NOR2_X1 U11965 ( .A1(n16912), .A2(n17139), .ZN(n10306) );
  NAND2_X1 U11966 ( .A1(n10054), .A2(n16919), .ZN(n10276) );
  NAND2_X1 U11967 ( .A1(n10277), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16624) );
  NAND2_X1 U11968 ( .A1(n16637), .A2(n16928), .ZN(n9993) );
  INV_X1 U11969 ( .A(n16661), .ZN(n10447) );
  NOR2_X1 U11970 ( .A1(n14893), .A2(n16939), .ZN(n10446) );
  INV_X1 U11971 ( .A(n10425), .ZN(n10424) );
  INV_X1 U11972 ( .A(n10337), .ZN(n10336) );
  OAI21_X1 U11973 ( .B1(n16533), .B2(n17134), .A(n13154), .ZN(n10337) );
  OAI21_X1 U11974 ( .B1(n16700), .B2(n9628), .A(n13148), .ZN(n16967) );
  NAND2_X1 U11975 ( .A1(n16775), .A2(n17056), .ZN(n9787) );
  INV_X1 U11976 ( .A(n16754), .ZN(n9788) );
  NAND2_X1 U11977 ( .A1(n11505), .A2(n11238), .ZN(n17116) );
  INV_X1 U11978 ( .A(n17116), .ZN(n17127) );
  INV_X1 U11979 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20291) );
  INV_X1 U11980 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20582) );
  INV_X1 U11981 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20574) );
  NAND2_X1 U11982 ( .A1(n19756), .A2(n18538), .ZN(n19754) );
  AOI21_X1 U11983 ( .B1(n19587), .B2(n19588), .A(n18576), .ZN(n19756) );
  OAI21_X1 U11984 ( .B1(n17691), .B2(n19704), .A(n10001), .ZN(n10000) );
  NAND2_X1 U11985 ( .A1(n17997), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n10001) );
  NOR2_X1 U11986 ( .A1(n17785), .A2(n18000), .ZN(n17777) );
  AND2_X1 U11987 ( .A1(n18102), .A2(n17361), .ZN(n18096) );
  NAND2_X1 U11988 ( .A1(n18317), .A2(n9755), .ZN(n18263) );
  AND2_X1 U11989 ( .A1(n10222), .A2(n10219), .ZN(n18383) );
  AND2_X1 U11990 ( .A1(n10220), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(n10219) );
  AND2_X1 U11991 ( .A1(n10222), .A2(n10221), .ZN(n18389) );
  AND2_X1 U11992 ( .A1(n10221), .A2(P3_EBX_REG_0__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U11993 ( .A1(n18413), .A2(n18600), .ZN(n18408) );
  NOR2_X1 U11994 ( .A1(n18431), .A2(n19171), .ZN(n18427) );
  NOR2_X1 U11995 ( .A1(n18443), .A2(n10058), .ZN(n10057) );
  NAND2_X1 U11996 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_16__SCAN_IN), 
        .ZN(n10058) );
  AOI21_X1 U11997 ( .B1(n18824), .B2(n13330), .A(n9810), .ZN(n9809) );
  INV_X1 U11998 ( .A(n14748), .ZN(n9810) );
  INV_X1 U11999 ( .A(n9811), .ZN(n14879) );
  NAND2_X1 U12000 ( .A1(n18780), .A2(n11712), .ZN(n18681) );
  NAND2_X1 U12001 ( .A1(n10321), .A2(n11716), .ZN(n17333) );
  NOR2_X1 U12002 ( .A1(n10245), .A2(n19089), .ZN(n18924) );
  NOR2_X1 U12003 ( .A1(n17338), .A2(n10246), .ZN(n10245) );
  OAI21_X1 U12004 ( .B1(n18971), .B2(n10247), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10246) );
  NOR2_X1 U12005 ( .A1(n17337), .A2(n17339), .ZN(n10247) );
  AND2_X1 U12006 ( .A1(n17301), .A2(n17282), .ZN(n19099) );
  INV_X1 U12007 ( .A(n19119), .ZN(n19044) );
  INV_X1 U12008 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18536) );
  NAND2_X1 U12009 ( .A1(n14861), .A2(n9585), .ZN(n12779) );
  OR2_X1 U12010 ( .A1(n12274), .A2(n12273), .ZN(n12903) );
  NAND2_X1 U12011 ( .A1(n12085), .A2(n10115), .ZN(n12959) );
  NAND2_X1 U12012 ( .A1(n10095), .A2(n12091), .ZN(n9907) );
  NAND2_X1 U12013 ( .A1(n10775), .A2(n10131), .ZN(n9871) );
  NAND2_X1 U12014 ( .A1(n20046), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10133) );
  NAND2_X1 U12015 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10161) );
  INV_X1 U12016 ( .A(n10778), .ZN(n9866) );
  NAND2_X1 U12017 ( .A1(n20209), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10162) );
  OAI21_X1 U12018 ( .B1(n20140), .B2(n10774), .A(n10130), .ZN(n9873) );
  NAND2_X1 U12019 ( .A1(n20324), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10130) );
  NAND2_X1 U12020 ( .A1(n10647), .A2(n9614), .ZN(n10279) );
  NAND2_X1 U12021 ( .A1(n10647), .A2(n9613), .ZN(n10278) );
  INV_X1 U12022 ( .A(n20324), .ZN(n10710) );
  NAND2_X1 U12023 ( .A1(n20237), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10147) );
  NAND2_X1 U12024 ( .A1(n10797), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10261) );
  NAND2_X1 U12025 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  NAND2_X1 U12026 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10263) );
  NAND2_X1 U12027 ( .A1(n10651), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10264) );
  NAND2_X1 U12028 ( .A1(n10647), .A2(n10159), .ZN(n10160) );
  AND2_X1 U12029 ( .A1(n9574), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10159) );
  NAND2_X1 U12030 ( .A1(n13684), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10206) );
  NAND2_X1 U12031 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10207) );
  NAND2_X1 U12032 ( .A1(n10668), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10208) );
  NAND2_X1 U12033 ( .A1(n9587), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10201) );
  NAND2_X1 U12034 ( .A1(n9575), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10200) );
  NAND2_X1 U12035 ( .A1(n13577), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10202) );
  NAND2_X1 U12036 ( .A1(n10668), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10197) );
  NAND2_X1 U12037 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10196) );
  NAND2_X1 U12038 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10198) );
  NAND2_X1 U12039 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10212) );
  NAND2_X1 U12040 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10211) );
  NAND2_X1 U12041 ( .A1(n13577), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10213) );
  AND2_X1 U12042 ( .A1(n21294), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12795) );
  AOI21_X1 U12043 ( .B1(n12814), .B2(n12813), .A(n12812), .ZN(n12824) );
  NOR2_X1 U12044 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20835), .ZN(
        n12827) );
  OR2_X1 U12045 ( .A1(n9604), .A2(n10441), .ZN(n10440) );
  NAND2_X1 U12046 ( .A1(n20854), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10441) );
  OR2_X1 U12047 ( .A1(n9600), .A2(n10025), .ZN(n10023) );
  INV_X1 U12048 ( .A(n10021), .ZN(n9888) );
  INV_X1 U12049 ( .A(n12899), .ZN(n12320) );
  AOI22_X1 U12050 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12154) );
  OR2_X1 U12051 ( .A1(n12250), .A2(n12249), .ZN(n12904) );
  NAND2_X1 U12052 ( .A1(n10192), .A2(n20859), .ZN(n9769) );
  NAND2_X1 U12053 ( .A1(n10050), .A2(n9620), .ZN(n10592) );
  INV_X1 U12054 ( .A(n10597), .ZN(n10049) );
  NOR2_X1 U12055 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13507) );
  CLKBUF_X1 U12056 ( .A(n13678), .Z(n13658) );
  NAND2_X1 U12057 ( .A1(n10662), .A2(n10669), .ZN(n13475) );
  NAND2_X1 U12058 ( .A1(n11193), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10597) );
  INV_X1 U12059 ( .A(n10460), .ZN(n10137) );
  INV_X1 U12060 ( .A(n13286), .ZN(n10364) );
  AOI22_X1 U12061 ( .A1(n19978), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U12062 ( .A1(n10796), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10164) );
  OR2_X1 U12063 ( .A1(n10696), .A2(n10695), .ZN(n10900) );
  NAND2_X1 U12064 ( .A1(n9798), .A2(n10604), .ZN(n11249) );
  AOI22_X1 U12065 ( .A1(n13577), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9596), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10562) );
  INV_X1 U12066 ( .A(n11659), .ZN(n9940) );
  AOI21_X1 U12067 ( .B1(n11659), .B2(n9939), .A(n9938), .ZN(n9936) );
  INV_X1 U12068 ( .A(n14170), .ZN(n9938) );
  AND2_X1 U12069 ( .A1(n21538), .A2(n11857), .ZN(n11867) );
  AND2_X1 U12070 ( .A1(n11865), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U12071 ( .A1(n12820), .A2(n12953), .ZN(n12830) );
  OR2_X1 U12072 ( .A1(n12568), .A2(n12486), .ZN(n12534) );
  NAND2_X1 U12073 ( .A1(n12468), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12732) );
  NAND2_X1 U12074 ( .A1(n12367), .A2(n12366), .ZN(n12391) );
  AND2_X1 U12075 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12366) );
  INV_X1 U12076 ( .A(n12231), .ZN(n10385) );
  NOR2_X1 U12077 ( .A1(n14995), .A2(n14903), .ZN(n10121) );
  NAND2_X1 U12078 ( .A1(n9912), .A2(n9909), .ZN(n10073) );
  INV_X1 U12079 ( .A(n15477), .ZN(n9763) );
  OR2_X1 U12080 ( .A1(n15583), .A2(n12943), .ZN(n15560) );
  NAND2_X1 U12081 ( .A1(n14522), .A2(n14521), .ZN(n12893) );
  NAND2_X1 U12082 ( .A1(n9819), .A2(n12902), .ZN(n9818) );
  AOI21_X1 U12083 ( .B1(n12278), .B2(n9726), .A(n9919), .ZN(n9916) );
  NOR2_X1 U12084 ( .A1(n12869), .A2(n10084), .ZN(n9919) );
  NAND2_X1 U12085 ( .A1(n14229), .A2(n12883), .ZN(n12888) );
  NAND2_X1 U12086 ( .A1(n9947), .A2(n12901), .ZN(n14522) );
  AND2_X1 U12087 ( .A1(n12253), .A2(n9583), .ZN(n9947) );
  NAND2_X1 U12088 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  NAND2_X1 U12089 ( .A1(n14114), .A2(n20832), .ZN(n12974) );
  OAI21_X1 U12090 ( .B1(n14336), .B2(n12951), .A(n9735), .ZN(n12952) );
  NAND2_X1 U12091 ( .A1(n12196), .A2(n10235), .ZN(n10234) );
  INV_X1 U12092 ( .A(n12107), .ZN(n12091) );
  AOI22_X1 U12093 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U12094 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12747), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U12095 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U12096 ( .A1(n14019), .A2(n14018), .ZN(n14367) );
  OAI21_X1 U12097 ( .B1(n10880), .B2(n13271), .A(n10879), .ZN(n10903) );
  NAND2_X1 U12098 ( .A1(n13271), .A2(n11186), .ZN(n10879) );
  NOR2_X1 U12099 ( .A1(n13241), .A2(n15979), .ZN(n13240) );
  AND2_X1 U12100 ( .A1(n10966), .A2(n10999), .ZN(n10378) );
  INV_X1 U12101 ( .A(n16419), .ZN(n10405) );
  NAND2_X1 U12102 ( .A1(n10050), .A2(n9619), .ZN(n10607) );
  AND2_X1 U12103 ( .A1(n10049), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n9619) );
  CLKBUF_X1 U12104 ( .A(n13577), .Z(n13683) );
  NOR2_X1 U12105 ( .A1(n16388), .A2(n16391), .ZN(n16375) );
  CLKBUF_X1 U12106 ( .A(n13505), .Z(n13679) );
  AND2_X1 U12107 ( .A1(n14046), .A2(n13352), .ZN(n14186) );
  AND2_X1 U12108 ( .A1(n17491), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13352) );
  NAND2_X1 U12109 ( .A1(n10283), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13241) );
  AND2_X1 U12110 ( .A1(n11139), .A2(n11138), .ZN(n11143) );
  NOR2_X1 U12111 ( .A1(n13236), .A2(n16600), .ZN(n10283) );
  AND2_X1 U12112 ( .A1(n13225), .A2(n9746), .ZN(n13237) );
  NAND2_X1 U12113 ( .A1(n13225), .A2(n9629), .ZN(n13234) );
  NOR2_X1 U12114 ( .A1(n13211), .A2(n10290), .ZN(n13217) );
  NAND2_X1 U12115 ( .A1(n10292), .A2(n10291), .ZN(n10290) );
  INV_X1 U12116 ( .A(n10294), .ZN(n10292) );
  NOR2_X1 U12117 ( .A1(n10293), .A2(n13219), .ZN(n10291) );
  INV_X1 U12118 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U12119 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10294) );
  NAND2_X1 U12120 ( .A1(n9774), .A2(n9773), .ZN(n10605) );
  NAND2_X1 U12121 ( .A1(n10591), .A2(n10586), .ZN(n9773) );
  INV_X1 U12122 ( .A(n9796), .ZN(n9774) );
  AND2_X1 U12123 ( .A1(n9637), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10416) );
  INV_X1 U12124 ( .A(n16024), .ZN(n10351) );
  INV_X1 U12125 ( .A(n16630), .ZN(n9963) );
  OR2_X1 U12126 ( .A1(n16057), .A2(n11513), .ZN(n11036) );
  NAND2_X1 U12127 ( .A1(n9660), .A2(n9615), .ZN(n16608) );
  AND2_X1 U12128 ( .A1(n11478), .A2(n14825), .ZN(n14887) );
  NAND2_X1 U12129 ( .A1(n9978), .A2(n13159), .ZN(n9977) );
  INV_X1 U12130 ( .A(n14811), .ZN(n9978) );
  AND2_X1 U12131 ( .A1(n9640), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10158) );
  AND2_X1 U12132 ( .A1(n13163), .A2(n9752), .ZN(n10448) );
  NOR2_X1 U12133 ( .A1(n16699), .A2(n17029), .ZN(n10415) );
  AND2_X1 U12134 ( .A1(n11075), .A2(n11074), .ZN(n14406) );
  INV_X1 U12135 ( .A(n14401), .ZN(n10394) );
  INV_X1 U12136 ( .A(n10852), .ZN(n9828) );
  NAND2_X1 U12137 ( .A1(n16791), .A2(n11265), .ZN(n10154) );
  NAND2_X1 U12138 ( .A1(n16833), .A2(n10828), .ZN(n9843) );
  NAND2_X1 U12139 ( .A1(n10829), .A2(n11513), .ZN(n16791) );
  AOI21_X1 U12140 ( .B1(n9795), .B2(n10937), .A(n13293), .ZN(n9794) );
  OR2_X1 U12141 ( .A1(n10793), .A2(n10792), .ZN(n11318) );
  INV_X1 U12142 ( .A(n17098), .ZN(n11526) );
  NAND2_X1 U12143 ( .A1(n14186), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13353) );
  CLKBUF_X1 U12144 ( .A(n11495), .Z(n11496) );
  NAND2_X1 U12145 ( .A1(n10574), .A2(n9727), .ZN(n10169) );
  NAND2_X1 U12146 ( .A1(n10578), .A2(n19862), .ZN(n10167) );
  AND2_X1 U12147 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13508) );
  INV_X1 U12148 ( .A(n10156), .ZN(n10442) );
  NAND2_X1 U12149 ( .A1(n13313), .A2(n9730), .ZN(n14729) );
  OR2_X1 U12150 ( .A1(n9996), .A2(n18740), .ZN(n9995) );
  NAND2_X1 U12151 ( .A1(n9997), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9996) );
  INV_X1 U12152 ( .A(n18774), .ZN(n9997) );
  OAI22_X1 U12153 ( .A1(n17189), .A2(n9638), .B1(n11722), .B2(n10312), .ZN(
        n14717) );
  NAND2_X1 U12154 ( .A1(n10317), .A2(n17316), .ZN(n10312) );
  INV_X1 U12155 ( .A(n11941), .ZN(n11942) );
  AOI21_X1 U12156 ( .B1(n11940), .B2(n11939), .A(n19153), .ZN(n11941) );
  INV_X1 U12157 ( .A(n19011), .ZN(n10251) );
  OR2_X1 U12158 ( .A1(n11872), .A2(n11871), .ZN(n11885) );
  INV_X1 U12159 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14064) );
  AOI21_X1 U12160 ( .B1(n19588), .B2(n10463), .A(n14026), .ZN(n14501) );
  AOI21_X1 U12161 ( .B1(n19739), .B2(n19127), .A(n19612), .ZN(n19138) );
  INV_X1 U12162 ( .A(n20674), .ZN(n20694) );
  NAND2_X1 U12163 ( .A1(n14114), .A2(n15637), .ZN(n13082) );
  INV_X1 U12164 ( .A(n10121), .ZN(n14905) );
  NAND2_X1 U12165 ( .A1(n14114), .A2(n15689), .ZN(n13066) );
  NOR2_X1 U12166 ( .A1(n15085), .A2(n13055), .ZN(n15056) );
  AND2_X1 U12167 ( .A1(n14343), .A2(n12841), .ZN(n14010) );
  NAND2_X1 U12168 ( .A1(n9580), .A2(n10079), .ZN(n13141) );
  AND2_X1 U12169 ( .A1(n12036), .A2(n10080), .ZN(n10079) );
  INV_X1 U12170 ( .A(n20838), .ZN(n20836) );
  INV_X1 U12171 ( .A(n12765), .ZN(n12772) );
  INV_X1 U12172 ( .A(n12734), .ZN(n12735) );
  INV_X1 U12173 ( .A(n12621), .ZN(n12620) );
  INV_X1 U12174 ( .A(n12552), .ZN(n12487) );
  NOR2_X2 U12175 ( .A1(n12534), .A2(n15505), .ZN(n12549) );
  AND2_X1 U12176 ( .A1(n10388), .A2(n15112), .ZN(n10387) );
  OR2_X1 U12177 ( .A1(n12425), .A2(n12424), .ZN(n12483) );
  INV_X1 U12178 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12482) );
  AND2_X1 U12179 ( .A1(n15220), .A2(n10388), .ZN(n15110) );
  NAND2_X1 U12180 ( .A1(n12440), .A2(n12393), .ZN(n12425) );
  AND2_X1 U12181 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12393) );
  INV_X1 U12182 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12424) );
  CLKBUF_X1 U12183 ( .A(n15220), .Z(n15221) );
  INV_X1 U12184 ( .A(n12330), .ZN(n12331) );
  INV_X1 U12185 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12298) );
  NAND2_X1 U12186 ( .A1(n14296), .A2(n14424), .ZN(n14529) );
  AOI21_X1 U12187 ( .B1(n12305), .B2(n12464), .A(n12304), .ZN(n14530) );
  INV_X1 U12188 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12254) );
  XNOR2_X1 U12189 ( .A(n12888), .B(n13129), .ZN(n14256) );
  INV_X1 U12190 ( .A(n14259), .ZN(n12230) );
  XNOR2_X1 U12191 ( .A(n12881), .B(n14107), .ZN(n14230) );
  OAI21_X1 U12192 ( .B1(n9943), .B2(n15646), .A(n9942), .ZN(n9822) );
  NAND2_X1 U12193 ( .A1(n10121), .A2(n10120), .ZN(n14977) );
  INV_X1 U12194 ( .A(n14859), .ZN(n10120) );
  NAND2_X1 U12195 ( .A1(n13079), .A2(n10093), .ZN(n14978) );
  NAND2_X1 U12196 ( .A1(n14114), .A2(n15642), .ZN(n10093) );
  NAND2_X1 U12197 ( .A1(n10070), .A2(n10069), .ZN(n10021) );
  NOR2_X1 U12198 ( .A1(n10432), .A2(n10075), .ZN(n10069) );
  INV_X1 U12199 ( .A(n10071), .ZN(n10022) );
  NAND2_X1 U12200 ( .A1(n10026), .A2(n12946), .ZN(n15432) );
  AND2_X1 U12201 ( .A1(n10125), .A2(n10123), .ZN(n10122) );
  INV_X1 U12202 ( .A(n13772), .ZN(n10123) );
  NAND2_X1 U12203 ( .A1(n10124), .A2(n10125), .ZN(n15045) );
  OAI21_X1 U12204 ( .B1(n10430), .B2(n9750), .A(n15595), .ZN(n10433) );
  NAND2_X1 U12205 ( .A1(n15496), .A2(n10066), .ZN(n15488) );
  AND2_X1 U12206 ( .A1(n15583), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10066) );
  NAND2_X1 U12207 ( .A1(n13043), .A2(n10091), .ZN(n15084) );
  NAND2_X1 U12208 ( .A1(n14114), .A2(n10092), .ZN(n10091) );
  AND2_X1 U12209 ( .A1(n13042), .A2(n13041), .ZN(n15104) );
  NAND2_X1 U12210 ( .A1(n14114), .A2(n10088), .ZN(n13032) );
  NAND2_X1 U12211 ( .A1(n15516), .A2(n9812), .ZN(n15524) );
  NAND2_X1 U12212 ( .A1(n9581), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9812) );
  AND2_X1 U12213 ( .A1(n13037), .A2(n13036), .ZN(n15137) );
  AND2_X1 U12214 ( .A1(n15549), .A2(n12942), .ZN(n15539) );
  NAND2_X1 U12215 ( .A1(n14114), .A2(n15797), .ZN(n13024) );
  NOR2_X1 U12216 ( .A1(n15565), .A2(n12938), .ZN(n15551) );
  NAND2_X1 U12217 ( .A1(n15593), .A2(n15514), .ZN(n15552) );
  AND2_X1 U12218 ( .A1(n13030), .A2(n13029), .ZN(n15168) );
  AND2_X1 U12219 ( .A1(n9611), .A2(n9699), .ZN(n10127) );
  NAND2_X1 U12220 ( .A1(n13013), .A2(n10089), .ZN(n15205) );
  NAND2_X1 U12221 ( .A1(n14114), .A2(n10090), .ZN(n10089) );
  NAND2_X1 U12222 ( .A1(n15224), .A2(n9611), .ZN(n15207) );
  NAND2_X1 U12223 ( .A1(n15224), .A2(n15223), .ZN(n15226) );
  NAND2_X1 U12224 ( .A1(n9821), .A2(n12935), .ZN(n10231) );
  CLKBUF_X1 U12225 ( .A(n17503), .Z(n17504) );
  NAND2_X1 U12226 ( .A1(n14114), .A2(n13129), .ZN(n12977) );
  NAND2_X1 U12227 ( .A1(n13102), .A2(n10085), .ZN(n13103) );
  INV_X1 U12228 ( .A(n9761), .ZN(n12468) );
  NAND2_X1 U12229 ( .A1(n14356), .A2(n9745), .ZN(n14358) );
  INV_X1 U12230 ( .A(n14367), .ZN(n15906) );
  AND2_X1 U12231 ( .A1(n21207), .A2(n21329), .ZN(n21175) );
  OAI21_X1 U12232 ( .B1(n21173), .B2(n21230), .A(n21235), .ZN(n21178) );
  AND2_X1 U12233 ( .A1(n9599), .A2(n20840), .ZN(n21203) );
  OR2_X1 U12234 ( .A1(n9599), .A2(n20840), .ZN(n21234) );
  INV_X1 U12235 ( .A(n21203), .ZN(n21086) );
  NOR2_X1 U12236 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21384) );
  AOI21_X1 U12237 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21294), .A(n21000), 
        .ZN(n21380) );
  AND2_X1 U12238 ( .A1(n15927), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13767) );
  INV_X1 U12239 ( .A(n15945), .ZN(n15927) );
  INV_X1 U12240 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15884) );
  OR2_X1 U12241 ( .A1(n10578), .A2(n11279), .ZN(n10583) );
  MUX2_X1 U12242 ( .A(n10873), .B(n10872), .S(n13271), .Z(n10899) );
  AND2_X1 U12243 ( .A1(n20598), .A2(n10891), .ZN(n14574) );
  NOR2_X1 U12244 ( .A1(n10580), .A2(n19862), .ZN(n10155) );
  AND2_X1 U12245 ( .A1(n15992), .A2(n15993), .ZN(n15983) );
  NAND2_X1 U12246 ( .A1(n16249), .A2(n13231), .ZN(n16054) );
  NOR2_X1 U12247 ( .A1(n10902), .A2(n10969), .ZN(n10970) );
  AND2_X1 U12248 ( .A1(n13225), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13229) );
  NOR2_X1 U12249 ( .A1(n10375), .A2(n10973), .ZN(n10374) );
  INV_X1 U12250 ( .A(n10470), .ZN(n10375) );
  INV_X1 U12251 ( .A(n11005), .ZN(n10998) );
  NOR2_X1 U12252 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20608) );
  AND2_X1 U12253 ( .A1(n10007), .A2(n10954), .ZN(n16251) );
  AND2_X1 U12254 ( .A1(n14574), .A2(n14601), .ZN(n13253) );
  NOR2_X1 U12255 ( .A1(n16423), .A2(n9740), .ZN(n9778) );
  AND2_X1 U12256 ( .A1(n11111), .A2(n11110), .ZN(n16090) );
  NOR2_X1 U12257 ( .A1(n10342), .A2(n15968), .ZN(n10341) );
  INV_X1 U12258 ( .A(n15972), .ZN(n10342) );
  NOR2_X1 U12259 ( .A1(n16376), .A2(n16375), .ZN(n16385) );
  NAND2_X1 U12260 ( .A1(n13609), .A2(n13593), .ZN(n16388) );
  AND2_X1 U12261 ( .A1(n11485), .A2(n11484), .ZN(n16013) );
  XNOR2_X1 U12262 ( .A(n9778), .B(n16408), .ZN(n16415) );
  NAND2_X1 U12263 ( .A1(n16415), .A2(n16414), .ZN(n16413) );
  AND2_X1 U12264 ( .A1(n11468), .A2(n11467), .ZN(n13146) );
  NAND2_X1 U12265 ( .A1(n10396), .A2(n14610), .ZN(n9777) );
  AND2_X1 U12266 ( .A1(n10398), .A2(n10397), .ZN(n10396) );
  INV_X1 U12267 ( .A(n14681), .ZN(n10397) );
  INV_X1 U12268 ( .A(n13836), .ZN(n13897) );
  AND2_X2 U12269 ( .A1(n13718), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19839)
         );
  INV_X1 U12270 ( .A(n11232), .ZN(n10401) );
  INV_X1 U12271 ( .A(n16627), .ZN(n9960) );
  OR2_X1 U12272 ( .A1(n16609), .A2(n16630), .ZN(n9957) );
  AND2_X1 U12273 ( .A1(n11127), .A2(n11126), .ZN(n16036) );
  AND2_X1 U12274 ( .A1(n9665), .A2(n11123), .ZN(n10408) );
  AND2_X1 U12275 ( .A1(n11122), .A2(n14843), .ZN(n11123) );
  NOR2_X1 U12276 ( .A1(n13208), .A2(n16747), .ZN(n13210) );
  INV_X1 U12277 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16747) );
  INV_X1 U12278 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13206) );
  OR2_X1 U12279 ( .A1(n13203), .A2(n13206), .ZN(n13208) );
  NOR2_X1 U12280 ( .A1(n13199), .A2(n16811), .ZN(n13201) );
  INV_X1 U12281 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16811) );
  NAND2_X1 U12282 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10296) );
  NAND2_X1 U12283 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13196) );
  NOR2_X1 U12284 ( .A1(n13196), .A2(n14637), .ZN(n13195) );
  INV_X1 U12285 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14637) );
  NAND2_X1 U12286 ( .A1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13739), .ZN(
        n9984) );
  NAND2_X1 U12287 ( .A1(n13190), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9985) );
  AND2_X1 U12288 ( .A1(n13283), .A2(n13282), .ZN(n13288) );
  AOI21_X1 U12289 ( .B1(n13273), .B2(n13293), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13281) );
  INV_X1 U12290 ( .A(n13273), .ZN(n11514) );
  NOR3_X1 U12291 ( .A1(n11173), .A2(n11513), .A3(n11504), .ZN(n13278) );
  AOI21_X1 U12292 ( .B1(n15950), .B2(n13293), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13280) );
  OR2_X1 U12293 ( .A1(n16887), .A2(n11502), .ZN(n16865) );
  AND2_X1 U12294 ( .A1(n15976), .A2(n15958), .ZN(n11233) );
  OAI21_X1 U12295 ( .B1(n9624), .B2(n9861), .A(n9860), .ZN(n9859) );
  NOR2_X1 U12296 ( .A1(n16597), .A2(n16595), .ZN(n9861) );
  NAND2_X1 U12297 ( .A1(n9624), .A2(n9864), .ZN(n9860) );
  OR2_X1 U12298 ( .A1(n16899), .A2(n11268), .ZN(n16887) );
  AND2_X1 U12299 ( .A1(n11135), .A2(n11134), .ZN(n16002) );
  NAND2_X1 U12300 ( .A1(n16103), .A2(n9718), .ZN(n16022) );
  OAI21_X1 U12301 ( .B1(n10429), .B2(n16663), .A(n10426), .ZN(n10425) );
  AOI21_X1 U12302 ( .B1(n14835), .B2(n10428), .A(n10427), .ZN(n10426) );
  INV_X1 U12303 ( .A(n16651), .ZN(n10428) );
  INV_X1 U12304 ( .A(n14837), .ZN(n10427) );
  INV_X1 U12305 ( .A(n14835), .ZN(n10429) );
  AND2_X1 U12306 ( .A1(n13151), .A2(n9665), .ZN(n16088) );
  AND2_X1 U12307 ( .A1(n11107), .A2(n11106), .ZN(n14689) );
  NAND2_X1 U12308 ( .A1(n13151), .A2(n9651), .ZN(n16089) );
  AND2_X1 U12309 ( .A1(n10421), .A2(n9682), .ZN(n10417) );
  AND2_X1 U12310 ( .A1(n16703), .A2(n16687), .ZN(n10421) );
  NAND2_X1 U12311 ( .A1(n11415), .A2(n10347), .ZN(n10345) );
  AND3_X1 U12312 ( .A1(n11414), .A2(n11413), .A3(n11412), .ZN(n14252) );
  NAND2_X1 U12313 ( .A1(n16754), .A2(n10415), .ZN(n16738) );
  CLKBUF_X1 U12314 ( .A(n14163), .Z(n14164) );
  AND2_X1 U12315 ( .A1(n11345), .A2(n14001), .ZN(n10340) );
  INV_X1 U12316 ( .A(n14041), .ZN(n11345) );
  INV_X1 U12317 ( .A(n14417), .ZN(n11064) );
  NOR2_X1 U12318 ( .A1(n17130), .A2(n11256), .ZN(n17078) );
  NAND2_X1 U12319 ( .A1(n14002), .A2(n14001), .ZN(n14000) );
  NAND2_X1 U12320 ( .A1(n16832), .A2(n10937), .ZN(n10270) );
  OR2_X1 U12321 ( .A1(n10933), .A2(n10934), .ZN(n9845) );
  NAND2_X1 U12322 ( .A1(n10913), .A2(n9847), .ZN(n9846) );
  OR2_X1 U12323 ( .A1(n14646), .A2(n14634), .ZN(n17130) );
  AND3_X1 U12324 ( .A1(n11315), .A2(n11314), .A3(n11313), .ZN(n16298) );
  NAND2_X1 U12325 ( .A1(n10913), .A2(n16313), .ZN(n16847) );
  AND2_X1 U12326 ( .A1(n11310), .A2(n11309), .ZN(n14643) );
  AND3_X1 U12327 ( .A1(n11261), .A2(n11260), .A3(n14785), .ZN(n17095) );
  CLKBUF_X1 U12328 ( .A(n11493), .Z(n11494) );
  XNOR2_X1 U12329 ( .A(n10642), .B(n10641), .ZN(n13359) );
  XNOR2_X1 U12330 ( .A(n10640), .B(n10639), .ZN(n10641) );
  NAND2_X1 U12331 ( .A1(n10643), .A2(n10638), .ZN(n10642) );
  INV_X1 U12332 ( .A(n11258), .ZN(n14786) );
  INV_X1 U12333 ( .A(n13164), .ZN(n14791) );
  AOI21_X1 U12334 ( .B1(n9574), .B2(n13360), .A(n13357), .ZN(n14004) );
  INV_X1 U12335 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U12336 ( .A1(n13190), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13191) );
  AND2_X2 U12337 ( .A1(n9825), .A2(n10651), .ZN(n19851) );
  INV_X1 U12338 ( .A(n10796), .ZN(n19947) );
  NAND2_X1 U12339 ( .A1(n10553), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10554) );
  AND2_X1 U12340 ( .A1(n20419), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19894) );
  NOR2_X2 U12341 ( .A1(n19837), .A2(n19838), .ZN(n19893) );
  AND3_X1 U12342 ( .A1(n14223), .A2(n14222), .A3(n14221), .ZN(n14582) );
  NOR2_X1 U12343 ( .A1(n18578), .A2(n19140), .ZN(n14710) );
  INV_X1 U12344 ( .A(n14023), .ZN(n9901) );
  NAND2_X1 U12345 ( .A1(n9994), .A2(n13324), .ZN(n17763) );
  NOR2_X1 U12346 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17921), .ZN(n17910) );
  NAND2_X1 U12347 ( .A1(n17934), .A2(n17923), .ZN(n17921) );
  NOR2_X1 U12348 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17950), .ZN(n17934) );
  NAND2_X1 U12349 ( .A1(n17962), .A2(n18371), .ZN(n17950) );
  NOR2_X1 U12350 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17978), .ZN(n17962) );
  NAND2_X1 U12351 ( .A1(n10226), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n10225) );
  INV_X1 U12352 ( .A(n18048), .ZN(n10226) );
  INV_X1 U12353 ( .A(n10229), .ZN(n10228) );
  OR2_X1 U12354 ( .A1(n10230), .A2(n17979), .ZN(n10229) );
  NAND2_X1 U12355 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .ZN(n10230) );
  NOR2_X1 U12356 ( .A1(n18596), .A2(n10061), .ZN(n10060) );
  OR2_X1 U12357 ( .A1(n11655), .A2(n11654), .ZN(n11896) );
  NOR2_X1 U12358 ( .A1(n11594), .A2(n10320), .ZN(n10319) );
  INV_X1 U12359 ( .A(n11586), .ZN(n10318) );
  NOR2_X1 U12360 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11563) );
  NOR2_X1 U12361 ( .A1(n19162), .A2(n19166), .ZN(n14508) );
  OAI21_X1 U12362 ( .B1(n14023), .B2(n19614), .A(n19735), .ZN(n18537) );
  NOR2_X1 U12363 ( .A1(n10217), .A2(n18576), .ZN(n18577) );
  NOR2_X1 U12364 ( .A1(n17212), .A2(n18774), .ZN(n18761) );
  INV_X1 U12365 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18803) );
  NAND2_X1 U12366 ( .A1(n14717), .A2(n10315), .ZN(n14720) );
  NOR2_X1 U12367 ( .A1(n10316), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10315) );
  NOR2_X1 U12368 ( .A1(n11944), .A2(n11950), .ZN(n13332) );
  NOR2_X1 U12369 ( .A1(n18652), .A2(n18712), .ZN(n18651) );
  INV_X1 U12370 ( .A(n17332), .ZN(n18653) );
  NAND2_X1 U12371 ( .A1(n10321), .A2(n11717), .ZN(n18710) );
  NAND2_X1 U12372 ( .A1(n19010), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18985) );
  OR2_X1 U12373 ( .A1(n10324), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10323) );
  OR2_X1 U12374 ( .A1(n18809), .A2(n9756), .ZN(n18782) );
  OR2_X1 U12375 ( .A1(n14385), .A2(n10316), .ZN(n18835) );
  OR2_X1 U12376 ( .A1(n18795), .A2(n18712), .ZN(n18833) );
  NOR2_X1 U12377 ( .A1(n14387), .A2(n21579), .ZN(n14386) );
  NOR2_X1 U12378 ( .A1(n14169), .A2(n14390), .ZN(n14168) );
  XNOR2_X1 U12379 ( .A(n11615), .B(n11613), .ZN(n14119) );
  INV_X1 U12380 ( .A(n11899), .ZN(n10237) );
  XNOR2_X1 U12381 ( .A(n14666), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14145) );
  INV_X1 U12382 ( .A(n17350), .ZN(n17348) );
  NAND2_X1 U12383 ( .A1(n17348), .A2(n13332), .ZN(n19588) );
  INV_X1 U12384 ( .A(n11731), .ZN(n10056) );
  INV_X1 U12385 ( .A(n18538), .ZN(n19140) );
  INV_X1 U12386 ( .A(n19384), .ZN(n19428) );
  AOI21_X1 U12387 ( .B1(n19585), .B2(n19592), .A(n14276), .ZN(n19582) );
  NAND2_X1 U12388 ( .A1(n13942), .A2(n10082), .ZN(n13943) );
  INV_X1 U12389 ( .A(n20681), .ZN(n15228) );
  INV_X1 U12390 ( .A(n13790), .ZN(n13771) );
  AND2_X1 U12391 ( .A1(n15270), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20674) );
  NAND2_X1 U12392 ( .A1(n13796), .A2(n13794), .ZN(n15287) );
  INV_X1 U12393 ( .A(n15228), .ZN(n20691) );
  AND2_X1 U12394 ( .A1(n13796), .A2(n13775), .ZN(n20693) );
  NAND2_X1 U12395 ( .A1(n15287), .A2(n15270), .ZN(n20673) );
  INV_X1 U12396 ( .A(n15328), .ZN(n20707) );
  AND2_X1 U12397 ( .A1(n14307), .A2(n14306), .ZN(n20721) );
  INV_X1 U12398 ( .A(n20721), .ZN(n20741) );
  INV_X1 U12399 ( .A(n15343), .ZN(n15420) );
  NOR2_X1 U12400 ( .A1(n15072), .A2(n9645), .ZN(n15503) );
  INV_X1 U12401 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15505) );
  OR2_X1 U12402 ( .A1(n14679), .A2(n14678), .ZN(n15325) );
  INV_X1 U12403 ( .A(n15530), .ZN(n20772) );
  AOI22_X1 U12404 ( .A1(n14934), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n10095), .ZN(n14935) );
  OAI22_X1 U12405 ( .A1(n13173), .A2(n9731), .B1(n13172), .B2(n12947), .ZN(
        n12948) );
  NAND2_X1 U12406 ( .A1(n10037), .A2(n10036), .ZN(n15650) );
  NAND2_X1 U12407 ( .A1(n10041), .A2(n10042), .ZN(n10036) );
  NAND2_X1 U12408 ( .A1(n10043), .A2(n10039), .ZN(n10038) );
  NAND2_X1 U12409 ( .A1(n15450), .A2(n10076), .ZN(n15442) );
  INV_X1 U12410 ( .A(n15496), .ZN(n15467) );
  OAI21_X1 U12411 ( .B1(n15525), .B2(n9814), .A(n9813), .ZN(n15517) );
  INV_X1 U12412 ( .A(n15516), .ZN(n9814) );
  NAND2_X1 U12413 ( .A1(n15525), .A2(n15515), .ZN(n9813) );
  AND2_X1 U12414 ( .A1(n17545), .A2(n15843), .ZN(n17535) );
  INV_X1 U12415 ( .A(n20771), .ZN(n20804) );
  NAND2_X1 U12416 ( .A1(n13115), .A2(n13090), .ZN(n20808) );
  INV_X1 U12417 ( .A(n15862), .ZN(n20828) );
  NAND2_X1 U12418 ( .A1(n10435), .A2(n12879), .ZN(n14108) );
  NAND2_X1 U12419 ( .A1(n12220), .A2(n9650), .ZN(n10435) );
  INV_X1 U12420 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21294) );
  INV_X1 U12421 ( .A(n21384), .ZN(n21382) );
  INV_X1 U12422 ( .A(n21382), .ZN(n21210) );
  CLKBUF_X1 U12423 ( .A(n14350), .Z(n21119) );
  INV_X1 U12424 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20835) );
  NOR2_X1 U12425 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14926) );
  NAND2_X1 U12426 ( .A1(n9762), .A2(n20995), .ZN(n14020) );
  INV_X1 U12427 ( .A(n12232), .ZN(n9762) );
  OAI211_X1 U12428 ( .C1(n20851), .C2(n20848), .A(n21182), .B(n20846), .ZN(
        n20890) );
  INV_X1 U12429 ( .A(n20913), .ZN(n20916) );
  INV_X1 U12430 ( .A(n21047), .ZN(n21038) );
  OAI211_X1 U12431 ( .C1(n21054), .C2(n21248), .A(n21336), .B(n21053), .ZN(
        n21082) );
  OAI211_X1 U12432 ( .C1(n10472), .C2(n21248), .A(n21182), .B(n21127), .ZN(
        n21144) );
  INV_X1 U12433 ( .A(n21107), .ZN(n21143) );
  INV_X1 U12434 ( .A(n21395), .ZN(n21259) );
  INV_X1 U12435 ( .A(n21401), .ZN(n21264) );
  INV_X1 U12436 ( .A(n21407), .ZN(n21269) );
  INV_X1 U12437 ( .A(n21415), .ZN(n21274) );
  INV_X1 U12438 ( .A(n21421), .ZN(n21279) );
  INV_X1 U12439 ( .A(n21427), .ZN(n21285) );
  OAI211_X1 U12440 ( .C1(n21249), .C2(n21248), .A(n21336), .B(n21247), .ZN(
        n21288) );
  OAI211_X1 U12441 ( .C1(n21360), .C2(n21337), .A(n21336), .B(n21335), .ZN(
        n21364) );
  INV_X1 U12442 ( .A(n20884), .ZN(n10087) );
  AND2_X1 U12443 ( .A1(n20854), .A2(n20884), .ZN(n21389) );
  AND2_X1 U12444 ( .A1(n20856), .A2(n20865), .ZN(n21390) );
  AND2_X1 U12445 ( .A1(n20859), .A2(n20884), .ZN(n21395) );
  INV_X1 U12446 ( .A(n21263), .ZN(n21396) );
  AND2_X1 U12447 ( .A1(n20866), .A2(n20865), .ZN(n21402) );
  INV_X1 U12448 ( .A(n21436), .ZN(n21410) );
  AND2_X1 U12449 ( .A1(n20869), .A2(n20884), .ZN(n21407) );
  INV_X1 U12450 ( .A(n21273), .ZN(n21408) );
  AND2_X1 U12451 ( .A1(n12084), .A2(n20884), .ZN(n21415) );
  AND2_X1 U12452 ( .A1(n20878), .A2(n20884), .ZN(n21421) );
  INV_X1 U12453 ( .A(n21283), .ZN(n21422) );
  INV_X1 U12454 ( .A(n21413), .ZN(n21432) );
  AND2_X1 U12455 ( .A1(n20885), .A2(n20884), .ZN(n21427) );
  INV_X1 U12456 ( .A(n21291), .ZN(n21429) );
  INV_X1 U12457 ( .A(n13767), .ZN(n15940) );
  INV_X1 U12458 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21248) );
  NAND2_X1 U12459 ( .A1(n13831), .A2(n16368), .ZN(n13823) );
  AND2_X1 U12460 ( .A1(n13291), .A2(n11044), .ZN(n15998) );
  NAND2_X1 U12461 ( .A1(n10367), .A2(n10473), .ZN(n16029) );
  NAND2_X1 U12462 ( .A1(n16351), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16340) );
  INV_X1 U12463 ( .A(n16358), .ZN(n16339) );
  INV_X1 U12464 ( .A(n16351), .ZN(n16288) );
  NAND2_X1 U12465 ( .A1(n10963), .A2(n10962), .ZN(n10982) );
  AND2_X1 U12466 ( .A1(n10961), .A2(n10949), .ZN(n16245) );
  INV_X1 U12467 ( .A(n16350), .ZN(n16337) );
  NAND2_X1 U12468 ( .A1(n13250), .A2(n13249), .ZN(n16345) );
  INV_X1 U12469 ( .A(n16304), .ZN(n16365) );
  INV_X1 U12470 ( .A(n9778), .ZN(n16406) );
  OR2_X1 U12471 ( .A1(n11461), .A2(n11460), .ZN(n14659) );
  NOR2_X1 U12472 ( .A1(n14441), .A2(n13385), .ZN(n14660) );
  OR2_X1 U12473 ( .A1(n11395), .A2(n11394), .ZN(n14329) );
  OAI21_X1 U12474 ( .B1(n14198), .B2(n9783), .A(n13384), .ZN(n9781) );
  OR2_X1 U12475 ( .A1(n11359), .A2(n11358), .ZN(n14266) );
  OR2_X1 U12476 ( .A1(n11341), .A2(n11340), .ZN(n14399) );
  NOR2_X1 U12477 ( .A1(n14237), .A2(n14236), .ZN(n14414) );
  INV_X1 U12478 ( .A(n16433), .ZN(n16435) );
  NAND2_X1 U12479 ( .A1(n10129), .A2(n9905), .ZN(n9904) );
  INV_X1 U12480 ( .A(n10189), .ZN(n10129) );
  NAND2_X1 U12481 ( .A1(n14044), .A2(n14047), .ZN(n21692) );
  NAND2_X1 U12482 ( .A1(n16430), .A2(n19895), .ZN(n16433) );
  INV_X1 U12483 ( .A(n21692), .ZN(n19840) );
  INV_X1 U12484 ( .A(n19795), .ZN(n19796) );
  OAI21_X1 U12485 ( .B1(n13929), .B2(n20618), .A(n13928), .ZN(n19826) );
  OR2_X1 U12486 ( .A1(n14220), .A2(n13927), .ZN(n13928) );
  INV_X1 U12487 ( .A(n13877), .ZN(n13918) );
  OR2_X1 U12488 ( .A1(n13831), .A2(n17491), .ZN(n13929) );
  NAND2_X1 U12489 ( .A1(n9985), .A2(n9984), .ZN(n9983) );
  NAND2_X1 U12490 ( .A1(n9857), .A2(n10857), .ZN(n11535) );
  INV_X1 U12491 ( .A(n14848), .ZN(n9897) );
  NAND2_X1 U12492 ( .A1(n10101), .A2(n9674), .ZN(n10100) );
  NAND2_X1 U12493 ( .A1(n14815), .A2(n16674), .ZN(n10101) );
  NAND2_X1 U12494 ( .A1(n16700), .A2(n16974), .ZN(n10216) );
  NAND2_X1 U12495 ( .A1(n10407), .A2(n11048), .ZN(n14191) );
  NAND2_X1 U12496 ( .A1(n10326), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10153) );
  NAND2_X1 U12497 ( .A1(n10326), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10325) );
  NAND2_X1 U12498 ( .A1(n10140), .A2(n10144), .ZN(n16907) );
  NAND2_X1 U12499 ( .A1(n10277), .A2(n9652), .ZN(n10140) );
  NAND2_X1 U12500 ( .A1(n16648), .A2(n16651), .ZN(n14836) );
  INV_X1 U12501 ( .A(n10157), .ZN(n16673) );
  AND2_X1 U12502 ( .A1(n16674), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10339) );
  NOR2_X1 U12503 ( .A1(n10176), .A2(n16966), .ZN(n10175) );
  NOR2_X1 U12504 ( .A1(n13148), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10176) );
  NAND2_X1 U12505 ( .A1(n16705), .A2(n16702), .ZN(n10422) );
  AND2_X1 U12506 ( .A1(n9758), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10414) );
  OAI21_X1 U12507 ( .B1(n16728), .B2(n16725), .A(n16726), .ZN(n9903) );
  NAND2_X1 U12508 ( .A1(n16606), .A2(n16772), .ZN(n16759) );
  INV_X1 U12509 ( .A(n10648), .ZN(n10052) );
  AND2_X1 U12510 ( .A1(n20606), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20587) );
  NAND2_X1 U12511 ( .A1(n14007), .A2(n14006), .ZN(n20585) );
  OR2_X1 U12512 ( .A1(n14005), .A2(n14004), .ZN(n14007) );
  INV_X1 U12513 ( .A(n14099), .ZN(n14100) );
  INV_X1 U12514 ( .A(n14198), .ZN(n14199) );
  INV_X1 U12515 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17496) );
  OR2_X1 U12516 ( .A1(n19908), .A2(n19906), .ZN(n19935) );
  OAI21_X1 U12517 ( .B1(n19943), .B2(n20326), .A(n19944), .ZN(n19965) );
  AND2_X1 U12518 ( .A1(n19947), .A2(n19946), .ZN(n19943) );
  OAI211_X1 U12519 ( .C1(n19977), .C2(n19975), .A(n19974), .B(n20419), .ZN(
        n20006) );
  INV_X1 U12520 ( .A(n20020), .ZN(n20038) );
  OAI21_X1 U12521 ( .B1(n20019), .B2(n20570), .A(n20013), .ZN(n20036) );
  OAI211_X1 U12522 ( .C1(n20049), .C2(n20044), .A(n20419), .B(n20043), .ZN(
        n20073) );
  OAI21_X1 U12523 ( .B1(n20079), .B2(n20211), .A(n20078), .ZN(n20103) );
  OAI211_X1 U12524 ( .C1(n20114), .C2(n20113), .A(n20419), .B(n20112), .ZN(
        n20132) );
  INV_X1 U12525 ( .A(n10806), .ZN(n20111) );
  OAI21_X1 U12526 ( .B1(n20109), .B2(n20570), .A(n20108), .ZN(n20130) );
  NAND2_X1 U12527 ( .A1(n9785), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20108) );
  OR2_X1 U12528 ( .A1(n10806), .A2(n20145), .ZN(n9785) );
  OAI21_X1 U12529 ( .B1(n20185), .B2(n20184), .A(n20183), .ZN(n20204) );
  OAI21_X1 U12530 ( .B1(n20238), .B2(n20211), .A(n20210), .ZN(n20230) );
  OAI211_X1 U12531 ( .C1(n20249), .C2(n20607), .A(n20248), .B(n20419), .ZN(
        n20287) );
  INV_X1 U12532 ( .A(n20295), .ZN(n20319) );
  OAI21_X1 U12533 ( .B1(n20294), .B2(n20326), .A(n20293), .ZN(n20318) );
  AOI21_X1 U12534 ( .B1(n20326), .B2(n20325), .A(n20327), .ZN(n20355) );
  INV_X1 U12535 ( .A(n20243), .ZN(n20412) );
  AND2_X1 U12536 ( .A1(n17491), .A2(n19894), .ZN(n20425) );
  AND2_X1 U12537 ( .A1(n19859), .A2(n20419), .ZN(n20426) );
  AND2_X1 U12538 ( .A1(n19864), .A2(n20419), .ZN(n20432) );
  INV_X1 U12539 ( .A(n20268), .ZN(n20444) );
  INV_X1 U12540 ( .A(n20472), .ZN(n20452) );
  AND2_X1 U12541 ( .A1(n19881), .A2(n20419), .ZN(n20450) );
  OAI21_X1 U12542 ( .B1(n20410), .B2(n20570), .A(n20409), .ZN(n20466) );
  AND2_X1 U12543 ( .A1(n19898), .A2(n20419), .ZN(n20465) );
  AND3_X1 U12544 ( .A1(n17141), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n14601) );
  OR3_X1 U12545 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20485), .A3(n20487), .ZN(
        n20618) );
  INV_X1 U12546 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n21590) );
  NAND2_X1 U12547 ( .A1(n19743), .A2(n19589), .ZN(n18576) );
  INV_X1 U12548 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19740) );
  XNOR2_X1 U12549 ( .A(n17674), .B(n17673), .ZN(n17678) );
  NOR2_X1 U12550 ( .A1(n19699), .A2(n17727), .ZN(n17703) );
  NAND2_X1 U12551 ( .A1(n17762), .A2(n18106), .ZN(n17759) );
  INV_X1 U12552 ( .A(n18731), .ZN(n10004) );
  INV_X1 U12553 ( .A(n10005), .ZN(n17786) );
  NOR2_X1 U12554 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17873), .ZN(n17861) );
  INV_X1 U12555 ( .A(n18034), .ZN(n18004) );
  AND2_X1 U12556 ( .A1(n19615), .A2(n13337), .ZN(n17997) );
  AND4_X1 U12557 ( .A1(n19055), .A2(n19751), .A3(n19621), .A4(n19631), .ZN(
        n17983) );
  INV_X1 U12558 ( .A(n18011), .ZN(n18038) );
  INV_X1 U12559 ( .A(n17997), .ZN(n18039) );
  AND2_X1 U12560 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18105), .ZN(n18101) );
  NOR3_X1 U12561 ( .A1(n18149), .A2(n10225), .A3(n10223), .ZN(n18105) );
  NAND2_X1 U12562 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .ZN(n10223) );
  NOR2_X1 U12563 ( .A1(n18201), .A2(n18204), .ZN(n18184) );
  NAND2_X1 U12564 ( .A1(n18205), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n18201) );
  NAND2_X1 U12565 ( .A1(n18317), .A2(n9635), .ZN(n18280) );
  AND2_X1 U12566 ( .A1(n18317), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n18301) );
  NAND2_X1 U12567 ( .A1(n18422), .A2(n9641), .ZN(n18413) );
  INV_X1 U12568 ( .A(n18426), .ZN(n18422) );
  NAND2_X1 U12569 ( .A1(n18422), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n18421) );
  NAND2_X1 U12570 ( .A1(n18427), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n18426) );
  NAND2_X1 U12571 ( .A1(n18475), .A2(n9642), .ZN(n18431) );
  NAND2_X1 U12572 ( .A1(n18475), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18471) );
  NOR2_X2 U12573 ( .A1(n18396), .A2(n18522), .ZN(n18469) );
  NOR2_X1 U12574 ( .A1(n18479), .A2(n18642), .ZN(n18475) );
  NOR2_X1 U12575 ( .A1(n18508), .A2(n10062), .ZN(n18480) );
  NAND2_X1 U12576 ( .A1(n18480), .A2(P3_EAX_REG_14__SCAN_IN), .ZN(n18479) );
  NAND2_X1 U12577 ( .A1(n18395), .A2(n18513), .ZN(n18508) );
  AND2_X1 U12578 ( .A1(n18395), .A2(n11836), .ZN(n18512) );
  OR2_X1 U12579 ( .A1(n11674), .A2(n11673), .ZN(n18518) );
  NAND2_X1 U12580 ( .A1(n14508), .A2(n18395), .ZN(n18525) );
  INV_X1 U12581 ( .A(n18531), .ZN(n18528) );
  INV_X1 U12582 ( .A(n18512), .ZN(n18438) );
  INV_X1 U12583 ( .A(n18525), .ZN(n18530) );
  INV_X1 U12584 ( .A(n18395), .ZN(n14663) );
  INV_X1 U12585 ( .A(n18565), .ZN(n18575) );
  NOR2_X1 U12586 ( .A1(n18578), .A2(n18638), .ZN(n18633) );
  INV_X1 U12587 ( .A(n18619), .ZN(n18638) );
  OR2_X1 U12589 ( .A1(n11722), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U12590 ( .A1(n18730), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14732) );
  NAND2_X1 U12591 ( .A1(n9898), .A2(n14875), .ZN(n17216) );
  INV_X1 U12592 ( .A(n18810), .ZN(n9898) );
  NAND2_X1 U12593 ( .A1(n9937), .A2(n11659), .ZN(n14171) );
  NAND2_X1 U12594 ( .A1(n14159), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9937) );
  INV_X1 U12595 ( .A(n19479), .ZN(n19515) );
  INV_X1 U12596 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18882) );
  INV_X1 U12597 ( .A(n17286), .ZN(n17302) );
  INV_X1 U12598 ( .A(n10314), .ZN(n17188) );
  NAND2_X1 U12599 ( .A1(n9928), .A2(n9927), .ZN(n17202) );
  NAND2_X1 U12600 ( .A1(n17335), .A2(n10248), .ZN(n17338) );
  NAND2_X1 U12601 ( .A1(n10249), .A2(n18978), .ZN(n10248) );
  INV_X1 U12602 ( .A(n18927), .ZN(n10249) );
  NOR2_X1 U12603 ( .A1(n14385), .A2(n10324), .ZN(n17219) );
  NAND2_X1 U12604 ( .A1(n14385), .A2(n18795), .ZN(n17254) );
  NAND2_X1 U12605 ( .A1(n10238), .A2(n10239), .ZN(n14151) );
  INV_X1 U12606 ( .A(n11919), .ZN(n10242) );
  AND2_X1 U12607 ( .A1(n11891), .A2(n19743), .ZN(n19053) );
  INV_X1 U12608 ( .A(n19053), .ZN(n19121) );
  NOR2_X1 U12609 ( .A1(n19077), .A2(n19121), .ZN(n19119) );
  INV_X1 U12610 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19583) );
  NOR2_X1 U12611 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19740), .ZN(n19628) );
  INV_X1 U12612 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19723) );
  OR2_X1 U12613 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19638), .ZN(n19731) );
  INV_X2 U12614 ( .A(n19731), .ZN(n19749) );
  NOR2_X1 U12615 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13761), .ZN(n17632)
         );
  NAND2_X1 U12617 ( .A1(n10118), .A2(n10117), .ZN(P1_U2842) );
  AOI21_X1 U12618 ( .B1(n14950), .B2(n20708), .A(n9733), .ZN(n10117) );
  INV_X1 U12619 ( .A(n14950), .ZN(n15337) );
  OAI21_X1 U12620 ( .B1(n15659), .B2(n20633), .A(n10308), .ZN(P1_U2972) );
  INV_X1 U12621 ( .A(n10309), .ZN(n10308) );
  INV_X1 U12622 ( .A(n15440), .ZN(n10380) );
  AND2_X1 U12623 ( .A1(n9926), .A2(n13755), .ZN(n13756) );
  NAND2_X1 U12624 ( .A1(n10068), .A2(n9724), .ZN(P1_U3011) );
  INV_X1 U12625 ( .A(n13275), .ZN(n13276) );
  NOR2_X1 U12626 ( .A1(n13266), .A2(n13265), .ZN(n13277) );
  OAI21_X1 U12627 ( .B1(n13707), .B2(n16353), .A(n13274), .ZN(n13275) );
  NAND2_X1 U12628 ( .A1(n15954), .A2(n10285), .ZN(P2_U2826) );
  AOI21_X1 U12629 ( .B1(n10289), .B2(n10288), .A(n10286), .ZN(n10285) );
  NOR2_X1 U12630 ( .A1(n13729), .A2(n13728), .ZN(n13730) );
  NOR2_X1 U12631 ( .A1(n13707), .A2(n16459), .ZN(n13729) );
  INV_X1 U12632 ( .A(n13306), .ZN(n13310) );
  OAI211_X1 U12633 ( .C1(n10030), .C2(n9983), .A(n13307), .B(n9982), .ZN(
        n13309) );
  OAI21_X1 U12634 ( .B1(n16369), .B2(n19838), .A(n13305), .ZN(n13306) );
  INV_X1 U12635 ( .A(n16572), .ZN(n10027) );
  NAND2_X1 U12636 ( .A1(n16573), .A2(n13307), .ZN(n10029) );
  AOI21_X1 U12637 ( .B1(n16874), .B2(n13307), .A(n16586), .ZN(n16587) );
  INV_X1 U12638 ( .A(n10009), .ZN(n10327) );
  OAI21_X1 U12639 ( .B1(n10326), .B2(n16592), .A(n10010), .ZN(n10009) );
  INV_X1 U12640 ( .A(n10143), .ZN(n10142) );
  NAND2_X1 U12641 ( .A1(n9652), .A2(n10138), .ZN(n10141) );
  AOI21_X1 U12642 ( .B1(n16913), .B2(n16827), .A(n16628), .ZN(n9964) );
  NAND2_X1 U12643 ( .A1(n16932), .A2(n13307), .ZN(n9800) );
  NOR2_X1 U12644 ( .A1(n16655), .A2(n16846), .ZN(n9824) );
  AOI21_X1 U12645 ( .B1(n16686), .B2(n16827), .A(n16685), .ZN(n10255) );
  NAND2_X1 U12646 ( .A1(n10258), .A2(n10257), .ZN(n10256) );
  NAND2_X1 U12647 ( .A1(n9786), .A2(n13307), .ZN(n16781) );
  OAI211_X1 U12648 ( .C1(n13731), .C2(n17139), .A(n13745), .B(n9688), .ZN(
        P2_U3015) );
  NAND2_X1 U12649 ( .A1(n13308), .A2(n17136), .ZN(n13745) );
  NAND2_X1 U12650 ( .A1(n16440), .A2(n17121), .ZN(n13747) );
  NAND2_X1 U12651 ( .A1(n11522), .A2(n17121), .ZN(n11534) );
  INV_X1 U12652 ( .A(n11501), .ZN(n11507) );
  NAND2_X1 U12653 ( .A1(n16573), .A2(n17136), .ZN(n11506) );
  NOR2_X1 U12654 ( .A1(n11546), .A2(n9646), .ZN(n11547) );
  OAI21_X1 U12655 ( .B1(n16922), .B2(n17124), .A(n10301), .ZN(P2_U3023) );
  NAND2_X1 U12656 ( .A1(n10304), .A2(n10303), .ZN(n10302) );
  INV_X1 U12657 ( .A(n16911), .ZN(n10305) );
  OR2_X1 U12658 ( .A1(n14900), .A2(n17136), .ZN(n9894) );
  NOR2_X1 U12659 ( .A1(n16655), .A2(n17124), .ZN(n9823) );
  NAND2_X1 U12660 ( .A1(n16967), .A2(n10339), .ZN(n10338) );
  NAND2_X1 U12661 ( .A1(n13169), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13170) );
  NAND2_X1 U12662 ( .A1(n9786), .A2(n17136), .ZN(n17063) );
  NAND2_X1 U12663 ( .A1(n10002), .A2(n9998), .ZN(P3_U2642) );
  AND2_X1 U12664 ( .A1(n17690), .A2(n9999), .ZN(n9998) );
  NOR2_X1 U12665 ( .A1(n17687), .A2(n10000), .ZN(n9999) );
  INV_X1 U12666 ( .A(n18096), .ZN(n17458) );
  NOR2_X1 U12667 ( .A1(n18149), .A2(n18049), .ZN(n18115) );
  AND2_X1 U12668 ( .A1(n18317), .A2(n9639), .ZN(n18264) );
  NAND2_X1 U12669 ( .A1(n10222), .A2(n10220), .ZN(n18391) );
  NOR2_X1 U12670 ( .A1(n14736), .A2(n9808), .ZN(n14737) );
  INV_X1 U12671 ( .A(n18681), .ZN(n18673) );
  AND2_X1 U12672 ( .A1(n11961), .A2(n11960), .ZN(n11962) );
  AOI21_X1 U12673 ( .B1(n18924), .B2(n18923), .A(n10244), .ZN(n18925) );
  AND2_X1 U12674 ( .A1(n19089), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n10244) );
  INV_X1 U12675 ( .A(n18054), .ZN(n18327) );
  INV_X1 U12676 ( .A(n17461), .ZN(n11735) );
  INV_X1 U12677 ( .A(n11628), .ZN(n18323) );
  AND2_X1 U12678 ( .A1(n15506), .A2(n9751), .ZN(n9600) );
  AND2_X1 U12679 ( .A1(n14033), .A2(n11562), .ZN(n17376) );
  INV_X1 U12680 ( .A(n11606), .ZN(n18253) );
  NAND2_X1 U12681 ( .A1(n9714), .A2(n11415), .ZN(n14250) );
  NAND2_X1 U12682 ( .A1(n10412), .A2(n14436), .ZN(n14435) );
  NAND3_X1 U12683 ( .A1(n9802), .A2(n10051), .A3(n9630), .ZN(n10939) );
  AND4_X1 U12684 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_8__SCAN_IN), .ZN(n9603) );
  INV_X1 U12685 ( .A(n18170), .ZN(n18321) );
  INV_X2 U12686 ( .A(n13475), .ZN(n10757) );
  NAND2_X1 U12687 ( .A1(n11709), .A2(n18712), .ZN(n18677) );
  INV_X1 U12688 ( .A(n12083), .ZN(n10083) );
  NOR2_X1 U12689 ( .A1(n10298), .A2(n10297), .ZN(n13197) );
  NOR2_X1 U12690 ( .A1(n10348), .A2(n10345), .ZN(n14382) );
  AND2_X1 U12691 ( .A1(n12196), .A2(n12872), .ZN(n9604) );
  INV_X1 U12692 ( .A(n20885), .ZN(n12036) );
  AND3_X1 U12693 ( .A1(n9594), .A2(n10096), .A3(n14580), .ZN(n9605) );
  INV_X1 U12694 ( .A(n15253), .ZN(n13101) );
  OR2_X1 U12695 ( .A1(n10944), .A2(n10372), .ZN(n9606) );
  AND2_X1 U12696 ( .A1(n10394), .A2(n14269), .ZN(n9607) );
  AND2_X1 U12697 ( .A1(n9607), .A2(n10392), .ZN(n9608) );
  NAND2_X1 U12698 ( .A1(n16103), .A2(n9716), .ZN(n16021) );
  NAND2_X1 U12699 ( .A1(n11029), .A2(n11031), .ZN(n11041) );
  INV_X1 U12700 ( .A(n14065), .ZN(n11564) );
  INV_X1 U12701 ( .A(n9844), .ZN(n9992) );
  AND2_X1 U12702 ( .A1(n13014), .A2(n15223), .ZN(n9611) );
  AND4_X1 U12703 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n9612) );
  AND2_X1 U12704 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n9613) );
  AND2_X1 U12705 ( .A1(n9574), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n9614) );
  AND2_X2 U12706 ( .A1(n10668), .A2(n10669), .ZN(n13534) );
  AND3_X1 U12707 ( .A1(n14832), .A2(n14838), .A3(n9698), .ZN(n9615) );
  AND2_X1 U12708 ( .A1(n18677), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9616) );
  NAND2_X1 U12709 ( .A1(n12946), .A2(n15583), .ZN(n10025) );
  NOR3_X1 U12710 ( .A1(n15975), .A2(n15974), .A3(n9732), .ZN(n10400) );
  AND4_X1 U12711 ( .A1(n11763), .A2(n11762), .A3(n11761), .A4(n11760), .ZN(
        n9618) );
  AND2_X1 U12712 ( .A1(n10049), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n9620) );
  INV_X1 U12713 ( .A(n19904), .ZN(n10797) );
  AND2_X1 U12714 ( .A1(n13700), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9621) );
  INV_X1 U12715 ( .A(n10070), .ZN(n15477) );
  INV_X1 U12716 ( .A(n15477), .ZN(n10430) );
  AND2_X1 U12717 ( .A1(n10378), .A2(n9725), .ZN(n9623) );
  AND2_X1 U12718 ( .A1(n11169), .A2(n11047), .ZN(n9624) );
  INV_X1 U12719 ( .A(n16830), .ZN(n9953) );
  AND2_X1 U12720 ( .A1(n11163), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9625) );
  NOR2_X1 U12721 ( .A1(n9604), .A2(n12094), .ZN(n9626) );
  AND2_X1 U12722 ( .A1(n10657), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n9627) );
  AND2_X1 U12723 ( .A1(n18389), .A2(n19171), .ZN(n18385) );
  NAND2_X1 U12724 ( .A1(n9805), .A2(n10589), .ZN(n11235) );
  INV_X1 U12725 ( .A(n15583), .ZN(n10434) );
  OR2_X1 U12726 ( .A1(n17124), .A2(n16974), .ZN(n9628) );
  NAND2_X1 U12727 ( .A1(n10393), .A2(n9607), .ZN(n14268) );
  OR2_X1 U12728 ( .A1(n18381), .A2(n10230), .ZN(n18376) );
  INV_X2 U12729 ( .A(n20708), .ZN(n15330) );
  AND2_X1 U12730 ( .A1(n9742), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9629) );
  NAND2_X1 U12731 ( .A1(n9782), .A2(n9780), .ZN(n14328) );
  AND2_X1 U12732 ( .A1(n10750), .A2(n10265), .ZN(n9630) );
  AND2_X1 U12733 ( .A1(n15595), .A2(n15642), .ZN(n9631) );
  NAND2_X1 U12734 ( .A1(n10393), .A2(n9608), .ZN(n10395) );
  OR2_X1 U12735 ( .A1(n13576), .A2(n9740), .ZN(n9632) );
  OR2_X1 U12736 ( .A1(n9628), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9633) );
  AND2_X1 U12737 ( .A1(n10416), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9634) );
  AND2_X1 U12738 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .ZN(n9635) );
  NAND2_X1 U12739 ( .A1(n11719), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9636) );
  AND2_X1 U12740 ( .A1(n10856), .A2(n9753), .ZN(n9637) );
  OR2_X1 U12741 ( .A1(n18712), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9638) );
  INV_X1 U12742 ( .A(n13868), .ZN(n10102) );
  AND2_X1 U12743 ( .A1(n9635), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n9639) );
  AND2_X1 U12744 ( .A1(n10448), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9640) );
  AND2_X1 U12745 ( .A1(n10060), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9641) );
  AND2_X1 U12746 ( .A1(n10057), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n9642) );
  AND2_X1 U12747 ( .A1(n9984), .A2(n13190), .ZN(n9643) );
  INV_X1 U12748 ( .A(n18218), .ZN(n18345) );
  AND2_X2 U12749 ( .A1(n13507), .A2(n10671), .ZN(n10686) );
  OR2_X1 U12750 ( .A1(n19582), .A2(n19623), .ZN(n9644) );
  AND2_X1 U12751 ( .A1(n17200), .A2(n10484), .ZN(n11722) );
  INV_X2 U12752 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10669) );
  NAND2_X1 U12753 ( .A1(n10990), .A2(n10378), .ZN(n10979) );
  INV_X1 U12754 ( .A(n18330), .ZN(n18352) );
  NOR2_X1 U12755 ( .A1(n15098), .A2(n15053), .ZN(n9645) );
  XNOR2_X1 U12756 ( .A(n13368), .B(n13366), .ZN(n14098) );
  INV_X1 U12757 ( .A(n10217), .ZN(n17647) );
  OR3_X1 U12758 ( .A1(n11946), .A2(n19140), .A3(n10218), .ZN(n10217) );
  NOR2_X1 U12759 ( .A1(n14679), .A2(n10011), .ZN(n15239) );
  OR2_X2 U12760 ( .A1(n11695), .A2(n18515), .ZN(n18712) );
  NAND2_X1 U12761 ( .A1(n14660), .A2(n14659), .ZN(n14658) );
  AND2_X1 U12762 ( .A1(n16469), .A2(n17121), .ZN(n9646) );
  NAND2_X1 U12763 ( .A1(n15220), .A2(n15222), .ZN(n15202) );
  INV_X1 U12764 ( .A(n10179), .ZN(n10826) );
  AND4_X1 U12765 ( .A1(n12969), .A2(n12094), .A3(n12084), .A4(n20885), .ZN(
        n9647) );
  AND2_X1 U12766 ( .A1(n15551), .A2(n12939), .ZN(n9648) );
  NOR2_X1 U12767 ( .A1(n13279), .A2(n13278), .ZN(n9649) );
  INV_X1 U12768 ( .A(n10254), .ZN(n18665) );
  NAND2_X1 U12769 ( .A1(n10334), .A2(n14784), .ZN(n10649) );
  AND2_X1 U12770 ( .A1(n10467), .A2(n9583), .ZN(n9650) );
  NOR2_X1 U12771 ( .A1(n16035), .A2(n16036), .ZN(n16018) );
  AND2_X1 U12772 ( .A1(n11103), .A2(n10410), .ZN(n9651) );
  AND2_X1 U12773 ( .A1(n10146), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9652) );
  NAND2_X1 U12774 ( .A1(n16661), .A2(n16939), .ZN(n9653) );
  NOR2_X1 U12775 ( .A1(n16423), .A2(n16424), .ZN(n16418) );
  AND2_X1 U12776 ( .A1(n10164), .A2(n10163), .ZN(n9654) );
  AND2_X1 U12777 ( .A1(n16103), .A2(n11480), .ZN(n9655) );
  NAND2_X1 U12778 ( .A1(n10968), .A2(n10376), .ZN(n9656) );
  AND4_X1 U12779 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(
        n9657) );
  OR3_X1 U12780 ( .A1(n18149), .A2(n10224), .A3(n18049), .ZN(n9658) );
  NAND2_X1 U12781 ( .A1(n10968), .A2(n10374), .ZN(n9659) );
  INV_X1 U12782 ( .A(n18730), .ZN(n18725) );
  AND2_X1 U12783 ( .A1(n18906), .A2(n18801), .ZN(n18730) );
  AOI21_X1 U12784 ( .B1(n12909), .B2(n12464), .A(n12326), .ZN(n14678) );
  AND4_X1 U12785 ( .A1(n16681), .A2(n14810), .A3(n11026), .A4(n16702), .ZN(
        n9660) );
  AND4_X1 U12786 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n9661) );
  OR2_X1 U12787 ( .A1(n13211), .A2(n16719), .ZN(n9662) );
  INV_X1 U12788 ( .A(n13359), .ZN(n14784) );
  CLKBUF_X3 U12789 ( .A(n13359), .Z(n13361) );
  AND2_X1 U12790 ( .A1(n16054), .A2(n16635), .ZN(n9663) );
  INV_X1 U12791 ( .A(n9593), .ZN(n20620) );
  NOR2_X1 U12792 ( .A1(n13196), .A2(n10296), .ZN(n13192) );
  AND2_X1 U12793 ( .A1(n11716), .A2(n17307), .ZN(n9664) );
  NAND2_X1 U12794 ( .A1(n9784), .A2(n10270), .ZN(n16823) );
  OAI21_X1 U12795 ( .B1(n9602), .B2(n10075), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10071) );
  AND2_X1 U12796 ( .A1(n9651), .A2(n10409), .ZN(n9665) );
  OR2_X1 U12797 ( .A1(n16171), .A2(n11513), .ZN(n9666) );
  OR2_X1 U12798 ( .A1(n11752), .A2(n11751), .ZN(n19166) );
  AND2_X1 U12799 ( .A1(n10268), .A2(n16595), .ZN(n9667) );
  AND2_X1 U12800 ( .A1(n12107), .A2(n10190), .ZN(n9668) );
  AND2_X1 U12801 ( .A1(n10520), .A2(n10521), .ZN(n9669) );
  AND3_X1 U12802 ( .A1(n10280), .A2(n10279), .A3(n10278), .ZN(n9670) );
  AND2_X1 U12803 ( .A1(n12085), .A2(n12113), .ZN(n9671) );
  AND2_X1 U12804 ( .A1(n10013), .A2(n15238), .ZN(n9672) );
  AND2_X1 U12805 ( .A1(n13700), .A2(n9590), .ZN(n9673) );
  NAND2_X1 U12806 ( .A1(n10116), .A2(n10334), .ZN(n20366) );
  OR3_X1 U12807 ( .A1(n10743), .A2(n10742), .A3(n10741), .ZN(n10880) );
  AND2_X1 U12808 ( .A1(n10157), .A2(n13307), .ZN(n9674) );
  OR2_X1 U12809 ( .A1(n11036), .A2(n16928), .ZN(n16631) );
  AND3_X1 U12810 ( .A1(n10648), .A2(n13361), .A3(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n9675) );
  OR2_X1 U12811 ( .A1(n14615), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9676) );
  NAND2_X1 U12812 ( .A1(n17833), .A2(n18697), .ZN(n9677) );
  AND4_X1 U12813 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n9679) );
  AND2_X1 U12814 ( .A1(n9960), .A2(n9957), .ZN(n9680) );
  AND2_X1 U12815 ( .A1(n19153), .A2(n19157), .ZN(n9681) );
  NAND2_X1 U12816 ( .A1(n14660), .A2(n10398), .ZN(n14673) );
  OR2_X1 U12817 ( .A1(n10418), .A2(n13157), .ZN(n9682) );
  INV_X1 U12818 ( .A(n10025), .ZN(n10024) );
  AND2_X1 U12819 ( .A1(n18710), .A2(n11719), .ZN(n9683) );
  AND2_X1 U12820 ( .A1(n11079), .A2(n11078), .ZN(n14326) );
  OR2_X1 U12821 ( .A1(n16903), .A2(n19838), .ZN(n9684) );
  AND3_X1 U12822 ( .A1(n13708), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10558), 
        .ZN(n9685) );
  INV_X1 U12823 ( .A(n9924), .ZN(n9923) );
  NOR2_X1 U12824 ( .A1(n13752), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9924) );
  INV_X1 U12825 ( .A(n16347), .ZN(n10646) );
  NAND2_X1 U12826 ( .A1(n10023), .A2(n10022), .ZN(n9686) );
  AND2_X1 U12827 ( .A1(n10806), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n9687) );
  AND2_X1 U12828 ( .A1(n13746), .A2(n13747), .ZN(n9688) );
  NAND2_X1 U12829 ( .A1(n10990), .A2(n9623), .ZN(n9689) );
  AND2_X1 U12830 ( .A1(n9684), .A2(n10145), .ZN(n9690) );
  OR2_X1 U12831 ( .A1(n16964), .A2(n16863), .ZN(n9691) );
  NAND2_X1 U12832 ( .A1(n9913), .A2(n9602), .ZN(n15459) );
  NOR2_X1 U12833 ( .A1(n11170), .A2(n16597), .ZN(n13284) );
  INV_X1 U12834 ( .A(n13284), .ZN(n9837) );
  AND2_X1 U12835 ( .A1(n11279), .A2(n11205), .ZN(n9692) );
  OAI21_X1 U12836 ( .B1(n16795), .B2(n17068), .A(n10154), .ZN(n10333) );
  INV_X1 U12837 ( .A(n10333), .ZN(n10853) );
  AND3_X1 U12838 ( .A1(n11733), .A2(n11732), .A3(n11734), .ZN(n9693) );
  INV_X1 U12839 ( .A(n10604), .ZN(n10166) );
  AND2_X1 U12840 ( .A1(n10334), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9694) );
  INV_X1 U12841 ( .A(n10825), .ZN(n9979) );
  AND2_X1 U12842 ( .A1(n13361), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9696) );
  NOR2_X1 U12843 ( .A1(n13112), .A2(n10190), .ZN(n9697) );
  AND2_X1 U12844 ( .A1(n16650), .A2(n16662), .ZN(n9698) );
  AND2_X1 U12845 ( .A1(n15182), .A2(n15194), .ZN(n9699) );
  NOR2_X1 U12846 ( .A1(n18809), .A2(n19024), .ZN(n9700) );
  AND2_X1 U12847 ( .A1(n12939), .A2(n12941), .ZN(n9701) );
  INV_X1 U12848 ( .A(n10937), .ZN(n9793) );
  AND2_X1 U12849 ( .A1(n12969), .A2(n20885), .ZN(n9702) );
  AND2_X1 U12850 ( .A1(n11305), .A2(n11311), .ZN(n9703) );
  AND2_X1 U12851 ( .A1(n9799), .A2(n16638), .ZN(n9704) );
  AND2_X1 U12852 ( .A1(n10310), .A2(n10128), .ZN(n9705) );
  AND2_X1 U12853 ( .A1(n9863), .A2(n11547), .ZN(n9706) );
  INV_X1 U12854 ( .A(n10054), .ZN(n10277) );
  NAND2_X1 U12855 ( .A1(n14841), .A2(n10053), .ZN(n10054) );
  AND2_X1 U12856 ( .A1(n9591), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U12857 ( .A1(n20859), .A2(n9585), .ZN(n9708) );
  AND2_X1 U12858 ( .A1(n9623), .A2(n10976), .ZN(n9709) );
  NAND2_X1 U12859 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11920), .ZN(
        n9710) );
  AND2_X1 U12860 ( .A1(n10658), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9711) );
  INV_X1 U12861 ( .A(n13930), .ZN(n20617) );
  AND2_X1 U12862 ( .A1(n10578), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13930) );
  NAND2_X1 U12863 ( .A1(n9706), .A2(n9853), .ZN(P2_U3020) );
  INV_X1 U12864 ( .A(n10663), .ZN(n13483) );
  NAND2_X1 U12865 ( .A1(n10281), .A2(n13191), .ZN(n13243) );
  NAND2_X1 U12867 ( .A1(n12094), .A2(n12083), .ZN(n10084) );
  INV_X2 U12868 ( .A(n16430), .ZN(n16438) );
  NAND2_X1 U12869 ( .A1(n10907), .A2(n10908), .ZN(n10945) );
  OR2_X1 U12870 ( .A1(n10346), .A2(n10348), .ZN(n9713) );
  NAND2_X1 U12871 ( .A1(n13045), .A2(n13044), .ZN(n15085) );
  INV_X1 U12872 ( .A(n15085), .ZN(n10124) );
  NOR2_X1 U12873 ( .A1(n18263), .A2(n17836), .ZN(n18205) );
  AND2_X1 U12874 ( .A1(n18364), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n18316) );
  AND2_X1 U12875 ( .A1(n14163), .A2(n14195), .ZN(n9714) );
  INV_X1 U12876 ( .A(n9714), .ZN(n10348) );
  NOR2_X1 U12877 ( .A1(n14400), .A2(n10390), .ZN(n14325) );
  NAND2_X1 U12878 ( .A1(n10412), .A2(n10411), .ZN(n14441) );
  NAND2_X1 U12879 ( .A1(n11495), .A2(n13700), .ZN(n11236) );
  INV_X1 U12880 ( .A(n17124), .ZN(n17136) );
  INV_X1 U12881 ( .A(n10007), .ZN(n10946) );
  NAND2_X1 U12882 ( .A1(n10907), .A2(n10008), .ZN(n10007) );
  AND2_X1 U12883 ( .A1(n18422), .A2(n10060), .ZN(n9715) );
  INV_X1 U12884 ( .A(n10907), .ZN(n10373) );
  INV_X1 U12885 ( .A(n12209), .ZN(n10386) );
  INV_X1 U12886 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n13189) );
  AND2_X1 U12887 ( .A1(n11480), .A2(n16046), .ZN(n9716) );
  AND2_X1 U12888 ( .A1(n10476), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13222) );
  NAND2_X1 U12889 ( .A1(n16626), .A2(n16635), .ZN(n10284) );
  NOR2_X1 U12890 ( .A1(n14441), .A2(n9777), .ZN(n14682) );
  NAND2_X1 U12891 ( .A1(n13151), .A2(n11103), .ZN(n13149) );
  NOR2_X1 U12892 ( .A1(n14400), .A2(n14401), .ZN(n14267) );
  INV_X1 U12893 ( .A(n16597), .ZN(n9864) );
  OR2_X2 U12894 ( .A1(n14304), .A2(n15918), .ZN(n20633) );
  INV_X1 U12895 ( .A(n20633), .ZN(n20779) );
  AND2_X1 U12896 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n9717) );
  AND2_X1 U12897 ( .A1(n9716), .A2(n10351), .ZN(n9718) );
  OAI21_X1 U12898 ( .B1(n16273), .B2(n16274), .A(n11323), .ZN(n13982) );
  NAND2_X1 U12899 ( .A1(n14800), .A2(n11305), .ZN(n14642) );
  AND2_X1 U12900 ( .A1(n13222), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13225) );
  NOR2_X1 U12901 ( .A1(n14189), .A2(n14238), .ZN(n14239) );
  AND2_X1 U12902 ( .A1(n16663), .A2(n16662), .ZN(n9719) );
  AND2_X1 U12903 ( .A1(n16713), .A2(n16712), .ZN(n9720) );
  XOR2_X1 U12904 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .Z(n9721) );
  AND2_X1 U12905 ( .A1(n12084), .A2(n20854), .ZN(n12953) );
  AND2_X1 U12906 ( .A1(n13244), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13246) );
  AND2_X1 U12907 ( .A1(n18184), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n18164) );
  AND2_X1 U12908 ( .A1(n13240), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13244) );
  OR3_X1 U12909 ( .A1(n13211), .A2(n10294), .A3(n10293), .ZN(n9722) );
  AND2_X1 U12910 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19628), .ZN(n19743) );
  AND2_X1 U12911 ( .A1(n10473), .A2(n10366), .ZN(n9723) );
  NOR2_X1 U12912 ( .A1(n15738), .A2(n10067), .ZN(n9724) );
  OR2_X1 U12913 ( .A1(n10902), .A2(n16135), .ZN(n9725) );
  OR2_X1 U12914 ( .A1(n10770), .A2(n10769), .ZN(n11312) );
  INV_X1 U12915 ( .A(n11312), .ZN(n10266) );
  AND2_X1 U12916 ( .A1(n9920), .A2(n9583), .ZN(n9726) );
  AND2_X1 U12917 ( .A1(n10572), .A2(n10573), .ZN(n9727) );
  AND2_X1 U12918 ( .A1(n10389), .A2(n15222), .ZN(n9728) );
  OR2_X1 U12919 ( .A1(n11428), .A2(n11427), .ZN(n14442) );
  AND2_X1 U12920 ( .A1(n18475), .A2(n10057), .ZN(n9729) );
  AND2_X1 U12921 ( .A1(n13311), .A2(n9717), .ZN(n9730) );
  NAND2_X1 U12922 ( .A1(n12957), .A2(n9769), .ZN(n13092) );
  INV_X1 U12923 ( .A(n13092), .ZN(n9768) );
  NAND2_X1 U12924 ( .A1(n9581), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9731) );
  OR2_X1 U12925 ( .A1(n10401), .A2(n10404), .ZN(n9732) );
  OR2_X1 U12926 ( .A1(n20869), .A2(n14376), .ZN(n12238) );
  NOR2_X1 U12927 ( .A1(n20712), .A2(n13145), .ZN(n9733) );
  INV_X1 U12928 ( .A(n14328), .ZN(n10412) );
  AND2_X1 U12929 ( .A1(n10168), .A2(n10167), .ZN(n9734) );
  AND2_X1 U12930 ( .A1(n12950), .A2(n9585), .ZN(n9735) );
  NAND2_X1 U12931 ( .A1(n9568), .A2(n11212), .ZN(n9736) );
  OR2_X1 U12932 ( .A1(n9977), .A2(n9976), .ZN(n9737) );
  INV_X1 U12933 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16719) );
  OR2_X1 U12934 ( .A1(n17116), .A2(n14784), .ZN(n9738) );
  INV_X1 U12935 ( .A(n10283), .ZN(n11149) );
  AND2_X1 U12936 ( .A1(n10376), .A2(n10969), .ZN(n9739) );
  INV_X1 U12937 ( .A(n12898), .ZN(n9920) );
  INV_X1 U12938 ( .A(n18294), .ZN(n18214) );
  NAND2_X1 U12939 ( .A1(n11552), .A2(n11564), .ZN(n11623) );
  NOR2_X1 U12940 ( .A1(n19752), .A2(n11947), .ZN(n19586) );
  NAND2_X1 U12941 ( .A1(n11146), .A2(n17491), .ZN(n16863) );
  NOR2_X1 U12942 ( .A1(n14729), .A2(n17685), .ZN(n13318) );
  NOR2_X1 U12943 ( .A1(n18381), .A2(n10229), .ZN(n14713) );
  OR2_X1 U12944 ( .A1(n16424), .A2(n10405), .ZN(n9740) );
  NOR2_X1 U12945 ( .A1(n18381), .A2(n18012), .ZN(n18379) );
  OR2_X1 U12946 ( .A1(n17212), .A2(n9996), .ZN(n9741) );
  AND2_X1 U12947 ( .A1(n13313), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14730) );
  AND2_X1 U12948 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9742) );
  OR3_X1 U12949 ( .A1(n19024), .A2(n19035), .A3(n18997), .ZN(n9743) );
  AND2_X1 U12950 ( .A1(n13570), .A2(n13569), .ZN(n16407) );
  NAND2_X1 U12951 ( .A1(n10577), .A2(n10576), .ZN(n13699) );
  AND2_X1 U12952 ( .A1(n13313), .A2(n9717), .ZN(n13312) );
  OR2_X1 U12953 ( .A1(n20878), .A2(n21373), .ZN(n12364) );
  INV_X1 U12954 ( .A(n12364), .ZN(n12464) );
  AND2_X1 U12955 ( .A1(n13942), .A2(n10104), .ZN(n9744) );
  OR2_X1 U12956 ( .A1(n14357), .A2(n10111), .ZN(n9745) );
  INV_X1 U12957 ( .A(n14610), .ZN(n13385) );
  OR2_X1 U12958 ( .A1(n11445), .A2(n11444), .ZN(n14610) );
  INV_X1 U12959 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18012) );
  AND2_X1 U12960 ( .A1(n12221), .A2(n12084), .ZN(n12106) );
  AND2_X1 U12961 ( .A1(n9629), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9746) );
  AND2_X1 U12962 ( .A1(n9634), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9747) );
  INV_X1 U12963 ( .A(n13941), .ZN(n10232) );
  AND2_X1 U12964 ( .A1(n10243), .A2(n10242), .ZN(n9748) );
  AND2_X1 U12965 ( .A1(n10228), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n9749) );
  INV_X1 U12966 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18388) );
  INV_X1 U12967 ( .A(n17465), .ZN(n18358) );
  INV_X1 U12968 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10088) );
  INV_X1 U12969 ( .A(n20837), .ZN(n20778) );
  NAND2_X1 U12970 ( .A1(n21210), .A2(n13179), .ZN(n20837) );
  NAND2_X1 U12971 ( .A1(n13317), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18696) );
  AND3_X1 U12972 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17946) );
  NAND4_X1 U12973 ( .A1(n15497), .A2(n15733), .A3(n10092), .A4(n15480), .ZN(
        n9750) );
  NOR2_X1 U12974 ( .A1(n17233), .A2(n18864), .ZN(n17248) );
  INV_X1 U12975 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U12976 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17990) );
  AND3_X1 U12977 ( .A1(n15711), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n9751) );
  NOR2_X1 U12978 ( .A1(n14065), .A2(n14074), .ZN(n17478) );
  NOR2_X1 U12979 ( .A1(n16974), .A2(n16969), .ZN(n9752) );
  NOR2_X1 U12980 ( .A1(n11502), .A2(n16864), .ZN(n9753) );
  AND2_X1 U12981 ( .A1(n10158), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9754) );
  AND2_X1 U12982 ( .A1(n9639), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n9755) );
  OR2_X1 U12983 ( .A1(n19024), .A2(n19035), .ZN(n9756) );
  NOR2_X1 U12984 ( .A1(n15422), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9757) );
  INV_X1 U12985 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10090) );
  INV_X1 U12986 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n10061) );
  AND2_X1 U12987 ( .A1(n10415), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9758) );
  AND2_X1 U12988 ( .A1(n15879), .A2(n15878), .ZN(n9759) );
  INV_X1 U12989 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9939) );
  INV_X1 U12990 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16674) );
  INV_X1 U12991 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10317) );
  AND2_X1 U12992 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9760) );
  INV_X1 U12993 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20326) );
  AOI211_X1 U12994 ( .C1(n17678), .C2(n18025), .A(n17677), .B(n17676), .ZN(
        n17681) );
  AOI22_X2 U12995 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19892), .ZN(n20436) );
  AOI22_X2 U12996 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19892), .ZN(n20392) );
  AOI22_X2 U12997 ( .A1(DATAI_20_), .A2(n20839), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20883), .ZN(n21414) );
  AOI22_X2 U12998 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20883), .B1(DATAI_16_), 
        .B2(n20839), .ZN(n21341) );
  NOR2_X2 U12999 ( .A1(n20837), .A2(n20836), .ZN(n20883) );
  AOI22_X2 U13000 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19892), .ZN(n20430) );
  NOR2_X2 U13001 ( .A1(n19839), .A2(n19838), .ZN(n19892) );
  OR2_X1 U13002 ( .A1(n12468), .A2(n9585), .ZN(n12837) );
  AND2_X1 U13003 ( .A1(n12468), .A2(n14930), .ZN(n14923) );
  AND2_X1 U13004 ( .A1(n12468), .A2(n9759), .ZN(n15880) );
  NAND3_X1 U13005 ( .A1(n9761), .A2(n12959), .A3(n20854), .ZN(n12118) );
  NAND2_X1 U13006 ( .A1(n9761), .A2(n12959), .ZN(n12089) );
  NAND3_X1 U13007 ( .A1(n10034), .A2(n10033), .A3(n10178), .ZN(n9906) );
  NAND2_X1 U13008 ( .A1(n15595), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12942) );
  XNOR2_X1 U13009 ( .A(n12232), .B(n20995), .ZN(n14350) );
  NAND2_X1 U13010 ( .A1(n12754), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12074) );
  NAND2_X1 U13011 ( .A1(n12754), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12052) );
  AOI22_X1 U13012 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12012) );
  NAND3_X1 U13013 ( .A1(n9880), .A2(n15551), .A3(n9879), .ZN(n9765) );
  NAND2_X2 U13014 ( .A1(n9572), .A2(n12306), .ZN(n14679) );
  XNOR2_X2 U13015 ( .A(n9770), .B(n12148), .ZN(n12223) );
  INV_X1 U13016 ( .A(n14855), .ZN(n9771) );
  INV_X1 U13017 ( .A(n12277), .ZN(n9772) );
  INV_X1 U13018 ( .A(n10178), .ZN(n15873) );
  OR2_X2 U13019 ( .A1(n12202), .A2(n12203), .ZN(n12277) );
  AND2_X2 U13020 ( .A1(n9776), .A2(n9775), .ZN(n9796) );
  NAND2_X1 U13021 ( .A1(n9840), .A2(n10575), .ZN(n9775) );
  INV_X1 U13022 ( .A(n9839), .ZN(n9776) );
  NAND2_X1 U13023 ( .A1(n14682), .A2(n14687), .ZN(n14686) );
  NAND2_X1 U13024 ( .A1(n9779), .A2(n13380), .ZN(n14185) );
  INV_X1 U13025 ( .A(n9781), .ZN(n9780) );
  OR2_X1 U13026 ( .A1(n14197), .A2(n9783), .ZN(n9782) );
  INV_X1 U13027 ( .A(n13380), .ZN(n9783) );
  NOR2_X2 U13028 ( .A1(n16824), .A2(n9828), .ZN(n9827) );
  NAND3_X1 U13029 ( .A1(n9950), .A2(n9952), .A3(n9949), .ZN(n9784) );
  NAND2_X1 U13030 ( .A1(n14841), .A2(n10416), .ZN(n11503) );
  NAND2_X1 U13031 ( .A1(n9790), .A2(n11513), .ZN(n10063) );
  NAND2_X1 U13032 ( .A1(n9790), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10828) );
  INV_X1 U13033 ( .A(n9791), .ZN(n10576) );
  NAND2_X1 U13034 ( .A1(n9791), .A2(n10096), .ZN(n9840) );
  AND2_X1 U13035 ( .A1(n11287), .A2(n9791), .ZN(n11209) );
  NAND2_X2 U13036 ( .A1(n9796), .A2(n10460), .ZN(n11212) );
  OAI21_X2 U13037 ( .B1(n16606), .B2(n16608), .A(n16607), .ZN(n16632) );
  NAND2_X2 U13038 ( .A1(n10960), .A2(n10959), .ZN(n16606) );
  NAND3_X1 U13039 ( .A1(n10941), .A2(n16819), .A3(n10940), .ZN(n16766) );
  INV_X1 U13040 ( .A(n10936), .ZN(n9795) );
  NAND3_X1 U13041 ( .A1(n9794), .A2(n9792), .A3(n10938), .ZN(n9831) );
  NAND3_X1 U13042 ( .A1(n9793), .A2(n10936), .A3(n10311), .ZN(n9792) );
  NAND2_X1 U13043 ( .A1(n9796), .A2(n10155), .ZN(n10858) );
  NAND2_X1 U13044 ( .A1(n9796), .A2(n10098), .ZN(n13251) );
  NAND3_X1 U13045 ( .A1(n10136), .A2(n9796), .A3(n13930), .ZN(n10135) );
  NAND2_X1 U13046 ( .A1(n9797), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10608) );
  NAND2_X1 U13047 ( .A1(n11249), .A2(n10606), .ZN(n9797) );
  INV_X1 U13048 ( .A(n10605), .ZN(n9798) );
  NAND2_X1 U13049 ( .A1(n9800), .A2(n9704), .ZN(P2_U2992) );
  NAND2_X1 U13050 ( .A1(n10204), .A2(n10193), .ZN(n9801) );
  AND2_X2 U13051 ( .A1(n9802), .A2(n10744), .ZN(n10215) );
  NAND2_X1 U13052 ( .A1(n9569), .A2(n9842), .ZN(n16790) );
  NAND3_X1 U13053 ( .A1(n9569), .A2(n9842), .A3(n10853), .ZN(n9807) );
  OAI21_X1 U13054 ( .B1(n9811), .B2(n14735), .A(n9809), .ZN(n9808) );
  NAND2_X2 U13055 ( .A1(n9644), .A2(n14280), .ZN(n18906) );
  NAND2_X2 U13056 ( .A1(n11560), .A2(n11561), .ZN(n18256) );
  AND2_X2 U13057 ( .A1(n17345), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11560) );
  NOR2_X2 U13058 ( .A1(n18995), .A2(n19736), .ZN(n19585) );
  INV_X1 U13059 ( .A(n15512), .ZN(n9820) );
  NAND2_X1 U13060 ( .A1(n12928), .A2(n9915), .ZN(n9821) );
  NAND3_X1 U13061 ( .A1(n9877), .A2(n9908), .A3(n13173), .ZN(n9876) );
  AND2_X1 U13062 ( .A1(n9832), .A2(n9825), .ZN(n9833) );
  NAND2_X1 U13063 ( .A1(n10097), .A2(n9825), .ZN(n10280) );
  OR2_X4 U13064 ( .A1(n9827), .A2(n9826), .ZN(n14841) );
  OAI21_X2 U13065 ( .B1(n9842), .B2(n9828), .A(n10853), .ZN(n9826) );
  XNOR2_X2 U13066 ( .A(n10215), .B(n9980), .ZN(n14635) );
  NAND2_X2 U13067 ( .A1(n9830), .A2(n10020), .ZN(n10825) );
  NAND3_X1 U13068 ( .A1(n9830), .A2(n10020), .A3(n16853), .ZN(n9990) );
  NAND2_X1 U13069 ( .A1(n9990), .A2(n9844), .ZN(n9988) );
  NAND2_X1 U13070 ( .A1(n14635), .A2(n14636), .ZN(n9829) );
  AND2_X1 U13071 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n9832)
         );
  NAND2_X1 U13072 ( .A1(n9834), .A2(n14580), .ZN(n10606) );
  NAND4_X1 U13073 ( .A1(n10574), .A2(n10572), .A3(n10166), .A4(n10573), .ZN(
        n9834) );
  NAND2_X1 U13074 ( .A1(n10570), .A2(n19862), .ZN(n9835) );
  NAND2_X1 U13075 ( .A1(n11205), .A2(n10580), .ZN(n9836) );
  OAI21_X1 U13076 ( .B1(n10605), .B2(n13271), .A(n10606), .ZN(n10579) );
  AOI21_X2 U13077 ( .B1(n10352), .B2(n9667), .A(n9837), .ZN(n16578) );
  NAND2_X2 U13078 ( .A1(n16606), .A2(n10355), .ZN(n10352) );
  NAND2_X2 U13079 ( .A1(n10634), .A2(n10189), .ZN(n9838) );
  NAND2_X1 U13080 ( .A1(n10644), .A2(n9838), .ZN(n10643) );
  OAI21_X1 U13081 ( .B1(n10637), .B2(n9838), .A(n10618), .ZN(n10622) );
  NAND2_X1 U13082 ( .A1(n9904), .A2(n9838), .ZN(n13350) );
  NAND2_X2 U13083 ( .A1(n9841), .A2(n10581), .ZN(n10629) );
  AND4_X1 U13084 ( .A1(n10608), .A2(n9841), .A3(n10607), .A4(n10609), .ZN(
        n10610) );
  NAND2_X2 U13085 ( .A1(n9843), .A2(n10826), .ZN(n9842) );
  XNOR2_X1 U13086 ( .A(n10825), .B(n9992), .ZN(n16854) );
  NAND3_X1 U13087 ( .A1(n9852), .A2(n13700), .A3(n9707), .ZN(n9849) );
  AND2_X2 U13088 ( .A1(n13701), .A2(n13708), .ZN(n9852) );
  NAND3_X1 U13089 ( .A1(n9856), .A2(n9855), .A3(n9854), .ZN(n9863) );
  NAND2_X1 U13090 ( .A1(n11040), .A2(n9858), .ZN(n9854) );
  NAND3_X1 U13091 ( .A1(n9857), .A2(n17136), .A3(n10857), .ZN(n9853) );
  NAND3_X1 U13092 ( .A1(n9856), .A2(n9859), .A3(n9854), .ZN(n11548) );
  NOR2_X1 U13093 ( .A1(n9866), .A2(n9865), .ZN(n9869) );
  NAND3_X1 U13094 ( .A1(n10162), .A2(n10132), .A3(n10773), .ZN(n9865) );
  AND2_X2 U13095 ( .A1(n9867), .A2(n10795), .ZN(n10936) );
  NAND4_X1 U13096 ( .A1(n9872), .A2(n9869), .A3(n9870), .A4(n9868), .ZN(n9867)
         );
  INV_X1 U13097 ( .A(n9873), .ZN(n9872) );
  NAND3_X1 U13098 ( .A1(n16691), .A2(n10216), .A3(n13307), .ZN(n16698) );
  NAND2_X2 U13099 ( .A1(n9874), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16691) );
  NAND3_X1 U13100 ( .A1(n14805), .A2(n14804), .A3(n9738), .ZN(P2_U3044) );
  NAND4_X1 U13101 ( .A1(n10517), .A2(n10518), .A3(n10516), .A4(n10515), .ZN(
        n10553) );
  NAND2_X1 U13102 ( .A1(n10352), .A2(n10353), .ZN(n16599) );
  NAND2_X1 U13103 ( .A1(n9876), .A2(n9875), .ZN(n13176) );
  NAND2_X1 U13104 ( .A1(n9877), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9875) );
  NAND2_X1 U13105 ( .A1(n9908), .A2(n13173), .ZN(n9878) );
  XNOR2_X1 U13106 ( .A(n9878), .B(n15416), .ZN(n15640) );
  INV_X1 U13107 ( .A(n12935), .ZN(n9879) );
  NAND2_X1 U13108 ( .A1(n9890), .A2(n9894), .ZN(n14901) );
  NAND2_X1 U13109 ( .A1(n10444), .A2(n9891), .ZN(n9890) );
  NAND2_X1 U13110 ( .A1(n9892), .A2(n9896), .ZN(n14849) );
  NAND2_X1 U13111 ( .A1(n10444), .A2(n9893), .ZN(n9892) );
  AND2_X1 U13112 ( .A1(n10443), .A2(n9897), .ZN(n9893) );
  NAND2_X1 U13113 ( .A1(n9897), .A2(n16846), .ZN(n9896) );
  NAND3_X1 U13114 ( .A1(n11810), .A2(n11809), .A3(n11811), .ZN(n9900) );
  AND2_X2 U13115 ( .A1(n17226), .A2(n17294), .ZN(n18780) );
  NOR2_X2 U13116 ( .A1(n18998), .A2(n19586), .ZN(n19029) );
  NAND2_X2 U13117 ( .A1(n14068), .A2(n9902), .ZN(n18998) );
  INV_X1 U13118 ( .A(n10634), .ZN(n9905) );
  XNOR2_X1 U13119 ( .A(n9906), .B(n12329), .ZN(n12915) );
  AND2_X1 U13120 ( .A1(n12323), .A2(n9906), .ZN(n12909) );
  NAND2_X1 U13121 ( .A1(n13172), .A2(n15595), .ZN(n9908) );
  INV_X1 U13122 ( .A(n9945), .ZN(n9911) );
  NAND2_X1 U13123 ( .A1(n10070), .A2(n9914), .ZN(n9913) );
  NAND2_X1 U13124 ( .A1(n12278), .A2(n9583), .ZN(n9917) );
  NAND2_X1 U13125 ( .A1(n12901), .A2(n12898), .ZN(n9918) );
  INV_X1 U13126 ( .A(n12892), .ZN(n20774) );
  NAND3_X1 U13127 ( .A1(n9925), .A2(n9923), .A3(n9921), .ZN(n15672) );
  NAND3_X1 U13128 ( .A1(n9925), .A2(n9922), .A3(n9921), .ZN(n9926) );
  NAND3_X1 U13129 ( .A1(n13753), .A2(n13752), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9925) );
  AND2_X2 U13130 ( .A1(n12839), .A2(n14335), .ZN(n10106) );
  NAND2_X1 U13131 ( .A1(n12949), .A2(n13080), .ZN(n12839) );
  NAND3_X1 U13132 ( .A1(n9928), .A2(n9927), .A3(n11721), .ZN(n17200) );
  AOI21_X2 U13133 ( .B1(n10322), .B2(n18677), .A(n9636), .ZN(n18652) );
  NAND2_X1 U13134 ( .A1(n9931), .A2(n11616), .ZN(n13809) );
  NAND2_X1 U13135 ( .A1(n14119), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9931) );
  OAI21_X1 U13136 ( .B1(n14119), .B2(n9935), .A(n9932), .ZN(n11639) );
  NAND2_X1 U13137 ( .A1(n11616), .A2(n9934), .ZN(n9933) );
  INV_X1 U13138 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n9934) );
  INV_X1 U13139 ( .A(n11616), .ZN(n9935) );
  OAI21_X1 U13140 ( .B1(n9940), .B2(n14159), .A(n9936), .ZN(n11678) );
  NAND2_X2 U13141 ( .A1(n9657), .A2(n9610), .ZN(n14666) );
  NAND4_X1 U13142 ( .A1(n10319), .A2(n9657), .A3(n9610), .A4(n10318), .ZN(
        n9944) );
  NAND2_X1 U13143 ( .A1(n11617), .A2(n9944), .ZN(n11595) );
  OR2_X2 U13144 ( .A1(n18795), .A2(n18985), .ZN(n18713) );
  NAND2_X2 U13145 ( .A1(n11707), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18795) );
  NAND2_X1 U13146 ( .A1(n9948), .A2(n11312), .ZN(n10020) );
  INV_X1 U13147 ( .A(n10215), .ZN(n9948) );
  NAND3_X1 U13148 ( .A1(n9988), .A2(n10827), .A3(n10179), .ZN(n9949) );
  NAND2_X1 U13149 ( .A1(n16830), .A2(n10179), .ZN(n9951) );
  NAND4_X1 U13150 ( .A1(n9954), .A2(n10826), .A3(n9953), .A4(n9990), .ZN(n9952) );
  NAND3_X1 U13151 ( .A1(n17013), .A2(n17012), .A3(n13307), .ZN(n16737) );
  NAND2_X1 U13152 ( .A1(n10777), .A2(n10133), .ZN(n9955) );
  INV_X2 U13153 ( .A(n11205), .ZN(n19862) );
  NAND3_X1 U13154 ( .A1(n10532), .A2(n10534), .A3(n10533), .ZN(n9968) );
  NAND3_X1 U13155 ( .A1(n10475), .A2(n10537), .A3(n10538), .ZN(n9969) );
  NAND4_X1 U13156 ( .A1(n10512), .A2(n10514), .A3(n10513), .A4(n10511), .ZN(
        n10556) );
  NOR2_X2 U13157 ( .A1(n9973), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14540) );
  NAND3_X2 U13158 ( .A1(n14559), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10496) );
  NAND2_X1 U13159 ( .A1(n13160), .A2(n13159), .ZN(n14812) );
  NAND2_X1 U13160 ( .A1(n13251), .A2(n17493), .ZN(n11493) );
  NAND2_X1 U13161 ( .A1(n10613), .A2(n10612), .ZN(n10640) );
  OR2_X2 U13162 ( .A1(n11212), .A2(n10597), .ZN(n10614) );
  NAND2_X1 U13163 ( .A1(n10825), .A2(n16853), .ZN(n9991) );
  INV_X1 U13164 ( .A(n9980), .ZN(n10019) );
  NAND2_X2 U13165 ( .A1(n10051), .A2(n10750), .ZN(n9980) );
  NAND2_X1 U13166 ( .A1(n9980), .A2(n11312), .ZN(n10017) );
  NAND2_X1 U13167 ( .A1(n9987), .A2(n9953), .ZN(n16833) );
  NAND2_X1 U13168 ( .A1(n9989), .A2(n9988), .ZN(n9987) );
  NAND3_X1 U13169 ( .A1(n9991), .A2(n9992), .A3(n10825), .ZN(n9989) );
  NAND2_X1 U13170 ( .A1(n9992), .A2(n9979), .ZN(n10771) );
  NAND2_X1 U13171 ( .A1(n16854), .A2(n16853), .ZN(n10108) );
  NOR2_X1 U13172 ( .A1(n17753), .A2(n17754), .ZN(n17752) );
  INV_X1 U13173 ( .A(n17765), .ZN(n9994) );
  NOR2_X2 U13174 ( .A1(n17212), .A2(n9995), .ZN(n13317) );
  NAND3_X1 U13175 ( .A1(n17684), .A2(n10003), .A3(n18025), .ZN(n10002) );
  NAND2_X1 U13176 ( .A1(n17683), .A2(n17682), .ZN(n10003) );
  INV_X2 U13177 ( .A(n13331), .ZN(n18000) );
  AND2_X1 U13178 ( .A1(n10005), .A2(n10004), .ZN(n17785) );
  NAND2_X1 U13179 ( .A1(n13331), .A2(n9677), .ZN(n10005) );
  MUX2_X1 U13180 ( .A(n9591), .B(n11006), .S(n11005), .Z(n11008) );
  NOR2_X4 U13181 ( .A1(n14988), .A2(n14989), .ZN(n13750) );
  OAI21_X2 U13182 ( .B1(n15870), .B2(n12364), .A(n12262), .ZN(n14297) );
  INV_X1 U13183 ( .A(n14679), .ZN(n14528) );
  NAND3_X1 U13184 ( .A1(n10019), .A2(n10215), .A3(n10266), .ZN(n10018) );
  NAND3_X1 U13185 ( .A1(n10029), .A2(n10028), .A3(n10027), .ZN(P2_U2985) );
  OR2_X1 U13186 ( .A1(n16574), .A2(n16863), .ZN(n10028) );
  NOR2_X1 U13187 ( .A1(n12202), .A2(n12898), .ZN(n10032) );
  NOR2_X1 U13188 ( .A1(n12202), .A2(n10035), .ZN(n10034) );
  NAND2_X1 U13189 ( .A1(n15426), .A2(n10434), .ZN(n10042) );
  OAI21_X1 U13190 ( .B1(n15650), .B2(n20633), .A(n15431), .ZN(P1_U2971) );
  AND2_X1 U13191 ( .A1(n10040), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U13192 ( .A1(n15425), .A2(n9760), .ZN(n10043) );
  NAND2_X2 U13193 ( .A1(n10602), .A2(n10601), .ZN(n10634) );
  XNOR2_X2 U13194 ( .A(n10046), .B(n10636), .ZN(n10644) );
  INV_X1 U13195 ( .A(n10045), .ZN(n10044) );
  INV_X1 U13196 ( .A(n10635), .ZN(n10046) );
  NAND2_X1 U13197 ( .A1(n10262), .A2(n10048), .ZN(n10260) );
  INV_X1 U13198 ( .A(n11212), .ZN(n10050) );
  NAND2_X1 U13199 ( .A1(n10052), .A2(n10658), .ZN(n10156) );
  AOI21_X1 U13200 ( .B1(n17127), .B2(n10052), .A(n14645), .ZN(n14648) );
  OAI21_X1 U13201 ( .B1(n16922), .B2(n16846), .A(n16629), .ZN(P2_U2991) );
  INV_X1 U13202 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n10059) );
  NAND3_X1 U13203 ( .A1(n9603), .A2(P3_EAX_REG_11__SCAN_IN), .A3(
        P3_EAX_REG_10__SCAN_IN), .ZN(n10062) );
  AND2_X2 U13204 ( .A1(n17346), .A2(n14074), .ZN(n11562) );
  OR2_X1 U13205 ( .A1(n15737), .A2(n15862), .ZN(n10068) );
  AOI21_X1 U13206 ( .B1(n10432), .B2(n10074), .A(n15583), .ZN(n10072) );
  INV_X1 U13207 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10076) );
  AND2_X2 U13208 ( .A1(n10078), .A2(n11979), .ZN(n12050) );
  AND2_X2 U13209 ( .A1(n10078), .A2(n10107), .ZN(n12063) );
  AND2_X2 U13210 ( .A1(n10111), .A2(n10078), .ZN(n12045) );
  AND2_X1 U13211 ( .A1(n10081), .A2(n20878), .ZN(n10080) );
  NAND2_X1 U13212 ( .A1(n20854), .A2(n10190), .ZN(n15260) );
  NAND2_X1 U13213 ( .A1(n10232), .A2(n9585), .ZN(n10082) );
  NOR2_X1 U13214 ( .A1(n15261), .A2(n10190), .ZN(n13796) );
  INV_X1 U13215 ( .A(n19875), .ZN(n10096) );
  AOI21_X1 U13216 ( .B1(n16676), .B2(n16827), .A(n16675), .ZN(n10099) );
  NAND2_X1 U13217 ( .A1(n10102), .A2(n9721), .ZN(n10103) );
  OAI21_X1 U13218 ( .B1(n13089), .B2(n12969), .A(n10106), .ZN(n10105) );
  NAND2_X1 U13219 ( .A1(n11974), .A2(n10107), .ZN(n10379) );
  NAND2_X1 U13220 ( .A1(n10108), .A2(n10771), .ZN(n16829) );
  OAI21_X1 U13221 ( .B1(n16854), .B2(n16853), .A(n10108), .ZN(n17137) );
  AND2_X4 U13222 ( .A1(n10111), .A2(n14341), .ZN(n12702) );
  NAND2_X1 U13223 ( .A1(n10111), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14352) );
  AND2_X1 U13224 ( .A1(n10111), .A2(n14365), .ZN(n12264) );
  AND2_X2 U13225 ( .A1(n11974), .A2(n10111), .ZN(n12160) );
  INV_X1 U13226 ( .A(n15283), .ZN(n10112) );
  NAND2_X1 U13227 ( .A1(n15283), .A2(n9626), .ZN(n10113) );
  NAND2_X1 U13228 ( .A1(n9694), .A2(n10116), .ZN(n10271) );
  OR2_X1 U13229 ( .A1(n14960), .A2(n15328), .ZN(n10118) );
  NOR2_X2 U13230 ( .A1(n14977), .A2(n14978), .ZN(n14976) );
  AOI22_X1 U13231 ( .A1(n20046), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n19851), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U13232 ( .A1(n10124), .A2(n10122), .ZN(n15034) );
  AND2_X2 U13233 ( .A1(n15224), .A2(n10127), .ZN(n15184) );
  NAND3_X2 U13234 ( .A1(n10135), .A2(n10600), .A3(n10134), .ZN(n10623) );
  OAI21_X1 U13235 ( .B1(n10710), .B2(n10652), .A(n10147), .ZN(n10656) );
  INV_X1 U13236 ( .A(n14764), .ZN(n14770) );
  NAND2_X1 U13237 ( .A1(n14841), .A2(n9747), .ZN(n10148) );
  AND2_X4 U13238 ( .A1(n10150), .A2(n14541), .ZN(n13678) );
  NOR2_X1 U13239 ( .A1(n10150), .A2(n14556), .ZN(n14558) );
  AND2_X1 U13240 ( .A1(n13507), .A2(n10150), .ZN(n13541) );
  MUX2_X1 U13241 ( .A(n13292), .B(n13291), .S(n9594), .Z(n14761) );
  NAND3_X1 U13242 ( .A1(n9793), .A2(n10311), .A3(n10936), .ZN(n10829) );
  NAND2_X1 U13243 ( .A1(n14841), .A2(n9640), .ZN(n10157) );
  NAND2_X1 U13244 ( .A1(n10160), .A2(n9678), .ZN(n10719) );
  NAND2_X1 U13245 ( .A1(n20209), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10163) );
  OAI21_X1 U13246 ( .B1(n20209), .B2(n20326), .A(n20607), .ZN(n10165) );
  NAND2_X1 U13247 ( .A1(n10169), .A2(n14580), .ZN(n10168) );
  NAND2_X1 U13248 ( .A1(n16677), .A2(n10170), .ZN(P2_U2997) );
  OR2_X1 U13249 ( .A1(n16678), .A2(n16863), .ZN(n10170) );
  XNOR2_X2 U13250 ( .A(n10171), .B(n10633), .ZN(n10648) );
  INV_X1 U13251 ( .A(n10171), .ZN(n10407) );
  NAND2_X1 U13252 ( .A1(n10622), .A2(n10621), .ZN(n10171) );
  INV_X1 U13253 ( .A(n9594), .ZN(n10173) );
  OAI21_X1 U13254 ( .B1(n16700), .B2(n9633), .A(n10175), .ZN(n10174) );
  NOR2_X1 U13255 ( .A1(n16965), .A2(n10174), .ZN(n16968) );
  NAND2_X1 U13256 ( .A1(n12133), .A2(n10177), .ZN(n12134) );
  NAND2_X1 U13257 ( .A1(n20893), .A2(n10177), .ZN(n15283) );
  NAND2_X1 U13258 ( .A1(n15871), .A2(n15873), .ZN(n21087) );
  NAND4_X1 U13259 ( .A1(n10508), .A2(n10509), .A3(n10510), .A4(n10507), .ZN(
        n10180) );
  NAND4_X1 U13260 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10182) );
  AND2_X1 U13261 ( .A1(n10801), .A2(n10800), .ZN(n10184) );
  INV_X1 U13262 ( .A(n10807), .ZN(n10188) );
  INV_X2 U13263 ( .A(n12108), .ZN(n10191) );
  OAI21_X1 U13264 ( .B1(n10199), .B2(n10194), .A(n10669), .ZN(n10193) );
  NAND4_X1 U13265 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10194) );
  NAND4_X1 U13266 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10199) );
  OAI21_X1 U13267 ( .B1(n10210), .B2(n10205), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10204) );
  NAND4_X1 U13268 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10205) );
  NAND2_X1 U13269 ( .A1(n13678), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10209) );
  NAND4_X1 U13270 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10210) );
  NOR2_X2 U13271 ( .A1(n18522), .A2(n10218), .ZN(n18470) );
  NOR3_X1 U13272 ( .A1(n18149), .A2(n18049), .A3(n10225), .ZN(n18102) );
  INV_X1 U13273 ( .A(n18381), .ZN(n10227) );
  NAND2_X1 U13274 ( .A1(n10227), .A2(n9749), .ZN(n18368) );
  XNOR2_X1 U13275 ( .A(n10231), .B(n15607), .ZN(n15863) );
  NAND2_X1 U13276 ( .A1(n12232), .A2(n12134), .ZN(n14332) );
  NAND3_X1 U13277 ( .A1(n12232), .A2(n12134), .A3(n14376), .ZN(n10236) );
  NOR2_X1 U13278 ( .A1(n11909), .A2(n10237), .ZN(n14118) );
  INV_X1 U13279 ( .A(n10243), .ZN(n13807) );
  OR2_X1 U13280 ( .A1(n18809), .A2(n9743), .ZN(n10254) );
  NAND2_X1 U13281 ( .A1(n18809), .A2(n10253), .ZN(n10252) );
  NAND3_X1 U13282 ( .A1(n10256), .A2(n10255), .A3(n9691), .ZN(P2_U2998) );
  NAND2_X1 U13283 ( .A1(n19851), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10259) );
  AND4_X2 U13284 ( .A1(n10269), .A2(n11247), .A3(n10585), .A4(n10588), .ZN(
        n11495) );
  INV_X2 U13285 ( .A(n10578), .ZN(n14580) );
  INV_X1 U13286 ( .A(n14841), .ZN(n16775) );
  AND2_X4 U13287 ( .A1(n14841), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16754) );
  NAND2_X1 U13288 ( .A1(n16624), .A2(n10276), .ZN(n16922) );
  NAND2_X1 U13289 ( .A1(n13303), .A2(n13189), .ZN(n10281) );
  NOR2_X1 U13290 ( .A1(n13211), .A2(n10294), .ZN(n13215) );
  AOI21_X1 U13291 ( .B1(n15992), .B2(n10295), .A(n13243), .ZN(n15959) );
  NAND2_X1 U13292 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10297) );
  NAND3_X1 U13293 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U13294 ( .A1(n10299), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16818) );
  XNOR2_X1 U13295 ( .A(n10935), .B(n17110), .ZN(n16834) );
  NAND2_X1 U13296 ( .A1(n12928), .A2(n10465), .ZN(n14614) );
  NAND2_X1 U13297 ( .A1(n10307), .A2(n12210), .ZN(n12201) );
  XNOR2_X1 U13298 ( .A(n10307), .B(n12210), .ZN(n15864) );
  NAND2_X1 U13299 ( .A1(n10442), .A2(n9696), .ZN(n10310) );
  INV_X1 U13300 ( .A(n10939), .ZN(n10311) );
  NAND2_X1 U13301 ( .A1(n10311), .A2(n10936), .ZN(n10823) );
  NAND3_X1 U13302 ( .A1(n11587), .A2(n11588), .A3(n11589), .ZN(n10320) );
  CLKBUF_X1 U13303 ( .A(n18677), .Z(n10321) );
  NAND2_X2 U13304 ( .A1(n17478), .A2(n14064), .ZN(n18218) );
  OAI21_X1 U13305 ( .B1(n10329), .B2(n10330), .A(n10327), .ZN(n16593) );
  NAND2_X1 U13306 ( .A1(n10653), .A2(n10334), .ZN(n20290) );
  NAND2_X1 U13307 ( .A1(n14800), .A2(n9703), .ZN(n16299) );
  INV_X1 U13308 ( .A(n16299), .ZN(n11317) );
  NAND2_X2 U13309 ( .A1(n14841), .A2(n13163), .ZN(n16700) );
  NAND3_X1 U13310 ( .A1(n13170), .A2(n10338), .A3(n10335), .ZN(P2_U3029) );
  NAND2_X1 U13311 ( .A1(n14002), .A2(n10340), .ZN(n14040) );
  INV_X1 U13312 ( .A(n14040), .ZN(n11364) );
  NAND2_X1 U13313 ( .A1(n15973), .A2(n15972), .ZN(n15971) );
  INV_X1 U13314 ( .A(n15966), .ZN(n15967) );
  NAND2_X1 U13315 ( .A1(n9714), .A2(n10343), .ZN(n16131) );
  NAND3_X1 U13316 ( .A1(n11415), .A2(n16157), .A3(n10347), .ZN(n10346) );
  AOI21_X1 U13317 ( .B1(n16575), .B2(n10361), .A(n10359), .ZN(n11509) );
  OR2_X1 U13318 ( .A1(n11163), .A2(n10364), .ZN(n10363) );
  INV_X2 U13319 ( .A(n10502), .ZN(n13577) );
  NAND2_X2 U13320 ( .A1(n14540), .A2(n14550), .ZN(n10502) );
  NAND2_X1 U13321 ( .A1(n10963), .A2(n10365), .ZN(n10992) );
  INV_X1 U13322 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U13323 ( .A1(n10907), .A2(n10368), .ZN(n10985) );
  INV_X1 U13324 ( .A(n10908), .ZN(n10371) );
  NAND2_X1 U13325 ( .A1(n10968), .A2(n9739), .ZN(n11030) );
  NAND2_X1 U13326 ( .A1(n10968), .A2(n10470), .ZN(n10972) );
  NAND2_X1 U13327 ( .A1(n10990), .A2(n9709), .ZN(n10975) );
  INV_X1 U13328 ( .A(n12204), .ZN(n10382) );
  AOI21_X1 U13329 ( .B1(n12209), .B2(n12364), .A(n10385), .ZN(n10384) );
  AND2_X1 U13330 ( .A1(n15220), .A2(n9728), .ZN(n15132) );
  INV_X1 U13331 ( .A(n10395), .ZN(n14324) );
  NOR2_X1 U13332 ( .A1(n15975), .A2(n15974), .ZN(n15976) );
  INV_X1 U13333 ( .A(n10400), .ZN(n10403) );
  INV_X1 U13334 ( .A(n15958), .ZN(n10404) );
  NAND2_X1 U13335 ( .A1(n10407), .A2(n10406), .ZN(n14189) );
  NAND2_X1 U13336 ( .A1(n13151), .A2(n10408), .ZN(n16035) );
  NAND2_X1 U13337 ( .A1(n16754), .A2(n10414), .ZN(n10413) );
  NAND2_X1 U13338 ( .A1(n16754), .A2(n9758), .ZN(n17012) );
  NAND2_X1 U13339 ( .A1(n16754), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16755) );
  NAND2_X1 U13340 ( .A1(n10413), .A2(n16989), .ZN(n16701) );
  NAND2_X1 U13341 ( .A1(n10960), .A2(n10419), .ZN(n10423) );
  OAI21_X2 U13342 ( .B1(n10423), .B2(n10418), .A(n10417), .ZN(n16679) );
  AND2_X1 U13343 ( .A1(n10422), .A2(n16703), .ZN(n16690) );
  INV_X1 U13344 ( .A(n10433), .ZN(n15468) );
  NAND2_X1 U13345 ( .A1(n10447), .A2(n10445), .ZN(n10444) );
  NAND2_X1 U13346 ( .A1(n14841), .A2(n10448), .ZN(n14815) );
  AOI21_X2 U13347 ( .B1(n15583), .B2(n15661), .A(n15450), .ZN(n15425) );
  AND2_X1 U13348 ( .A1(n15975), .A2(n11144), .ZN(n11536) );
  INV_X1 U13349 ( .A(n11532), .ZN(n11533) );
  INV_X1 U13350 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11963) );
  NAND2_X1 U13351 ( .A1(n16428), .A2(n16429), .ZN(n16423) );
  AOI22_X1 U13352 ( .A1(n10636), .A2(n10635), .B1(n10640), .B2(n10619), .ZN(
        n10618) );
  AND2_X1 U13353 ( .A1(n10600), .A2(n10599), .ZN(n10601) );
  INV_X1 U13354 ( .A(n20290), .ZN(n10803) );
  NAND2_X1 U13355 ( .A1(n10629), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10582) );
  AOI22_X1 U13356 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10539) );
  OAI22_X2 U13357 ( .A1(n18770), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n18713), .B2(n11708), .ZN(n18766) );
  INV_X1 U13358 ( .A(n13371), .ZN(n13360) );
  OR2_X1 U13359 ( .A1(n11535), .A2(n16846), .ZN(n10449) );
  INV_X1 U13360 ( .A(n16846), .ZN(n13307) );
  OR2_X1 U13361 ( .A1(n13346), .A2(n13345), .ZN(P3_U2640) );
  OR2_X1 U13362 ( .A1(n14922), .A2(n20837), .ZN(n10451) );
  AND4_X1 U13363 ( .A1(n12467), .A2(n15136), .A3(n15179), .A4(n12466), .ZN(
        n10452) );
  INV_X1 U13364 ( .A(n12769), .ZN(n12713) );
  INV_X1 U13365 ( .A(n11346), .ZN(n13485) );
  INV_X1 U13366 ( .A(n13610), .ZN(n13593) );
  AND2_X1 U13367 ( .A1(n14427), .A2(n14426), .ZN(n10453) );
  INV_X1 U13368 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18371) );
  AND2_X1 U13369 ( .A1(n14839), .A2(n14838), .ZN(n10454) );
  AND2_X1 U13370 ( .A1(n16681), .A2(n16688), .ZN(n10455) );
  AND2_X1 U13371 ( .A1(n10715), .A2(n10714), .ZN(n10456) );
  AND2_X1 U13372 ( .A1(n18805), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10457) );
  AND2_X1 U13373 ( .A1(n15413), .A2(n12036), .ZN(n10458) );
  NAND2_X2 U13374 ( .A1(n15413), .A2(n14127), .ZN(n15415) );
  NOR2_X1 U13375 ( .A1(n17539), .A2(n14617), .ZN(n10459) );
  AND2_X1 U13376 ( .A1(n11205), .A2(n13719), .ZN(n10460) );
  OR2_X1 U13377 ( .A1(n11513), .A2(n13739), .ZN(n10461) );
  AND2_X1 U13378 ( .A1(n18997), .A2(n19035), .ZN(n10462) );
  OR2_X1 U13379 ( .A1(n10217), .A2(n18578), .ZN(n10463) );
  OR2_X1 U13380 ( .A1(n10631), .A2(n20591), .ZN(n10464) );
  OR2_X1 U13381 ( .A1(n17509), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10465) );
  INV_X1 U13382 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n11859) );
  INV_X1 U13383 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n14376) );
  OR2_X1 U13384 ( .A1(n13671), .A2(n13670), .ZN(n10466) );
  NAND2_X1 U13385 ( .A1(n12219), .A2(n12218), .ZN(n10467) );
  AND2_X1 U13386 ( .A1(n10316), .A2(n17309), .ZN(n10468) );
  OR2_X1 U13387 ( .A1(n18712), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10469) );
  INV_X1 U13388 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11720) );
  INV_X1 U13389 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19660) );
  INV_X1 U13390 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16164) );
  INV_X1 U13391 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16225) );
  INV_X1 U13392 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10964) );
  INV_X1 U13393 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19165) );
  INV_X1 U13394 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11721) );
  INV_X1 U13395 ( .A(n11299), .ZN(n11432) );
  INV_X1 U13396 ( .A(n15098), .ZN(n15070) );
  INV_X1 U13397 ( .A(n17283), .ZN(n11724) );
  OR2_X1 U13398 ( .A1(n10902), .A2(n10967), .ZN(n10470) );
  NAND2_X1 U13399 ( .A1(n9583), .A2(n12899), .ZN(n10471) );
  NOR2_X1 U13400 ( .A1(n21240), .A2(n21205), .ZN(n10472) );
  NOR2_X1 U13401 ( .A1(n15978), .A2(n11513), .ZN(n16577) );
  OR2_X1 U13402 ( .A1(n10902), .A2(n16038), .ZN(n10473) );
  INV_X1 U13403 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11865) );
  INV_X1 U13404 ( .A(n13351), .ZN(n14044) );
  OAI21_X1 U13405 ( .B1(n13350), .B2(n13371), .A(n13349), .ZN(n13351) );
  INV_X1 U13406 ( .A(n18025), .ZN(n19631) );
  NOR2_X1 U13407 ( .A1(n18536), .A2(n19633), .ZN(n18025) );
  INV_X1 U13408 ( .A(n17708), .ZN(n13329) );
  AND2_X1 U13409 ( .A1(n10540), .A2(n10539), .ZN(n10474) );
  AND3_X1 U13410 ( .A1(n10536), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10535), .ZN(n10475) );
  AND2_X1 U13411 ( .A1(n13217), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10476) );
  NOR2_X1 U13412 ( .A1(n21240), .A2(n21048), .ZN(n10477) );
  INV_X1 U13413 ( .A(n14493), .ZN(n14500) );
  NAND2_X1 U13414 ( .A1(n12850), .A2(n13767), .ZN(n15400) );
  INV_X2 U13415 ( .A(n15400), .ZN(n15413) );
  INV_X1 U13416 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20607) );
  NAND2_X1 U13417 ( .A1(n21384), .A2(n15884), .ZN(n10478) );
  AND2_X1 U13418 ( .A1(n13180), .A2(n21373), .ZN(n20666) );
  OR2_X1 U13419 ( .A1(n18015), .A2(n14734), .ZN(n10479) );
  XNOR2_X1 U13420 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13294), .ZN(
        n10480) );
  AND2_X1 U13421 ( .A1(n11462), .A2(n13293), .ZN(n10481) );
  OR2_X1 U13422 ( .A1(n13280), .A2(n13278), .ZN(n10482) );
  OR2_X1 U13423 ( .A1(n11411), .A2(n11410), .ZN(n14436) );
  INV_X2 U13424 ( .A(n19171), .ZN(n11836) );
  INV_X1 U13425 ( .A(n11141), .ZN(n11142) );
  AND2_X1 U13426 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10483) );
  NOR2_X1 U13427 ( .A1(n18651), .A2(n10468), .ZN(n10484) );
  AND2_X1 U13428 ( .A1(n13652), .A2(n16378), .ZN(n10485) );
  AND2_X1 U13429 ( .A1(n11999), .A2(n11998), .ZN(n10486) );
  AND4_X1 U13430 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n10487) );
  OAI211_X1 U13431 ( .C1(n12815), .C2(n12173), .A(n12174), .B(n12172), .ZN(
        n12217) );
  INV_X1 U13432 ( .A(n12217), .ZN(n12218) );
  INV_X2 U13433 ( .A(n12111), .ZN(n12094) );
  AND3_X1 U13434 ( .A1(n12776), .A2(n12775), .A3(n12784), .ZN(n12789) );
  AOI22_X1 U13435 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13528), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10723) );
  INV_X1 U13436 ( .A(n10889), .ZN(n10860) );
  OAI21_X1 U13437 ( .B1(n13092), .B2(n12096), .A(n12189), .ZN(n12097) );
  INV_X1 U13438 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11969) );
  OR2_X1 U13439 ( .A1(n12294), .A2(n12293), .ZN(n12917) );
  AND3_X1 U13440 ( .A1(n12118), .A2(n12117), .A3(n12116), .ZN(n12119) );
  NAND2_X1 U13441 ( .A1(n12808), .A2(n12807), .ZN(n12814) );
  NAND2_X1 U13442 ( .A1(n13719), .A2(n19869), .ZN(n10587) );
  OR2_X1 U13443 ( .A1(n11837), .A2(n11847), .ZN(n11839) );
  INV_X1 U13444 ( .A(n12391), .ZN(n12392) );
  AND2_X1 U13445 ( .A1(n12276), .A2(n12275), .ZN(n12898) );
  OR2_X1 U13446 ( .A1(n12199), .A2(n12198), .ZN(n12200) );
  NAND2_X1 U13447 ( .A1(n12969), .A2(n12932), .ZN(n12174) );
  OR2_X1 U13448 ( .A1(n12316), .A2(n12315), .ZN(n12916) );
  AND2_X1 U13449 ( .A1(n12215), .A2(n12176), .ZN(n12177) );
  INV_X1 U13450 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10962) );
  INV_X1 U13451 ( .A(n10880), .ZN(n11308) );
  AND2_X1 U13452 ( .A1(n12392), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12446) );
  AND2_X1 U13453 ( .A1(n12318), .A2(n12317), .ZN(n12319) );
  OR2_X1 U13454 ( .A1(n12188), .A2(n12187), .ZN(n12872) );
  AOI22_X1 U13455 ( .A1(n17515), .A2(n12925), .B1(n17505), .B2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U13456 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9554), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11992) );
  AND3_X1 U13457 ( .A1(n12192), .A2(n12191), .A3(n12190), .ZN(n12197) );
  NAND2_X1 U13458 ( .A1(n9590), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10904) );
  AND2_X1 U13459 ( .A1(n17496), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10881) );
  AND2_X2 U13460 ( .A1(n11288), .A2(n11273), .ZN(n11297) );
  INV_X1 U13461 ( .A(n14190), .ZN(n11053) );
  AND2_X1 U13462 ( .A1(n11479), .A2(n14887), .ZN(n11480) );
  INV_X1 U13463 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11856) );
  NAND2_X1 U13464 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17177) );
  NAND2_X1 U13465 ( .A1(n11678), .A2(n11677), .ZN(n11699) );
  INV_X1 U13466 ( .A(n15024), .ZN(n12619) );
  NAND2_X1 U13467 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12048) );
  NAND2_X1 U13468 ( .A1(n12735), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12737) );
  INV_X1 U13469 ( .A(n14131), .ZN(n12229) );
  NAND2_X1 U13470 ( .A1(n10905), .A2(n10904), .ZN(n10911) );
  OR2_X1 U13471 ( .A1(n16408), .A2(n13574), .ZN(n13575) );
  AND2_X1 U13472 ( .A1(n11491), .A2(n11490), .ZN(n11517) );
  AND2_X1 U13473 ( .A1(n13152), .A2(n13150), .ZN(n11103) );
  INV_X1 U13474 ( .A(n14252), .ZN(n11415) );
  INV_X1 U13475 ( .A(n14079), .ZN(n11363) );
  INV_X1 U13476 ( .A(n16298), .ZN(n11316) );
  INV_X1 U13477 ( .A(n10873), .ZN(n11296) );
  NAND2_X1 U13478 ( .A1(n11856), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n21538) );
  OAI21_X1 U13479 ( .B1(n11286), .B2(n11285), .A(n11284), .ZN(n11290) );
  NAND2_X1 U13480 ( .A1(n14044), .A2(n13353), .ZN(n13358) );
  XNOR2_X1 U13481 ( .A(n13379), .B(n13377), .ZN(n14198) );
  INV_X1 U13482 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11853) );
  INV_X1 U13483 ( .A(n17177), .ZN(n13311) );
  NAND2_X1 U13484 ( .A1(n18843), .A2(n11703), .ZN(n11704) );
  AND2_X1 U13485 ( .A1(n11914), .A2(n11895), .ZN(n11916) );
  INV_X1 U13486 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18207) );
  NAND2_X1 U13487 ( .A1(n12237), .A2(n12236), .ZN(n20995) );
  AND2_X1 U13488 ( .A1(n13065), .A2(n13064), .ZN(n15033) );
  OR2_X1 U13489 ( .A1(n15052), .A2(n15053), .ZN(n15039) );
  INV_X1 U13490 ( .A(n12713), .ZN(n12451) );
  OR2_X1 U13491 ( .A1(n14304), .A2(n14339), .ZN(n14305) );
  OR2_X1 U13492 ( .A1(n12737), .A2(n12736), .ZN(n13182) );
  NAND2_X1 U13493 ( .A1(n12620), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12640) );
  AND2_X1 U13494 ( .A1(n12380), .A2(n12379), .ZN(n15203) );
  OR2_X1 U13495 ( .A1(n15583), .A2(n15842), .ZN(n15512) );
  OR2_X1 U13496 ( .A1(n13114), .A2(n13113), .ZN(n14344) );
  INV_X1 U13497 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14342) );
  AND2_X1 U13498 ( .A1(n12235), .A2(n21368), .ZN(n20845) );
  INV_X1 U13499 ( .A(n21293), .ZN(n21370) );
  INV_X1 U13500 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21120) );
  INV_X1 U13501 ( .A(n13229), .ZN(n13227) );
  NAND2_X1 U13502 ( .A1(n10868), .A2(n10867), .ZN(n20598) );
  AND2_X1 U13503 ( .A1(n11057), .A2(n11056), .ZN(n14238) );
  OR2_X1 U13504 ( .A1(n13611), .A2(n16389), .ZN(n13629) );
  AND2_X1 U13505 ( .A1(n13563), .A2(n13562), .ZN(n13571) );
  AND2_X1 U13506 ( .A1(n17078), .A2(n11265), .ZN(n17031) );
  INV_X1 U13507 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14550) );
  INV_X1 U13508 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14559) );
  AND2_X1 U13509 ( .A1(n19904), .A2(n19903), .ZN(n19908) );
  NAND2_X1 U13510 ( .A1(n11943), .A2(n11942), .ZN(n11950) );
  NAND2_X1 U13511 ( .A1(n13340), .A2(n10479), .ZN(n13341) );
  AOI22_X1 U13512 ( .A1(n11684), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11628), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11591) );
  INV_X1 U13513 ( .A(n14877), .ZN(n11723) );
  INV_X1 U13514 ( .A(n19024), .ZN(n19032) );
  INV_X1 U13515 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17346) );
  AND2_X1 U13516 ( .A1(n14926), .A2(n14376), .ZN(n13180) );
  OR2_X1 U13517 ( .A1(n15287), .A2(n15246), .ZN(n20700) );
  INV_X1 U13518 ( .A(n15205), .ZN(n13014) );
  NOR2_X1 U13519 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12769) );
  OR2_X1 U13520 ( .A1(n12861), .A2(n20836), .ZN(n15387) );
  OAI21_X1 U13521 ( .B1(n14013), .B2(n14010), .A(n12849), .ZN(n12850) );
  AOI21_X1 U13522 ( .B1(n15533), .B2(n14906), .A(n13754), .ZN(n13755) );
  NAND2_X1 U13523 ( .A1(n12549), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12552) );
  OR2_X1 U13524 ( .A1(n12483), .A2(n12482), .ZN(n12568) );
  NAND2_X1 U13525 ( .A1(n14133), .A2(n14132), .ZN(n14131) );
  OR2_X1 U13526 ( .A1(n15583), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12947) );
  INV_X1 U13527 ( .A(n20666), .ZN(n20771) );
  NOR2_X1 U13528 ( .A1(n13946), .A2(n12094), .ZN(n14925) );
  INV_X1 U13529 ( .A(n14013), .ZN(n14374) );
  AND2_X1 U13530 ( .A1(n20962), .A2(n20988), .ZN(n20966) );
  NOR2_X1 U13531 ( .A1(n21239), .A2(n21000), .ZN(n21182) );
  INV_X1 U13532 ( .A(n21389), .ZN(n21254) );
  INV_X1 U13533 ( .A(n12880), .ZN(n20840) );
  INV_X1 U13534 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21373) );
  INV_X1 U13535 ( .A(n16340), .ZN(n16359) );
  NAND2_X1 U13536 ( .A1(n11141), .A2(n11140), .ZN(n15975) );
  INV_X1 U13537 ( .A(n16357), .ZN(n16335) );
  AND2_X1 U13538 ( .A1(n11102), .A2(n11101), .ZN(n14608) );
  OR2_X1 U13539 ( .A1(n13629), .A2(n13631), .ZN(n16377) );
  INV_X1 U13540 ( .A(n16407), .ZN(n16408) );
  AND2_X1 U13541 ( .A1(n19795), .A2(n13720), .ZN(n16543) );
  NAND2_X1 U13542 ( .A1(n13288), .A2(n13287), .ZN(n13289) );
  AOI21_X1 U13543 ( .B1(n11536), .B2(n16827), .A(n11153), .ZN(n11154) );
  AND2_X1 U13544 ( .A1(n11098), .A2(n11097), .ZN(n14657) );
  NAND2_X1 U13545 ( .A1(n13828), .A2(n11147), .ZN(n16839) );
  INV_X1 U13546 ( .A(n16973), .ZN(n13166) );
  AND3_X1 U13547 ( .A1(n11381), .A2(n11380), .A3(n11379), .ZN(n14165) );
  AND3_X1 U13548 ( .A1(n11321), .A2(n11320), .A3(n11319), .ZN(n16274) );
  AND2_X1 U13549 ( .A1(n20608), .A2(n20606), .ZN(n16837) );
  NAND2_X1 U13550 ( .A1(n14005), .A2(n14004), .ZN(n14006) );
  NAND2_X1 U13551 ( .A1(n11199), .A2(n11198), .ZN(n14570) );
  INV_X1 U13552 ( .A(n19912), .ZN(n19934) );
  OR2_X1 U13553 ( .A1(n20245), .A2(n20241), .ZN(n20284) );
  NOR2_X1 U13554 ( .A1(n20177), .A2(n20615), .ZN(n20331) );
  INV_X1 U13555 ( .A(n19893), .ZN(n19889) );
  AND2_X1 U13556 ( .A1(n19584), .A2(n19593), .ZN(n14276) );
  NOR2_X1 U13557 ( .A1(n13342), .A2(n13341), .ZN(n13343) );
  NOR2_X1 U13558 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17800), .ZN(n17787) );
  NOR2_X1 U13559 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17897), .ZN(n17882) );
  NAND2_X1 U13560 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .ZN(n14712) );
  OR2_X1 U13561 ( .A1(n18713), .A2(n17315), .ZN(n17287) );
  INV_X1 U13562 ( .A(n19736), .ZN(n18578) );
  INV_X1 U13563 ( .A(n11957), .ZN(n17160) );
  NOR2_X1 U13564 ( .A1(n19121), .A2(n18947), .ZN(n19000) );
  AND2_X1 U13565 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19032), .ZN(
        n19010) );
  AND2_X1 U13566 ( .A1(n11894), .A2(n11893), .ZN(n19584) );
  AND4_X1 U13567 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n11832) );
  INV_X1 U13568 ( .A(n19641), .ZN(n19735) );
  AND2_X1 U13569 ( .A1(n13796), .A2(n13795), .ZN(n20681) );
  AND2_X1 U13570 ( .A1(n15270), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13789) );
  INV_X1 U13571 ( .A(n9573), .ZN(n14934) );
  AND2_X1 U13572 ( .A1(n15413), .A2(n14128), .ZN(n15401) );
  INV_X2 U13573 ( .A(n14498), .ZN(n20768) );
  NAND2_X1 U13574 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n12331), .ZN(
        n12359) );
  NAND2_X1 U13575 ( .A1(n20633), .A2(n13181), .ZN(n15530) );
  OR2_X1 U13576 ( .A1(n14013), .A2(n15940), .ZN(n14304) );
  NOR2_X1 U13577 ( .A1(n15758), .A2(n13132), .ZN(n15698) );
  NOR2_X1 U13578 ( .A1(n13129), .A2(n20819), .ZN(n14628) );
  OR2_X1 U13579 ( .A1(n14628), .A2(n20811), .ZN(n17545) );
  AND2_X1 U13580 ( .A1(n13115), .A2(n13944), .ZN(n20811) );
  NAND2_X1 U13581 ( .A1(n14374), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15931) );
  OAI22_X1 U13582 ( .A1(n20851), .A2(n20850), .B1(n21123), .B2(n20997), .ZN(
        n20889) );
  INV_X1 U13583 ( .A(n20954), .ZN(n20921) );
  OAI22_X1 U13584 ( .A1(n20927), .A2(n20926), .B1(n21123), .B2(n21056), .ZN(
        n20950) );
  OAI211_X1 U13585 ( .C1(n20927), .C2(n20925), .A(n21182), .B(n20924), .ZN(
        n20951) );
  OAI21_X1 U13586 ( .B1(n10477), .B2(n21001), .A(n21336), .ZN(n21018) );
  NAND2_X1 U13587 ( .A1(n15870), .A2(n15867), .ZN(n20958) );
  OAI22_X1 U13588 ( .A1(n21058), .A2(n21057), .B1(n21331), .B2(n21056), .ZN(
        n21081) );
  INV_X1 U13589 ( .A(n21234), .ZN(n21118) );
  NOR2_X2 U13590 ( .A1(n21211), .A2(n21301), .ZN(n21198) );
  NOR2_X2 U13591 ( .A1(n21211), .A2(n21328), .ZN(n21230) );
  INV_X1 U13592 ( .A(n21250), .ZN(n21287) );
  NAND2_X1 U13593 ( .A1(n14376), .A2(n14375), .ZN(n21000) );
  OAI21_X1 U13594 ( .B1(n21300), .B2(n21299), .A(n21380), .ZN(n21324) );
  NOR2_X2 U13595 ( .A1(n21379), .A2(n21301), .ZN(n21363) );
  INV_X1 U13596 ( .A(n21253), .ZN(n21376) );
  AND2_X1 U13597 ( .A1(n12107), .A2(n20884), .ZN(n21401) );
  INV_X1 U13598 ( .A(n21278), .ZN(n21416) );
  NAND2_X1 U13599 ( .A1(n9599), .A2(n12880), .ZN(n21328) );
  INV_X1 U13600 ( .A(n17555), .ZN(n14378) );
  INV_X1 U13601 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21442) );
  INV_X1 U13602 ( .A(n21500), .ZN(n21501) );
  AND2_X1 U13603 ( .A1(n13823), .A2(n13272), .ZN(n16357) );
  OR2_X1 U13604 ( .A1(n11378), .A2(n11377), .ZN(n14410) );
  OR2_X1 U13605 ( .A1(n14571), .A2(n14570), .ZN(n14218) );
  INV_X1 U13606 ( .A(n13693), .ZN(n13694) );
  OR3_X1 U13607 ( .A1(n13428), .A2(n13427), .A3(n13426), .ZN(n14687) );
  INV_X1 U13608 ( .A(n19803), .ZN(n19793) );
  INV_X1 U13609 ( .A(n13929), .ZN(n13905) );
  NAND2_X1 U13610 ( .A1(n13252), .A2(n13253), .ZN(n13831) );
  INV_X1 U13611 ( .A(n17018), .ZN(n16735) );
  INV_X1 U13612 ( .A(n16863), .ZN(n16836) );
  NOR2_X1 U13613 ( .A1(n11220), .A2(n10898), .ZN(n11146) );
  NAND2_X1 U13614 ( .A1(n16649), .A2(n16662), .ZN(n16653) );
  NAND2_X1 U13615 ( .A1(n13166), .A2(n13165), .ZN(n13167) );
  AND2_X1 U13616 ( .A1(n11505), .A2(n11498), .ZN(n17121) );
  INV_X1 U13617 ( .A(n17121), .ZN(n17134) );
  OAI211_X1 U13618 ( .C1(n19912), .C2(n20607), .A(n19911), .B(n20419), .ZN(
        n19937) );
  INV_X1 U13619 ( .A(n19945), .ZN(n19966) );
  OAI21_X1 U13620 ( .B1(n19981), .B2(n19980), .A(n19979), .ZN(n20005) );
  OAI21_X1 U13621 ( .B1(n20049), .B2(n20048), .A(n20047), .ZN(n20072) );
  INV_X1 U13622 ( .A(n20087), .ZN(n20104) );
  INV_X1 U13623 ( .A(n20176), .ZN(n20131) );
  NAND2_X1 U13624 ( .A1(n20148), .A2(n20147), .ZN(n20172) );
  OR2_X1 U13625 ( .A1(n20567), .A2(n21692), .ZN(n20115) );
  INV_X1 U13626 ( .A(n20562), .ZN(n20250) );
  INV_X1 U13627 ( .A(n20329), .ZN(n20365) );
  NOR2_X2 U13628 ( .A1(n20335), .A2(n20334), .ZN(n20397) );
  INV_X1 U13629 ( .A(n20264), .ZN(n20438) );
  AND2_X1 U13630 ( .A1(n19886), .A2(n20419), .ZN(n20458) );
  INV_X1 U13631 ( .A(n16345), .ZN(n16292) );
  INV_X1 U13632 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20493) );
  AND2_X1 U13633 ( .A1(n11881), .A2(n11884), .ZN(n19589) );
  NAND2_X1 U13634 ( .A1(n13344), .A2(n13343), .ZN(n13345) );
  NOR2_X1 U13635 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17759), .ZN(n17728) );
  NOR2_X1 U13636 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17826), .ZN(n17812) );
  NOR2_X1 U13637 ( .A1(n19681), .A2(n17819), .ZN(n17794) );
  NAND2_X1 U13638 ( .A1(n17861), .A2(n17857), .ZN(n17854) );
  NOR2_X1 U13639 ( .A1(n19670), .A2(n17892), .ZN(n17885) );
  INV_X1 U13640 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17979) );
  NOR2_X2 U13641 ( .A1(n19754), .A2(n19615), .ZN(n18034) );
  INV_X1 U13642 ( .A(n17983), .ZN(n18042) );
  NOR2_X1 U13643 ( .A1(n19171), .A2(n18471), .ZN(n18465) );
  OR2_X1 U13644 ( .A1(n11694), .A2(n11693), .ZN(n17282) );
  INV_X1 U13645 ( .A(n18801), .ZN(n18737) );
  NOR2_X1 U13646 ( .A1(n18576), .A2(n18537), .ZN(n18565) );
  OAI21_X1 U13647 ( .B1(n18578), .B2(n19617), .A(n18577), .ZN(n18622) );
  AND2_X1 U13648 ( .A1(n18578), .A2(n18577), .ZN(n18617) );
  NOR2_X2 U13649 ( .A1(n18860), .A2(n18536), .ZN(n18824) );
  AND2_X1 U13650 ( .A1(n14728), .A2(n17282), .ZN(n18846) );
  NOR2_X1 U13651 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19138), .ZN(n19384) );
  INV_X1 U13652 ( .A(n19114), .ZN(n19008) );
  INV_X1 U13653 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19088) );
  AND2_X1 U13654 ( .A1(n19053), .A2(n19584), .ZN(n17301) );
  NOR3_X1 U13655 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n17653), .ZN(n19291) );
  NOR2_X1 U13656 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19723), .ZN(
        n19612) );
  INV_X1 U13657 ( .A(n19216), .ZN(n19241) );
  INV_X1 U13658 ( .A(n19259), .ZN(n19263) );
  INV_X1 U13659 ( .A(n19306), .ZN(n19332) );
  INV_X1 U13660 ( .A(n19344), .ZN(n19355) );
  INV_X1 U13661 ( .A(n19397), .ZN(n19401) );
  INV_X1 U13662 ( .A(n19413), .ZN(n19423) );
  INV_X1 U13663 ( .A(n19443), .ZN(n19447) );
  INV_X1 U13664 ( .A(n19551), .ZN(n19495) );
  INV_X1 U13665 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19638) );
  INV_X1 U13666 ( .A(n19839), .ZN(n19837) );
  INV_X1 U13667 ( .A(U212), .ZN(n17600) );
  NAND2_X1 U13668 ( .A1(n14448), .A2(n13866), .ZN(n21521) );
  INV_X1 U13669 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21050) );
  AOI21_X1 U13670 ( .B1(n15627), .B2(n20693), .A(n14947), .ZN(n14948) );
  AND2_X1 U13671 ( .A1(n15242), .A2(n15114), .ZN(n15217) );
  NAND2_X1 U13672 ( .A1(n13771), .A2(n13789), .ZN(n15255) );
  AND2_X1 U13673 ( .A1(n15255), .A2(n15254), .ZN(n20672) );
  AND2_X2 U13674 ( .A1(n13144), .A2(n13767), .ZN(n20712) );
  INV_X1 U13675 ( .A(n15401), .ZN(n15412) );
  INV_X1 U13676 ( .A(n20736), .ZN(n20732) );
  NOR2_X1 U13677 ( .A1(n14448), .A2(n14447), .ZN(n14498) );
  OR2_X1 U13678 ( .A1(n13137), .A2(n13136), .ZN(n13138) );
  NAND2_X1 U13679 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15823), .ZN(
        n20819) );
  OAI21_X1 U13680 ( .B1(n14377), .B2(n17560), .A(n21000), .ZN(n20834) );
  OR2_X1 U13681 ( .A1(n20958), .A2(n21234), .ZN(n20913) );
  OR2_X1 U13682 ( .A1(n20958), .A2(n21301), .ZN(n20954) );
  OR2_X1 U13683 ( .A1(n20958), .A2(n21328), .ZN(n20994) );
  OR2_X1 U13684 ( .A1(n20958), .A2(n21086), .ZN(n21021) );
  OR2_X1 U13685 ( .A1(n21087), .A2(n21234), .ZN(n21047) );
  OR2_X1 U13686 ( .A1(n21087), .A2(n21301), .ZN(n21085) );
  OR2_X1 U13687 ( .A1(n21087), .A2(n21086), .ZN(n21107) );
  OR2_X1 U13688 ( .A1(n21087), .A2(n21328), .ZN(n21117) );
  NAND2_X1 U13689 ( .A1(n21204), .A2(n21118), .ZN(n21171) );
  AOI22_X1 U13690 ( .A1(n21178), .A2(n21175), .B1(n21174), .B2(n21330), .ZN(
        n21202) );
  NAND2_X1 U13691 ( .A1(n21204), .A2(n21203), .ZN(n21250) );
  AOI22_X1 U13692 ( .A1(n21246), .A2(n21243), .B1(n21239), .B2(n21238), .ZN(
        n21292) );
  OR2_X1 U13693 ( .A1(n21379), .A2(n21234), .ZN(n21327) );
  OR2_X1 U13694 ( .A1(n21379), .A2(n21086), .ZN(n21413) );
  OR2_X1 U13695 ( .A1(n21379), .A2(n21328), .ZN(n21436) );
  NAND2_X1 U13696 ( .A1(n15884), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15945) );
  INV_X1 U13697 ( .A(n21510), .ZN(n21507) );
  INV_X1 U13698 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20628) );
  OR2_X1 U13699 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20628), .ZN(n21532) );
  INV_X1 U13700 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20615) );
  AOI211_X1 U13701 ( .C1(n14761), .C2(n16357), .A(n14760), .B(n14759), .ZN(
        n14763) );
  INV_X1 U13702 ( .A(n11536), .ZN(n16394) );
  OR2_X1 U13703 ( .A1(n16105), .A2(n16104), .ZN(n16948) );
  NAND2_X1 U13704 ( .A1(n13823), .A2(n13264), .ZN(n16304) );
  INV_X1 U13705 ( .A(n16342), .ZN(n16353) );
  OR2_X1 U13706 ( .A1(n14672), .A2(n14671), .ZN(n16963) );
  AOI21_X2 U13707 ( .B1(n14218), .B2(n14203), .A(n14226), .ZN(n16430) );
  INV_X1 U13708 ( .A(n20585), .ZN(n20009) );
  NAND2_X1 U13709 ( .A1(n19795), .A2(n13705), .ZN(n16562) );
  AND2_X1 U13710 ( .A1(n16459), .A2(n16562), .ZN(n16565) );
  AND2_X1 U13711 ( .A1(n13987), .A2(n13986), .ZN(n19803) );
  NAND2_X1 U13712 ( .A1(n19826), .A2(n13930), .ZN(n13980) );
  OR2_X1 U13713 ( .A1(n19833), .A2(n19826), .ZN(n19828) );
  INV_X1 U13714 ( .A(n19826), .ZN(n19836) );
  OR2_X1 U13715 ( .A1(n13831), .A2(n13830), .ZN(n13836) );
  NAND2_X1 U13716 ( .A1(n11146), .A2(n9593), .ZN(n16846) );
  XNOR2_X1 U13717 ( .A(n16653), .B(n16652), .ZN(n16946) );
  NAND2_X1 U13718 ( .A1(n11505), .A2(n20595), .ZN(n17124) );
  INV_X1 U13719 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20591) );
  INV_X1 U13720 ( .A(n17497), .ZN(n17156) );
  NAND2_X1 U13721 ( .A1(n20136), .A2(n20077), .ZN(n19940) );
  OR2_X1 U13722 ( .A1(n20010), .A2(n20562), .ZN(n20003) );
  OR2_X1 U13723 ( .A1(n20115), .A2(n20334), .ZN(n20087) );
  OR2_X1 U13724 ( .A1(n20010), .A2(n20334), .ZN(n20076) );
  NAND2_X1 U13725 ( .A1(n20361), .A2(n20077), .ZN(n20135) );
  OR2_X1 U13726 ( .A1(n20115), .A2(n20414), .ZN(n20176) );
  NAND2_X1 U13727 ( .A1(n20362), .A2(n20136), .ZN(n20208) );
  NAND2_X1 U13728 ( .A1(n20251), .A2(n20250), .ZN(n20295) );
  INV_X1 U13729 ( .A(n20427), .ZN(n20341) );
  INV_X1 U13730 ( .A(n20459), .ZN(n20354) );
  INV_X1 U13731 ( .A(n20433), .ZN(n20381) );
  INV_X1 U13732 ( .A(n20309), .ZN(n20448) );
  NAND2_X1 U13733 ( .A1(n20362), .A2(n20361), .ZN(n20455) );
  INV_X1 U13734 ( .A(n20560), .ZN(n20474) );
  INV_X1 U13735 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n17653) );
  INV_X1 U13736 ( .A(n19089), .ZN(n19120) );
  NAND2_X1 U13737 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18042), .ZN(n18015) );
  NAND2_X1 U13738 ( .A1(n18096), .A2(P3_EBX_REG_28__SCAN_IN), .ZN(n18093) );
  AND3_X1 U13739 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(n18465), .ZN(n18463) );
  INV_X1 U13740 ( .A(n17282), .ZN(n18515) );
  INV_X1 U13741 ( .A(n11896), .ZN(n18524) );
  AND2_X1 U13742 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n14515), .ZN(n14518) );
  OR2_X1 U13743 ( .A1(n18536), .A2(n18737), .ZN(n19744) );
  INV_X1 U13744 ( .A(n18622), .ZN(n18619) );
  INV_X1 U13745 ( .A(n18846), .ZN(n18829) );
  NAND2_X1 U13746 ( .A1(n19384), .A2(n19291), .ZN(n19479) );
  OR2_X1 U13747 ( .A1(n18945), .A2(n18948), .ZN(n18969) );
  NAND2_X1 U13748 ( .A1(n19753), .A2(n19740), .ZN(n19055) );
  INV_X1 U13749 ( .A(n19099), .ZN(n19058) );
  OR2_X1 U13750 ( .A1(n19053), .A2(n19089), .ZN(n19114) );
  INV_X1 U13751 ( .A(n17489), .ZN(n14076) );
  INV_X1 U13752 ( .A(n19528), .ZN(n19464) );
  INV_X1 U13753 ( .A(n19482), .ZN(n19519) );
  INV_X1 U13754 ( .A(n19187), .ZN(n19537) );
  INV_X1 U13755 ( .A(n19743), .ZN(n19623) );
  INV_X1 U13756 ( .A(n19720), .ZN(n19717) );
  INV_X1 U13757 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19656) );
  AND2_X2 U13758 ( .A1(n12860), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20838)
         );
  INV_X1 U13759 ( .A(n17605), .ZN(n17603) );
  INV_X1 U13760 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20499) );
  NAND2_X1 U13761 ( .A1(n10451), .A2(n13756), .ZN(P1_U2973) );
  OAI211_X1 U13762 ( .C1(n13731), .C2(n16863), .A(n13310), .B(n13309), .ZN(
        P2_U2983) );
  OAI211_X1 U13763 ( .C1(n16574), .C2(n17139), .A(n11507), .B(n11506), .ZN(
        P2_U3017) );
  INV_X2 U13764 ( .A(n10496), .ZN(n10564) );
  AOI22_X1 U13765 ( .A1(n13577), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9596), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10494) );
  AND2_X4 U13766 ( .A1(n10670), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13505) );
  AND3_X4 U13767 ( .A1(n10490), .A2(n10489), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13684) );
  AOI22_X1 U13768 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13684), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10493) );
  AND2_X4 U13769 ( .A1(n10670), .A2(n14541), .ZN(n13506) );
  AOI22_X1 U13770 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13771 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10491) );
  NAND4_X1 U13772 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10495) );
  AOI22_X1 U13773 ( .A1(n9575), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9576), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10500) );
  INV_X2 U13774 ( .A(n10496), .ZN(n10545) );
  AOI22_X1 U13775 ( .A1(n13577), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9596), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13776 ( .A1(n9587), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9589), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13777 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9592), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10497) );
  NAND4_X1 U13778 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10501) );
  INV_X2 U13779 ( .A(n10502), .ZN(n10662) );
  AOI22_X1 U13780 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10662), .B1(
        n10564), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13781 ( .A1(n9575), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n13684), .ZN(n10505) );
  AOI22_X1 U13782 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13783 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13784 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9576), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13785 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13786 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13787 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10564), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13788 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13684), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13789 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13790 ( .A1(n13682), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13791 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10564), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13792 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13793 ( .A1(n9575), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9576), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13794 ( .A1(n13682), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10515) );
  NAND3_X1 U13795 ( .A1(n10556), .A2(n10553), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13796 ( .A1(n13577), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U13797 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13684), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13798 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13799 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13800 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13801 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9576), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13802 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13803 ( .A1(n13682), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10523) );
  NAND4_X1 U13804 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10552) );
  NAND3_X1 U13805 ( .A1(n10557), .A2(n10552), .A3(n10669), .ZN(n10527) );
  NAND2_X1 U13806 ( .A1(n10528), .A2(n10527), .ZN(n10529) );
  AOI22_X1 U13807 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10564), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13808 ( .A1(n9587), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13809 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13684), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13810 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13811 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13812 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13813 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13814 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13684), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10537) );
  NAND2_X1 U13815 ( .A1(n13577), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10540) );
  NAND2_X1 U13816 ( .A1(n10564), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10543) );
  AOI22_X1 U13817 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13818 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13684), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10541) );
  NAND4_X1 U13819 ( .A1(n10474), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10544) );
  AOI22_X1 U13820 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10564), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13821 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13822 ( .A1(n9575), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13684), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13823 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10546) );
  NAND4_X1 U13824 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10550) );
  NAND2_X1 U13825 ( .A1(n10550), .A2(n10669), .ZN(n10551) );
  NAND2_X1 U13826 ( .A1(n10552), .A2(n10669), .ZN(n10555) );
  NAND2_X1 U13827 ( .A1(n19895), .A2(n13347), .ZN(n10571) );
  INV_X2 U13828 ( .A(n10596), .ZN(n13700) );
  AOI22_X1 U13829 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9576), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13830 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13831 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10559) );
  NAND4_X1 U13832 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        n10563) );
  AOI22_X1 U13833 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9596), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13834 ( .A1(n9575), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13684), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13835 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13836 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10565) );
  NAND4_X1 U13837 ( .A1(n10568), .A2(n10567), .A3(n10566), .A4(n10565), .ZN(
        n10569) );
  NOR2_X1 U13838 ( .A1(n13719), .A2(n19875), .ZN(n10570) );
  NAND2_X1 U13839 ( .A1(n19875), .A2(n19895), .ZN(n11239) );
  NAND2_X1 U13840 ( .A1(n11239), .A2(n10571), .ZN(n10573) );
  NAND2_X1 U13841 ( .A1(n11287), .A2(n19869), .ZN(n10572) );
  NAND2_X1 U13842 ( .A1(n10575), .A2(n16405), .ZN(n10604) );
  NOR2_X1 U13843 ( .A1(n19875), .A2(n19895), .ZN(n10577) );
  NAND2_X1 U13844 ( .A1(n10579), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10581) );
  INV_X1 U13845 ( .A(n20608), .ZN(n10631) );
  NAND2_X1 U13846 ( .A1(n10583), .A2(n13271), .ZN(n11247) );
  INV_X1 U13847 ( .A(n11239), .ZN(n10585) );
  NAND2_X1 U13848 ( .A1(n10604), .A2(n10586), .ZN(n10588) );
  NAND2_X1 U13849 ( .A1(n10623), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10595) );
  INV_X1 U13850 ( .A(n13699), .ZN(n10591) );
  AOI22_X1 U13851 ( .A1(n9547), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10593) );
  INV_X1 U13852 ( .A(n13271), .ZN(n11193) );
  AND2_X1 U13853 ( .A1(n10593), .A2(n10592), .ZN(n10594) );
  NOR2_X1 U13854 ( .A1(n10636), .A2(n10635), .ZN(n10637) );
  NOR2_X1 U13855 ( .A1(n10597), .A2(n10596), .ZN(n10598) );
  OAI22_X1 U13856 ( .A1(n10629), .A2(n10598), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10624), .ZN(n10602) );
  NAND2_X1 U13857 ( .A1(n20608), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10599) );
  NAND2_X1 U13858 ( .A1(n10623), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10611) );
  MUX2_X1 U13859 ( .A(n13189), .B(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .S(
        P2_STATE2_REG_1__SCAN_IN), .Z(n10603) );
  AOI21_X1 U13860 ( .B1(n9547), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10603), .ZN(
        n10609) );
  NAND2_X1 U13861 ( .A1(n10629), .A2(n17154), .ZN(n10613) );
  AOI21_X1 U13862 ( .B1(n13189), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13863 ( .A1(n11084), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U13864 ( .A1(n10623), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10615) );
  NAND3_X1 U13865 ( .A1(n10617), .A2(n10616), .A3(n10615), .ZN(n10619) );
  INV_X1 U13866 ( .A(n10640), .ZN(n10620) );
  NAND2_X1 U13867 ( .A1(n10620), .A2(n10639), .ZN(n10621) );
  NAND2_X1 U13868 ( .A1(n10623), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10628) );
  AOI22_X1 U13869 ( .A1(n10624), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10626) );
  NAND2_X1 U13870 ( .A1(n11084), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10625) );
  NAND2_X1 U13871 ( .A1(n10629), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10630) );
  OAI21_X1 U13872 ( .B1(n20574), .B2(n10631), .A(n10630), .ZN(n10632) );
  INV_X1 U13873 ( .A(n10637), .ZN(n10638) );
  BUF_X1 U13874 ( .A(n10643), .Z(n10645) );
  NOR2_X1 U13875 ( .A1(n9574), .A2(n16366), .ZN(n10651) );
  INV_X1 U13876 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n21605) );
  INV_X1 U13877 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10652) );
  INV_X1 U13878 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13406) );
  INV_X1 U13879 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10654) );
  OAI22_X1 U13880 ( .A1(n20290), .A2(n13406), .B1(n20417), .B2(n10654), .ZN(
        n10655) );
  NOR2_X1 U13881 ( .A1(n10656), .A2(n10655), .ZN(n10661) );
  AND2_X2 U13882 ( .A1(n10659), .A2(n14784), .ZN(n20182) );
  AOI21_X1 U13883 ( .B1(n20182), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(n9593), .ZN(n10660) );
  AND2_X2 U13884 ( .A1(n9575), .A2(n10669), .ZN(n13528) );
  AOI22_X1 U13885 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11346), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10667) );
  AND2_X2 U13886 ( .A1(n9595), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11327) );
  AOI22_X1 U13887 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10666) );
  AND2_X2 U13888 ( .A1(n13506), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10780) );
  AOI22_X1 U13889 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13542), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10665) );
  AND2_X2 U13890 ( .A1(n13678), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10663) );
  AOI22_X1 U13891 ( .A1(n10757), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10664) );
  NAND4_X1 U13892 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10681) );
  AOI22_X1 U13893 ( .A1(n13534), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10679) );
  INV_X1 U13894 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10674) );
  AND2_X2 U13895 ( .A1(n10670), .A2(n13507), .ZN(n13535) );
  NAND2_X1 U13896 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10673) );
  AND2_X1 U13897 ( .A1(n14559), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10671) );
  NAND2_X1 U13898 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10672) );
  OAI211_X1 U13899 ( .C1(n10727), .C2(n10674), .A(n10673), .B(n10672), .ZN(
        n10675) );
  INV_X1 U13900 ( .A(n10675), .ZN(n10678) );
  AOI22_X1 U13901 ( .A1(n13541), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10677) );
  NAND2_X1 U13902 ( .A1(n13527), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10676) );
  NAND4_X1 U13903 ( .A1(n10679), .A2(n10678), .A3(n10677), .A4(n10676), .ZN(
        n10680) );
  AND2_X1 U13904 ( .A1(n11277), .A2(n9593), .ZN(n10745) );
  AOI22_X1 U13905 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13528), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13906 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10780), .B1(
        n11346), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13907 ( .A1(n10757), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13526), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10682) );
  NAND4_X1 U13909 ( .A1(n10685), .A2(n10684), .A3(n10683), .A4(n10682), .ZN(
        n10696) );
  AOI22_X1 U13910 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n13533), .B1(
        n13534), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10694) );
  INV_X1 U13911 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10689) );
  NAND2_X1 U13912 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10688) );
  NAND2_X1 U13913 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10687) );
  OAI211_X1 U13914 ( .C1(n10727), .C2(n10689), .A(n10688), .B(n10687), .ZN(
        n10690) );
  INV_X1 U13915 ( .A(n10690), .ZN(n10693) );
  AOI22_X1 U13916 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13540), .B1(
        n13541), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10692) );
  NAND2_X1 U13917 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10691) );
  NAND4_X1 U13918 ( .A1(n10694), .A2(n10693), .A3(n10692), .A4(n10691), .ZN(
        n10695) );
  NAND2_X1 U13919 ( .A1(n10745), .A2(n10900), .ZN(n10751) );
  AOI22_X1 U13920 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13528), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13921 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13526), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13922 ( .A1(n10757), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13923 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11346), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10697) );
  NAND4_X1 U13924 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n10709) );
  AOI22_X1 U13925 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n13533), .B1(
        n13534), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10707) );
  INV_X1 U13926 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13425) );
  NAND2_X1 U13927 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10702) );
  NAND2_X1 U13928 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10701) );
  OAI211_X1 U13929 ( .C1(n10727), .C2(n13425), .A(n10702), .B(n10701), .ZN(
        n10703) );
  INV_X1 U13930 ( .A(n10703), .ZN(n10706) );
  AOI22_X1 U13931 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13540), .B1(
        n13541), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U13932 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10704) );
  NAND4_X1 U13933 ( .A1(n10707), .A2(n10706), .A3(n10705), .A4(n10704), .ZN(
        n10708) );
  NAND2_X1 U13934 ( .A1(n10751), .A2(n11296), .ZN(n10750) );
  AOI22_X1 U13935 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20016), .B1(
        n10806), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13936 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20182), .B1(
        n20237), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10712) );
  NAND2_X1 U13937 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10711) );
  AOI22_X1 U13938 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10796), .B1(
        n20046), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13939 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19978), .B1(
        n19851), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10714) );
  INV_X1 U13940 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10732) );
  NAND2_X1 U13941 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10718) );
  INV_X1 U13942 ( .A(n20366), .ZN(n10716) );
  NAND2_X1 U13943 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10717) );
  OAI211_X1 U13944 ( .C1(n20140), .C2(n10732), .A(n10718), .B(n10717), .ZN(
        n10720) );
  INV_X1 U13945 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13434) );
  INV_X1 U13946 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13436) );
  NOR2_X1 U13947 ( .A1(n10720), .A2(n10719), .ZN(n10721) );
  INV_X1 U13948 ( .A(n10723), .ZN(n10726) );
  INV_X1 U13949 ( .A(n11327), .ZN(n13480) );
  INV_X1 U13950 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13433) );
  INV_X1 U13951 ( .A(n13527), .ZN(n13487) );
  INV_X1 U13952 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10724) );
  OAI22_X1 U13953 ( .A1(n13480), .A2(n13433), .B1(n13487), .B2(n10724), .ZN(
        n10725) );
  OR2_X1 U13954 ( .A1(n10726), .A2(n10725), .ZN(n10743) );
  AOI22_X1 U13955 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13535), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13956 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n13541), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10730) );
  OR2_X1 U13957 ( .A1(n10727), .A2(n13434), .ZN(n10729) );
  NAND2_X1 U13958 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10728) );
  NAND4_X1 U13959 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10735) );
  INV_X1 U13960 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13439) );
  OAI22_X1 U13961 ( .A1(n13439), .A2(n13465), .B1(n10733), .B2(n10732), .ZN(
        n10734) );
  OR2_X1 U13962 ( .A1(n10735), .A2(n10734), .ZN(n10742) );
  INV_X1 U13963 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11388) );
  INV_X1 U13964 ( .A(n10780), .ZN(n13477) );
  INV_X1 U13965 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10736) );
  OAI22_X1 U13966 ( .A1(n11388), .A2(n13477), .B1(n13475), .B2(n10736), .ZN(
        n10740) );
  INV_X1 U13967 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10738) );
  INV_X1 U13968 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10737) );
  OAI22_X1 U13969 ( .A1(n13485), .A2(n10738), .B1(n13483), .B2(n10737), .ZN(
        n10739) );
  NAND2_X1 U13970 ( .A1(n11308), .A2(n9593), .ZN(n10744) );
  INV_X1 U13971 ( .A(n10745), .ZN(n13872) );
  NAND2_X1 U13972 ( .A1(n13872), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13871) );
  INV_X1 U13973 ( .A(n13871), .ZN(n10747) );
  INV_X1 U13974 ( .A(n10900), .ZN(n10746) );
  XNOR2_X1 U13975 ( .A(n11277), .B(n10746), .ZN(n10748) );
  NAND2_X1 U13976 ( .A1(n10747), .A2(n10748), .ZN(n10749) );
  XNOR2_X1 U13977 ( .A(n13871), .B(n10748), .ZN(n13954) );
  NAND2_X1 U13978 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13954), .ZN(
        n13955) );
  NAND2_X1 U13979 ( .A1(n10749), .A2(n13955), .ZN(n10752) );
  XOR2_X1 U13980 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10752), .Z(
        n14776) );
  OAI21_X1 U13981 ( .B1(n10751), .B2(n11296), .A(n10750), .ZN(n14775) );
  NAND2_X1 U13982 ( .A1(n14776), .A2(n14775), .ZN(n10754) );
  NAND2_X1 U13983 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10752), .ZN(
        n10753) );
  NAND2_X1 U13984 ( .A1(n10754), .A2(n10753), .ZN(n10755) );
  INV_X1 U13985 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14634) );
  XNOR2_X1 U13986 ( .A(n10755), .B(n14634), .ZN(n14636) );
  NAND2_X1 U13987 ( .A1(n10755), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10756) );
  AOI22_X1 U13988 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13528), .B1(
        n11346), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13989 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13526), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13990 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13991 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10757), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10758) );
  NAND4_X1 U13992 ( .A1(n10761), .A2(n10760), .A3(n10759), .A4(n10758), .ZN(
        n10770) );
  AOI22_X1 U13993 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13533), .B1(
        n13534), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10768) );
  INV_X1 U13994 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13455) );
  NAND2_X1 U13995 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10763) );
  NAND2_X1 U13996 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10762) );
  OAI211_X1 U13997 ( .C1(n10727), .C2(n13455), .A(n10763), .B(n10762), .ZN(
        n10764) );
  INV_X1 U13998 ( .A(n10764), .ZN(n10767) );
  AOI22_X1 U13999 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13540), .B1(
        n13541), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10766) );
  NAND2_X1 U14000 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10765) );
  NAND4_X1 U14001 ( .A1(n10768), .A2(n10767), .A3(n10766), .A4(n10765), .ZN(
        n10769) );
  INV_X1 U14002 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16853) );
  INV_X1 U14003 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U14004 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10773) );
  NAND2_X1 U14005 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10772) );
  INV_X1 U14006 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13466) );
  INV_X1 U14007 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13644) );
  AOI22_X1 U14008 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19851), .B1(
        n19978), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U14009 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10775) );
  AOI22_X1 U14010 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U14011 ( .A1(n11346), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U14012 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13542), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U14013 ( .A1(n13526), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10781) );
  NAND4_X1 U14014 ( .A1(n10784), .A2(n10783), .A3(n10782), .A4(n10781), .ZN(
        n10793) );
  AOI22_X1 U14015 ( .A1(n13534), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10791) );
  NAND2_X1 U14016 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10786) );
  NAND2_X1 U14017 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10785) );
  OAI211_X1 U14018 ( .C1(n10727), .C2(n13466), .A(n10786), .B(n10785), .ZN(
        n10787) );
  INV_X1 U14019 ( .A(n10787), .ZN(n10790) );
  AOI22_X1 U14020 ( .A1(n13541), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10789) );
  NAND2_X1 U14021 ( .A1(n13527), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10788) );
  NAND4_X1 U14022 ( .A1(n10791), .A2(n10790), .A3(n10789), .A4(n10788), .ZN(
        n10792) );
  INV_X1 U14023 ( .A(n11318), .ZN(n10794) );
  NAND2_X1 U14024 ( .A1(n10794), .A2(n9593), .ZN(n10795) );
  INV_X1 U14025 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17110) );
  INV_X1 U14026 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10808) );
  INV_X1 U14027 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13486) );
  AOI22_X1 U14028 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20182), .B1(
        n20237), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U14029 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10779), .B1(
        n20324), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10800) );
  NAND2_X1 U14030 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10799) );
  INV_X1 U14031 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13478) );
  NAND2_X1 U14032 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10805) );
  NAND2_X1 U14033 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10804) );
  OAI211_X1 U14034 ( .C1(n20140), .C2(n13478), .A(n10805), .B(n10804), .ZN(
        n10807) );
  AOI22_X1 U14035 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U14036 ( .A1(n13541), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10811) );
  OR2_X1 U14037 ( .A1(n10727), .A2(n10808), .ZN(n10810) );
  NAND2_X1 U14038 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10809) );
  NAND4_X1 U14039 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(
        n10814) );
  INV_X1 U14040 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13499) );
  OAI22_X1 U14041 ( .A1(n10733), .A2(n13478), .B1(n13465), .B2(n13499), .ZN(
        n10813) );
  NOR2_X1 U14042 ( .A1(n10814), .A2(n10813), .ZN(n10820) );
  INV_X1 U14043 ( .A(n13528), .ZN(n13489) );
  INV_X1 U14044 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13474) );
  INV_X1 U14045 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13481) );
  OAI22_X1 U14046 ( .A1(n13489), .A2(n13474), .B1(n13487), .B2(n13481), .ZN(
        n10816) );
  INV_X1 U14047 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13476) );
  INV_X1 U14048 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13488) );
  OAI22_X1 U14049 ( .A1(n13485), .A2(n13476), .B1(n13483), .B2(n13488), .ZN(
        n10815) );
  NOR2_X1 U14050 ( .A1(n10816), .A2(n10815), .ZN(n10819) );
  AOI22_X1 U14051 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U14052 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10817) );
  NAND4_X1 U14053 ( .A1(n10820), .A2(n10819), .A3(n10818), .A4(n10817), .ZN(
        n11322) );
  INV_X1 U14054 ( .A(n11322), .ZN(n10821) );
  NAND2_X1 U14055 ( .A1(n10821), .A2(n9593), .ZN(n10822) );
  NAND2_X1 U14056 ( .A1(n10823), .A2(n10937), .ZN(n10824) );
  INV_X1 U14057 ( .A(n10829), .ZN(n10850) );
  NAND2_X1 U14058 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10833) );
  NAND2_X1 U14059 ( .A1(n10757), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10832) );
  NAND2_X1 U14060 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10831) );
  NAND2_X1 U14061 ( .A1(n13526), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10830) );
  NAND2_X1 U14062 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10837) );
  NAND2_X1 U14063 ( .A1(n11346), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10836) );
  NAND2_X1 U14064 ( .A1(n13527), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10835) );
  NAND2_X1 U14065 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10834) );
  AOI22_X1 U14066 ( .A1(n13534), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10847) );
  INV_X1 U14067 ( .A(n13542), .ZN(n13437) );
  INV_X1 U14068 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10840) );
  NAND2_X1 U14069 ( .A1(n13541), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10839) );
  NAND2_X1 U14070 ( .A1(n13540), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10838) );
  OAI211_X1 U14071 ( .C1(n13437), .C2(n10840), .A(n10839), .B(n10838), .ZN(
        n10845) );
  INV_X1 U14072 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10843) );
  NAND2_X1 U14073 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10842) );
  NAND2_X1 U14074 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10841) );
  OAI211_X1 U14075 ( .C1(n10727), .C2(n10843), .A(n10842), .B(n10841), .ZN(
        n10844) );
  NOR2_X1 U14076 ( .A1(n10845), .A2(n10844), .ZN(n10846) );
  INV_X1 U14077 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17080) );
  OAI21_X1 U14078 ( .B1(n16791), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10851) );
  OAI21_X1 U14079 ( .B1(n16795), .B2(n17080), .A(n10851), .ZN(n10852) );
  AND2_X1 U14080 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11265) );
  NAND2_X1 U14081 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17024) );
  INV_X1 U14082 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16699) );
  NOR2_X1 U14083 ( .A1(n17024), .A2(n16699), .ZN(n16984) );
  NAND2_X1 U14084 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13147) );
  INV_X1 U14085 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16989) );
  NOR2_X1 U14086 ( .A1(n13147), .A2(n16989), .ZN(n10854) );
  AND2_X1 U14087 ( .A1(n16984), .A2(n10854), .ZN(n13163) );
  AND3_X1 U14088 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10855) );
  AND2_X1 U14089 ( .A1(n13163), .A2(n10855), .ZN(n16949) );
  NAND2_X1 U14090 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16949), .ZN(
        n14820) );
  INV_X1 U14091 ( .A(n14820), .ZN(n14818) );
  NAND4_X1 U14092 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(n14818), .ZN(n11267) );
  NAND3_X1 U14093 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11268) );
  NOR2_X1 U14094 ( .A1(n11267), .A2(n11268), .ZN(n10856) );
  INV_X1 U14095 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11538) );
  INV_X1 U14096 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11539) );
  NAND2_X1 U14097 ( .A1(n16594), .A2(n11539), .ZN(n10857) );
  AND2_X1 U14098 ( .A1(n9593), .A2(n10578), .ZN(n13268) );
  INV_X1 U14099 ( .A(n13268), .ZN(n10859) );
  NOR2_X1 U14100 ( .A1(n10858), .A2(n10859), .ZN(n20595) );
  XNOR2_X1 U14101 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11176) );
  NAND2_X1 U14102 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20291), .ZN(
        n10889) );
  NAND2_X1 U14103 ( .A1(n11176), .A2(n10860), .ZN(n10862) );
  NAND2_X1 U14104 ( .A1(n20591), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10861) );
  NAND2_X1 U14105 ( .A1(n10862), .A2(n10861), .ZN(n10871) );
  XNOR2_X1 U14106 ( .A(n17154), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10870) );
  NAND2_X1 U14107 ( .A1(n10871), .A2(n10870), .ZN(n10869) );
  NAND2_X1 U14108 ( .A1(n20582), .A2(n17154), .ZN(n10863) );
  NAND2_X1 U14109 ( .A1(n10869), .A2(n10863), .ZN(n10878) );
  XNOR2_X1 U14110 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10877) );
  NOR2_X1 U14111 ( .A1(n10669), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10864) );
  AOI21_X1 U14112 ( .B1(n10878), .B2(n10877), .A(n10864), .ZN(n10882) );
  INV_X1 U14113 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n10865) );
  NAND2_X1 U14114 ( .A1(n10865), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10866) );
  NAND2_X1 U14115 ( .A1(n10882), .A2(n10866), .ZN(n10868) );
  INV_X1 U14116 ( .A(n10881), .ZN(n10867) );
  OAI21_X1 U14117 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20291), .A(
        n10889), .ZN(n11177) );
  INV_X1 U14118 ( .A(n11177), .ZN(n11179) );
  MUX2_X1 U14119 ( .A(n11277), .B(n11179), .S(n13271), .Z(n10919) );
  INV_X1 U14120 ( .A(n10919), .ZN(n10876) );
  INV_X1 U14121 ( .A(n11176), .ZN(n10875) );
  OAI21_X1 U14122 ( .B1(n10871), .B2(n10870), .A(n10869), .ZN(n11182) );
  INV_X1 U14123 ( .A(n11182), .ZN(n10872) );
  INV_X1 U14124 ( .A(n10899), .ZN(n10874) );
  OAI21_X1 U14125 ( .B1(n10876), .B2(n10875), .A(n10874), .ZN(n10886) );
  XNOR2_X1 U14126 ( .A(n10878), .B(n10877), .ZN(n11186) );
  INV_X1 U14127 ( .A(n10903), .ZN(n10884) );
  AND2_X1 U14128 ( .A1(n10882), .A2(n10881), .ZN(n11192) );
  INV_X1 U14129 ( .A(n11192), .ZN(n10883) );
  MUX2_X1 U14130 ( .A(n11312), .B(n10883), .S(n13271), .Z(n10906) );
  NAND2_X1 U14131 ( .A1(n10884), .A2(n10906), .ZN(n11174) );
  INV_X1 U14132 ( .A(n11174), .ZN(n10885) );
  NAND2_X1 U14133 ( .A1(n10886), .A2(n10885), .ZN(n20597) );
  NAND3_X1 U14134 ( .A1(n20595), .A2(n20598), .A3(n20597), .ZN(n10897) );
  INV_X1 U14135 ( .A(n10858), .ZN(n10895) );
  INV_X1 U14136 ( .A(n14202), .ZN(n10887) );
  AND2_X1 U14137 ( .A1(n10887), .A2(n17496), .ZN(n17492) );
  NAND2_X1 U14138 ( .A1(n13480), .A2(n17492), .ZN(n10888) );
  INV_X1 U14139 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n17498) );
  NAND2_X1 U14140 ( .A1(n10888), .A2(n17498), .ZN(n21688) );
  NOR3_X1 U14141 ( .A1(n11186), .A2(n11182), .A3(n11192), .ZN(n10890) );
  INV_X1 U14142 ( .A(n10890), .ZN(n10892) );
  XNOR2_X1 U14143 ( .A(n11176), .B(n10889), .ZN(n11178) );
  NAND2_X1 U14144 ( .A1(n11178), .A2(n10890), .ZN(n10891) );
  OAI21_X1 U14145 ( .B1(n11177), .B2(n10892), .A(n14574), .ZN(n10893) );
  INV_X1 U14146 ( .A(n10893), .ZN(n10894) );
  MUX2_X1 U14147 ( .A(n21688), .B(n10894), .S(n17141), .Z(n17499) );
  NAND3_X1 U14148 ( .A1(n10895), .A2(n17491), .A3(n17499), .ZN(n10896) );
  NAND2_X1 U14149 ( .A1(n10578), .A2(n14601), .ZN(n10898) );
  INV_X1 U14150 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n16321) );
  MUX2_X1 U14151 ( .A(n10899), .B(n16321), .S(n9590), .Z(n10914) );
  INV_X1 U14152 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14008) );
  INV_X1 U14153 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n16349) );
  NAND3_X1 U14154 ( .A1(n9590), .A2(n14008), .A3(n16349), .ZN(n10901) );
  NAND2_X1 U14155 ( .A1(n10900), .A2(n10902), .ZN(n11286) );
  NAND2_X1 U14156 ( .A1(n10901), .A2(n11286), .ZN(n10915) );
  NAND2_X1 U14157 ( .A1(n10914), .A2(n10915), .ZN(n10918) );
  NAND2_X1 U14158 ( .A1(n10903), .A2(n10902), .ZN(n10905) );
  INV_X1 U14159 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n16290) );
  MUX2_X1 U14160 ( .A(n10906), .B(n16290), .S(n9590), .Z(n10926) );
  INV_X1 U14161 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14241) );
  MUX2_X1 U14162 ( .A(n14241), .B(n11318), .S(n10902), .Z(n10908) );
  NAND2_X1 U14163 ( .A1(n10373), .A2(n10371), .ZN(n10909) );
  NAND2_X1 U14164 ( .A1(n10945), .A2(n10909), .ZN(n16284) );
  NAND2_X1 U14165 ( .A1(n14635), .A2(n11513), .ZN(n10913) );
  INV_X1 U14166 ( .A(n10910), .ZN(n10928) );
  NAND2_X1 U14167 ( .A1(n10918), .A2(n10911), .ZN(n10912) );
  NAND2_X1 U14168 ( .A1(n10928), .A2(n10912), .ZN(n16313) );
  INV_X1 U14169 ( .A(n10914), .ZN(n10916) );
  INV_X1 U14170 ( .A(n10915), .ZN(n10921) );
  NAND2_X1 U14171 ( .A1(n10916), .A2(n10921), .ZN(n10917) );
  NAND2_X1 U14172 ( .A1(n10918), .A2(n10917), .ZN(n16322) );
  XNOR2_X1 U14173 ( .A(n16322), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14774) );
  MUX2_X1 U14174 ( .A(n10919), .B(P2_EBX_REG_0__SCAN_IN), .S(n9590), .Z(n16356) );
  NAND2_X1 U14175 ( .A1(n16356), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13953) );
  NAND3_X1 U14176 ( .A1(n9590), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U14177 ( .A1(n10921), .A2(n10920), .ZN(n16334) );
  INV_X1 U14178 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14056) );
  AND2_X1 U14179 ( .A1(n16334), .A2(n14056), .ZN(n10922) );
  OAI22_X1 U14180 ( .A1(n13953), .A2(n10922), .B1(n14056), .B2(n16334), .ZN(
        n14773) );
  NAND2_X1 U14181 ( .A1(n14774), .A2(n14773), .ZN(n10925) );
  INV_X1 U14182 ( .A(n16322), .ZN(n10923) );
  NAND2_X1 U14183 ( .A1(n10923), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10924) );
  NAND2_X1 U14184 ( .A1(n10925), .A2(n10924), .ZN(n16848) );
  INV_X1 U14185 ( .A(n10926), .ZN(n10927) );
  NAND2_X1 U14186 ( .A1(n10928), .A2(n10927), .ZN(n10929) );
  NAND2_X1 U14187 ( .A1(n10373), .A2(n10929), .ZN(n16850) );
  NAND2_X1 U14188 ( .A1(n16850), .A2(n16853), .ZN(n10931) );
  OAI21_X1 U14189 ( .B1(n16848), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10931), .ZN(n10930) );
  INV_X1 U14190 ( .A(n10930), .ZN(n10934) );
  NAND3_X1 U14191 ( .A1(n10931), .A2(n16848), .A3(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10932) );
  OAI21_X1 U14192 ( .B1(n16850), .B2(n16853), .A(n10932), .ZN(n10933) );
  NAND2_X1 U14193 ( .A1(n16818), .A2(n16835), .ZN(n10941) );
  NAND2_X1 U14194 ( .A1(n10939), .A2(n10937), .ZN(n10938) );
  INV_X1 U14195 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n16262) );
  MUX2_X1 U14196 ( .A(n16262), .B(n11322), .S(n10902), .Z(n10943) );
  INV_X1 U14197 ( .A(n10943), .ZN(n10953) );
  XNOR2_X1 U14198 ( .A(n10945), .B(n10953), .ZN(n16269) );
  INV_X1 U14199 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17100) );
  NAND2_X1 U14200 ( .A1(n10942), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16767) );
  INV_X1 U14201 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14419) );
  MUX2_X1 U14202 ( .A(n14419), .B(n13293), .S(n10902), .Z(n10951) );
  NAND2_X1 U14203 ( .A1(n10943), .A2(n10951), .ZN(n10944) );
  NAND2_X1 U14204 ( .A1(n9591), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10947) );
  INV_X1 U14205 ( .A(n10947), .ZN(n10948) );
  NAND2_X1 U14206 ( .A1(n10007), .A2(n10948), .ZN(n10949) );
  AND2_X1 U14207 ( .A1(n13293), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10950) );
  NAND2_X1 U14208 ( .A1(n16245), .A2(n10950), .ZN(n16782) );
  INV_X1 U14209 ( .A(n10951), .ZN(n10952) );
  OAI21_X1 U14210 ( .B1(n10945), .B2(n10953), .A(n10952), .ZN(n10954) );
  NAND2_X1 U14211 ( .A1(n16251), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16808) );
  AND2_X1 U14212 ( .A1(n16782), .A2(n16808), .ZN(n16768) );
  INV_X1 U14213 ( .A(n16245), .ZN(n10956) );
  INV_X1 U14214 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17068) );
  OAI21_X1 U14215 ( .B1(n10956), .B2(n11513), .A(n17068), .ZN(n16783) );
  INV_X1 U14216 ( .A(n16251), .ZN(n10957) );
  NAND2_X1 U14217 ( .A1(n10957), .A2(n17080), .ZN(n16806) );
  AND2_X1 U14218 ( .A1(n16783), .A2(n16806), .ZN(n16769) );
  NAND2_X1 U14219 ( .A1(n9590), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10958) );
  XNOR2_X1 U14220 ( .A(n10961), .B(n10958), .ZN(n16223) );
  NAND2_X1 U14221 ( .A1(n16223), .A2(n13293), .ZN(n10989) );
  INV_X1 U14222 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17056) );
  NAND2_X1 U14223 ( .A1(n10989), .A2(n17056), .ZN(n16771) );
  AND2_X1 U14224 ( .A1(n16769), .A2(n16771), .ZN(n10959) );
  INV_X1 U14225 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n14272) );
  INV_X1 U14226 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n16191) );
  NOR2_X1 U14227 ( .A1(n10902), .A2(n16191), .ZN(n10991) );
  INV_X1 U14228 ( .A(n10991), .ZN(n10965) );
  NAND2_X1 U14229 ( .A1(n9591), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10999) );
  OAI21_X1 U14230 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n9590), .ZN(n10966) );
  INV_X1 U14231 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n16135) );
  NAND2_X1 U14232 ( .A1(n9591), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10976) );
  INV_X1 U14233 ( .A(n10975), .ZN(n10968) );
  INV_X1 U14234 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10967) );
  INV_X1 U14235 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n16095) );
  NOR2_X1 U14236 ( .A1(n10902), .A2(n16095), .ZN(n10973) );
  INV_X1 U14237 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n16431) );
  INV_X1 U14238 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10969) );
  AND2_X1 U14239 ( .A1(n9656), .A2(n10970), .ZN(n10971) );
  OR2_X1 U14240 ( .A1(n11029), .A2(n10971), .ZN(n16069) );
  NAND2_X1 U14241 ( .A1(n11013), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14839) );
  INV_X1 U14242 ( .A(n10973), .ZN(n10974) );
  XNOR2_X1 U14243 ( .A(n10972), .B(n10974), .ZN(n16093) );
  NAND2_X1 U14244 ( .A1(n16093), .A2(n13293), .ZN(n11015) );
  INV_X1 U14245 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16939) );
  INV_X1 U14246 ( .A(n10976), .ZN(n10977) );
  NAND2_X1 U14247 ( .A1(n9689), .A2(n10977), .ZN(n10978) );
  NAND2_X1 U14248 ( .A1(n10975), .A2(n10978), .ZN(n16126) );
  NOR2_X1 U14249 ( .A1(n11019), .A2(n16674), .ZN(n14811) );
  NAND3_X1 U14250 ( .A1(n10979), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n9590), .ZN(
        n10980) );
  OAI211_X1 U14251 ( .C1(n10979), .C2(P2_EBX_REG_16__SCAN_IN), .A(n10980), .B(
        n11043), .ZN(n16133) );
  NOR2_X1 U14252 ( .A1(n16133), .A2(n11513), .ZN(n11017) );
  NAND2_X1 U14253 ( .A1(n11017), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13159) );
  NOR2_X1 U14254 ( .A1(n10902), .A2(n10964), .ZN(n10981) );
  AND2_X1 U14255 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  NOR2_X1 U14256 ( .A1(n10984), .A2(n10983), .ZN(n16202) );
  NAND2_X1 U14257 ( .A1(n16202), .A2(n13293), .ZN(n11022) );
  OR2_X1 U14258 ( .A1(n11022), .A2(n16699), .ZN(n16743) );
  NAND2_X1 U14259 ( .A1(n9591), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10986) );
  MUX2_X1 U14260 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n10986), .S(n10985), .Z(
        n10987) );
  NAND2_X1 U14261 ( .A1(n10987), .A2(n11043), .ZN(n16211) );
  NAND2_X1 U14262 ( .A1(n13293), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10988) );
  OR2_X1 U14263 ( .A1(n16211), .A2(n10988), .ZN(n16756) );
  OR2_X1 U14264 ( .A1(n10989), .A2(n17056), .ZN(n16772) );
  AND2_X1 U14265 ( .A1(n16756), .A2(n16772), .ZN(n16740) );
  NAND2_X1 U14266 ( .A1(n16743), .A2(n16740), .ZN(n16715) );
  INV_X1 U14267 ( .A(n10990), .ZN(n11001) );
  NAND2_X1 U14268 ( .A1(n10992), .A2(n10991), .ZN(n10993) );
  NAND2_X1 U14269 ( .A1(n11001), .A2(n10993), .ZN(n16188) );
  NAND2_X1 U14270 ( .A1(n13293), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10994) );
  NOR2_X1 U14271 ( .A1(n16188), .A2(n10994), .ZN(n16725) );
  NOR2_X1 U14272 ( .A1(n16715), .A2(n16725), .ZN(n11003) );
  INV_X1 U14273 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10995) );
  NAND2_X1 U14274 ( .A1(n10998), .A2(n10995), .ZN(n11007) );
  NAND3_X1 U14275 ( .A1(n11007), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n9590), .ZN(
        n10996) );
  AND2_X1 U14276 ( .A1(n10996), .A2(n10979), .ZN(n16153) );
  AND2_X1 U14277 ( .A1(n13293), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10997) );
  NAND2_X1 U14278 ( .A1(n16153), .A2(n10997), .ZN(n16687) );
  INV_X1 U14279 ( .A(n10999), .ZN(n11000) );
  NAND2_X1 U14280 ( .A1(n11001), .A2(n11000), .ZN(n11002) );
  NAND2_X1 U14281 ( .A1(n11005), .A2(n11002), .ZN(n16171) );
  INV_X1 U14282 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17002) );
  NOR3_X1 U14283 ( .A1(n16171), .A2(n11513), .A3(n17002), .ZN(n13156) );
  INV_X1 U14284 ( .A(n13156), .ZN(n16713) );
  NAND4_X1 U14285 ( .A1(n13159), .A2(n11003), .A3(n16687), .A4(n16713), .ZN(
        n11004) );
  NOR2_X1 U14286 ( .A1(n14811), .A2(n11004), .ZN(n11009) );
  XNOR2_X1 U14287 ( .A(n10975), .B(n10470), .ZN(n16114) );
  NAND2_X1 U14288 ( .A1(n16114), .A2(n13293), .ZN(n11016) );
  INV_X1 U14289 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16952) );
  OR2_X1 U14290 ( .A1(n11016), .A2(n16952), .ZN(n16663) );
  NAND2_X1 U14291 ( .A1(n9591), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U14292 ( .A1(n11008), .A2(n11007), .ZN(n16168) );
  NOR2_X1 U14293 ( .A1(n16168), .A2(n11513), .ZN(n11024) );
  NAND2_X1 U14294 ( .A1(n11024), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16703) );
  AND4_X1 U14295 ( .A1(n16651), .A2(n11009), .A3(n16663), .A4(n16703), .ZN(
        n11012) );
  NAND2_X1 U14296 ( .A1(n9659), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11010) );
  MUX2_X1 U14297 ( .A(n9659), .B(n11010), .S(n9591), .Z(n11011) );
  NAND2_X1 U14298 ( .A1(n11027), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14837) );
  AND3_X1 U14299 ( .A1(n14839), .A2(n11012), .A3(n14837), .ZN(n16607) );
  INV_X1 U14300 ( .A(n11013), .ZN(n11014) );
  INV_X1 U14301 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14892) );
  NAND2_X1 U14302 ( .A1(n11014), .A2(n14892), .ZN(n14838) );
  NAND2_X1 U14303 ( .A1(n11015), .A2(n16939), .ZN(n16650) );
  NAND2_X1 U14304 ( .A1(n11016), .A2(n16952), .ZN(n16662) );
  INV_X1 U14305 ( .A(n11017), .ZN(n11018) );
  XNOR2_X1 U14306 ( .A(n11018), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16681) );
  NAND2_X1 U14307 ( .A1(n11019), .A2(n16674), .ZN(n14810) );
  INV_X1 U14308 ( .A(n16153), .ZN(n11020) );
  INV_X1 U14309 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16974) );
  NAND2_X1 U14310 ( .A1(n9666), .A2(n17002), .ZN(n16712) );
  INV_X1 U14311 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16730) );
  OAI21_X1 U14312 ( .B1(n16188), .B2(n11513), .A(n16730), .ZN(n16726) );
  OR2_X1 U14313 ( .A1(n16211), .A2(n11513), .ZN(n11021) );
  INV_X1 U14314 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17029) );
  NAND2_X1 U14315 ( .A1(n11021), .A2(n17029), .ZN(n16757) );
  NAND2_X1 U14316 ( .A1(n11022), .A2(n16699), .ZN(n16742) );
  AND3_X1 U14317 ( .A1(n16726), .A2(n16757), .A3(n16742), .ZN(n11023) );
  AND2_X1 U14318 ( .A1(n16712), .A2(n11023), .ZN(n13155) );
  AND2_X1 U14319 ( .A1(n16688), .A2(n13155), .ZN(n11026) );
  INV_X1 U14320 ( .A(n11024), .ZN(n11025) );
  NAND2_X1 U14321 ( .A1(n11025), .A2(n16989), .ZN(n16702) );
  INV_X1 U14322 ( .A(n11027), .ZN(n11028) );
  INV_X1 U14323 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14893) );
  NAND2_X1 U14324 ( .A1(n11028), .A2(n14893), .ZN(n14832) );
  NAND2_X1 U14325 ( .A1(n9590), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11031) );
  INV_X1 U14326 ( .A(n11031), .ZN(n11032) );
  NAND2_X1 U14327 ( .A1(n11030), .A2(n11032), .ZN(n11033) );
  NAND2_X1 U14328 ( .A1(n11041), .A2(n11033), .ZN(n16057) );
  INV_X1 U14329 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16928) );
  NAND2_X1 U14330 ( .A1(n11036), .A2(n16928), .ZN(n16630) );
  INV_X1 U14331 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16038) );
  XNOR2_X1 U14332 ( .A(n11041), .B(n10473), .ZN(n16045) );
  NAND2_X1 U14333 ( .A1(n16045), .A2(n13293), .ZN(n16610) );
  INV_X1 U14334 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16919) );
  NAND2_X1 U14335 ( .A1(n16610), .A2(n16919), .ZN(n11034) );
  NAND2_X1 U14336 ( .A1(n16631), .A2(n16919), .ZN(n11037) );
  INV_X1 U14337 ( .A(n16610), .ZN(n16611) );
  NAND2_X1 U14338 ( .A1(n11043), .A2(n13293), .ZN(n11039) );
  INV_X1 U14339 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16618) );
  NOR2_X1 U14340 ( .A1(n11039), .A2(n16618), .ZN(n16612) );
  AOI21_X1 U14341 ( .B1(n11037), .B2(n16611), .A(n16612), .ZN(n11038) );
  NAND2_X1 U14342 ( .A1(n11039), .A2(n16618), .ZN(n16613) );
  INV_X1 U14343 ( .A(n16599), .ZN(n11040) );
  NAND2_X1 U14344 ( .A1(n11039), .A2(n11538), .ZN(n16595) );
  NOR2_X1 U14345 ( .A1(n11039), .A2(n11538), .ZN(n16597) );
  NOR2_X1 U14346 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n11042) );
  NAND2_X1 U14347 ( .A1(n16028), .A2(n11042), .ZN(n11160) );
  INV_X1 U14348 ( .A(n11157), .ZN(n13291) );
  OAI211_X1 U14349 ( .C1(n16008), .C2(P2_EBX_REG_25__SCAN_IN), .A(
        P2_EBX_REG_26__SCAN_IN), .B(n9591), .ZN(n11044) );
  AND2_X1 U14350 ( .A1(n13293), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11045) );
  NAND2_X1 U14351 ( .A1(n15998), .A2(n11045), .ZN(n11169) );
  INV_X1 U14352 ( .A(n15998), .ZN(n11046) );
  OAI21_X1 U14353 ( .B1(n11046), .B2(n11513), .A(n11539), .ZN(n11047) );
  NAND2_X1 U14354 ( .A1(n13299), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11052) );
  AOI22_X1 U14355 ( .A1(n11523), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11050) );
  NAND2_X1 U14356 ( .A1(n11084), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11049) );
  AND2_X1 U14357 ( .A1(n11050), .A2(n11049), .ZN(n11051) );
  NAND2_X1 U14358 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11057) );
  AOI22_X1 U14359 ( .A1(n11523), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11055) );
  NAND2_X1 U14360 ( .A1(n11084), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11054) );
  AND2_X1 U14361 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  INV_X1 U14362 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20503) );
  NAND2_X1 U14363 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11059) );
  AOI22_X1 U14364 ( .A1(n11523), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11058) );
  OAI211_X1 U14365 ( .C1(n20503), .C2(n13297), .A(n11059), .B(n11058), .ZN(
        n14286) );
  NAND2_X1 U14366 ( .A1(n14239), .A2(n14286), .ZN(n14285) );
  INV_X1 U14367 ( .A(n14285), .ZN(n11065) );
  NAND2_X1 U14368 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11063) );
  AOI22_X1 U14369 ( .A1(n11523), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11061) );
  NAND2_X1 U14370 ( .A1(n11084), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11060) );
  AND2_X1 U14371 ( .A1(n11061), .A2(n11060), .ZN(n11062) );
  NAND2_X1 U14372 ( .A1(n11065), .A2(n11064), .ZN(n14400) );
  NAND2_X1 U14373 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11069) );
  AOI22_X1 U14374 ( .A1(n11523), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11067) );
  NAND2_X1 U14375 ( .A1(n11084), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11066) );
  AND2_X1 U14376 ( .A1(n11067), .A2(n11066), .ZN(n11068) );
  INV_X1 U14377 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20508) );
  NAND2_X1 U14378 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11071) );
  AOI22_X1 U14379 ( .A1(n11523), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11070) );
  OAI211_X1 U14380 ( .C1(n20508), .C2(n13297), .A(n11071), .B(n11070), .ZN(
        n14269) );
  NAND2_X1 U14381 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11075) );
  AOI22_X1 U14382 ( .A1(n11523), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11073) );
  NAND2_X1 U14383 ( .A1(n11084), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11072) );
  AND2_X1 U14384 ( .A1(n11073), .A2(n11072), .ZN(n11074) );
  NAND2_X1 U14385 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11079) );
  AOI22_X1 U14386 ( .A1(n11523), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11077) );
  NAND2_X1 U14387 ( .A1(n11084), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11076) );
  AND2_X1 U14388 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  NAND2_X1 U14389 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11083) );
  AOI22_X1 U14390 ( .A1(n10624), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11081) );
  NAND2_X1 U14391 ( .A1(n11084), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11080) );
  AND2_X1 U14392 ( .A1(n11081), .A2(n11080), .ZN(n11082) );
  NAND2_X1 U14393 ( .A1(n11083), .A2(n11082), .ZN(n14433) );
  AND2_X2 U14394 ( .A1(n14325), .A2(n14433), .ZN(n14440) );
  NAND2_X1 U14395 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11088) );
  AOI22_X1 U14396 ( .A1(n10624), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11086) );
  NAND2_X1 U14397 ( .A1(n11084), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11085) );
  AND2_X1 U14398 ( .A1(n11086), .A2(n11085), .ZN(n11087) );
  NAND2_X1 U14399 ( .A1(n11088), .A2(n11087), .ZN(n14439) );
  AND2_X2 U14400 ( .A1(n14440), .A2(n14439), .ZN(n13151) );
  INV_X1 U14401 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20519) );
  NAND2_X1 U14402 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11090) );
  AOI22_X1 U14403 ( .A1(n11523), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11089) );
  OAI211_X1 U14404 ( .C1(n20519), .C2(n13297), .A(n11090), .B(n11089), .ZN(
        n13152) );
  NAND2_X1 U14405 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11094) );
  AOI22_X1 U14406 ( .A1(n11523), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11092) );
  NAND2_X1 U14407 ( .A1(n11223), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11091) );
  AND2_X1 U14408 ( .A1(n11092), .A2(n11091), .ZN(n11093) );
  AND2_X1 U14409 ( .A1(n11094), .A2(n11093), .ZN(n14669) );
  NAND2_X1 U14410 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11098) );
  AOI22_X1 U14411 ( .A1(n11523), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11096) );
  NAND2_X1 U14412 ( .A1(n11223), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11095) );
  AND2_X1 U14413 ( .A1(n11096), .A2(n11095), .ZN(n11097) );
  NAND2_X1 U14414 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11102) );
  AOI22_X1 U14415 ( .A1(n11523), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11100) );
  NAND2_X1 U14416 ( .A1(n11223), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11099) );
  AND2_X1 U14417 ( .A1(n11100), .A2(n11099), .ZN(n11101) );
  NOR2_X1 U14418 ( .A1(n14669), .A2(n14653), .ZN(n13150) );
  NAND2_X1 U14419 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11107) );
  AOI22_X1 U14420 ( .A1(n11523), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11105) );
  NAND2_X1 U14421 ( .A1(n11223), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11104) );
  AND2_X1 U14422 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  NAND2_X1 U14423 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11111) );
  AOI22_X1 U14424 ( .A1(n10624), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11109) );
  NAND2_X1 U14425 ( .A1(n11223), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11108) );
  AND2_X1 U14426 ( .A1(n11109), .A2(n11108), .ZN(n11110) );
  NAND2_X1 U14427 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11115) );
  AOI22_X1 U14428 ( .A1(n10624), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11113) );
  NAND2_X1 U14429 ( .A1(n11223), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11112) );
  AND2_X1 U14430 ( .A1(n11113), .A2(n11112), .ZN(n11114) );
  INV_X1 U14431 ( .A(n16053), .ZN(n11122) );
  INV_X1 U14432 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20527) );
  NAND2_X1 U14433 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11117) );
  AOI22_X1 U14434 ( .A1(n10624), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11116) );
  OAI211_X1 U14435 ( .C1(n20527), .C2(n13297), .A(n11117), .B(n11116), .ZN(
        n14844) );
  NAND2_X1 U14436 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11121) );
  AOI22_X1 U14437 ( .A1(n11523), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11119) );
  NAND2_X1 U14438 ( .A1(n11223), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11118) );
  AND2_X1 U14439 ( .A1(n11119), .A2(n11118), .ZN(n11120) );
  NAND2_X1 U14440 ( .A1(n11121), .A2(n11120), .ZN(n14817) );
  NAND2_X1 U14441 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11127) );
  AOI22_X1 U14442 ( .A1(n10624), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11125) );
  NAND2_X1 U14443 ( .A1(n11223), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11124) );
  AND2_X1 U14444 ( .A1(n11125), .A2(n11124), .ZN(n11126) );
  NAND2_X1 U14445 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11131) );
  AOI22_X1 U14446 ( .A1(n10624), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11129) );
  NAND2_X1 U14447 ( .A1(n11223), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11128) );
  AND2_X1 U14448 ( .A1(n11129), .A2(n11128), .ZN(n11130) );
  NAND2_X1 U14449 ( .A1(n11131), .A2(n11130), .ZN(n16019) );
  NAND2_X1 U14450 ( .A1(n16018), .A2(n16019), .ZN(n16001) );
  NAND2_X1 U14451 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11135) );
  AOI22_X1 U14452 ( .A1(n10624), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11133) );
  NAND2_X1 U14453 ( .A1(n11223), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11132) );
  AND2_X1 U14454 ( .A1(n11133), .A2(n11132), .ZN(n11134) );
  NOR2_X2 U14455 ( .A1(n16001), .A2(n16002), .ZN(n11141) );
  NAND2_X1 U14456 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11139) );
  AOI22_X1 U14457 ( .A1(n10624), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11137) );
  NAND2_X1 U14458 ( .A1(n11223), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11136) );
  AND2_X1 U14459 ( .A1(n11137), .A2(n11136), .ZN(n11138) );
  INV_X1 U14460 ( .A(n11143), .ZN(n11140) );
  NAND2_X1 U14461 ( .A1(n11142), .A2(n11143), .ZN(n11144) );
  NOR2_X1 U14462 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14591) );
  NAND2_X1 U14463 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n21689) );
  INV_X1 U14464 ( .A(n21689), .ZN(n13817) );
  OAI22_X1 U14465 ( .A1(n14591), .A2(n13817), .B1(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20607), .ZN(n11145) );
  INV_X1 U14466 ( .A(n19838), .ZN(n16827) );
  INV_X1 U14467 ( .A(n11146), .ZN(n13828) );
  NOR2_X1 U14468 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17490) );
  OR2_X1 U14469 ( .A1(n20606), .A2(n17490), .ZN(n20583) );
  NAND2_X1 U14470 ( .A1(n20583), .A2(n13189), .ZN(n11147) );
  NAND2_X1 U14471 ( .A1(n13189), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13371) );
  NAND2_X1 U14472 ( .A1(n20615), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13248) );
  NAND2_X1 U14473 ( .A1(n13371), .A2(n13248), .ZN(n13874) );
  NAND2_X1 U14474 ( .A1(n13197), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13199) );
  NAND2_X1 U14475 ( .A1(n13201), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13204) );
  INV_X1 U14476 ( .A(n13204), .ZN(n11148) );
  NAND2_X1 U14477 ( .A1(n11148), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13203) );
  NAND2_X1 U14478 ( .A1(n13210), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13211) );
  INV_X1 U14479 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n13219) );
  INV_X1 U14480 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16121) );
  INV_X1 U14481 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13233) );
  NAND2_X1 U14482 ( .A1(n13237), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13236) );
  INV_X1 U14483 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16600) );
  INV_X1 U14484 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11150) );
  NAND2_X1 U14485 ( .A1(n11149), .A2(n11150), .ZN(n11151) );
  NAND2_X1 U14486 ( .A1(n13241), .A2(n11151), .ZN(n15993) );
  INV_X2 U14487 ( .A(n16837), .ZN(n16810) );
  INV_X1 U14488 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20536) );
  NOR2_X1 U14489 ( .A1(n16810), .A2(n20536), .ZN(n11541) );
  AOI21_X1 U14490 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n11541), .ZN(n11152) );
  OAI21_X1 U14491 ( .B1(n16856), .B2(n15993), .A(n11152), .ZN(n11153) );
  OAI21_X1 U14492 ( .B1(n11548), .B2(n16863), .A(n11154), .ZN(n11155) );
  INV_X1 U14493 ( .A(n11155), .ZN(n11156) );
  NAND2_X1 U14494 ( .A1(n10449), .A2(n11156), .ZN(P2_U2988) );
  NAND2_X1 U14495 ( .A1(n9591), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11158) );
  INV_X1 U14496 ( .A(n11158), .ZN(n11159) );
  NAND2_X1 U14497 ( .A1(n11160), .A2(n11159), .ZN(n11161) );
  NAND2_X1 U14498 ( .A1(n11165), .A2(n11161), .ZN(n15978) );
  INV_X1 U14499 ( .A(n11162), .ZN(n11163) );
  NOR2_X1 U14500 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13286) );
  INV_X1 U14501 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11164) );
  NOR2_X1 U14502 ( .A1(n10902), .A2(n11164), .ZN(n11166) );
  INV_X1 U14503 ( .A(n11511), .ZN(n11168) );
  NAND2_X1 U14504 ( .A1(n11165), .A2(n11166), .ZN(n11167) );
  NAND2_X1 U14505 ( .A1(n11168), .A2(n11167), .ZN(n15962) );
  INV_X1 U14506 ( .A(n16579), .ZN(n11171) );
  INV_X1 U14507 ( .A(n11169), .ZN(n11170) );
  NAND2_X1 U14508 ( .A1(n9591), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11510) );
  INV_X1 U14509 ( .A(n11510), .ZN(n11172) );
  INV_X1 U14510 ( .A(n15950), .ZN(n11173) );
  INV_X1 U14511 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11504) );
  XNOR2_X1 U14512 ( .A(n11509), .B(n10482), .ZN(n16574) );
  NAND2_X1 U14513 ( .A1(n19875), .A2(n10578), .ZN(n11200) );
  NAND2_X1 U14514 ( .A1(n9593), .A2(n19875), .ZN(n11202) );
  NAND2_X1 U14515 ( .A1(n11174), .A2(n13271), .ZN(n11190) );
  NAND2_X1 U14516 ( .A1(n20617), .A2(n20620), .ZN(n11175) );
  MUX2_X1 U14517 ( .A(n13271), .B(n11175), .S(n11182), .Z(n11185) );
  INV_X1 U14518 ( .A(n13701), .ZN(n11183) );
  OAI21_X1 U14519 ( .B1(n10875), .B2(n11177), .A(n11193), .ZN(n11181) );
  OAI211_X1 U14520 ( .C1(n17491), .C2(n11179), .A(n14580), .B(n11178), .ZN(
        n11180) );
  OAI211_X1 U14521 ( .C1(n11183), .C2(n11182), .A(n11181), .B(n11180), .ZN(
        n11184) );
  NAND2_X1 U14522 ( .A1(n11185), .A2(n11184), .ZN(n11188) );
  INV_X1 U14523 ( .A(n11186), .ZN(n11187) );
  NAND2_X1 U14524 ( .A1(n11188), .A2(n11187), .ZN(n11189) );
  NAND2_X1 U14525 ( .A1(n11190), .A2(n11189), .ZN(n11195) );
  NAND2_X1 U14526 ( .A1(n20598), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11191) );
  AOI21_X1 U14527 ( .B1(n11193), .B2(n11192), .A(n11191), .ZN(n11194) );
  NAND2_X1 U14528 ( .A1(n11195), .A2(n11194), .ZN(n11199) );
  INV_X1 U14529 ( .A(n20598), .ZN(n11197) );
  NOR2_X1 U14530 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11196) );
  AOI21_X1 U14531 ( .B1(n13930), .B2(n11197), .A(n11196), .ZN(n11198) );
  MUX2_X1 U14532 ( .A(n11200), .B(n11202), .S(n14570), .Z(n11221) );
  NAND2_X1 U14533 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20613) );
  AND2_X1 U14534 ( .A1(n14574), .A2(n20613), .ZN(n11214) );
  MUX2_X1 U14535 ( .A(n19862), .B(n10050), .S(n17491), .Z(n11213) );
  INV_X1 U14536 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20475) );
  NOR2_X1 U14537 ( .A1(n20475), .A2(n20493), .ZN(n20485) );
  NOR2_X1 U14538 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20487) );
  INV_X1 U14539 ( .A(n20618), .ZN(n11215) );
  NAND3_X1 U14540 ( .A1(n14574), .A2(n20613), .A3(n11215), .ZN(n11211) );
  NAND2_X1 U14541 ( .A1(n11209), .A2(n19895), .ZN(n11201) );
  NAND2_X1 U14542 ( .A1(n11201), .A2(n13268), .ZN(n11246) );
  NAND2_X1 U14543 ( .A1(n11202), .A2(n14580), .ZN(n11203) );
  NAND2_X1 U14544 ( .A1(n11203), .A2(n19895), .ZN(n11204) );
  AOI21_X1 U14545 ( .B1(n11204), .B2(n11205), .A(n13700), .ZN(n11208) );
  NAND2_X1 U14546 ( .A1(n11287), .A2(n19875), .ZN(n11243) );
  NAND2_X1 U14547 ( .A1(n11243), .A2(n11205), .ZN(n11206) );
  NAND2_X1 U14548 ( .A1(n17493), .A2(n11206), .ZN(n11207) );
  INV_X1 U14549 ( .A(n11209), .ZN(n11210) );
  NAND2_X1 U14550 ( .A1(n11210), .A2(n10096), .ZN(n11244) );
  OAI211_X1 U14551 ( .C1(n11212), .C2(n11211), .A(n11241), .B(n11244), .ZN(
        n14216) );
  AOI21_X1 U14552 ( .B1(n11214), .B2(n11213), .A(n14216), .ZN(n11219) );
  AND2_X1 U14553 ( .A1(n11215), .A2(n20620), .ZN(n11216) );
  NAND2_X1 U14554 ( .A1(n14570), .A2(n11216), .ZN(n14220) );
  NAND2_X1 U14555 ( .A1(n19862), .A2(n20613), .ZN(n11217) );
  OR2_X1 U14556 ( .A1(n14220), .A2(n11217), .ZN(n11218) );
  NAND4_X1 U14557 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11222) );
  AND2_X2 U14558 ( .A1(n11222), .A2(n14601), .ZN(n11505) );
  NOR2_X1 U14559 ( .A1(n10858), .A2(n13271), .ZN(n20602) );
  NAND2_X1 U14560 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11227) );
  AOI22_X1 U14561 ( .A1(n10624), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11225) );
  NAND2_X1 U14562 ( .A1(n11223), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11224) );
  AND2_X1 U14563 ( .A1(n11225), .A2(n11224), .ZN(n11226) );
  INV_X1 U14564 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20539) );
  NAND2_X1 U14565 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11229) );
  AOI22_X1 U14566 ( .A1(n10624), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11228) );
  OAI211_X1 U14567 ( .C1(n20539), .C2(n13297), .A(n11229), .B(n11228), .ZN(
        n15958) );
  INV_X1 U14568 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20541) );
  NAND2_X1 U14569 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11231) );
  AOI22_X1 U14570 ( .A1(n10624), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11230) );
  OAI211_X1 U14571 ( .C1(n20541), .C2(n13297), .A(n11231), .B(n11230), .ZN(
        n11232) );
  NAND2_X1 U14572 ( .A1(n11235), .A2(n9593), .ZN(n11237) );
  NAND2_X1 U14573 ( .A1(n11237), .A2(n11236), .ZN(n11238) );
  NOR2_X1 U14574 ( .A1(n11239), .A2(n20620), .ZN(n11240) );
  NAND2_X1 U14575 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14790) );
  INV_X1 U14576 ( .A(n14790), .ZN(n14788) );
  NAND2_X1 U14577 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14788), .ZN(
        n14789) );
  INV_X1 U14578 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11242) );
  NAND2_X1 U14579 ( .A1(n11242), .A2(n14790), .ZN(n14787) );
  INV_X1 U14580 ( .A(n14787), .ZN(n11257) );
  AOI21_X1 U14581 ( .B1(n14786), .B2(n14789), .A(n11257), .ZN(n11255) );
  NAND3_X1 U14582 ( .A1(n11244), .A2(n19895), .A3(n11243), .ZN(n11245) );
  NAND2_X1 U14583 ( .A1(n11245), .A2(n20620), .ZN(n14548) );
  NAND2_X1 U14584 ( .A1(n14548), .A2(n11246), .ZN(n11248) );
  INV_X1 U14585 ( .A(n11247), .ZN(n20619) );
  AOI22_X1 U14586 ( .A1(n11248), .A2(n19869), .B1(n20619), .B2(n19875), .ZN(
        n11252) );
  NAND2_X1 U14587 ( .A1(n11249), .A2(n11247), .ZN(n11250) );
  NAND2_X1 U14588 ( .A1(n11250), .A2(n13700), .ZN(n11251) );
  INV_X1 U14589 ( .A(n11253), .ZN(n14203) );
  NAND2_X1 U14590 ( .A1(n14535), .A2(n14203), .ZN(n11254) );
  NAND2_X1 U14591 ( .A1(n11255), .A2(n11526), .ZN(n14646) );
  NOR2_X1 U14592 ( .A1(n17110), .A2(n16853), .ZN(n17111) );
  NAND2_X1 U14593 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17111), .ZN(
        n11256) );
  INV_X1 U14594 ( .A(n11267), .ZN(n14842) );
  NAND2_X1 U14595 ( .A1(n17031), .A2(n14842), .ZN(n16899) );
  AND2_X1 U14596 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11537) );
  INV_X1 U14597 ( .A(n11537), .ZN(n11502) );
  NOR2_X1 U14598 ( .A1(n16865), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16878) );
  NAND2_X1 U14599 ( .A1(n13164), .A2(n14789), .ZN(n11261) );
  NAND2_X1 U14600 ( .A1(n11258), .A2(n11257), .ZN(n11260) );
  INV_X1 U14601 ( .A(n11505), .ZN(n11259) );
  NAND2_X1 U14602 ( .A1(n11259), .A2(n16810), .ZN(n14785) );
  NAND2_X1 U14603 ( .A1(n17095), .A2(n17098), .ZN(n17097) );
  INV_X1 U14604 ( .A(n17097), .ZN(n17032) );
  INV_X1 U14605 ( .A(n17095), .ZN(n11263) );
  NAND3_X1 U14606 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n17111), .ZN(n11262) );
  OR2_X1 U14607 ( .A1(n11263), .A2(n11262), .ZN(n11264) );
  NAND2_X1 U14608 ( .A1(n17097), .A2(n11264), .ZN(n17081) );
  INV_X1 U14609 ( .A(n11265), .ZN(n17065) );
  NAND2_X1 U14610 ( .A1(n11526), .A2(n17065), .ZN(n11266) );
  NAND2_X1 U14611 ( .A1(n17081), .A2(n11266), .ZN(n17028) );
  NOR2_X1 U14612 ( .A1(n17028), .A2(n11267), .ZN(n14891) );
  INV_X1 U14613 ( .A(n11268), .ZN(n11269) );
  NAND2_X1 U14614 ( .A1(n14891), .A2(n11269), .ZN(n11270) );
  NAND2_X1 U14615 ( .A1(n11270), .A2(n17097), .ZN(n16901) );
  OAI21_X1 U14616 ( .B1(n11537), .B2(n17032), .A(n16901), .ZN(n16880) );
  OR2_X1 U14617 ( .A1(n16878), .A2(n16880), .ZN(n16868) );
  NOR2_X1 U14618 ( .A1(n16810), .A2(n20541), .ZN(n16569) );
  INV_X1 U14619 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16582) );
  AOI21_X1 U14620 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n11504), .A(
        n16582), .ZN(n11271) );
  AOI211_X1 U14621 ( .C1(n11504), .C2(n16582), .A(n11271), .B(n16865), .ZN(
        n11272) );
  AOI211_X1 U14622 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16868), .A(
        n16569), .B(n11272), .ZN(n11500) );
  NAND2_X1 U14623 ( .A1(n11297), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11276) );
  AOI21_X1 U14624 ( .B1(n17491), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11275) );
  INV_X1 U14625 ( .A(n19895), .ZN(n13706) );
  NAND2_X1 U14626 ( .A1(n13706), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11274) );
  NAND3_X1 U14627 ( .A1(n11276), .A2(n11275), .A3(n11274), .ZN(n13992) );
  NAND3_X1 U14628 ( .A1(n9593), .A2(n10902), .A3(n20607), .ZN(n11307) );
  INV_X1 U14629 ( .A(n11277), .ZN(n11281) );
  INV_X1 U14630 ( .A(n11288), .ZN(n11278) );
  OAI21_X1 U14631 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20607), .A(
        n11278), .ZN(n11280) );
  INV_X1 U14632 ( .A(n11287), .ZN(n13705) );
  AND2_X1 U14633 ( .A1(n11279), .A2(n20607), .ZN(n11299) );
  NAND2_X1 U14634 ( .A1(n13705), .A2(n11299), .ZN(n11295) );
  OAI211_X1 U14635 ( .C1(n11307), .C2(n11281), .A(n11280), .B(n11295), .ZN(
        n13991) );
  NAND2_X1 U14636 ( .A1(n13992), .A2(n13991), .ZN(n13993) );
  INV_X1 U14637 ( .A(n11297), .ZN(n11283) );
  INV_X1 U14638 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20494) );
  AND2_X2 U14639 ( .A1(n13706), .A2(n20607), .ZN(n11298) );
  AOI22_X1 U14640 ( .A1(n11298), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11299), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11282) );
  OAI21_X1 U14641 ( .B1(n11283), .B2(n20494), .A(n11282), .ZN(n11291) );
  XNOR2_X1 U14642 ( .A(n13993), .B(n11291), .ZN(n14051) );
  NAND2_X1 U14643 ( .A1(n9593), .A2(n20607), .ZN(n11285) );
  NAND2_X1 U14644 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11284) );
  AND2_X1 U14645 ( .A1(n11288), .A2(n11287), .ZN(n11289) );
  NOR2_X1 U14646 ( .A1(n11290), .A2(n11289), .ZN(n14050) );
  NAND2_X1 U14647 ( .A1(n14051), .A2(n14050), .ZN(n14049) );
  INV_X1 U14648 ( .A(n11291), .ZN(n11292) );
  NAND2_X1 U14649 ( .A1(n13993), .A2(n11292), .ZN(n11293) );
  NAND2_X1 U14650 ( .A1(n14049), .A2(n11293), .ZN(n11304) );
  NAND2_X1 U14651 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11294) );
  OAI211_X1 U14652 ( .C1(n11307), .C2(n11296), .A(n11295), .B(n11294), .ZN(
        n11302) );
  XNOR2_X1 U14653 ( .A(n11304), .B(n11302), .ZN(n14798) );
  NAND2_X1 U14654 ( .A1(n11297), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14655 ( .A1(n11298), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13732), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11300) );
  AND2_X1 U14656 ( .A1(n11301), .A2(n11300), .ZN(n14797) );
  INV_X1 U14657 ( .A(n11302), .ZN(n11303) );
  NAND2_X1 U14658 ( .A1(n11304), .A2(n11303), .ZN(n11305) );
  OAI22_X1 U14659 ( .A1(n11432), .A2(n14634), .B1(n20574), .B2(n20607), .ZN(
        n11306) );
  AOI21_X1 U14660 ( .B1(n11297), .B2(P2_REIP_REG_3__SCAN_IN), .A(n11306), .ZN(
        n11310) );
  AOI22_X1 U14661 ( .A1(n11462), .A2(n10880), .B1(n11298), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n11309) );
  INV_X1 U14662 ( .A(n14643), .ZN(n11311) );
  NAND2_X1 U14663 ( .A1(n11297), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14664 ( .A1(n11298), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13732), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U14665 ( .A1(n11462), .A2(n11312), .ZN(n11313) );
  NAND2_X1 U14666 ( .A1(n11317), .A2(n11316), .ZN(n16273) );
  NAND2_X1 U14667 ( .A1(n11297), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14668 ( .A1(n11298), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13732), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11320) );
  NAND2_X1 U14669 ( .A1(n11462), .A2(n11318), .ZN(n11319) );
  NAND2_X1 U14670 ( .A1(n11462), .A2(n11322), .ZN(n11323) );
  AOI22_X1 U14671 ( .A1(n11298), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13732), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11324) );
  OAI21_X1 U14672 ( .B1(n13734), .B2(n20503), .A(n11324), .ZN(n13983) );
  AOI21_X1 U14673 ( .B1(n13982), .B2(n13983), .A(n10481), .ZN(n11325) );
  INV_X1 U14674 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20505) );
  AOI22_X1 U14675 ( .A1(n11298), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13732), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11326) );
  OAI21_X1 U14676 ( .B1(n13734), .B2(n20505), .A(n11326), .ZN(n14001) );
  NAND2_X1 U14677 ( .A1(n11297), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14678 ( .A1(n11298), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13732), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14679 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14680 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14681 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14682 ( .A1(n11346), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11328) );
  NAND4_X1 U14683 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n11341) );
  AOI22_X1 U14684 ( .A1(n13534), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11339) );
  INV_X1 U14685 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11334) );
  NAND2_X1 U14686 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U14687 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11332) );
  OAI211_X1 U14688 ( .C1(n10727), .C2(n11334), .A(n11333), .B(n11332), .ZN(
        n11335) );
  INV_X1 U14689 ( .A(n11335), .ZN(n11338) );
  AOI22_X1 U14690 ( .A1(n13541), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11337) );
  NAND2_X1 U14691 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11336) );
  NAND4_X1 U14692 ( .A1(n11339), .A2(n11338), .A3(n11337), .A4(n11336), .ZN(
        n11340) );
  NAND2_X1 U14693 ( .A1(n11462), .A2(n14399), .ZN(n11342) );
  NAND2_X1 U14694 ( .A1(n11297), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14695 ( .A1(n11298), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13732), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14696 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11346), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14697 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10757), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14698 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14699 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11347) );
  NAND4_X1 U14700 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n11359) );
  AOI22_X1 U14701 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n13534), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11357) );
  NAND2_X1 U14702 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11352) );
  NAND2_X1 U14703 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11351) );
  OAI211_X1 U14704 ( .C1(n10727), .C2(n21605), .A(n11352), .B(n11351), .ZN(
        n11353) );
  INV_X1 U14705 ( .A(n11353), .ZN(n11356) );
  AOI22_X1 U14706 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13541), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U14707 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11354) );
  NAND4_X1 U14708 ( .A1(n11357), .A2(n11356), .A3(n11355), .A4(n11354), .ZN(
        n11358) );
  NAND2_X1 U14709 ( .A1(n11462), .A2(n14266), .ZN(n11360) );
  NAND2_X1 U14710 ( .A1(n11364), .A2(n11363), .ZN(n14078) );
  NAND2_X1 U14711 ( .A1(n11297), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14712 ( .A1(n11298), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14713 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10780), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14714 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13526), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14715 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14716 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n11346), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11365) );
  NAND4_X1 U14717 ( .A1(n11368), .A2(n11367), .A3(n11366), .A4(n11365), .ZN(
        n11378) );
  AOI22_X1 U14718 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n13534), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11376) );
  INV_X1 U14719 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11371) );
  NAND2_X1 U14720 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11370) );
  NAND2_X1 U14721 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11369) );
  OAI211_X1 U14722 ( .C1(n10727), .C2(n11371), .A(n11370), .B(n11369), .ZN(
        n11372) );
  INV_X1 U14723 ( .A(n11372), .ZN(n11375) );
  AOI22_X1 U14724 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13541), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11374) );
  NAND2_X1 U14725 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11373) );
  NAND4_X1 U14726 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11377) );
  NAND2_X1 U14727 ( .A1(n11462), .A2(n14410), .ZN(n11379) );
  INV_X1 U14728 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16746) );
  AOI22_X1 U14729 ( .A1(n11298), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14730 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n13528), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14731 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10757), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14732 ( .A1(n11346), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14733 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11382) );
  NAND4_X1 U14734 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11395) );
  AOI22_X1 U14735 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n13534), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11393) );
  NAND2_X1 U14736 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11387) );
  NAND2_X1 U14737 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11386) );
  OAI211_X1 U14738 ( .C1(n10727), .C2(n11388), .A(n11387), .B(n11386), .ZN(
        n11389) );
  INV_X1 U14739 ( .A(n11389), .ZN(n11392) );
  AOI22_X1 U14740 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13541), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11391) );
  NAND2_X1 U14741 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11390) );
  NAND4_X1 U14742 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n11394) );
  NAND2_X1 U14743 ( .A1(n11462), .A2(n14329), .ZN(n11396) );
  OAI211_X1 U14744 ( .C1(n13734), .C2(n16746), .A(n11397), .B(n11396), .ZN(
        n14195) );
  NAND2_X1 U14745 ( .A1(n11297), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14746 ( .A1(n11298), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14747 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10780), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14748 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13526), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14749 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U14750 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11346), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U14751 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11411) );
  AOI22_X1 U14752 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13534), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11409) );
  INV_X1 U14753 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11404) );
  NAND2_X1 U14754 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11403) );
  NAND2_X1 U14755 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11402) );
  OAI211_X1 U14756 ( .C1(n10727), .C2(n11404), .A(n11403), .B(n11402), .ZN(
        n11405) );
  INV_X1 U14757 ( .A(n11405), .ZN(n11408) );
  AOI22_X1 U14758 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13541), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11407) );
  NAND2_X1 U14759 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11406) );
  NAND4_X1 U14760 ( .A1(n11409), .A2(n11408), .A3(n11407), .A4(n11406), .ZN(
        n11410) );
  NAND2_X1 U14761 ( .A1(n11462), .A2(n14436), .ZN(n11412) );
  NAND2_X1 U14762 ( .A1(n11297), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14763 ( .A1(n11298), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14764 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10780), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14765 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14766 ( .A1(n11346), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14767 ( .A1(n10757), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11416) );
  NAND4_X1 U14768 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n11428) );
  AOI22_X1 U14769 ( .A1(n13534), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11426) );
  INV_X1 U14770 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13634) );
  NAND2_X1 U14771 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11421) );
  NAND2_X1 U14772 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11420) );
  OAI211_X1 U14773 ( .C1(n10727), .C2(n13634), .A(n11421), .B(n11420), .ZN(
        n11422) );
  INV_X1 U14774 ( .A(n11422), .ZN(n11425) );
  AOI22_X1 U14775 ( .A1(n13541), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11424) );
  NAND2_X1 U14776 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11423) );
  NAND4_X1 U14777 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(
        n11427) );
  NAND2_X1 U14778 ( .A1(n11462), .A2(n14442), .ZN(n11429) );
  INV_X1 U14779 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n16706) );
  INV_X2 U14780 ( .A(n11432), .ZN(n13732) );
  AOI22_X1 U14781 ( .A1(n11298), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14782 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14783 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14784 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14785 ( .A1(n11346), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U14786 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n11445) );
  AOI22_X1 U14787 ( .A1(n13534), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11443) );
  INV_X1 U14788 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13482) );
  NAND2_X1 U14789 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11438) );
  NAND2_X1 U14790 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11437) );
  OAI211_X1 U14791 ( .C1(n10727), .C2(n13482), .A(n11438), .B(n11437), .ZN(
        n11439) );
  INV_X1 U14792 ( .A(n11439), .ZN(n11442) );
  AOI22_X1 U14793 ( .A1(n13541), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U14794 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11440) );
  NAND4_X1 U14795 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(
        n11444) );
  NAND2_X1 U14796 ( .A1(n11462), .A2(n14610), .ZN(n11446) );
  OAI211_X1 U14797 ( .C1(n13734), .C2(n16706), .A(n11447), .B(n11446), .ZN(
        n16157) );
  INV_X1 U14798 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n16692) );
  AOI22_X1 U14799 ( .A1(n11298), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14800 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14801 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n11346), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14802 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14803 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n11327), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11448) );
  NAND4_X1 U14804 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11461) );
  AOI22_X1 U14805 ( .A1(n13534), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11459) );
  INV_X1 U14806 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U14807 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11453) );
  NAND2_X1 U14808 ( .A1(n13540), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11452) );
  OAI211_X1 U14809 ( .C1(n10727), .C2(n11454), .A(n11453), .B(n11452), .ZN(
        n11455) );
  INV_X1 U14810 ( .A(n11455), .ZN(n11458) );
  AOI22_X1 U14811 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13541), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U14812 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11456) );
  NAND4_X1 U14813 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11460) );
  NAND2_X1 U14814 ( .A1(n11462), .A2(n14659), .ZN(n11463) );
  OAI211_X1 U14815 ( .C1(n13734), .C2(n16692), .A(n11464), .B(n11463), .ZN(
        n16154) );
  NAND2_X1 U14816 ( .A1(n11297), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U14817 ( .A1(n11298), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11465) );
  OR2_X2 U14818 ( .A1(n16131), .A2(n16132), .ZN(n16129) );
  NAND2_X1 U14819 ( .A1(n11297), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14820 ( .A1(n11298), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11467) );
  NOR2_X4 U14821 ( .A1(n16129), .A2(n13146), .ZN(n16103) );
  NAND2_X1 U14822 ( .A1(n11297), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14823 ( .A1(n11298), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11469) );
  AND2_X1 U14824 ( .A1(n11470), .A2(n11469), .ZN(n16062) );
  INV_X1 U14825 ( .A(n16062), .ZN(n11479) );
  NAND2_X1 U14826 ( .A1(n11297), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14827 ( .A1(n11298), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11471) );
  AND2_X1 U14828 ( .A1(n11472), .A2(n11471), .ZN(n14890) );
  INV_X1 U14829 ( .A(n14890), .ZN(n11478) );
  NAND2_X1 U14830 ( .A1(n11297), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14831 ( .A1(n11298), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11473) );
  AND2_X1 U14832 ( .A1(n11474), .A2(n11473), .ZN(n14827) );
  INV_X1 U14833 ( .A(n14827), .ZN(n11477) );
  INV_X1 U14834 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20523) );
  AOI22_X1 U14835 ( .A1(n11298), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11475) );
  OAI21_X1 U14836 ( .B1(n13734), .B2(n20523), .A(n11475), .ZN(n16087) );
  INV_X1 U14837 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20521) );
  AOI22_X1 U14838 ( .A1(n11298), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11476) );
  OAI21_X1 U14839 ( .B1(n13734), .B2(n20521), .A(n11476), .ZN(n16102) );
  AND2_X1 U14840 ( .A1(n16087), .A2(n16102), .ZN(n14824) );
  INV_X1 U14841 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20531) );
  AOI22_X1 U14842 ( .A1(n11298), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11481) );
  OAI21_X1 U14843 ( .B1(n13734), .B2(n20531), .A(n11481), .ZN(n16046) );
  NAND2_X1 U14844 ( .A1(n11297), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14845 ( .A1(n11298), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11482) );
  AND2_X1 U14846 ( .A1(n11483), .A2(n11482), .ZN(n16024) );
  NAND2_X1 U14847 ( .A1(n11297), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14848 ( .A1(n11298), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14849 ( .A1(n11298), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11486) );
  OAI21_X1 U14850 ( .B1(n13734), .B2(n20536), .A(n11486), .ZN(n11543) );
  AND2_X2 U14851 ( .A1(n16015), .A2(n11543), .ZN(n15973) );
  INV_X1 U14852 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20538) );
  AOI22_X1 U14853 ( .A1(n11298), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11487) );
  OAI21_X1 U14854 ( .B1(n13734), .B2(n20538), .A(n11487), .ZN(n15972) );
  NAND2_X1 U14855 ( .A1(n11297), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14856 ( .A1(n11298), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11488) );
  AND2_X1 U14857 ( .A1(n11489), .A2(n11488), .ZN(n15968) );
  NAND2_X1 U14858 ( .A1(n11297), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14859 ( .A1(n11298), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11490) );
  INV_X1 U14860 ( .A(n11517), .ZN(n11492) );
  NAND2_X1 U14861 ( .A1(n11494), .A2(n17491), .ZN(n11497) );
  NAND2_X1 U14862 ( .A1(n9736), .A2(n11496), .ZN(n14571) );
  NAND2_X1 U14863 ( .A1(n11497), .A2(n14571), .ZN(n11498) );
  NAND2_X1 U14864 ( .A1(n15955), .A2(n17121), .ZN(n11499) );
  OAI211_X1 U14865 ( .C1(n16571), .C2(n17116), .A(n11500), .B(n11499), .ZN(
        n11501) );
  INV_X1 U14866 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16864) );
  INV_X1 U14867 ( .A(n13278), .ZN(n11508) );
  OAI21_X1 U14868 ( .B1(n11509), .B2(n13280), .A(n11508), .ZN(n11516) );
  NAND2_X1 U14869 ( .A1(n9590), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11512) );
  INV_X1 U14870 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13739) );
  NOR2_X1 U14871 ( .A1(n11514), .A2(n10461), .ZN(n13279) );
  NOR2_X1 U14872 ( .A1(n13279), .A2(n13281), .ZN(n11515) );
  XNOR2_X1 U14873 ( .A(n11516), .B(n11515), .ZN(n14772) );
  INV_X1 U14874 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20546) );
  AOI22_X1 U14875 ( .A1(n11298), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11518) );
  OAI21_X1 U14876 ( .B1(n13734), .B2(n20546), .A(n11518), .ZN(n11519) );
  INV_X1 U14877 ( .A(n13707), .ZN(n11522) );
  NAND2_X1 U14878 ( .A1(n9548), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11525) );
  AOI22_X1 U14879 ( .A1(n10624), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11524) );
  OAI211_X1 U14880 ( .C1(n20546), .C2(n13297), .A(n11525), .B(n11524), .ZN(
        n13295) );
  NAND3_X1 U14881 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13738) );
  AOI21_X1 U14882 ( .B1(n11526), .B2(n13738), .A(n16880), .ZN(n13737) );
  INV_X1 U14883 ( .A(n13737), .ZN(n11528) );
  NOR2_X1 U14884 ( .A1(n16810), .A2(n20546), .ZN(n14765) );
  NOR3_X1 U14885 ( .A1(n16865), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n13738), .ZN(n11527) );
  AOI211_X1 U14886 ( .C1(n11528), .C2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14765), .B(n11527), .ZN(n11529) );
  OAI21_X1 U14887 ( .B1(n14806), .B2(n17116), .A(n11529), .ZN(n11530) );
  INV_X1 U14888 ( .A(n11530), .ZN(n11531) );
  OAI21_X1 U14889 ( .B1(n14764), .B2(n17124), .A(n11531), .ZN(n11532) );
  OAI211_X1 U14890 ( .C1(n14772), .C2(n17139), .A(n11534), .B(n11533), .ZN(
        P2_U3016) );
  INV_X1 U14891 ( .A(n16901), .ZN(n16890) );
  AOI211_X1 U14892 ( .C1(n11539), .C2(n11538), .A(n11537), .B(n16887), .ZN(
        n11540) );
  AOI211_X1 U14893 ( .C1(n16890), .C2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11541), .B(n11540), .ZN(n11542) );
  OAI21_X1 U14894 ( .B1(n16394), .B2(n17116), .A(n11542), .ZN(n11546) );
  INV_X1 U14895 ( .A(n11543), .ZN(n11545) );
  INV_X1 U14896 ( .A(n16015), .ZN(n11544) );
  AOI21_X1 U14897 ( .B1(n11545), .B2(n11544), .A(n15973), .ZN(n16469) );
  INV_X1 U14898 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18354) );
  NAND2_X1 U14899 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11550) );
  NAND2_X1 U14900 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11549) );
  OAI211_X1 U14901 ( .C1(n18218), .C2(n18354), .A(n11550), .B(n11549), .ZN(
        n11551) );
  INV_X1 U14902 ( .A(n11551), .ZN(n11556) );
  AOI22_X1 U14903 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11555) );
  AND2_X2 U14904 ( .A1(n11557), .A2(n17351), .ZN(n17461) );
  AOI22_X1 U14905 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11554) );
  NAND2_X1 U14906 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11553) );
  AOI22_X1 U14907 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11568) );
  AND2_X2 U14908 ( .A1(n11558), .A2(n11559), .ZN(n18330) );
  NAND2_X2 U14909 ( .A1(n11558), .A2(n11562), .ZN(n17408) );
  AOI22_X1 U14910 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14911 ( .A1(n11649), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11566) );
  AND2_X4 U14912 ( .A1(n11564), .A2(n11563), .ZN(n18170) );
  AOI22_X1 U14913 ( .A1(n11628), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11565) );
  INV_X1 U14914 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18228) );
  NAND2_X1 U14915 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11570) );
  NAND2_X1 U14916 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11569) );
  OAI211_X1 U14917 ( .C1(n18218), .C2(n18228), .A(n11570), .B(n11569), .ZN(
        n11571) );
  INV_X1 U14918 ( .A(n11571), .ZN(n11575) );
  AOI22_X1 U14919 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14920 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11573) );
  NAND2_X1 U14921 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11572) );
  NAND4_X1 U14922 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11581) );
  AOI22_X1 U14923 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14924 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14925 ( .A1(n11649), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14926 ( .A1(n11628), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11576) );
  NAND4_X1 U14927 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11580) );
  NAND2_X1 U14928 ( .A1(n14512), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14277) );
  INV_X1 U14929 ( .A(n14277), .ZN(n14144) );
  NAND2_X1 U14930 ( .A1(n14145), .A2(n14144), .ZN(n11583) );
  INV_X1 U14931 ( .A(n14666), .ZN(n11906) );
  NAND2_X1 U14932 ( .A1(n11906), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11582) );
  NAND2_X1 U14933 ( .A1(n11583), .A2(n11582), .ZN(n14093) );
  INV_X1 U14934 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17379) );
  NAND2_X1 U14935 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11585) );
  NAND2_X1 U14936 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11584) );
  OAI211_X1 U14937 ( .C1(n18218), .C2(n17379), .A(n11585), .B(n11584), .ZN(
        n11586) );
  AOI22_X1 U14938 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14939 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11588) );
  NAND2_X1 U14940 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11587) );
  AOI22_X1 U14941 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11649), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14942 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11590) );
  NAND4_X1 U14943 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n11594) );
  XNOR2_X1 U14944 ( .A(n11595), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14092) );
  NAND2_X1 U14945 ( .A1(n14093), .A2(n14092), .ZN(n11598) );
  INV_X1 U14946 ( .A(n11595), .ZN(n11596) );
  NAND2_X1 U14947 ( .A1(n11596), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11597) );
  INV_X1 U14948 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17432) );
  NAND2_X1 U14949 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U14950 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11599) );
  OAI211_X1 U14951 ( .C1(n18218), .C2(n17432), .A(n11600), .B(n11599), .ZN(
        n11601) );
  INV_X1 U14952 ( .A(n11601), .ZN(n11605) );
  AOI22_X1 U14953 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14954 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11603) );
  NAND2_X1 U14955 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11602) );
  NAND4_X1 U14956 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11612) );
  AOI22_X1 U14957 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14958 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14959 ( .A1(n11649), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14960 ( .A1(n11628), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11607) );
  NAND4_X1 U14961 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11611) );
  INV_X1 U14962 ( .A(n14509), .ZN(n11910) );
  XNOR2_X1 U14963 ( .A(n11617), .B(n11910), .ZN(n11613) );
  INV_X1 U14964 ( .A(n11613), .ZN(n11614) );
  NAND2_X1 U14965 ( .A1(n11615), .A2(n11614), .ZN(n11616) );
  INV_X1 U14966 ( .A(n11617), .ZN(n11618) );
  NAND2_X1 U14967 ( .A1(n11618), .A2(n14509), .ZN(n11640) );
  INV_X1 U14968 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11621) );
  NAND2_X1 U14969 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11620) );
  NAND2_X1 U14970 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11619) );
  OAI211_X1 U14971 ( .C1(n18218), .C2(n11621), .A(n11620), .B(n11619), .ZN(
        n11622) );
  INV_X1 U14972 ( .A(n11622), .ZN(n11627) );
  AOI22_X1 U14973 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14974 ( .A1(n11784), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U14975 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11624) );
  NAND4_X1 U14976 ( .A1(n11627), .A2(n11626), .A3(n11625), .A4(n11624), .ZN(
        n11634) );
  AOI22_X1 U14977 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14978 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14979 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9559), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14980 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11629) );
  NAND4_X1 U14981 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11633) );
  INV_X1 U14982 ( .A(n18529), .ZN(n11635) );
  XNOR2_X1 U14983 ( .A(n11640), .B(n11635), .ZN(n11636) );
  XNOR2_X1 U14984 ( .A(n11636), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13810) );
  INV_X1 U14985 ( .A(n11636), .ZN(n11637) );
  NAND2_X1 U14986 ( .A1(n11637), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11638) );
  INV_X1 U14987 ( .A(n11640), .ZN(n11641) );
  NAND2_X1 U14988 ( .A1(n11641), .A2(n18529), .ZN(n11660) );
  INV_X1 U14989 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17471) );
  NAND2_X1 U14990 ( .A1(n9556), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11643) );
  NAND2_X1 U14991 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11642) );
  OAI211_X1 U14992 ( .C1(n18218), .C2(n17471), .A(n11643), .B(n11642), .ZN(
        n11644) );
  INV_X1 U14993 ( .A(n11644), .ZN(n11648) );
  AOI22_X1 U14994 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14995 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11646) );
  NAND2_X1 U14996 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11645) );
  NAND4_X1 U14997 ( .A1(n11648), .A2(n11647), .A3(n11646), .A4(n11645), .ZN(
        n11655) );
  AOI22_X1 U14998 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14999 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U15000 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11651) );
  INV_X1 U15001 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n21563) );
  AOI22_X1 U15002 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11650) );
  NAND4_X1 U15003 ( .A1(n11653), .A2(n11652), .A3(n11651), .A4(n11650), .ZN(
        n11654) );
  XNOR2_X1 U15004 ( .A(n11660), .B(n18524), .ZN(n11656) );
  INV_X1 U15005 ( .A(n11656), .ZN(n11657) );
  NAND2_X1 U15006 ( .A1(n11658), .A2(n11657), .ZN(n11659) );
  INV_X1 U15007 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11663) );
  NAND2_X1 U15008 ( .A1(n11606), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11662) );
  NAND2_X1 U15009 ( .A1(n18170), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11661) );
  OAI211_X1 U15010 ( .C1(n18218), .C2(n11663), .A(n11662), .B(n11661), .ZN(
        n11664) );
  INV_X1 U15011 ( .A(n11664), .ZN(n11668) );
  AOI22_X1 U15012 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U15013 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9559), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U15014 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11665) );
  NAND4_X1 U15015 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n11674) );
  AOI22_X1 U15016 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U15017 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U15018 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U15019 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U15020 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  XNOR2_X1 U15021 ( .A(n11675), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14170) );
  INV_X1 U15022 ( .A(n11675), .ZN(n11676) );
  NAND2_X1 U15023 ( .A1(n11676), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11677) );
  INV_X1 U15024 ( .A(n11679), .ZN(n11680) );
  INV_X1 U15025 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18255) );
  NAND2_X1 U15026 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11682) );
  NAND2_X1 U15027 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11681) );
  OAI211_X1 U15028 ( .C1(n18218), .C2(n18255), .A(n11682), .B(n11681), .ZN(
        n11683) );
  INV_X1 U15029 ( .A(n11683), .ZN(n11688) );
  AOI22_X1 U15030 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U15031 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11686) );
  NAND2_X1 U15032 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11685) );
  NAND4_X1 U15033 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n11694) );
  AOI22_X1 U15034 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U15035 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11691) );
  INV_X1 U15036 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n21652) );
  AOI22_X1 U15037 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U15038 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U15039 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11693) );
  NAND2_X1 U15040 ( .A1(n11695), .A2(n18515), .ZN(n11696) );
  NAND2_X1 U15041 ( .A1(n18712), .A2(n11696), .ZN(n11697) );
  XNOR2_X1 U15042 ( .A(n11699), .B(n11697), .ZN(n18854) );
  NAND2_X1 U15043 ( .A1(n18854), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11701) );
  INV_X1 U15044 ( .A(n11697), .ZN(n11698) );
  NAND2_X1 U15045 ( .A1(n11699), .A2(n11698), .ZN(n11700) );
  NAND2_X1 U15046 ( .A1(n11701), .A2(n11700), .ZN(n11707) );
  INV_X1 U15047 ( .A(n11707), .ZN(n11702) );
  NOR2_X1 U15048 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18843) );
  INV_X1 U15049 ( .A(n18843), .ZN(n17224) );
  NOR2_X1 U15050 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11703) );
  INV_X1 U15051 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11705) );
  INV_X1 U15052 ( .A(n18788), .ZN(n11706) );
  INV_X1 U15053 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18997) );
  INV_X1 U15054 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n19035) );
  INV_X1 U15055 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n19102) );
  NOR2_X1 U15056 ( .A1(n19102), .A2(n19088), .ZN(n17227) );
  NAND2_X1 U15057 ( .A1(n17227), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19060) );
  NOR2_X1 U15058 ( .A1(n19060), .A2(n11705), .ZN(n19021) );
  NAND2_X1 U15059 ( .A1(n19021), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n19024) );
  NAND2_X1 U15060 ( .A1(n10316), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11708) );
  INV_X1 U15061 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18979) );
  NAND2_X1 U15062 ( .A1(n18766), .A2(n18979), .ZN(n11709) );
  AND2_X1 U15063 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18952) );
  AND2_X1 U15064 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11710) );
  AND2_X1 U15065 ( .A1(n18952), .A2(n11710), .ZN(n11718) );
  NAND2_X1 U15066 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18973) );
  INV_X1 U15067 ( .A(n18973), .ZN(n11711) );
  AND2_X1 U15068 ( .A1(n11718), .A2(n11711), .ZN(n18937) );
  NAND2_X1 U15069 ( .A1(n18937), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17339) );
  INV_X1 U15070 ( .A(n17339), .ZN(n11712) );
  NAND2_X1 U15071 ( .A1(n11712), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18669) );
  INV_X1 U15072 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11713) );
  NAND2_X1 U15073 ( .A1(n18712), .A2(n11713), .ZN(n18754) );
  INV_X1 U15074 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18968) );
  INV_X1 U15075 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18935) );
  NAND2_X1 U15076 ( .A1(n18968), .A2(n18935), .ZN(n11714) );
  NOR2_X1 U15077 ( .A1(n18754), .A2(n11714), .ZN(n18711) );
  INV_X1 U15078 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18716) );
  INV_X1 U15079 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18921) );
  INV_X1 U15080 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18692) );
  NAND4_X1 U15081 ( .A1(n18711), .A2(n18716), .A3(n18921), .A4(n18692), .ZN(
        n11715) );
  AND2_X1 U15082 ( .A1(n11718), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11719) );
  NAND2_X1 U15083 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17309) );
  INV_X1 U15084 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17316) );
  INV_X1 U15085 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17300) );
  NAND2_X1 U15086 ( .A1(n11722), .A2(n10316), .ZN(n17283) );
  AND2_X1 U15087 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17290) );
  NAND2_X1 U15088 ( .A1(n17290), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14877) );
  NAND2_X1 U15089 ( .A1(n11724), .A2(n11723), .ZN(n11725) );
  NAND2_X1 U15090 ( .A1(n14720), .A2(n11725), .ZN(n11726) );
  XNOR2_X1 U15091 ( .A(n11726), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14886) );
  INV_X1 U15092 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11730) );
  NAND2_X1 U15093 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11729) );
  NAND2_X1 U15094 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11728) );
  OAI211_X1 U15095 ( .C1(n18218), .C2(n11730), .A(n11729), .B(n11728), .ZN(
        n11731) );
  AOI22_X1 U15096 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U15097 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11733) );
  NAND2_X1 U15098 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11732) );
  AOI22_X1 U15099 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11649), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11739) );
  INV_X2 U15100 ( .A(n18256), .ZN(n11784) );
  AOI22_X1 U15101 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U15102 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U15103 ( .A1(n11628), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11736) );
  INV_X1 U15104 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18062) );
  NAND2_X1 U15105 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11741) );
  NAND2_X1 U15106 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11740) );
  OAI211_X1 U15107 ( .C1(n18218), .C2(n18062), .A(n11741), .B(n11740), .ZN(
        n11742) );
  INV_X1 U15108 ( .A(n11742), .ZN(n11746) );
  AOI22_X1 U15109 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U15110 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11744) );
  NAND2_X1 U15111 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11743) );
  NAND4_X1 U15112 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n11752) );
  AOI22_X1 U15113 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U15114 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U15115 ( .A1(n11649), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U15116 ( .A1(n11628), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11747) );
  NAND4_X1 U15117 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11751) );
  INV_X1 U15118 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18134) );
  NAND2_X1 U15119 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11754) );
  NAND2_X1 U15120 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11753) );
  OAI211_X1 U15121 ( .C1(n18218), .C2(n18134), .A(n11754), .B(n11753), .ZN(
        n11755) );
  INV_X1 U15122 ( .A(n11755), .ZN(n11759) );
  AOI22_X1 U15123 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U15124 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U15125 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11756) );
  AOI22_X1 U15126 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U15127 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U15128 ( .A1(n11649), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U15129 ( .A1(n11628), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U15130 ( .A1(n19166), .A2(n19162), .ZN(n11936) );
  INV_X1 U15131 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18188) );
  NAND2_X1 U15132 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11765) );
  NAND2_X1 U15133 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11764) );
  OAI211_X1 U15134 ( .C1(n18218), .C2(n18188), .A(n11765), .B(n11764), .ZN(
        n11766) );
  INV_X1 U15135 ( .A(n11766), .ZN(n11770) );
  AOI22_X1 U15136 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U15137 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11768) );
  NAND2_X1 U15138 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11767) );
  NAND4_X1 U15139 ( .A1(n11770), .A2(n11769), .A3(n11768), .A4(n11767), .ZN(
        n11776) );
  AOI22_X1 U15140 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U15141 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U15142 ( .A1(n11649), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U15143 ( .A1(n11628), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11771) );
  NAND4_X1 U15144 ( .A1(n11774), .A2(n11773), .A3(n11772), .A4(n11771), .ZN(
        n11775) );
  INV_X1 U15145 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18252) );
  NAND2_X1 U15146 ( .A1(n18294), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U15147 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11777) );
  OAI211_X1 U15148 ( .C1(n18218), .C2(n18252), .A(n11778), .B(n11777), .ZN(
        n11779) );
  INV_X1 U15149 ( .A(n11779), .ZN(n11783) );
  AOI22_X1 U15150 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18054), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U15151 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17461), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11781) );
  NAND2_X1 U15152 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11780) );
  NAND4_X1 U15153 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11790) );
  AOI22_X1 U15154 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U15155 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U15156 ( .A1(n9582), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U15157 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11785) );
  NAND4_X1 U15158 ( .A1(n11788), .A2(n11787), .A3(n11786), .A4(n11785), .ZN(
        n11789) );
  INV_X1 U15159 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11793) );
  NAND2_X1 U15160 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11792) );
  NAND2_X1 U15161 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11791) );
  OAI211_X1 U15162 ( .C1(n18218), .C2(n11793), .A(n11792), .B(n11791), .ZN(
        n11794) );
  INV_X1 U15163 ( .A(n11794), .ZN(n11798) );
  AOI22_X1 U15164 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17450), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U15165 ( .A1(n11784), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U15166 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11795) );
  NAND4_X1 U15167 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11805) );
  AOI22_X1 U15168 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9556), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U15169 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U15170 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9559), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U15171 ( .A1(n18349), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11800) );
  NAND4_X1 U15172 ( .A1(n11803), .A2(n11802), .A3(n11801), .A4(n11800), .ZN(
        n11804) );
  INV_X1 U15173 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17399) );
  NAND2_X1 U15174 ( .A1(n9556), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11807) );
  NAND2_X1 U15175 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11806) );
  OAI211_X1 U15176 ( .C1(n18218), .C2(n17399), .A(n11807), .B(n11806), .ZN(
        n11808) );
  AOI22_X1 U15177 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U15178 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U15179 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11809) );
  AOI22_X1 U15180 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U15181 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U15182 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U15183 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U15184 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U15185 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U15186 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11817) );
  NAND2_X1 U15187 ( .A1(n11784), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U15188 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11823) );
  NAND2_X1 U15189 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11822) );
  NAND2_X1 U15190 ( .A1(n9556), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11821) );
  NAND2_X1 U15191 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11820) );
  NAND2_X1 U15192 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U15193 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11826) );
  NAND2_X1 U15194 ( .A1(n11684), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11825) );
  NAND2_X1 U15195 ( .A1(n18349), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11824) );
  NAND2_X1 U15196 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11829) );
  NAND2_X1 U15197 ( .A1(n11606), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11828) );
  OAI211_X1 U15198 ( .C1(n18218), .C2(n18207), .A(n11829), .B(n11828), .ZN(
        n11830) );
  INV_X1 U15199 ( .A(n11830), .ZN(n11831) );
  NAND2_X1 U15200 ( .A1(n19140), .A2(n19736), .ZN(n11935) );
  OAI21_X1 U15201 ( .B1(n18396), .B2(n19157), .A(n11935), .ZN(n11835) );
  NOR2_X1 U15202 ( .A1(n11946), .A2(n11835), .ZN(n11894) );
  NOR2_X1 U15203 ( .A1(n11836), .A2(n11846), .ZN(n11840) );
  INV_X1 U15204 ( .A(n19153), .ZN(n11837) );
  NAND2_X1 U15205 ( .A1(n19157), .A2(n14508), .ZN(n11838) );
  OAI211_X1 U15206 ( .C1(n19157), .C2(n11840), .A(n11839), .B(n11838), .ZN(
        n11842) );
  AOI21_X1 U15207 ( .B1(n9695), .B2(n11935), .A(n11846), .ZN(n11841) );
  NOR2_X1 U15208 ( .A1(n11842), .A2(n11841), .ZN(n11845) );
  NAND2_X1 U15209 ( .A1(n11843), .A2(n19140), .ZN(n11844) );
  NAND2_X1 U15210 ( .A1(n11894), .A2(n11943), .ZN(n11851) );
  INV_X1 U15211 ( .A(n14508), .ZN(n11848) );
  NAND2_X1 U15212 ( .A1(n19171), .A2(n11848), .ZN(n11849) );
  NAND3_X1 U15213 ( .A1(n18578), .A2(n18538), .A3(n11849), .ZN(n11939) );
  INV_X1 U15214 ( .A(n11939), .ZN(n11850) );
  AOI21_X1 U15215 ( .B1(n11851), .B2(n17657), .A(n11850), .ZN(n14025) );
  AND2_X1 U15216 ( .A1(n9695), .A2(n19736), .ZN(n11870) );
  INV_X1 U15217 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19647) );
  NAND2_X2 U15218 ( .A1(n19749), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19708) );
  OAI211_X1 U15219 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19647), .B(n19708), .ZN(n19641) );
  OAI21_X1 U15220 ( .B1(n9695), .B2(n19736), .A(n19641), .ZN(n11852) );
  NAND2_X1 U15221 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19617) );
  OAI21_X1 U15222 ( .B1(n11870), .B2(n11852), .A(n19617), .ZN(n17654) );
  MUX2_X1 U15223 ( .A(n11853), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11882) );
  NAND2_X1 U15224 ( .A1(n11882), .A2(n11864), .ZN(n11855) );
  NAND2_X1 U15225 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n11853), .ZN(
        n11854) );
  NAND2_X1 U15226 ( .A1(n11855), .A2(n11854), .ZN(n11868) );
  NAND2_X1 U15227 ( .A1(n17346), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11857) );
  NAND2_X1 U15228 ( .A1(n11868), .A2(n11867), .ZN(n11858) );
  NAND2_X1 U15229 ( .A1(n11858), .A2(n21538), .ZN(n11860) );
  OAI22_X1 U15230 ( .A1(n11860), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n11859), .ZN(n11876) );
  NAND2_X1 U15231 ( .A1(n11876), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11863) );
  NAND2_X1 U15232 ( .A1(n11860), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11877) );
  AND2_X1 U15233 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19583), .ZN(
        n11861) );
  NAND2_X1 U15234 ( .A1(n11877), .A2(n11861), .ZN(n11862) );
  NAND2_X1 U15235 ( .A1(n11863), .A2(n11862), .ZN(n11872) );
  INV_X1 U15236 ( .A(n11864), .ZN(n11873) );
  OAI21_X1 U15237 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11865), .A(
        n11873), .ZN(n11866) );
  NOR2_X1 U15238 ( .A1(n11872), .A2(n11866), .ZN(n11883) );
  XNOR2_X1 U15239 ( .A(n11868), .B(n11867), .ZN(n11871) );
  INV_X1 U15240 ( .A(n11871), .ZN(n11869) );
  AND2_X1 U15241 ( .A1(n11883), .A2(n11869), .ZN(n14275) );
  NAND2_X1 U15242 ( .A1(n11870), .A2(n19166), .ZN(n11892) );
  OAI22_X1 U15243 ( .A1(n17654), .A2(n11888), .B1(n14275), .B2(n11892), .ZN(
        n11889) );
  INV_X1 U15244 ( .A(n11885), .ZN(n11875) );
  XNOR2_X1 U15245 ( .A(n11882), .B(n11873), .ZN(n11874) );
  NAND2_X1 U15246 ( .A1(n11875), .A2(n11874), .ZN(n11881) );
  INV_X1 U15247 ( .A(n11876), .ZN(n11880) );
  NAND2_X1 U15248 ( .A1(n11877), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11879) );
  NOR2_X1 U15249 ( .A1(n19583), .A2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11878) );
  AOI21_X1 U15250 ( .B1(n11880), .B2(n11879), .A(n11878), .ZN(n11884) );
  NAND2_X1 U15251 ( .A1(n11883), .A2(n11882), .ZN(n11887) );
  AND2_X1 U15252 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  AOI22_X1 U15253 ( .A1(n11889), .A2(n19589), .B1(n19592), .B2(n11888), .ZN(
        n11890) );
  NAND2_X1 U15254 ( .A1(n14025), .A2(n11890), .ZN(n11891) );
  INV_X1 U15255 ( .A(n11892), .ZN(n11893) );
  NAND2_X1 U15256 ( .A1(n11904), .A2(n11898), .ZN(n11914) );
  AND2_X1 U15257 ( .A1(n14509), .A2(n18529), .ZN(n11895) );
  NAND2_X1 U15258 ( .A1(n11916), .A2(n11896), .ZN(n11921) );
  NOR2_X1 U15259 ( .A1(n11897), .A2(n11921), .ZN(n11925) );
  NAND2_X1 U15260 ( .A1(n11925), .A2(n17282), .ZN(n11926) );
  XNOR2_X1 U15261 ( .A(n11916), .B(n18524), .ZN(n11920) );
  XNOR2_X1 U15262 ( .A(n11904), .B(n11898), .ZN(n11900) );
  OAI21_X1 U15263 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n11900), .A(
        n11899), .ZN(n14085) );
  INV_X1 U15264 ( .A(n14512), .ZN(n11901) );
  INV_X1 U15265 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19020) );
  NAND2_X1 U15266 ( .A1(n11901), .A2(n19020), .ZN(n14278) );
  NAND2_X1 U15267 ( .A1(n14278), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11907) );
  INV_X1 U15268 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11902) );
  NAND2_X1 U15269 ( .A1(n19020), .A2(n11902), .ZN(n11903) );
  NAND2_X1 U15270 ( .A1(n11904), .A2(n11903), .ZN(n11905) );
  AOI21_X1 U15271 ( .B1(n11907), .B2(n11906), .A(n11905), .ZN(n14084) );
  INV_X1 U15272 ( .A(n14084), .ZN(n11908) );
  NOR2_X1 U15273 ( .A1(n14085), .A2(n11908), .ZN(n11909) );
  XNOR2_X1 U15274 ( .A(n11914), .B(n11910), .ZN(n11912) );
  INV_X1 U15275 ( .A(n11913), .ZN(n11911) );
  OAI21_X1 U15276 ( .B1(n11912), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11911), .ZN(n14117) );
  NOR2_X1 U15277 ( .A1(n14118), .A2(n14117), .ZN(n14116) );
  NOR2_X2 U15278 ( .A1(n14116), .A2(n11913), .ZN(n11918) );
  AOI21_X1 U15279 ( .B1(n11914), .B2(n14509), .A(n18529), .ZN(n11915) );
  NOR2_X1 U15280 ( .A1(n11918), .A2(n11917), .ZN(n11919) );
  INV_X1 U15281 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14157) );
  XNOR2_X1 U15282 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11920), .ZN(
        n14152) );
  XOR2_X1 U15283 ( .A(n11921), .B(n18518), .Z(n11923) );
  NOR2_X1 U15284 ( .A1(n11922), .A2(n11923), .ZN(n11924) );
  XNOR2_X1 U15285 ( .A(n11923), .B(n11922), .ZN(n14169) );
  INV_X1 U15286 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14390) );
  NOR2_X1 U15287 ( .A1(n11924), .A2(n14168), .ZN(n11927) );
  XNOR2_X1 U15288 ( .A(n11925), .B(n17282), .ZN(n11928) );
  NAND2_X1 U15289 ( .A1(n11927), .A2(n11928), .ZN(n18851) );
  NOR2_X1 U15290 ( .A1(n11926), .A2(n11930), .ZN(n11932) );
  INV_X1 U15291 ( .A(n11926), .ZN(n11931) );
  OR2_X1 U15292 ( .A1(n11928), .A2(n11927), .ZN(n18852) );
  OAI21_X1 U15293 ( .B1(n11931), .B2(n11930), .A(n18852), .ZN(n11929) );
  AOI21_X1 U15294 ( .B1(n11931), .B2(n11930), .A(n11929), .ZN(n14387) );
  INV_X1 U15295 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21579) );
  NOR2_X1 U15296 ( .A1(n11932), .A2(n14386), .ZN(n18809) );
  NAND3_X1 U15297 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17323) );
  INV_X1 U15298 ( .A(n17323), .ZN(n11933) );
  NAND2_X1 U15299 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n11933), .ZN(
        n11934) );
  NOR2_X1 U15300 ( .A1(n17339), .A2(n11934), .ZN(n17176) );
  INV_X1 U15301 ( .A(n17176), .ZN(n17315) );
  NAND2_X1 U15302 ( .A1(n17267), .A2(n11723), .ZN(n11957) );
  NOR2_X1 U15303 ( .A1(n19736), .A2(n18538), .ZN(n14505) );
  NAND2_X1 U15304 ( .A1(n9695), .A2(n19153), .ZN(n14069) );
  NOR2_X1 U15305 ( .A1(n11936), .A2(n14069), .ZN(n14502) );
  AND2_X1 U15306 ( .A1(n14505), .A2(n14502), .ZN(n11937) );
  NAND2_X1 U15307 ( .A1(n11937), .A2(n19171), .ZN(n11938) );
  INV_X1 U15308 ( .A(n13332), .ZN(n11945) );
  NOR2_X1 U15309 ( .A1(n14505), .A2(n14710), .ZN(n19752) );
  INV_X1 U15310 ( .A(n14024), .ZN(n11947) );
  NOR3_X1 U15311 ( .A1(n11949), .A2(n18578), .A3(n11948), .ZN(n11951) );
  NOR2_X1 U15312 ( .A1(n11951), .A2(n11950), .ZN(n14068) );
  NOR2_X1 U15313 ( .A1(n17287), .A2(n14877), .ZN(n17159) );
  NAND2_X1 U15314 ( .A1(n17301), .A2(n18515), .ZN(n19037) );
  OAI22_X1 U15315 ( .A1(n17160), .A2(n19044), .B1(n17159), .B2(n19037), .ZN(
        n17278) );
  NAND2_X1 U15316 ( .A1(n18995), .A2(n19053), .ZN(n17276) );
  INV_X1 U15317 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19113) );
  NOR3_X1 U15318 ( .A1(n19113), .A2(n14390), .A3(n21579), .ZN(n18982) );
  NAND3_X1 U15319 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18980) );
  NAND2_X1 U15320 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13803) );
  NOR2_X1 U15321 ( .A1(n18980), .A2(n13803), .ZN(n14153) );
  NAND2_X1 U15322 ( .A1(n18982), .A2(n14153), .ZN(n19023) );
  NOR2_X1 U15323 ( .A1(n18985), .A2(n19023), .ZN(n18928) );
  NAND4_X1 U15324 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17176), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A4(n18928), .ZN(n11953) );
  AOI21_X1 U15325 ( .B1(n17176), .B2(n18928), .A(n17314), .ZN(n11952) );
  AOI21_X1 U15326 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14082) );
  NOR2_X1 U15327 ( .A1(n14082), .A2(n18980), .ZN(n14155) );
  NAND2_X1 U15328 ( .A1(n14155), .A2(n18982), .ZN(n19025) );
  NOR2_X1 U15329 ( .A1(n18985), .A2(n19025), .ZN(n18972) );
  INV_X1 U15330 ( .A(n19586), .ZN(n18971) );
  AOI21_X1 U15331 ( .B1(n17176), .B2(n18972), .A(n18971), .ZN(n17310) );
  AOI211_X1 U15332 ( .C1(n18998), .C2(n11953), .A(n11952), .B(n17310), .ZN(
        n17273) );
  OR2_X1 U15333 ( .A1(n17273), .A2(n19121), .ZN(n11954) );
  NAND2_X1 U15334 ( .A1(n18536), .A2(n19723), .ZN(n18043) );
  NOR2_X1 U15335 ( .A1(n18043), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19753) );
  INV_X2 U15336 ( .A(n19055), .ZN(n19089) );
  OAI211_X1 U15337 ( .C1(n11723), .C2(n17276), .A(n11954), .B(n19114), .ZN(
        n14740) );
  OAI21_X1 U15338 ( .B1(n17278), .B2(n14740), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11961) );
  NAND2_X1 U15339 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18928), .ZN(
        n18999) );
  INV_X1 U15340 ( .A(n18999), .ZN(n11955) );
  AOI222_X1 U15341 ( .A1(n19586), .A2(n18972), .B1(n19122), .B2(n18928), .C1(
        n11955), .C2(n18998), .ZN(n18909) );
  NAND2_X1 U15342 ( .A1(n19584), .A2(n18515), .ZN(n19048) );
  OAI22_X1 U15343 ( .A1(n18909), .A2(n17315), .B1(n17287), .B2(n19048), .ZN(
        n17266) );
  NAND3_X1 U15344 ( .A1(n17266), .A2(n11723), .A3(n19053), .ZN(n11956) );
  OAI21_X1 U15345 ( .B1(n11957), .B2(n19044), .A(n11956), .ZN(n11959) );
  INV_X1 U15346 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14741) );
  INV_X1 U15347 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n11958) );
  NOR2_X1 U15348 ( .A1(n19120), .A2(n11958), .ZN(n14878) );
  AOI21_X1 U15349 ( .B1(n11959), .B2(n14741), .A(n14878), .ZN(n11960) );
  OAI21_X1 U15350 ( .B1(n14886), .B2(n19058), .A(n11962), .ZN(P3_U2832) );
  AND2_X2 U15351 ( .A1(n14355), .A2(n14365), .ZN(n12719) );
  NAND2_X1 U15352 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11968) );
  NAND2_X1 U15353 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11967) );
  INV_X1 U15354 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U15355 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11966) );
  NAND2_X1 U15356 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11965) );
  AND2_X4 U15357 ( .A1(n11974), .A2(n14355), .ZN(n12745) );
  NAND2_X1 U15358 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11973) );
  NAND2_X1 U15359 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11972) );
  NAND2_X1 U15360 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11971) );
  NAND2_X1 U15361 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11970) );
  NAND2_X1 U15362 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11978) );
  NAND2_X1 U15363 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11977) );
  AND2_X4 U15364 ( .A1(n11974), .A2(n11979), .ZN(n12755) );
  NAND2_X1 U15365 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11976) );
  NAND2_X1 U15366 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11975) );
  NAND2_X1 U15367 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11983) );
  NAND2_X1 U15368 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11982) );
  NAND2_X1 U15369 ( .A1(n12754), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U15370 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11980) );
  AOI22_X1 U15371 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15372 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15373 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12063), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15374 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9549), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15375 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11994) );
  NAND2_X2 U15376 ( .A1(n11997), .A2(n11996), .ZN(n12084) );
  AOI22_X1 U15377 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15378 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15379 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U15380 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12149), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15381 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15382 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15383 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15384 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15385 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15386 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15387 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12063), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15388 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15389 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15390 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15391 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12063), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15392 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U15393 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12025) );
  AOI22_X1 U15394 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15395 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15396 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15397 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12244), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12020) );
  NAND4_X1 U15398 ( .A1(n12023), .A2(n12022), .A3(n12021), .A4(n12020), .ZN(
        n12024) );
  AOI22_X1 U15399 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12264), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15400 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12160), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15401 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12063), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15402 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12026) );
  NAND4_X1 U15403 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12035) );
  AOI22_X1 U15404 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15405 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15406 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12031) );
  NAND4_X1 U15407 ( .A1(n12033), .A2(n12032), .A3(n12031), .A4(n12030), .ZN(
        n12034) );
  NAND2_X1 U15408 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12040) );
  NAND2_X1 U15409 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12039) );
  NAND2_X1 U15410 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12038) );
  NAND2_X1 U15411 ( .A1(n9550), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12037) );
  NAND2_X1 U15412 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12044) );
  NAND2_X1 U15413 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12043) );
  NAND2_X1 U15414 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12042) );
  NAND2_X1 U15415 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12041) );
  NAND2_X1 U15416 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12049) );
  NAND2_X1 U15417 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12047) );
  NAND2_X1 U15418 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12046) );
  NAND2_X1 U15419 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12053) );
  NAND2_X1 U15420 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12051) );
  NAND2_X1 U15421 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12062) );
  NAND2_X1 U15422 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12061) );
  NAND2_X1 U15423 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12060) );
  NAND2_X1 U15424 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12059) );
  NAND2_X1 U15425 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12067) );
  NAND2_X1 U15426 ( .A1(n12160), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12066) );
  NAND2_X1 U15427 ( .A1(n12149), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12065) );
  NAND2_X1 U15428 ( .A1(n12063), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12064) );
  NAND2_X1 U15429 ( .A1(n12264), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12071) );
  NAND2_X1 U15430 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12070) );
  NAND2_X1 U15431 ( .A1(n12068), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12069) );
  NAND2_X1 U15432 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12076) );
  NAND2_X1 U15433 ( .A1(n12244), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12075) );
  NAND2_X1 U15434 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12073) );
  NOR2_X1 U15435 ( .A1(n12083), .A2(n12111), .ZN(n12109) );
  NAND3_X1 U15436 ( .A1(n12093), .A2(n12109), .A3(n14861), .ZN(n14334) );
  NAND2_X1 U15437 ( .A1(n12106), .A2(n12969), .ZN(n12085) );
  NAND2_X1 U15438 ( .A1(n12112), .A2(n20869), .ZN(n12088) );
  NAND3_X1 U15439 ( .A1(n13096), .A2(n12089), .A3(n12117), .ZN(n12090) );
  OAI21_X1 U15440 ( .B1(n12101), .B2(n12090), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12098) );
  NAND2_X1 U15441 ( .A1(n13111), .A2(n12084), .ZN(n12874) );
  INV_X1 U15442 ( .A(n12950), .ZN(n12205) );
  NAND3_X1 U15443 ( .A1(n12874), .A2(n12205), .A3(n12091), .ZN(n12092) );
  INV_X1 U15444 ( .A(n9580), .ZN(n12095) );
  NAND2_X1 U15445 ( .A1(n12095), .A2(n12094), .ZN(n12096) );
  NAND2_X1 U15446 ( .A1(n12098), .A2(n12097), .ZN(n12126) );
  NAND2_X1 U15447 ( .A1(n12126), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12100) );
  NAND2_X1 U15448 ( .A1(n21372), .A2(n21294), .ZN(n21240) );
  NAND2_X1 U15449 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21206) );
  NAND2_X1 U15450 ( .A1(n21240), .A2(n21206), .ZN(n21179) );
  INV_X1 U15451 ( .A(n21179), .ZN(n21121) );
  AND2_X1 U15452 ( .A1(n15945), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12122) );
  AOI21_X1 U15453 ( .B1(n21121), .B2(n13180), .A(n12122), .ZN(n12099) );
  NAND2_X1 U15454 ( .A1(n12100), .A2(n12099), .ZN(n12102) );
  NAND2_X1 U15455 ( .A1(n12101), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12121) );
  XNOR2_X2 U15456 ( .A(n12102), .B(n12121), .ZN(n20959) );
  NAND2_X1 U15457 ( .A1(n12126), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12105) );
  INV_X1 U15458 ( .A(n13180), .ZN(n12103) );
  MUX2_X1 U15459 ( .A(n15927), .B(n12103), .S(n21294), .Z(n12104) );
  INV_X1 U15460 ( .A(n12106), .ZN(n14126) );
  AOI21_X1 U15461 ( .B1(n14126), .B2(n12107), .A(n10191), .ZN(n12110) );
  INV_X1 U15462 ( .A(n12113), .ZN(n12115) );
  NAND4_X1 U15463 ( .A1(n15260), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14926), 
        .A4(n9708), .ZN(n12114) );
  AOI21_X1 U15464 ( .B1(n14446), .B2(n12115), .A(n12114), .ZN(n12116) );
  INV_X1 U15465 ( .A(n12121), .ZN(n12125) );
  INV_X1 U15466 ( .A(n12122), .ZN(n12123) );
  NAND2_X1 U15467 ( .A1(n12123), .A2(n10077), .ZN(n12124) );
  NAND2_X1 U15468 ( .A1(n12125), .A2(n12124), .ZN(n12132) );
  NAND2_X1 U15469 ( .A1(n12126), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12128) );
  XNOR2_X1 U15470 ( .A(n21206), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20849) );
  AOI22_X1 U15471 ( .A1(n13180), .A2(n20849), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15945), .ZN(n12127) );
  INV_X1 U15472 ( .A(n12130), .ZN(n12131) );
  AND2_X1 U15473 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  AOI22_X1 U15474 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15475 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15476 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15477 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12135) );
  NAND4_X1 U15478 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12144) );
  AOI22_X1 U15479 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15480 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15481 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12140) );
  INV_X1 U15482 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n21645) );
  AOI22_X1 U15483 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12139) );
  NAND4_X1 U15484 ( .A1(n12142), .A2(n12141), .A3(n12140), .A4(n12139), .ZN(
        n12143) );
  NOR2_X1 U15485 ( .A1(n12144), .A2(n12143), .ZN(n12884) );
  OAI22_X1 U15486 ( .A1(n12815), .A2(n21645), .B1(n12239), .B2(n12884), .ZN(
        n12145) );
  INV_X1 U15487 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15488 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15489 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15490 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12063), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15491 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12150) );
  NAND4_X1 U15492 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12159) );
  AOI22_X1 U15493 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15494 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15495 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12155) );
  NAND4_X1 U15496 ( .A1(n12157), .A2(n12156), .A3(n12155), .A4(n12154), .ZN(
        n12158) );
  AOI22_X1 U15497 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15498 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n9551), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15499 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15500 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12161) );
  NAND4_X1 U15501 ( .A1(n12164), .A2(n12163), .A3(n12162), .A4(n12161), .ZN(
        n12170) );
  AOI22_X1 U15502 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15503 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12063), .B1(
        n12744), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15504 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15505 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n12745), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12165) );
  NAND4_X1 U15506 ( .A1(n12168), .A2(n12167), .A3(n12166), .A4(n12165), .ZN(
        n12169) );
  INV_X1 U15507 ( .A(n12171), .ZN(n12781) );
  OAI21_X1 U15508 ( .B1(n12877), .B2(n14376), .A(n12781), .ZN(n12172) );
  NOR2_X1 U15509 ( .A1(n12238), .A2(n12932), .ZN(n12178) );
  MUX2_X1 U15510 ( .A(n12929), .B(n12178), .S(n12877), .Z(n12175) );
  INV_X1 U15511 ( .A(n12175), .ZN(n12219) );
  INV_X1 U15512 ( .A(n12929), .ZN(n12176) );
  NAND2_X1 U15513 ( .A1(n12820), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12192) );
  INV_X1 U15514 ( .A(n12178), .ZN(n12191) );
  AOI22_X1 U15515 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12755), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15516 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15517 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15518 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12179) );
  NAND4_X1 U15519 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12188) );
  AOI22_X1 U15520 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15521 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15522 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15523 ( .A1(n12664), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12183) );
  NAND4_X1 U15524 ( .A1(n12186), .A2(n12185), .A3(n12184), .A4(n12183), .ZN(
        n12187) );
  NAND2_X1 U15525 ( .A1(n12189), .A2(n12872), .ZN(n12190) );
  INV_X1 U15526 ( .A(n20959), .ZN(n12195) );
  INV_X1 U15527 ( .A(n12193), .ZN(n12194) );
  INV_X1 U15528 ( .A(n12238), .ZN(n12196) );
  INV_X1 U15529 ( .A(n12197), .ZN(n12198) );
  NAND2_X1 U15530 ( .A1(n12203), .A2(n12202), .ZN(n12204) );
  AND2_X1 U15531 ( .A1(n12205), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12261) );
  INV_X1 U15532 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n12207) );
  XNOR2_X1 U15533 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20696) );
  AOI21_X1 U15534 ( .B1(n12769), .B2(n20696), .A(n12771), .ZN(n12206) );
  OAI21_X1 U15535 ( .B1(n12765), .B2(n12207), .A(n12206), .ZN(n12208) );
  AOI21_X1 U15536 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n12261), .A(
        n12208), .ZN(n12209) );
  NAND2_X1 U15537 ( .A1(n12771), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12231) );
  NAND2_X1 U15538 ( .A1(n15864), .A2(n12464), .ZN(n12214) );
  INV_X1 U15539 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12211) );
  INV_X1 U15540 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14233) );
  OAI22_X1 U15541 ( .A1(n12765), .A2(n12211), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14233), .ZN(n12212) );
  AOI21_X1 U15542 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12261), .A(
        n12212), .ZN(n12213) );
  NAND2_X1 U15543 ( .A1(n12880), .A2(n12221), .ZN(n12222) );
  NAND2_X1 U15544 ( .A1(n12222), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14103) );
  INV_X1 U15545 ( .A(n12261), .ZN(n12282) );
  INV_X1 U15546 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14930) );
  NAND2_X1 U15547 ( .A1(n21373), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12225) );
  NAND2_X1 U15548 ( .A1(n12772), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12224) );
  OAI211_X1 U15549 ( .C1(n12282), .C2(n14930), .A(n12225), .B(n12224), .ZN(
        n12226) );
  AOI21_X1 U15550 ( .B1(n12223), .B2(n12464), .A(n12226), .ZN(n12227) );
  OR2_X1 U15551 ( .A1(n14103), .A2(n12227), .ZN(n14104) );
  INV_X1 U15552 ( .A(n12227), .ZN(n14105) );
  OR2_X1 U15553 ( .A1(n14105), .A2(n12713), .ZN(n12228) );
  NAND2_X1 U15554 ( .A1(n14104), .A2(n12228), .ZN(n14132) );
  NAND2_X1 U15555 ( .A1(n12230), .A2(n12229), .ZN(n14257) );
  NAND2_X1 U15556 ( .A1(n12126), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12237) );
  INV_X1 U15557 ( .A(n21206), .ZN(n20955) );
  INV_X1 U15558 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21180) );
  NAND2_X1 U15559 ( .A1(n21180), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21048) );
  INV_X1 U15560 ( .A(n21048), .ZN(n12233) );
  NAND2_X1 U15561 ( .A1(n20955), .A2(n12233), .ZN(n21088) );
  NAND2_X1 U15562 ( .A1(n21088), .A2(n21180), .ZN(n12235) );
  NAND2_X1 U15563 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21371) );
  INV_X1 U15564 ( .A(n21371), .ZN(n12234) );
  NAND2_X1 U15565 ( .A1(n20955), .A2(n12234), .ZN(n21368) );
  AOI22_X1 U15566 ( .A1(n20845), .A2(n13180), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15945), .ZN(n12236) );
  NAND2_X1 U15567 ( .A1(n14350), .A2(n14376), .ZN(n12252) );
  AOI22_X1 U15568 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15569 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15570 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15571 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U15572 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12250) );
  AOI22_X1 U15573 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15574 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15575 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15576 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12245) );
  NAND4_X1 U15577 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n12245), .ZN(
        n12249) );
  AOI22_X1 U15578 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12820), .B1(
        n12834), .B2(n12904), .ZN(n12251) );
  NAND2_X1 U15579 ( .A1(n12277), .A2(n15873), .ZN(n12253) );
  INV_X1 U15580 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n12259) );
  INV_X1 U15581 ( .A(n12255), .ZN(n12257) );
  NOR2_X2 U15582 ( .A1(n12255), .A2(n12254), .ZN(n12279) );
  INV_X1 U15583 ( .A(n12279), .ZN(n12256) );
  OAI21_X1 U15584 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12257), .A(
        n12256), .ZN(n15274) );
  AOI22_X1 U15585 ( .A1(n12451), .A2(n15274), .B1(n12771), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12258) );
  OAI21_X1 U15586 ( .B1(n12765), .B2(n12259), .A(n12258), .ZN(n12260) );
  AOI21_X1 U15587 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12261), .A(
        n12260), .ZN(n12262) );
  AOI22_X1 U15588 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15589 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15590 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15591 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12265) );
  NAND4_X1 U15592 ( .A1(n12268), .A2(n12267), .A3(n12266), .A4(n12265), .ZN(
        n12274) );
  AOI22_X1 U15593 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15594 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15595 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15596 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12269) );
  NAND4_X1 U15597 ( .A1(n12272), .A2(n12271), .A3(n12270), .A4(n12269), .ZN(
        n12273) );
  NAND2_X1 U15598 ( .A1(n12834), .A2(n12903), .ZN(n12276) );
  NAND2_X1 U15599 ( .A1(n12820), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12275) );
  INV_X1 U15600 ( .A(n12322), .ZN(n12278) );
  OAI21_X1 U15601 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12279), .A(
        n12299), .ZN(n20782) );
  INV_X1 U15602 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14369) );
  OAI21_X1 U15603 ( .B1(n21050), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21373), .ZN(n12281) );
  NAND2_X1 U15604 ( .A1(n12772), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12280) );
  OAI211_X1 U15605 ( .C1(n12282), .C2(n14369), .A(n12281), .B(n12280), .ZN(
        n12283) );
  OAI21_X1 U15606 ( .B1(n12713), .B2(n20782), .A(n12283), .ZN(n12284) );
  NAND2_X1 U15607 ( .A1(n12820), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12296) );
  AOI22_X1 U15608 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15609 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15610 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15611 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12285) );
  NAND4_X1 U15612 ( .A1(n12288), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(
        n12294) );
  AOI22_X1 U15613 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15614 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15615 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15616 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12289) );
  NAND4_X1 U15617 ( .A1(n12292), .A2(n12291), .A3(n12290), .A4(n12289), .ZN(
        n12293) );
  NAND2_X1 U15618 ( .A1(n12834), .A2(n12917), .ZN(n12295) );
  NAND2_X1 U15619 ( .A1(n12322), .A2(n12899), .ZN(n12902) );
  OR2_X1 U15620 ( .A1(n12322), .A2(n12899), .ZN(n12297) );
  AND2_X1 U15621 ( .A1(n12902), .A2(n12297), .ZN(n12305) );
  INV_X1 U15622 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12303) );
  INV_X1 U15623 ( .A(n12299), .ZN(n12301) );
  NOR2_X2 U15624 ( .A1(n12299), .A2(n12298), .ZN(n12324) );
  INV_X1 U15625 ( .A(n12324), .ZN(n12300) );
  OAI21_X1 U15626 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12301), .A(
        n12300), .ZN(n20676) );
  AOI22_X1 U15627 ( .A1(n12451), .A2(n20676), .B1(n12771), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12302) );
  OAI21_X1 U15628 ( .B1(n12765), .B2(n12303), .A(n12302), .ZN(n12304) );
  INV_X1 U15629 ( .A(n14530), .ZN(n12306) );
  NAND2_X1 U15630 ( .A1(n12820), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12318) );
  AOI22_X1 U15631 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15632 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15633 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15634 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12307) );
  NAND4_X1 U15635 ( .A1(n12310), .A2(n12309), .A3(n12308), .A4(n12307), .ZN(
        n12316) );
  AOI22_X1 U15636 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15637 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15638 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15639 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12311) );
  NAND4_X1 U15640 ( .A1(n12314), .A2(n12313), .A3(n12312), .A4(n12311), .ZN(
        n12315) );
  NAND2_X1 U15641 ( .A1(n12834), .A2(n12916), .ZN(n12317) );
  NAND2_X1 U15642 ( .A1(n12902), .A2(n12319), .ZN(n12323) );
  INV_X1 U15643 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n21595) );
  OAI21_X1 U15644 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12324), .A(
        n12330), .ZN(n20671) );
  AOI22_X1 U15645 ( .A1(n12451), .A2(n20671), .B1(n12771), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12325) );
  OAI21_X1 U15646 ( .B1(n12765), .B2(n21595), .A(n12325), .ZN(n12326) );
  INV_X1 U15647 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U15648 ( .A1(n12834), .A2(n12932), .ZN(n12327) );
  OAI21_X1 U15649 ( .B1(n12328), .B2(n12815), .A(n12327), .ZN(n12329) );
  INV_X1 U15650 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12333) );
  OAI21_X1 U15651 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12331), .A(
        n12359), .ZN(n20661) );
  AOI22_X1 U15652 ( .A1(n12451), .A2(n20661), .B1(n12771), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12332) );
  OAI21_X1 U15653 ( .B1(n12765), .B2(n12333), .A(n12332), .ZN(n12334) );
  AOI22_X1 U15654 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n12756), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15655 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n9551), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15656 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12592), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15657 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n12755), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12335) );
  NAND4_X1 U15658 ( .A1(n12338), .A2(n12337), .A3(n12336), .A4(n12335), .ZN(
        n12344) );
  AOI22_X1 U15659 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15660 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12744), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12341) );
  AOI22_X1 U15661 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15662 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12745), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12339) );
  NAND4_X1 U15663 ( .A1(n12342), .A2(n12341), .A3(n12340), .A4(n12339), .ZN(
        n12343) );
  NOR2_X1 U15664 ( .A1(n12344), .A2(n12343), .ZN(n12348) );
  NAND2_X1 U15665 ( .A1(n12772), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12347) );
  INV_X1 U15666 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12345) );
  XNOR2_X1 U15667 ( .A(n12359), .B(n12345), .ZN(n15616) );
  AOI22_X1 U15668 ( .A1(n15616), .A2(n12451), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12771), .ZN(n12346) );
  OAI211_X1 U15669 ( .C1(n12348), .C2(n12364), .A(n12347), .B(n12346), .ZN(
        n15238) );
  AOI22_X1 U15670 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12755), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15671 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15672 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15673 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12349) );
  NAND4_X1 U15674 ( .A1(n12352), .A2(n12351), .A3(n12350), .A4(n12349), .ZN(
        n12358) );
  AOI22_X1 U15675 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9597), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15676 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15677 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15678 ( .A1(n12664), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12353) );
  NAND4_X1 U15679 ( .A1(n12356), .A2(n12355), .A3(n12354), .A4(n12353), .ZN(
        n12357) );
  NOR2_X1 U15680 ( .A1(n12358), .A2(n12357), .ZN(n12365) );
  NAND2_X1 U15681 ( .A1(n12772), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12363) );
  NAND2_X1 U15682 ( .A1(n12367), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12360) );
  INV_X1 U15683 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15231) );
  XNOR2_X1 U15684 ( .A(n12360), .B(n15231), .ZN(n15610) );
  INV_X1 U15685 ( .A(n12771), .ZN(n12581) );
  NOR2_X1 U15686 ( .A1(n12581), .A2(n15231), .ZN(n12361) );
  AOI21_X1 U15687 ( .B1(n15610), .B2(n12451), .A(n12361), .ZN(n12362) );
  OAI211_X1 U15688 ( .C1(n12365), .C2(n12364), .A(n12363), .B(n12362), .ZN(
        n15222) );
  XNOR2_X1 U15689 ( .A(n12391), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15600) );
  INV_X1 U15690 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15210) );
  OAI22_X1 U15691 ( .A1(n15600), .A2(n12713), .B1(n15210), .B2(n12581), .ZN(
        n12368) );
  AOI21_X1 U15692 ( .B1(n12772), .B2(P1_EAX_REG_10__SCAN_IN), .A(n12368), .ZN(
        n12380) );
  AOI22_X1 U15693 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15694 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12744), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15695 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15696 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9549), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U15697 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12378) );
  AOI22_X1 U15698 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15699 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15700 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15701 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12373) );
  NAND4_X1 U15702 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(
        n12377) );
  OAI21_X1 U15703 ( .B1(n12378), .B2(n12377), .A(n12464), .ZN(n12379) );
  AOI22_X1 U15704 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9551), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15705 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15706 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15707 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12381) );
  NAND4_X1 U15708 ( .A1(n12384), .A2(n12383), .A3(n12382), .A4(n12381), .ZN(
        n12390) );
  AOI22_X1 U15709 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15710 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15711 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15712 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12385) );
  NAND4_X1 U15713 ( .A1(n12388), .A2(n12387), .A3(n12386), .A4(n12385), .ZN(
        n12389) );
  OAI21_X1 U15714 ( .B1(n12390), .B2(n12389), .A(n12464), .ZN(n12397) );
  NAND2_X1 U15715 ( .A1(n12772), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12396) );
  AND2_X2 U15716 ( .A1(n12446), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12440) );
  XNOR2_X1 U15717 ( .A(n12425), .B(n12424), .ZN(n15556) );
  NAND2_X1 U15718 ( .A1(n15556), .A2(n12451), .ZN(n12395) );
  NAND2_X1 U15719 ( .A1(n12771), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12394) );
  NAND4_X1 U15720 ( .A1(n12397), .A2(n12396), .A3(n12395), .A4(n12394), .ZN(
        n15147) );
  AOI22_X1 U15721 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15722 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15723 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15724 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12398) );
  NAND4_X1 U15725 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n12398), .ZN(
        n12407) );
  AOI22_X1 U15726 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12405) );
  AOI22_X1 U15727 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15728 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15729 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12402) );
  NAND4_X1 U15730 ( .A1(n12405), .A2(n12404), .A3(n12403), .A4(n12402), .ZN(
        n12406) );
  OAI21_X1 U15731 ( .B1(n12407), .B2(n12406), .A(n12464), .ZN(n12413) );
  NAND2_X1 U15732 ( .A1(n12772), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U15733 ( .A1(n12440), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12409) );
  INV_X1 U15734 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12408) );
  XNOR2_X1 U15735 ( .A(n12409), .B(n12408), .ZN(n15568) );
  NAND2_X1 U15736 ( .A1(n15568), .A2(n12451), .ZN(n12411) );
  NAND2_X1 U15737 ( .A1(n12771), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12410) );
  NAND4_X1 U15738 ( .A1(n12413), .A2(n12412), .A3(n12411), .A4(n12410), .ZN(
        n15165) );
  AND2_X1 U15739 ( .A1(n15147), .A2(n15165), .ZN(n12467) );
  AOI22_X1 U15740 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12755), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15741 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15742 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15743 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12414) );
  NAND4_X1 U15744 ( .A1(n12417), .A2(n12416), .A3(n12415), .A4(n12414), .ZN(
        n12423) );
  AOI22_X1 U15745 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15746 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15747 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U15748 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12418) );
  NAND4_X1 U15749 ( .A1(n12421), .A2(n12420), .A3(n12419), .A4(n12418), .ZN(
        n12422) );
  OAI21_X1 U15750 ( .B1(n12423), .B2(n12422), .A(n12464), .ZN(n12429) );
  NAND2_X1 U15751 ( .A1(n12772), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12428) );
  XNOR2_X1 U15752 ( .A(n12483), .B(n12482), .ZN(n15545) );
  NAND2_X1 U15753 ( .A1(n15545), .A2(n12451), .ZN(n12427) );
  NAND2_X1 U15754 ( .A1(n12771), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12426) );
  NAND4_X1 U15755 ( .A1(n12429), .A2(n12428), .A3(n12427), .A4(n12426), .ZN(
        n15136) );
  AOI22_X1 U15756 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15757 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12755), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15758 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15759 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12430) );
  NAND4_X1 U15760 ( .A1(n12433), .A2(n12432), .A3(n12431), .A4(n12430), .ZN(
        n12439) );
  AOI22_X1 U15761 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15762 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15763 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15764 ( .A1(n12664), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12434) );
  NAND4_X1 U15765 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n12434), .ZN(
        n12438) );
  OAI21_X1 U15766 ( .B1(n12439), .B2(n12438), .A(n12464), .ZN(n12445) );
  NAND2_X1 U15767 ( .A1(n12772), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12444) );
  INV_X1 U15768 ( .A(n12440), .ZN(n12450) );
  INV_X1 U15769 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12441) );
  XNOR2_X1 U15770 ( .A(n12450), .B(n12441), .ZN(n15578) );
  NAND2_X1 U15771 ( .A1(n15578), .A2(n12769), .ZN(n12443) );
  NAND2_X1 U15772 ( .A1(n12771), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12442) );
  NAND4_X1 U15773 ( .A1(n12445), .A2(n12444), .A3(n12443), .A4(n12442), .ZN(
        n15179) );
  INV_X1 U15774 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n21575) );
  INV_X1 U15775 ( .A(n12446), .ZN(n12448) );
  INV_X1 U15776 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12447) );
  NAND2_X1 U15777 ( .A1(n12448), .A2(n12447), .ZN(n12449) );
  NAND2_X1 U15778 ( .A1(n12450), .A2(n12449), .ZN(n15589) );
  AOI22_X1 U15779 ( .A1(n15589), .A2(n12451), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12771), .ZN(n12452) );
  OAI21_X1 U15780 ( .B1(n12765), .B2(n21575), .A(n12452), .ZN(n15163) );
  INV_X1 U15781 ( .A(n15163), .ZN(n12465) );
  AOI22_X1 U15782 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15783 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15784 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15785 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12453) );
  NAND4_X1 U15786 ( .A1(n12456), .A2(n12455), .A3(n12454), .A4(n12453), .ZN(
        n12462) );
  AOI22_X1 U15787 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15788 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15789 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15790 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12457) );
  NAND4_X1 U15791 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12461) );
  OR2_X1 U15792 ( .A1(n12462), .A2(n12461), .ZN(n12463) );
  NAND2_X1 U15793 ( .A1(n12464), .A2(n12463), .ZN(n15193) );
  NAND2_X1 U15794 ( .A1(n12465), .A2(n15193), .ZN(n12466) );
  AOI22_X1 U15795 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12752), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15796 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n9551), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15797 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15798 ( .A1(n12664), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12469) );
  NAND4_X1 U15799 ( .A1(n12472), .A2(n12471), .A3(n12470), .A4(n12469), .ZN(
        n12478) );
  AOI22_X1 U15800 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12755), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15801 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n12745), .B1(
        n12045), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15802 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12744), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15803 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12473) );
  NAND4_X1 U15804 ( .A1(n12476), .A2(n12475), .A3(n12474), .A4(n12473), .ZN(
        n12477) );
  NOR2_X1 U15805 ( .A1(n12478), .A2(n12477), .ZN(n12481) );
  INV_X1 U15806 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15529) );
  AOI21_X1 U15807 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15529), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12479) );
  AOI21_X1 U15808 ( .B1(n12772), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12479), .ZN(
        n12480) );
  OAI21_X1 U15809 ( .B1(n12732), .B2(n12481), .A(n12480), .ZN(n12485) );
  XNOR2_X1 U15810 ( .A(n12568), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15532) );
  NAND2_X1 U15811 ( .A1(n15532), .A2(n12769), .ZN(n12484) );
  NAND2_X1 U15812 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12486) );
  AND2_X2 U15813 ( .A1(n12487), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12514) );
  NAND2_X2 U15814 ( .A1(n12514), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12589) );
  XNOR2_X1 U15815 ( .A(n12589), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15475) );
  INV_X1 U15816 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15471) );
  AOI21_X1 U15817 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15471), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12488) );
  AOI21_X1 U15818 ( .B1(n12772), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12488), .ZN(
        n12500) );
  AOI22_X1 U15819 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15820 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15821 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15822 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9549), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12489) );
  NAND4_X1 U15823 ( .A1(n12492), .A2(n12491), .A3(n12490), .A4(n12489), .ZN(
        n12498) );
  AOI22_X1 U15824 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9597), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15825 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U15826 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15827 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12493) );
  NAND4_X1 U15828 ( .A1(n12496), .A2(n12495), .A3(n12494), .A4(n12493), .ZN(
        n12497) );
  INV_X1 U15829 ( .A(n12732), .ZN(n12767) );
  OAI21_X1 U15830 ( .B1(n12498), .B2(n12497), .A(n12767), .ZN(n12499) );
  AOI22_X1 U15831 ( .A1(n15475), .A2(n12769), .B1(n12500), .B2(n12499), .ZN(
        n13765) );
  AOI22_X1 U15832 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9551), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15833 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U15834 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12755), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15835 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12501) );
  NAND4_X1 U15836 ( .A1(n12504), .A2(n12503), .A3(n12502), .A4(n12501), .ZN(
        n12510) );
  AOI22_X1 U15837 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U15838 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U15839 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15840 ( .A1(n12664), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12505) );
  NAND4_X1 U15841 ( .A1(n12508), .A2(n12507), .A3(n12506), .A4(n12505), .ZN(
        n12509) );
  NOR2_X1 U15842 ( .A1(n12510), .A2(n12509), .ZN(n12513) );
  INV_X1 U15843 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15369) );
  INV_X1 U15844 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15046) );
  OAI22_X1 U15845 ( .A1(n12765), .A2(n15369), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15046), .ZN(n12511) );
  INV_X1 U15846 ( .A(n12511), .ZN(n12512) );
  OAI21_X1 U15847 ( .B1(n12732), .B2(n12513), .A(n12512), .ZN(n12517) );
  INV_X1 U15848 ( .A(n12514), .ZN(n12515) );
  NAND2_X1 U15849 ( .A1(n12515), .A2(n15046), .ZN(n12516) );
  NAND2_X1 U15850 ( .A1(n12589), .A2(n12516), .ZN(n15483) );
  MUX2_X1 U15851 ( .A(n12517), .B(n15483), .S(n12769), .Z(n12518) );
  INV_X1 U15852 ( .A(n12518), .ZN(n15042) );
  XNOR2_X1 U15853 ( .A(n12552), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15494) );
  NAND2_X1 U15854 ( .A1(n15494), .A2(n12769), .ZN(n12533) );
  AOI22_X1 U15855 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12522) );
  AOI22_X1 U15856 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12521) );
  AOI22_X1 U15857 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U15858 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12519) );
  NAND4_X1 U15859 ( .A1(n12522), .A2(n12521), .A3(n12520), .A4(n12519), .ZN(
        n12528) );
  AOI22_X1 U15860 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12526) );
  AOI22_X1 U15861 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15862 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U15863 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12523) );
  NAND4_X1 U15864 ( .A1(n12526), .A2(n12525), .A3(n12524), .A4(n12523), .ZN(
        n12527) );
  NOR2_X1 U15865 ( .A1(n12528), .A2(n12527), .ZN(n12531) );
  INV_X1 U15866 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15490) );
  AOI21_X1 U15867 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15490), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12529) );
  AOI21_X1 U15868 ( .B1(n12772), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12529), .ZN(
        n12530) );
  OAI21_X1 U15869 ( .B1(n12732), .B2(n12531), .A(n12530), .ZN(n12532) );
  NAND2_X1 U15870 ( .A1(n12533), .A2(n12532), .ZN(n15052) );
  XNOR2_X1 U15871 ( .A(n12534), .B(n15505), .ZN(n15089) );
  AOI22_X1 U15872 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U15873 ( .A1(n12743), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15874 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U15875 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12535) );
  NAND4_X1 U15876 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12544) );
  AOI22_X1 U15877 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9552), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U15878 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12744), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12541) );
  AOI22_X1 U15879 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U15880 ( .A1(n9598), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12539) );
  NAND4_X1 U15881 ( .A1(n12542), .A2(n12541), .A3(n12540), .A4(n12539), .ZN(
        n12543) );
  NOR2_X1 U15882 ( .A1(n12544), .A2(n12543), .ZN(n12547) );
  INV_X1 U15883 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15381) );
  OAI22_X1 U15884 ( .A1(n12765), .A2(n15381), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15505), .ZN(n12545) );
  INV_X1 U15885 ( .A(n12545), .ZN(n12546) );
  OAI21_X1 U15886 ( .B1(n12732), .B2(n12547), .A(n12546), .ZN(n12548) );
  MUX2_X1 U15887 ( .A(n15089), .B(n12548), .S(n12713), .Z(n15087) );
  INV_X1 U15888 ( .A(n12549), .ZN(n12550) );
  INV_X1 U15889 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15073) );
  NAND2_X1 U15890 ( .A1(n12550), .A2(n15073), .ZN(n12551) );
  NAND2_X1 U15891 ( .A1(n12552), .A2(n12551), .ZN(n15501) );
  AOI22_X1 U15892 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12719), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15893 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15894 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15895 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12553) );
  NAND4_X1 U15896 ( .A1(n12556), .A2(n12555), .A3(n12554), .A4(n12553), .ZN(
        n12562) );
  AOI22_X1 U15897 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U15898 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15899 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15900 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12557) );
  NAND4_X1 U15901 ( .A1(n12560), .A2(n12559), .A3(n12558), .A4(n12557), .ZN(
        n12561) );
  NOR2_X1 U15902 ( .A1(n12562), .A2(n12561), .ZN(n12566) );
  INV_X1 U15903 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12563) );
  OAI22_X1 U15904 ( .A1(n12765), .A2(n12563), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15073), .ZN(n12564) );
  INV_X1 U15905 ( .A(n12564), .ZN(n12565) );
  OAI21_X1 U15906 ( .B1(n12732), .B2(n12566), .A(n12565), .ZN(n12567) );
  MUX2_X1 U15907 ( .A(n15501), .B(n12567), .S(n12713), .Z(n15071) );
  NAND2_X1 U15908 ( .A1(n15087), .A2(n15071), .ZN(n15053) );
  NOR2_X1 U15909 ( .A1(n15042), .A2(n15039), .ZN(n13763) );
  AND2_X1 U15910 ( .A1(n13765), .A2(n13763), .ZN(n12586) );
  OR2_X1 U15911 ( .A1(n12568), .A2(n15529), .ZN(n12569) );
  XNOR2_X1 U15912 ( .A(n12569), .B(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15522) );
  AOI22_X1 U15913 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12755), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15914 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15915 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U15916 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12570) );
  NAND4_X1 U15917 ( .A1(n12573), .A2(n12572), .A3(n12571), .A4(n12570), .ZN(
        n12579) );
  AOI22_X1 U15918 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U15919 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15920 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9549), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15921 ( .A1(n9554), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12574) );
  NAND4_X1 U15922 ( .A1(n12577), .A2(n12576), .A3(n12575), .A4(n12574), .ZN(
        n12578) );
  OR2_X1 U15923 ( .A1(n12579), .A2(n12578), .ZN(n12580) );
  NAND2_X1 U15924 ( .A1(n12767), .A2(n12580), .ZN(n12585) );
  INV_X1 U15925 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12582) );
  INV_X1 U15926 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15518) );
  OAI22_X1 U15927 ( .A1(n12765), .A2(n12582), .B1(n15518), .B2(n12581), .ZN(
        n12583) );
  INV_X1 U15928 ( .A(n12583), .ZN(n12584) );
  OAI211_X1 U15929 ( .C1(n15522), .C2(n12713), .A(n12585), .B(n12584), .ZN(
        n15099) );
  INV_X1 U15930 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12614) );
  OAI21_X1 U15931 ( .B1(n12589), .B2(n15471), .A(n12614), .ZN(n12590) );
  NAND2_X1 U15932 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12588) );
  OR2_X2 U15933 ( .A1(n12589), .A2(n12588), .ZN(n12621) );
  NAND2_X1 U15934 ( .A1(n12590), .A2(n12621), .ZN(n15463) );
  AOI22_X1 U15935 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n12603), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15936 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15937 ( .A1(n12592), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15938 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12593) );
  NAND4_X1 U15939 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12602) );
  AOI22_X1 U15940 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n9551), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U15941 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n12745), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15942 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12720), .B1(
        n12744), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15943 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12597) );
  NAND4_X1 U15944 ( .A1(n12600), .A2(n12599), .A3(n12598), .A4(n12597), .ZN(
        n12601) );
  NOR2_X1 U15945 ( .A1(n12602), .A2(n12601), .ZN(n12623) );
  AOI22_X1 U15946 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9598), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15947 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15948 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U15949 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12604) );
  NAND4_X1 U15950 ( .A1(n12607), .A2(n12606), .A3(n12605), .A4(n12604), .ZN(
        n12613) );
  AOI22_X1 U15951 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12611) );
  AOI22_X1 U15952 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15953 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U15954 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12608) );
  NAND4_X1 U15955 ( .A1(n12611), .A2(n12610), .A3(n12609), .A4(n12608), .ZN(
        n12612) );
  NOR2_X1 U15956 ( .A1(n12613), .A2(n12612), .ZN(n12624) );
  XNOR2_X1 U15957 ( .A(n12623), .B(n12624), .ZN(n12617) );
  INV_X1 U15958 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n15361) );
  OAI22_X1 U15959 ( .A1(n12765), .A2(n15361), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12614), .ZN(n12615) );
  INV_X1 U15960 ( .A(n12615), .ZN(n12616) );
  OAI21_X1 U15961 ( .B1(n12732), .B2(n12617), .A(n12616), .ZN(n12618) );
  MUX2_X1 U15962 ( .A(n15463), .B(n12618), .S(n12713), .Z(n15024) );
  INV_X1 U15963 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21640) );
  NAND2_X1 U15964 ( .A1(n12621), .A2(n21640), .ZN(n12622) );
  NAND2_X1 U15965 ( .A1(n12640), .A2(n12622), .ZN(n15455) );
  NOR2_X1 U15966 ( .A1(n12624), .A2(n12623), .ZN(n12643) );
  AOI22_X1 U15967 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U15968 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U15969 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U15970 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12625) );
  NAND4_X1 U15971 ( .A1(n12628), .A2(n12627), .A3(n12626), .A4(n12625), .ZN(
        n12634) );
  AOI22_X1 U15972 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U15973 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15974 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15975 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12629) );
  NAND4_X1 U15976 ( .A1(n12632), .A2(n12631), .A3(n12630), .A4(n12629), .ZN(
        n12633) );
  OR2_X1 U15977 ( .A1(n12634), .A2(n12633), .ZN(n12642) );
  XNOR2_X1 U15978 ( .A(n12643), .B(n12642), .ZN(n12637) );
  INV_X1 U15979 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15356) );
  OAI22_X1 U15980 ( .A1(n12765), .A2(n15356), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21640), .ZN(n12635) );
  INV_X1 U15981 ( .A(n12635), .ZN(n12636) );
  OAI21_X1 U15982 ( .B1(n12637), .B2(n12732), .A(n12636), .ZN(n12638) );
  MUX2_X1 U15983 ( .A(n15455), .B(n12638), .S(n12713), .Z(n15012) );
  INV_X1 U15984 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12639) );
  OR2_X2 U15985 ( .A1(n12640), .A2(n12639), .ZN(n12676) );
  NAND2_X1 U15986 ( .A1(n12640), .A2(n12639), .ZN(n12641) );
  NAND2_X1 U15987 ( .A1(n12676), .A2(n12641), .ZN(n15446) );
  NAND2_X1 U15988 ( .A1(n12643), .A2(n12642), .ZN(n12658) );
  AOI22_X1 U15989 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U15990 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15991 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12645) );
  AOI22_X1 U15992 ( .A1(n12743), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9549), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12644) );
  NAND4_X1 U15993 ( .A1(n12647), .A2(n12646), .A3(n12645), .A4(n12644), .ZN(
        n12653) );
  AOI22_X1 U15994 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U15995 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15996 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12744), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15997 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12648) );
  NAND4_X1 U15998 ( .A1(n12651), .A2(n12650), .A3(n12649), .A4(n12648), .ZN(
        n12652) );
  NOR2_X1 U15999 ( .A1(n12653), .A2(n12652), .ZN(n12659) );
  XNOR2_X1 U16000 ( .A(n12658), .B(n12659), .ZN(n12656) );
  OAI21_X1 U16001 ( .B1(n21050), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n21373), .ZN(n12655) );
  NAND2_X1 U16002 ( .A1(n12772), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n12654) );
  OAI211_X1 U16003 ( .C1(n12656), .C2(n12732), .A(n12655), .B(n12654), .ZN(
        n12657) );
  OAI21_X1 U16004 ( .B1(n15446), .B2(n12713), .A(n12657), .ZN(n14989) );
  XNOR2_X1 U16005 ( .A(n12676), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14906) );
  NAND2_X1 U16006 ( .A1(n14906), .A2(n12769), .ZN(n12675) );
  NOR2_X1 U16007 ( .A1(n12659), .A2(n12658), .ZN(n12681) );
  AOI22_X1 U16008 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U16009 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U16010 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U16011 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12660) );
  NAND4_X1 U16012 ( .A1(n12663), .A2(n12662), .A3(n12661), .A4(n12660), .ZN(
        n12670) );
  AOI22_X1 U16013 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U16014 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U16015 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12664), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U16016 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12665) );
  NAND4_X1 U16017 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n12665), .ZN(
        n12669) );
  OR2_X1 U16018 ( .A1(n12670), .A2(n12669), .ZN(n12680) );
  XNOR2_X1 U16019 ( .A(n12681), .B(n12680), .ZN(n12673) );
  NAND2_X1 U16020 ( .A1(n12772), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n12672) );
  OAI21_X1 U16021 ( .B1(n21050), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n21373), .ZN(n12671) );
  OAI211_X1 U16022 ( .C1(n12673), .C2(n12732), .A(n12672), .B(n12671), .ZN(
        n12674) );
  NAND2_X1 U16023 ( .A1(n12675), .A2(n12674), .ZN(n13748) );
  INV_X1 U16024 ( .A(n12676), .ZN(n12677) );
  NAND2_X1 U16025 ( .A1(n12677), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12678) );
  INV_X1 U16026 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14869) );
  OR2_X2 U16027 ( .A1(n12678), .A2(n14869), .ZN(n12734) );
  NAND2_X1 U16028 ( .A1(n12678), .A2(n14869), .ZN(n12679) );
  NAND2_X1 U16029 ( .A1(n12734), .A2(n12679), .ZN(n15439) );
  NAND2_X1 U16030 ( .A1(n12681), .A2(n12680), .ZN(n12696) );
  AOI22_X1 U16031 ( .A1(n12603), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U16032 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U16033 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U16034 ( .A1(n12664), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12682) );
  NAND4_X1 U16035 ( .A1(n12685), .A2(n12684), .A3(n12683), .A4(n12682), .ZN(
        n12691) );
  AOI22_X1 U16036 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12755), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U16037 ( .A1(n12743), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12744), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U16038 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U16039 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9549), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12686) );
  NAND4_X1 U16040 ( .A1(n12689), .A2(n12688), .A3(n12687), .A4(n12686), .ZN(
        n12690) );
  NOR2_X1 U16041 ( .A1(n12691), .A2(n12690), .ZN(n12697) );
  XNOR2_X1 U16042 ( .A(n12696), .B(n12697), .ZN(n12694) );
  OAI21_X1 U16043 ( .B1(n21050), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n21373), .ZN(n12693) );
  NAND2_X1 U16044 ( .A1(n12772), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12692) );
  OAI211_X1 U16045 ( .C1(n12694), .C2(n12732), .A(n12693), .B(n12692), .ZN(
        n12695) );
  OAI21_X1 U16046 ( .B1(n15439), .B2(n12713), .A(n12695), .ZN(n14856) );
  NOR2_X1 U16047 ( .A1(n13748), .A2(n14856), .ZN(n14857) );
  INV_X1 U16048 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14981) );
  XNOR2_X1 U16049 ( .A(n12734), .B(n14981), .ZN(n15428) );
  NOR2_X1 U16050 ( .A1(n12697), .A2(n12696), .ZN(n12728) );
  AOI22_X1 U16051 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U16052 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U16053 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U16054 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12068), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12698) );
  NAND4_X1 U16055 ( .A1(n12701), .A2(n12700), .A3(n12699), .A4(n12698), .ZN(
        n12708) );
  AOI22_X1 U16056 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9554), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U16057 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U16058 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U16059 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12703) );
  NAND4_X1 U16060 ( .A1(n12706), .A2(n12705), .A3(n12704), .A4(n12703), .ZN(
        n12707) );
  OR2_X1 U16061 ( .A1(n12708), .A2(n12707), .ZN(n12727) );
  XNOR2_X1 U16062 ( .A(n12728), .B(n12727), .ZN(n12711) );
  NAND2_X1 U16063 ( .A1(n12772), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n12710) );
  OAI21_X1 U16064 ( .B1(n21050), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n21373), .ZN(n12709) );
  OAI211_X1 U16065 ( .C1(n12711), .C2(n12732), .A(n12710), .B(n12709), .ZN(
        n12712) );
  OAI21_X1 U16066 ( .B1(n15428), .B2(n12713), .A(n12712), .ZN(n14975) );
  INV_X1 U16067 ( .A(n14975), .ZN(n12714) );
  AND2_X1 U16068 ( .A1(n14857), .A2(n12714), .ZN(n14961) );
  AOI22_X1 U16069 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12745), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U16070 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U16071 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9549), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U16072 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12715) );
  NAND4_X1 U16073 ( .A1(n12718), .A2(n12717), .A3(n12716), .A4(n12715), .ZN(
        n12726) );
  AOI22_X1 U16074 ( .A1(n12719), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12755), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U16075 ( .A1(n9552), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U16076 ( .A1(n12744), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U16077 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12721) );
  NAND4_X1 U16078 ( .A1(n12724), .A2(n12723), .A3(n12722), .A4(n12721), .ZN(
        n12725) );
  NOR2_X1 U16079 ( .A1(n12726), .A2(n12725), .ZN(n12742) );
  NAND2_X1 U16080 ( .A1(n12728), .A2(n12727), .ZN(n12741) );
  XNOR2_X1 U16081 ( .A(n12742), .B(n12741), .ZN(n12733) );
  INV_X1 U16082 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12729) );
  INV_X1 U16083 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12736) );
  OAI22_X1 U16084 ( .A1(n12765), .A2(n12729), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12736), .ZN(n12730) );
  INV_X1 U16085 ( .A(n12730), .ZN(n12731) );
  OAI21_X1 U16086 ( .B1(n12733), .B2(n12732), .A(n12731), .ZN(n12739) );
  NAND2_X1 U16087 ( .A1(n12737), .A2(n12736), .ZN(n12738) );
  NAND2_X1 U16088 ( .A1(n13182), .A2(n12738), .ZN(n15418) );
  MUX2_X1 U16089 ( .A(n12739), .B(n15418), .S(n12769), .Z(n14963) );
  AND2_X1 U16090 ( .A1(n14961), .A2(n14963), .ZN(n12740) );
  NOR2_X1 U16091 ( .A1(n12742), .A2(n12741), .ZN(n12764) );
  AOI22_X1 U16092 ( .A1(n12045), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U16093 ( .A1(n9551), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12743), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U16094 ( .A1(n12745), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12744), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U16095 ( .A1(n12747), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12746), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12748) );
  NAND4_X1 U16096 ( .A1(n12751), .A2(n12750), .A3(n12749), .A4(n12748), .ZN(
        n12762) );
  AOI22_X1 U16097 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12720), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U16098 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U16099 ( .A1(n12755), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12754), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U16100 ( .A1(n12756), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9550), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12757) );
  NAND4_X1 U16101 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12761) );
  NOR2_X1 U16102 ( .A1(n12762), .A2(n12761), .ZN(n12763) );
  XNOR2_X1 U16103 ( .A(n12764), .B(n12763), .ZN(n12768) );
  INV_X1 U16104 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15333) );
  INV_X1 U16105 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14952) );
  OAI22_X1 U16106 ( .A1(n12765), .A2(n15333), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14952), .ZN(n12766) );
  AOI21_X1 U16107 ( .B1(n12768), .B2(n12767), .A(n12766), .ZN(n12770) );
  XNOR2_X1 U16108 ( .A(n13182), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14951) );
  MUX2_X1 U16109 ( .A(n12770), .B(n14951), .S(n12769), .Z(n13140) );
  AOI22_X1 U16110 ( .A1(n12772), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12771), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12773) );
  XNOR2_X1 U16111 ( .A(n12774), .B(n12773), .ZN(n14931) );
  XNOR2_X1 U16112 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12794) );
  XNOR2_X1 U16113 ( .A(n12794), .B(n12795), .ZN(n12844) );
  NAND2_X1 U16114 ( .A1(n12820), .A2(n12844), .ZN(n12776) );
  NAND2_X1 U16115 ( .A1(n12834), .A2(n20854), .ZN(n12775) );
  NAND2_X1 U16116 ( .A1(n14861), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12784) );
  AND2_X1 U16117 ( .A1(n14930), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12777) );
  NOR2_X1 U16118 ( .A1(n12795), .A2(n12777), .ZN(n12780) );
  NAND2_X1 U16119 ( .A1(n12834), .A2(n12780), .ZN(n12778) );
  NAND2_X1 U16120 ( .A1(n12830), .A2(n12778), .ZN(n12783) );
  NAND2_X1 U16121 ( .A1(n12779), .A2(n12094), .ZN(n12799) );
  NAND2_X1 U16122 ( .A1(n12783), .A2(n12782), .ZN(n12788) );
  NAND2_X1 U16123 ( .A1(n12789), .A2(n12788), .ZN(n12787) );
  INV_X1 U16124 ( .A(n12834), .ZN(n12785) );
  NAND3_X1 U16125 ( .A1(n12785), .A2(n20854), .A3(n12784), .ZN(n12819) );
  NAND2_X1 U16126 ( .A1(n12819), .A2(n12844), .ZN(n12786) );
  NAND2_X1 U16127 ( .A1(n12787), .A2(n12786), .ZN(n12793) );
  INV_X1 U16128 ( .A(n12788), .ZN(n12791) );
  INV_X1 U16129 ( .A(n12789), .ZN(n12790) );
  NAND2_X1 U16130 ( .A1(n12791), .A2(n12790), .ZN(n12792) );
  NAND2_X1 U16131 ( .A1(n12793), .A2(n12792), .ZN(n12804) );
  NAND2_X1 U16132 ( .A1(n12795), .A2(n12794), .ZN(n12797) );
  NAND2_X1 U16133 ( .A1(n21372), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12796) );
  NAND2_X1 U16134 ( .A1(n12797), .A2(n12796), .ZN(n12806) );
  XNOR2_X1 U16135 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12805) );
  XNOR2_X1 U16136 ( .A(n12806), .B(n12805), .ZN(n12843) );
  INV_X1 U16137 ( .A(n12843), .ZN(n12800) );
  NAND2_X1 U16138 ( .A1(n12834), .A2(n12800), .ZN(n12798) );
  OAI211_X1 U16139 ( .C1(n12800), .C2(n12815), .A(n12798), .B(n12799), .ZN(
        n12803) );
  INV_X1 U16140 ( .A(n12799), .ZN(n12801) );
  AND3_X1 U16141 ( .A1(n12801), .A2(n12800), .A3(n12834), .ZN(n12802) );
  AOI21_X1 U16142 ( .B1(n12804), .B2(n12803), .A(n12802), .ZN(n12810) );
  NAND2_X1 U16143 ( .A1(n12806), .A2(n12805), .ZN(n12808) );
  NAND2_X1 U16144 ( .A1(n21120), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12807) );
  XNOR2_X1 U16145 ( .A(n12814), .B(n12813), .ZN(n12842) );
  AND2_X1 U16146 ( .A1(n12815), .A2(n12842), .ZN(n12809) );
  INV_X1 U16147 ( .A(n12830), .ZN(n12811) );
  NAND2_X1 U16148 ( .A1(n12811), .A2(n12842), .ZN(n12817) );
  NOR2_X1 U16149 ( .A1(n11964), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12812) );
  AND2_X1 U16150 ( .A1(n12824), .A2(n12827), .ZN(n12845) );
  AND2_X1 U16151 ( .A1(n12815), .A2(n12845), .ZN(n12816) );
  INV_X1 U16152 ( .A(n12819), .ZN(n12821) );
  NAND3_X1 U16153 ( .A1(n12821), .A2(n12820), .A3(n12845), .ZN(n12823) );
  NAND2_X1 U16154 ( .A1(n14376), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12822) );
  NAND2_X1 U16155 ( .A1(n12823), .A2(n12822), .ZN(n12831) );
  INV_X1 U16156 ( .A(n12824), .ZN(n12826) );
  NOR2_X1 U16157 ( .A1(n14369), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12825) );
  INV_X1 U16158 ( .A(n12827), .ZN(n12828) );
  AND2_X1 U16159 ( .A1(n13111), .A2(n12107), .ZN(n12838) );
  NAND2_X1 U16160 ( .A1(n13178), .A2(n15253), .ZN(n14343) );
  INV_X1 U16161 ( .A(n12839), .ZN(n12840) );
  NAND2_X1 U16162 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21523) );
  NAND2_X1 U16163 ( .A1(n12840), .A2(n21523), .ZN(n12841) );
  OR4_X1 U16164 ( .A1(n12845), .A2(n12844), .A3(n12843), .A4(n12842), .ZN(
        n12846) );
  AND2_X1 U16165 ( .A1(n12847), .A2(n12846), .ZN(n13945) );
  NAND2_X1 U16166 ( .A1(n13945), .A2(n21523), .ZN(n12961) );
  OR2_X1 U16167 ( .A1(n14335), .A2(n12961), .ZN(n14015) );
  OAI21_X1 U16168 ( .B1(n13101), .B2(n13141), .A(n14015), .ZN(n12848) );
  INV_X1 U16169 ( .A(n12848), .ZN(n12849) );
  NAND2_X1 U16170 ( .A1(n14931), .A2(n10458), .ZN(n12866) );
  NOR2_X1 U16171 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n21542) );
  NOR3_X1 U16172 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n12853) );
  NOR4_X1 U16173 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12852) );
  NOR4_X1 U16174 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12851) );
  AND4_X1 U16175 ( .A1(n21542), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n12859) );
  NOR4_X1 U16176 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12857) );
  NOR4_X1 U16177 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12856) );
  NOR4_X1 U16178 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12855) );
  NOR4_X1 U16179 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12854) );
  AND4_X1 U16180 ( .A1(n12857), .A2(n12856), .A3(n12855), .A4(n12854), .ZN(
        n12858) );
  NAND2_X1 U16181 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  INV_X1 U16182 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17565) );
  NOR2_X1 U16183 ( .A1(n15387), .A2(n17565), .ZN(n12864) );
  AOI22_X1 U16184 ( .A1(n15393), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15400), .ZN(n12862) );
  INV_X1 U16185 ( .A(n12862), .ZN(n12863) );
  NOR2_X1 U16186 ( .A1(n12864), .A2(n12863), .ZN(n12865) );
  NAND2_X1 U16187 ( .A1(n12866), .A2(n12865), .ZN(P1_U2873) );
  INV_X1 U16188 ( .A(n9583), .ZN(n12897) );
  NAND2_X1 U16189 ( .A1(n12872), .A2(n12877), .ZN(n12885) );
  NAND2_X1 U16190 ( .A1(n12885), .A2(n12884), .ZN(n12906) );
  NAND2_X1 U16191 ( .A1(n12906), .A2(n12904), .ZN(n12868) );
  INV_X1 U16192 ( .A(n12903), .ZN(n12867) );
  XNOR2_X1 U16193 ( .A(n12868), .B(n12867), .ZN(n12869) );
  INV_X1 U16194 ( .A(n12904), .ZN(n12870) );
  XNOR2_X1 U16195 ( .A(n12906), .B(n12870), .ZN(n12871) );
  NAND2_X1 U16196 ( .A1(n12871), .A2(n14446), .ZN(n14521) );
  AOI21_X1 U16197 ( .B1(n12893), .B2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12896) );
  OAI21_X1 U16198 ( .B1(n12872), .B2(n12877), .A(n12885), .ZN(n12873) );
  INV_X1 U16199 ( .A(n12873), .ZN(n12875) );
  AOI21_X1 U16200 ( .B1(n12875), .B2(n14446), .A(n12874), .ZN(n12876) );
  INV_X1 U16201 ( .A(n12877), .ZN(n12878) );
  AOI21_X1 U16202 ( .B1(n12878), .B2(n14446), .A(n9668), .ZN(n12879) );
  NAND2_X1 U16203 ( .A1(n14230), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14229) );
  INV_X1 U16204 ( .A(n12881), .ZN(n12882) );
  OR2_X1 U16205 ( .A1(n14107), .A2(n12882), .ZN(n12883) );
  INV_X1 U16206 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13129) );
  XNOR2_X1 U16207 ( .A(n12885), .B(n12884), .ZN(n12886) );
  AOI21_X1 U16208 ( .B1(n12886), .B2(n14446), .A(n9668), .ZN(n12887) );
  NAND2_X1 U16209 ( .A1(n14256), .A2(n14255), .ZN(n14254) );
  NAND2_X1 U16210 ( .A1(n12888), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12889) );
  INV_X1 U16211 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20785) );
  AND2_X1 U16212 ( .A1(n20785), .A2(n14521), .ZN(n12890) );
  NAND2_X1 U16213 ( .A1(n14522), .A2(n12890), .ZN(n12891) );
  OAI211_X1 U16214 ( .C1(n12892), .C2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n14520), .B(n12891), .ZN(n12895) );
  NAND3_X1 U16215 ( .A1(n12893), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12894) );
  OAI211_X1 U16216 ( .C1(n20774), .C2(n12896), .A(n12895), .B(n12894), .ZN(
        n17521) );
  OR2_X1 U16217 ( .A1(n12898), .A2(n12897), .ZN(n12900) );
  AND2_X1 U16218 ( .A1(n12904), .A2(n12903), .ZN(n12905) );
  NAND2_X1 U16219 ( .A1(n12906), .A2(n12905), .ZN(n12919) );
  XNOR2_X1 U16220 ( .A(n12919), .B(n12917), .ZN(n12907) );
  NAND2_X1 U16221 ( .A1(n12907), .A2(n14446), .ZN(n12908) );
  INV_X1 U16222 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14622) );
  XNOR2_X1 U16223 ( .A(n12923), .B(n14622), .ZN(n17522) );
  NAND2_X1 U16224 ( .A1(n17521), .A2(n17522), .ZN(n17503) );
  NAND2_X1 U16225 ( .A1(n12909), .A2(n9583), .ZN(n12914) );
  INV_X1 U16226 ( .A(n12919), .ZN(n12910) );
  NAND2_X1 U16227 ( .A1(n12910), .A2(n12917), .ZN(n12911) );
  XNOR2_X1 U16228 ( .A(n12911), .B(n12916), .ZN(n12912) );
  NAND2_X1 U16229 ( .A1(n12912), .A2(n14446), .ZN(n12913) );
  NAND2_X1 U16230 ( .A1(n12914), .A2(n12913), .ZN(n17515) );
  NOR2_X1 U16231 ( .A1(n17515), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17508) );
  NAND2_X1 U16232 ( .A1(n12915), .A2(n9583), .ZN(n12922) );
  NAND2_X1 U16233 ( .A1(n12917), .A2(n12916), .ZN(n12918) );
  OR2_X1 U16234 ( .A1(n12919), .A2(n12918), .ZN(n12931) );
  XNOR2_X1 U16235 ( .A(n12931), .B(n12932), .ZN(n12920) );
  NAND2_X1 U16236 ( .A1(n12920), .A2(n14446), .ZN(n12921) );
  NAND2_X1 U16237 ( .A1(n12922), .A2(n12921), .ZN(n17509) );
  NAND2_X1 U16238 ( .A1(n17509), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12927) );
  INV_X1 U16239 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17514) );
  NAND2_X1 U16240 ( .A1(n12924), .A2(n17514), .ZN(n12925) );
  INV_X1 U16241 ( .A(n12924), .ZN(n17505) );
  AND2_X1 U16242 ( .A1(n12929), .A2(n9583), .ZN(n12930) );
  INV_X1 U16243 ( .A(n12931), .ZN(n12933) );
  NAND3_X1 U16244 ( .A1(n12933), .A2(n14446), .A3(n12932), .ZN(n12934) );
  NAND2_X1 U16245 ( .A1(n14615), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12935) );
  INV_X1 U16246 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15803) );
  NAND2_X1 U16247 ( .A1(n9581), .A2(n15803), .ZN(n12936) );
  NAND2_X1 U16248 ( .A1(n15549), .A2(n12936), .ZN(n15565) );
  INV_X1 U16249 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15821) );
  NAND2_X1 U16250 ( .A1(n9581), .A2(n15821), .ZN(n15564) );
  NAND2_X1 U16251 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12937) );
  NAND2_X1 U16252 ( .A1(n15583), .A2(n12937), .ZN(n15562) );
  NAND2_X1 U16253 ( .A1(n15564), .A2(n15562), .ZN(n12938) );
  INV_X1 U16254 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15797) );
  NAND2_X1 U16255 ( .A1(n15583), .A2(n15797), .ZN(n12939) );
  INV_X1 U16256 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15784) );
  NAND2_X1 U16257 ( .A1(n15583), .A2(n15784), .ZN(n15537) );
  NAND2_X1 U16258 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U16259 ( .A1(n15583), .A2(n12940), .ZN(n12941) );
  OR2_X1 U16260 ( .A1(n15583), .A2(n15821), .ZN(n15563) );
  NOR2_X1 U16261 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12943) );
  INV_X1 U16262 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15842) );
  INV_X1 U16263 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15764) );
  AND3_X1 U16264 ( .A1(n15764), .A2(n15784), .A3(n10088), .ZN(n12944) );
  OR2_X1 U16265 ( .A1(n9581), .A2(n12944), .ZN(n12945) );
  XNOR2_X1 U16266 ( .A(n9581), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15506) );
  AND2_X1 U16267 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15711) );
  INV_X1 U16268 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15716) );
  INV_X1 U16269 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15497) );
  INV_X1 U16270 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15733) );
  INV_X1 U16271 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15480) );
  INV_X1 U16272 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15666) );
  INV_X1 U16273 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15689) );
  NAND2_X1 U16274 ( .A1(n15666), .A2(n15689), .ZN(n15422) );
  AND2_X1 U16275 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15667) );
  NAND2_X1 U16276 ( .A1(n15667), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15661) );
  INV_X1 U16277 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13133) );
  INV_X1 U16278 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15652) );
  INV_X1 U16279 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15642) );
  NAND2_X1 U16280 ( .A1(n15652), .A2(n15642), .ZN(n15645) );
  AND2_X1 U16281 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13126) );
  INV_X1 U16282 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15637) );
  XNOR2_X1 U16283 ( .A(n12948), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14854) );
  INV_X1 U16284 ( .A(n12949), .ZN(n14336) );
  NAND2_X1 U16285 ( .A1(n9721), .A2(n21442), .ZN(n15925) );
  NAND2_X1 U16286 ( .A1(n12094), .A2(n15925), .ZN(n13776) );
  NAND2_X1 U16287 ( .A1(n13776), .A2(n21523), .ZN(n12951) );
  NAND2_X1 U16288 ( .A1(n12952), .A2(n13111), .ZN(n12955) );
  AND2_X1 U16289 ( .A1(n9583), .A2(n12221), .ZN(n13112) );
  INV_X1 U16290 ( .A(n13112), .ZN(n12954) );
  MUX2_X1 U16291 ( .A(n12955), .B(n12954), .S(n14013), .Z(n12966) );
  NAND2_X1 U16292 ( .A1(n12957), .A2(n12956), .ZN(n13946) );
  INV_X1 U16293 ( .A(n13946), .ZN(n12958) );
  NAND2_X1 U16294 ( .A1(n12959), .A2(n9697), .ZN(n13098) );
  NAND2_X1 U16295 ( .A1(n12960), .A2(n13098), .ZN(n14017) );
  INV_X1 U16296 ( .A(n14017), .ZN(n12965) );
  NAND2_X1 U16297 ( .A1(n20854), .A2(n15925), .ZN(n12963) );
  INV_X1 U16298 ( .A(n12961), .ZN(n12962) );
  NAND3_X1 U16299 ( .A1(n12963), .A2(n20859), .A3(n12962), .ZN(n12964) );
  NAND3_X1 U16300 ( .A1(n12966), .A2(n12965), .A3(n12964), .ZN(n12967) );
  INV_X1 U16301 ( .A(n13115), .ZN(n12970) );
  NAND2_X1 U16302 ( .A1(n13178), .A2(n12968), .ZN(n13942) );
  CLKBUF_X3 U16303 ( .A(n12971), .Z(n12972) );
  INV_X1 U16304 ( .A(n12972), .ZN(n12973) );
  MUX2_X1 U16305 ( .A(n10191), .B(n12973), .S(P1_EBX_REG_0__SCAN_IN), .Z(
        n14113) );
  NAND2_X2 U16306 ( .A1(n9565), .A2(n13080), .ZN(n13078) );
  MUX2_X1 U16307 ( .A(n13078), .B(n9565), .S(P1_EBX_REG_1__SCAN_IN), .Z(n12975) );
  XNOR2_X1 U16308 ( .A(n14113), .B(n12976), .ZN(n14142) );
  AOI21_X1 U16309 ( .B1(n14142), .B2(n9573), .A(n12976), .ZN(n14292) );
  MUX2_X1 U16310 ( .A(n13078), .B(n9577), .S(P1_EBX_REG_2__SCAN_IN), .Z(n12978) );
  AND2_X1 U16311 ( .A1(n12978), .A2(n12977), .ZN(n14291) );
  NAND2_X1 U16312 ( .A1(n14292), .A2(n14291), .ZN(n14430) );
  INV_X1 U16313 ( .A(n14430), .ZN(n12988) );
  INV_X1 U16314 ( .A(n13078), .ZN(n13046) );
  INV_X1 U16315 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14432) );
  NAND2_X1 U16316 ( .A1(n13046), .A2(n14432), .ZN(n12982) );
  NAND2_X1 U16317 ( .A1(n9573), .A2(n14432), .ZN(n12980) );
  NAND2_X1 U16318 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12979) );
  NAND3_X1 U16319 ( .A1(n12980), .A2(n12972), .A3(n12979), .ZN(n12981) );
  AND2_X1 U16320 ( .A1(n12982), .A2(n12981), .ZN(n14427) );
  NAND2_X1 U16321 ( .A1(n12972), .A2(n20785), .ZN(n12985) );
  INV_X1 U16322 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12983) );
  NAND2_X1 U16323 ( .A1(n9573), .A2(n12983), .ZN(n12984) );
  NAND3_X1 U16324 ( .A1(n12985), .A2(n9577), .A3(n12984), .ZN(n12987) );
  OR2_X1 U16325 ( .A1(n9577), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U16326 ( .A1(n12987), .A2(n12986), .ZN(n14426) );
  INV_X1 U16327 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20711) );
  NAND2_X1 U16328 ( .A1(n13046), .A2(n20711), .ZN(n12992) );
  NAND2_X1 U16329 ( .A1(n9573), .A2(n20711), .ZN(n12990) );
  NAND2_X1 U16330 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12989) );
  NAND3_X1 U16331 ( .A1(n12990), .A2(n12972), .A3(n12989), .ZN(n12991) );
  AND2_X1 U16332 ( .A1(n12992), .A2(n12991), .ZN(n17536) );
  NAND2_X1 U16333 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12993) );
  NAND2_X1 U16334 ( .A1(n12972), .A2(n12993), .ZN(n12995) );
  INV_X1 U16335 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14532) );
  NAND2_X1 U16336 ( .A1(n9573), .A2(n14532), .ZN(n12994) );
  NAND2_X1 U16337 ( .A1(n12995), .A2(n12994), .ZN(n12997) );
  OR2_X1 U16338 ( .A1(n9577), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U16339 ( .A1(n12997), .A2(n12996), .ZN(n17537) );
  NAND2_X1 U16340 ( .A1(n17536), .A2(n17537), .ZN(n12998) );
  NAND2_X1 U16341 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12999) );
  NAND2_X1 U16342 ( .A1(n12972), .A2(n12999), .ZN(n13001) );
  INV_X1 U16343 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n15329) );
  NAND2_X1 U16344 ( .A1(n9573), .A2(n15329), .ZN(n13000) );
  NAND2_X1 U16345 ( .A1(n13001), .A2(n13000), .ZN(n13003) );
  OR2_X1 U16346 ( .A1(n9577), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n13002) );
  AND2_X1 U16347 ( .A1(n13003), .A2(n13002), .ZN(n14618) );
  INV_X1 U16348 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15324) );
  NAND2_X1 U16349 ( .A1(n9573), .A2(n15324), .ZN(n13005) );
  NAND2_X1 U16350 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13004) );
  NAND3_X1 U16351 ( .A1(n13005), .A2(n12972), .A3(n13004), .ZN(n13006) );
  OAI21_X1 U16352 ( .B1(n13078), .B2(P1_EBX_REG_8__SCAN_IN), .A(n13006), .ZN(
        n14619) );
  NOR2_X1 U16353 ( .A1(n14618), .A2(n14619), .ZN(n13007) );
  AND2_X2 U16354 ( .A1(n14617), .A2(n13007), .ZN(n15224) );
  NAND2_X1 U16355 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13008) );
  NAND2_X1 U16356 ( .A1(n12972), .A2(n13008), .ZN(n13010) );
  INV_X1 U16357 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15227) );
  NAND2_X1 U16358 ( .A1(n9573), .A2(n15227), .ZN(n13009) );
  NAND2_X1 U16359 ( .A1(n13010), .A2(n13009), .ZN(n13012) );
  OR2_X1 U16360 ( .A1(n9577), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n13011) );
  NAND2_X1 U16361 ( .A1(n13012), .A2(n13011), .ZN(n15223) );
  MUX2_X1 U16362 ( .A(n13078), .B(n9577), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13013) );
  INV_X1 U16363 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15319) );
  NAND2_X1 U16364 ( .A1(n13046), .A2(n15319), .ZN(n13018) );
  NAND2_X1 U16365 ( .A1(n9573), .A2(n15319), .ZN(n13016) );
  NAND2_X1 U16366 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13015) );
  NAND3_X1 U16367 ( .A1(n13016), .A2(n12972), .A3(n13015), .ZN(n13017) );
  AND2_X1 U16368 ( .A1(n13018), .A2(n13017), .ZN(n15182) );
  INV_X1 U16369 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15822) );
  NAND2_X1 U16370 ( .A1(n12972), .A2(n15822), .ZN(n13021) );
  INV_X1 U16371 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n13019) );
  NAND2_X1 U16372 ( .A1(n9573), .A2(n13019), .ZN(n13020) );
  NAND3_X1 U16373 ( .A1(n13021), .A2(n9577), .A3(n13020), .ZN(n13023) );
  OR2_X1 U16374 ( .A1(n9577), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n13022) );
  NAND2_X1 U16375 ( .A1(n13023), .A2(n13022), .ZN(n15194) );
  MUX2_X1 U16376 ( .A(n13078), .B(n9577), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13025) );
  NAND2_X1 U16377 ( .A1(n13025), .A2(n13024), .ZN(n15152) );
  NAND2_X1 U16378 ( .A1(n12972), .A2(n15803), .ZN(n13028) );
  INV_X1 U16379 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n13026) );
  NAND2_X1 U16380 ( .A1(n9573), .A2(n13026), .ZN(n13027) );
  NAND3_X1 U16381 ( .A1(n13028), .A2(n9577), .A3(n13027), .ZN(n13030) );
  OR2_X1 U16382 ( .A1(n9577), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n13029) );
  NOR2_X1 U16383 ( .A1(n15152), .A2(n15168), .ZN(n13031) );
  MUX2_X1 U16384 ( .A(n13078), .B(n9577), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13033) );
  NAND2_X1 U16385 ( .A1(n13033), .A2(n13032), .ZN(n15120) );
  NAND2_X1 U16386 ( .A1(n12972), .A2(n15784), .ZN(n13035) );
  INV_X1 U16387 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n21557) );
  NAND2_X1 U16388 ( .A1(n9573), .A2(n21557), .ZN(n13034) );
  NAND3_X1 U16389 ( .A1(n13035), .A2(n9577), .A3(n13034), .ZN(n13037) );
  OR2_X1 U16390 ( .A1(n9577), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n13036) );
  NOR2_X1 U16391 ( .A1(n15120), .A2(n15137), .ZN(n13038) );
  NAND2_X1 U16392 ( .A1(n12972), .A2(n15764), .ZN(n13040) );
  INV_X1 U16393 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15315) );
  NAND2_X1 U16394 ( .A1(n9573), .A2(n15315), .ZN(n13039) );
  NAND3_X1 U16395 ( .A1(n13040), .A2(n9577), .A3(n13039), .ZN(n13042) );
  OR2_X1 U16396 ( .A1(n9577), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n13041) );
  MUX2_X1 U16397 ( .A(n13078), .B(n9577), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n13043) );
  INV_X1 U16398 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U16399 ( .A1(n13046), .A2(n15312), .ZN(n13050) );
  NAND2_X1 U16400 ( .A1(n9573), .A2(n15312), .ZN(n13048) );
  NAND2_X1 U16401 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13047) );
  NAND3_X1 U16402 ( .A1(n13048), .A2(n12972), .A3(n13047), .ZN(n13049) );
  AND2_X1 U16403 ( .A1(n13050), .A2(n13049), .ZN(n15055) );
  NAND2_X1 U16404 ( .A1(n12972), .A2(n15497), .ZN(n13052) );
  INV_X1 U16405 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15313) );
  NAND2_X1 U16406 ( .A1(n9573), .A2(n15313), .ZN(n13051) );
  NAND3_X1 U16407 ( .A1(n13052), .A2(n9577), .A3(n13051), .ZN(n13054) );
  OR2_X1 U16408 ( .A1(n9577), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n13053) );
  NAND2_X1 U16409 ( .A1(n13054), .A2(n13053), .ZN(n15069) );
  NAND2_X1 U16410 ( .A1(n15055), .A2(n15069), .ZN(n13055) );
  NAND2_X1 U16411 ( .A1(n12972), .A2(n15480), .ZN(n13057) );
  INV_X1 U16412 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15311) );
  NAND2_X1 U16413 ( .A1(n9573), .A2(n15311), .ZN(n13056) );
  NAND3_X1 U16414 ( .A1(n13057), .A2(n9577), .A3(n13056), .ZN(n13059) );
  OR2_X1 U16415 ( .A1(n9577), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n13058) );
  NAND2_X1 U16416 ( .A1(n13059), .A2(n13058), .ZN(n15043) );
  MUX2_X1 U16417 ( .A(n13078), .B(n9577), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13060) );
  NAND2_X1 U16418 ( .A1(n12972), .A2(n10076), .ZN(n13063) );
  INV_X1 U16419 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n13061) );
  NAND2_X1 U16420 ( .A1(n9573), .A2(n13061), .ZN(n13062) );
  NAND3_X1 U16421 ( .A1(n13063), .A2(n9577), .A3(n13062), .ZN(n13065) );
  OR2_X1 U16422 ( .A1(n9577), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n13064) );
  NOR2_X2 U16423 ( .A1(n15034), .A2(n15033), .ZN(n15036) );
  MUX2_X1 U16424 ( .A(n13078), .B(n9577), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n13067) );
  AND2_X1 U16425 ( .A1(n13067), .A2(n13066), .ZN(n15007) );
  NAND2_X1 U16426 ( .A1(n12972), .A2(n15666), .ZN(n13069) );
  INV_X1 U16427 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15306) );
  NAND2_X1 U16428 ( .A1(n9573), .A2(n15306), .ZN(n13068) );
  NAND3_X1 U16429 ( .A1(n13069), .A2(n9577), .A3(n13068), .ZN(n13071) );
  OR2_X1 U16430 ( .A1(n9577), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n13070) );
  NAND2_X1 U16431 ( .A1(n13071), .A2(n13070), .ZN(n14993) );
  INV_X1 U16432 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21666) );
  NAND2_X1 U16433 ( .A1(n9573), .A2(n21666), .ZN(n13073) );
  NAND2_X1 U16434 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13072) );
  NAND3_X1 U16435 ( .A1(n13073), .A2(n12972), .A3(n13072), .ZN(n13074) );
  OAI21_X1 U16436 ( .B1(n13078), .B2(P1_EBX_REG_26__SCAN_IN), .A(n13074), .ZN(
        n14903) );
  NAND2_X1 U16437 ( .A1(n9577), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13075) );
  NAND2_X1 U16438 ( .A1(n12972), .A2(n13075), .ZN(n13077) );
  INV_X1 U16439 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n21565) );
  NAND2_X1 U16440 ( .A1(n9573), .A2(n21565), .ZN(n13076) );
  AOI22_X1 U16441 ( .A1(n13077), .A2(n13076), .B1(n10191), .B2(n21565), .ZN(
        n14859) );
  MUX2_X1 U16442 ( .A(n13078), .B(n9565), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13079) );
  INV_X1 U16443 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15304) );
  NAND2_X1 U16444 ( .A1(n9573), .A2(n15304), .ZN(n13081) );
  NAND2_X1 U16445 ( .A1(n13082), .A2(n13081), .ZN(n13084) );
  OR2_X1 U16446 ( .A1(n9577), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n13083) );
  OAI21_X1 U16447 ( .B1(n13084), .B2(n10191), .A(n13083), .ZN(n14964) );
  NAND2_X1 U16448 ( .A1(n14932), .A2(n10191), .ZN(n13085) );
  NAND2_X1 U16449 ( .A1(n13085), .A2(n13084), .ZN(n13087) );
  OR2_X1 U16450 ( .A1(n14976), .A2(n10191), .ZN(n13086) );
  OR2_X1 U16451 ( .A1(n13868), .A2(n20854), .ZN(n15926) );
  OAI21_X1 U16452 ( .B1(n13089), .B2(n20869), .A(n15926), .ZN(n13090) );
  NAND2_X1 U16453 ( .A1(n20666), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14850) );
  OAI21_X1 U16454 ( .B1(n14960), .B2(n20808), .A(n14850), .ZN(n13091) );
  INV_X1 U16455 ( .A(n13091), .ZN(n13139) );
  OR2_X1 U16456 ( .A1(n9580), .A2(n12036), .ZN(n13094) );
  INV_X1 U16457 ( .A(n15260), .ZN(n13093) );
  OAI211_X1 U16458 ( .C1(n9671), .C2(n9577), .A(n13096), .B(n13095), .ZN(
        n13114) );
  INV_X1 U16459 ( .A(n13114), .ZN(n13100) );
  NAND2_X1 U16460 ( .A1(n12221), .A2(n20859), .ZN(n13097) );
  AND2_X1 U16461 ( .A1(n13098), .A2(n13097), .ZN(n13099) );
  OAI211_X1 U16462 ( .C1(n9768), .C2(n13101), .A(n13100), .B(n13099), .ZN(
        n14338) );
  NAND2_X1 U16463 ( .A1(n9580), .A2(n12221), .ZN(n13102) );
  OR2_X1 U16464 ( .A1(n14338), .A2(n13103), .ZN(n13104) );
  NAND2_X1 U16465 ( .A1(n13115), .A2(n13104), .ZN(n15703) );
  NAND2_X2 U16466 ( .A1(n13115), .A2(n14925), .ZN(n15802) );
  NAND2_X1 U16467 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15841) );
  NOR2_X1 U16468 ( .A1(n15841), .A2(n17514), .ZN(n15844) );
  AND2_X1 U16469 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13105) );
  NAND2_X1 U16470 ( .A1(n15844), .A2(n13105), .ZN(n15833) );
  INV_X1 U16471 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21660) );
  NOR2_X1 U16472 ( .A1(n21660), .A2(n20785), .ZN(n20784) );
  NAND4_X1 U16473 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A4(n20784), .ZN(n13106) );
  OR2_X1 U16474 ( .A1(n15833), .A2(n13106), .ZN(n15815) );
  NAND2_X1 U16475 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13107) );
  NOR2_X1 U16476 ( .A1(n15815), .A2(n13107), .ZN(n15702) );
  NAND2_X1 U16477 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15702), .ZN(
        n15709) );
  AND2_X1 U16478 ( .A1(n15816), .A2(n15709), .ZN(n13110) );
  OR2_X1 U16479 ( .A1(n15703), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13109) );
  OR2_X1 U16480 ( .A1(n13115), .A2(n20804), .ZN(n13108) );
  NAND2_X1 U16481 ( .A1(n13109), .A2(n13108), .ZN(n15817) );
  NOR2_X1 U16482 ( .A1(n13110), .A2(n15817), .ZN(n15752) );
  NAND2_X1 U16483 ( .A1(n13112), .A2(n13111), .ZN(n13113) );
  INV_X1 U16484 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15883) );
  INV_X1 U16485 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20832) );
  OAI21_X1 U16486 ( .B1(n15883), .B2(n20832), .A(n13129), .ZN(n20790) );
  AND2_X1 U16487 ( .A1(n20790), .A2(n20784), .ZN(n13116) );
  NAND2_X1 U16488 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13116), .ZN(
        n14625) );
  INV_X1 U16489 ( .A(n14625), .ZN(n15843) );
  NAND2_X1 U16490 ( .A1(n15843), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13117) );
  OR2_X1 U16491 ( .A1(n15833), .A2(n13117), .ZN(n15814) );
  NOR2_X1 U16492 ( .A1(n15814), .A2(n15821), .ZN(n15749) );
  AND2_X1 U16493 ( .A1(n15749), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13130) );
  NAND3_X1 U16494 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15759) );
  INV_X1 U16495 ( .A(n15759), .ZN(n15754) );
  AND3_X1 U16496 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n15754), .ZN(n15707) );
  NAND2_X1 U16497 ( .A1(n13130), .A2(n15707), .ZN(n13118) );
  NAND2_X1 U16498 ( .A1(n20826), .A2(n13118), .ZN(n13119) );
  NAND2_X1 U16499 ( .A1(n15752), .A2(n13119), .ZN(n15746) );
  INV_X1 U16500 ( .A(n15711), .ZN(n13120) );
  OR2_X1 U16501 ( .A1(n15746), .A2(n13120), .ZN(n13121) );
  NAND2_X1 U16502 ( .A1(n13121), .A2(n17528), .ZN(n15721) );
  NOR2_X1 U16503 ( .A1(n15480), .A2(n15716), .ZN(n13131) );
  INV_X1 U16504 ( .A(n13131), .ZN(n15712) );
  NAND2_X1 U16505 ( .A1(n20826), .A2(n15712), .ZN(n13122) );
  NAND2_X1 U16506 ( .A1(n15721), .A2(n13122), .ZN(n15684) );
  INV_X1 U16507 ( .A(n15667), .ZN(n13123) );
  AND2_X1 U16508 ( .A1(n20826), .A2(n13123), .ZN(n13124) );
  OR2_X2 U16509 ( .A1(n15684), .A2(n13124), .ZN(n15675) );
  NAND2_X1 U16510 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13125) );
  INV_X1 U16511 ( .A(n20826), .ZN(n15755) );
  NAND2_X1 U16512 ( .A1(n15721), .A2(n15755), .ZN(n15622) );
  INV_X1 U16513 ( .A(n13126), .ZN(n15646) );
  NAND2_X1 U16514 ( .A1(n15622), .A2(n15646), .ZN(n13127) );
  NAND2_X1 U16515 ( .A1(n15653), .A2(n13127), .ZN(n15632) );
  AND2_X1 U16516 ( .A1(n20826), .A2(n15637), .ZN(n13128) );
  INV_X1 U16517 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15621) );
  OR3_X2 U16518 ( .A1(n15632), .A2(n13128), .A3(n15621), .ZN(n15623) );
  INV_X1 U16519 ( .A(n15623), .ZN(n13137) );
  NAND2_X1 U16520 ( .A1(n15802), .A2(n15883), .ZN(n20825) );
  NAND2_X1 U16521 ( .A1(n17545), .A2(n13130), .ZN(n15758) );
  NAND3_X1 U16522 ( .A1(n15707), .A2(n15711), .A3(n13131), .ZN(n13132) );
  NOR2_X1 U16523 ( .A1(n15661), .A2(n13133), .ZN(n13134) );
  NAND2_X1 U16524 ( .A1(n15698), .A2(n13134), .ZN(n15654) );
  OAI21_X1 U16525 ( .B1(n15631), .B2(n15637), .A(n15621), .ZN(n13135) );
  INV_X1 U16526 ( .A(n13135), .ZN(n13136) );
  OAI211_X1 U16527 ( .C1(n14854), .C2(n15862), .A(n13139), .B(n13138), .ZN(
        P1_U3001) );
  NAND2_X1 U16528 ( .A1(n14013), .A2(n13944), .ZN(n13143) );
  NAND2_X1 U16529 ( .A1(n13143), .A2(n13142), .ZN(n13144) );
  AND2_X1 U16530 ( .A1(n20712), .A2(n20885), .ZN(n20708) );
  INV_X1 U16531 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13145) );
  XNOR2_X1 U16532 ( .A(n16129), .B(n13146), .ZN(n16533) );
  NAND2_X1 U16533 ( .A1(n17031), .A2(n16984), .ZN(n16985) );
  NOR2_X1 U16534 ( .A1(n16985), .A2(n13147), .ZN(n16990) );
  NAND3_X1 U16535 ( .A1(n16990), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13148) );
  AND2_X1 U16536 ( .A1(n13151), .A2(n13150), .ZN(n14671) );
  OR2_X1 U16537 ( .A1(n14671), .A2(n13152), .ZN(n13153) );
  AND2_X1 U16538 ( .A1(n13149), .A2(n13153), .ZN(n16676) );
  NOR2_X1 U16539 ( .A1(n16810), .A2(n20519), .ZN(n16670) );
  AOI21_X1 U16540 ( .B1(n16676), .B2(n17127), .A(n16670), .ZN(n13154) );
  INV_X1 U16541 ( .A(n13155), .ZN(n13158) );
  NOR3_X1 U16542 ( .A1(n13156), .A2(n16715), .A3(n16725), .ZN(n13157) );
  NAND2_X1 U16543 ( .A1(n16679), .A2(n10455), .ZN(n13160) );
  INV_X1 U16544 ( .A(n14810), .ZN(n13161) );
  NOR2_X1 U16545 ( .A1(n14811), .A2(n13161), .ZN(n13162) );
  XNOR2_X1 U16546 ( .A(n14812), .B(n13162), .ZN(n16678) );
  OR2_X1 U16547 ( .A1(n16678), .A2(n17139), .ZN(n13171) );
  INV_X1 U16548 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16969) );
  NAND2_X1 U16549 ( .A1(n14786), .A2(n17124), .ZN(n13168) );
  INV_X1 U16550 ( .A(n17028), .ZN(n17057) );
  OAI21_X1 U16551 ( .B1(n17098), .B2(n13163), .A(n17057), .ZN(n16973) );
  NAND2_X1 U16552 ( .A1(n13164), .A2(n16974), .ZN(n13165) );
  OAI21_X1 U16553 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17098), .A(
        n16970), .ZN(n13169) );
  XNOR2_X1 U16554 ( .A(n9581), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15416) );
  NAND2_X1 U16555 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15637), .ZN(
        n13174) );
  AND2_X1 U16556 ( .A1(n15416), .A2(n13174), .ZN(n13175) );
  XNOR2_X1 U16557 ( .A(n13176), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15630) );
  NAND2_X1 U16558 ( .A1(n13178), .A2(n13177), .ZN(n15918) );
  AND3_X1 U16559 ( .A1(n14376), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n13179) );
  NAND2_X1 U16560 ( .A1(n14931), .A2(n20778), .ZN(n13188) );
  OR2_X1 U16561 ( .A1(n13180), .A2(n21384), .ZN(n21522) );
  NAND2_X1 U16562 ( .A1(n21522), .A2(n14376), .ZN(n13181) );
  INV_X1 U16563 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14946) );
  NOR2_X1 U16564 ( .A1(n20771), .A2(n14946), .ZN(n15625) );
  OR2_X2 U16565 ( .A1(n13182), .A2(n14952), .ZN(n13184) );
  INV_X1 U16566 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13183) );
  XNOR2_X2 U16567 ( .A(n13184), .B(n13183), .ZN(n13790) );
  NAND2_X1 U16568 ( .A1(n14376), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15944) );
  NAND2_X1 U16569 ( .A1(n21050), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13185) );
  NAND2_X1 U16570 ( .A1(n15944), .A2(n13185), .ZN(n14109) );
  NOR2_X1 U16571 ( .A1(n13790), .A2(n20783), .ZN(n13186) );
  AOI211_X1 U16572 ( .C1(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n20772), .A(
        n15625), .B(n13186), .ZN(n13187) );
  OAI211_X1 U16573 ( .C1(n15630), .C2(n20633), .A(n13188), .B(n13187), .ZN(
        P1_U2968) );
  INV_X1 U16574 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15979) );
  INV_X1 U16575 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14758) );
  INV_X1 U16576 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13190) );
  OR2_X1 U16577 ( .A1(n13195), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13194) );
  INV_X1 U16578 ( .A(n13192), .ZN(n13193) );
  NAND2_X1 U16579 ( .A1(n13194), .A2(n13193), .ZN(n16855) );
  AOI21_X1 U16580 ( .B1(n14637), .B2(n13196), .A(n13195), .ZN(n16308) );
  MUX2_X1 U16581 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16331) );
  INV_X1 U16582 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16338) );
  MUX2_X1 U16583 ( .A(n16338), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n16330) );
  NOR2_X1 U16584 ( .A1(n16331), .A2(n16330), .ZN(n16319) );
  OAI21_X1 U16585 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13196), .ZN(n16320) );
  NAND2_X1 U16586 ( .A1(n16319), .A2(n16320), .ZN(n16306) );
  NOR2_X1 U16587 ( .A1(n16308), .A2(n16306), .ZN(n16293) );
  NAND2_X1 U16588 ( .A1(n16855), .A2(n16293), .ZN(n16275) );
  NOR2_X1 U16589 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n13192), .ZN(
        n13198) );
  NOR2_X1 U16590 ( .A1(n13197), .A2(n13198), .ZN(n16843) );
  NOR2_X1 U16591 ( .A1(n16275), .A2(n16843), .ZN(n16260) );
  OAI21_X1 U16592 ( .B1(n13197), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13199), .ZN(n16822) );
  NAND2_X1 U16593 ( .A1(n16260), .A2(n16822), .ZN(n16248) );
  AND2_X1 U16594 ( .A1(n13199), .A2(n16811), .ZN(n13200) );
  NOR2_X1 U16595 ( .A1(n13201), .A2(n13200), .ZN(n16813) );
  OR2_X1 U16596 ( .A1(n16248), .A2(n16813), .ZN(n16238) );
  OR2_X1 U16597 ( .A1(n13201), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13202) );
  AND2_X1 U16598 ( .A1(n13204), .A2(n13202), .ZN(n16789) );
  NOR2_X1 U16599 ( .A1(n16238), .A2(n16789), .ZN(n16227) );
  NAND2_X1 U16600 ( .A1(n13204), .A2(n16225), .ZN(n13205) );
  NAND2_X1 U16601 ( .A1(n13203), .A2(n13205), .ZN(n16777) );
  AND2_X1 U16602 ( .A1(n16227), .A2(n16777), .ZN(n16216) );
  NAND2_X1 U16603 ( .A1(n13203), .A2(n13206), .ZN(n13207) );
  NAND2_X1 U16604 ( .A1(n13208), .A2(n13207), .ZN(n16763) );
  NAND2_X1 U16605 ( .A1(n16216), .A2(n16763), .ZN(n16200) );
  AND2_X1 U16606 ( .A1(n13208), .A2(n16747), .ZN(n13209) );
  NOR2_X1 U16607 ( .A1(n13210), .A2(n13209), .ZN(n16749) );
  OR2_X1 U16608 ( .A1(n16200), .A2(n16749), .ZN(n16193) );
  OR2_X1 U16609 ( .A1(n13210), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13212) );
  AND2_X1 U16610 ( .A1(n13212), .A2(n13211), .ZN(n16187) );
  OR2_X1 U16611 ( .A1(n16193), .A2(n16187), .ZN(n16174) );
  NAND2_X1 U16612 ( .A1(n13211), .A2(n16719), .ZN(n13213) );
  AND2_X1 U16613 ( .A1(n9662), .A2(n13213), .ZN(n16721) );
  NOR2_X1 U16614 ( .A1(n16174), .A2(n16721), .ZN(n16161) );
  AND2_X1 U16615 ( .A1(n9662), .A2(n16164), .ZN(n13214) );
  OR2_X1 U16616 ( .A1(n13214), .A2(n13215), .ZN(n16709) );
  AND2_X1 U16617 ( .A1(n16161), .A2(n16709), .ZN(n16146) );
  OR2_X1 U16618 ( .A1(n13215), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13216) );
  NAND2_X1 U16619 ( .A1(n9722), .A2(n13216), .ZN(n16694) );
  AND2_X1 U16620 ( .A1(n16146), .A2(n16694), .ZN(n16137) );
  INV_X1 U16621 ( .A(n13217), .ZN(n13218) );
  NAND2_X1 U16622 ( .A1(n9722), .A2(n13219), .ZN(n13220) );
  NAND2_X1 U16623 ( .A1(n13218), .A2(n13220), .ZN(n16683) );
  NAND2_X1 U16624 ( .A1(n16137), .A2(n16683), .ZN(n16118) );
  AND2_X1 U16625 ( .A1(n13218), .A2(n16121), .ZN(n13221) );
  OR2_X1 U16626 ( .A1(n13221), .A2(n10476), .ZN(n16672) );
  INV_X1 U16627 ( .A(n16672), .ZN(n16124) );
  OR2_X1 U16628 ( .A1(n16118), .A2(n16124), .ZN(n16109) );
  NOR2_X1 U16629 ( .A1(n10476), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13223) );
  OR2_X1 U16630 ( .A1(n13222), .A2(n13223), .ZN(n16666) );
  INV_X1 U16631 ( .A(n16666), .ZN(n13224) );
  NOR2_X1 U16632 ( .A1(n16109), .A2(n13224), .ZN(n16091) );
  NOR2_X1 U16633 ( .A1(n13222), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13226) );
  OR2_X1 U16634 ( .A1(n13225), .A2(n13226), .ZN(n16658) );
  AND2_X1 U16635 ( .A1(n16091), .A2(n16658), .ZN(n16075) );
  OR2_X1 U16636 ( .A1(n13225), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13228) );
  NAND2_X1 U16637 ( .A1(n13228), .A2(n13227), .ZN(n16639) );
  NAND2_X1 U16638 ( .A1(n16075), .A2(n16639), .ZN(n16065) );
  NOR2_X1 U16639 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13229), .ZN(
        n13230) );
  NOR2_X1 U16640 ( .A1(n13232), .A2(n13230), .ZN(n16066) );
  OR2_X1 U16641 ( .A1(n16065), .A2(n16066), .ZN(n13231) );
  OAI21_X1 U16642 ( .B1(n13232), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n13234), .ZN(n16635) );
  AND2_X1 U16643 ( .A1(n13234), .A2(n13233), .ZN(n13235) );
  OR2_X1 U16644 ( .A1(n13235), .A2(n13237), .ZN(n16626) );
  OR2_X1 U16645 ( .A1(n13237), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13238) );
  NAND2_X1 U16646 ( .A1(n13236), .A2(n13238), .ZN(n16621) );
  NAND2_X1 U16647 ( .A1(n16025), .A2(n16621), .ZN(n16004) );
  NAND2_X1 U16648 ( .A1(n13236), .A2(n16600), .ZN(n13239) );
  AND2_X1 U16649 ( .A1(n11149), .A2(n13239), .ZN(n16602) );
  INV_X1 U16650 ( .A(n13240), .ZN(n13245) );
  NAND2_X1 U16651 ( .A1(n13241), .A2(n15979), .ZN(n13242) );
  NAND2_X1 U16652 ( .A1(n13245), .A2(n13242), .ZN(n16589) );
  INV_X1 U16653 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15961) );
  AOI21_X1 U16654 ( .B1(n15961), .B2(n13245), .A(n13244), .ZN(n16583) );
  NOR2_X1 U16655 ( .A1(n13244), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13247) );
  OR2_X1 U16656 ( .A1(n13246), .A2(n13247), .ZN(n16567) );
  XOR2_X1 U16657 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n13246), .Z(
        n14766) );
  XNOR2_X1 U16658 ( .A(n14756), .B(n14766), .ZN(n13263) );
  INV_X1 U16659 ( .A(n13248), .ZN(n13250) );
  NOR2_X1 U16660 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13249) );
  INV_X1 U16661 ( .A(n13251), .ZN(n13252) );
  INV_X1 U16662 ( .A(n17493), .ZN(n14577) );
  NAND2_X1 U16663 ( .A1(n14577), .A2(n13253), .ZN(n16368) );
  AND2_X1 U16664 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U16665 ( .A1(n14591), .A2(n13254), .ZN(n14593) );
  NAND3_X1 U16666 ( .A1(n16345), .A2(n16810), .A3(n14593), .ZN(n13255) );
  NAND2_X1 U16667 ( .A1(n20613), .A2(n20615), .ZN(n13269) );
  NOR2_X1 U16668 ( .A1(n20618), .A2(n13269), .ZN(n13267) );
  INV_X1 U16669 ( .A(n13267), .ZN(n13256) );
  NAND2_X1 U16670 ( .A1(n13268), .A2(n13256), .ZN(n13259) );
  INV_X1 U16671 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13257) );
  NAND3_X1 U16672 ( .A1(n10578), .A2(n13257), .A3(n13269), .ZN(n13258) );
  NAND2_X1 U16673 ( .A1(n13259), .A2(n13258), .ZN(n13260) );
  NAND2_X1 U16674 ( .A1(n13823), .A2(n13260), .ZN(n16350) );
  AOI22_X1 U16675 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n16288), .B1(n16337), 
        .B2(P2_EBX_REG_30__SCAN_IN), .ZN(n13262) );
  NAND2_X1 U16676 ( .A1(n16359), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13261) );
  OAI211_X1 U16677 ( .C1(n13263), .C2(n16345), .A(n13262), .B(n13261), .ZN(
        n13266) );
  NOR2_X1 U16678 ( .A1(n13271), .A2(n13269), .ZN(n13264) );
  NOR2_X1 U16679 ( .A1(n14806), .A2(n16304), .ZN(n13265) );
  AND2_X1 U16680 ( .A1(n13268), .A2(n13267), .ZN(n14587) );
  NAND2_X1 U16681 ( .A1(n13269), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13270) );
  NOR2_X1 U16682 ( .A1(n13271), .A2(n13270), .ZN(n13272) );
  NAND2_X1 U16683 ( .A1(n13277), .A2(n13276), .ZN(P2_U2825) );
  INV_X1 U16684 ( .A(n13281), .ZN(n13282) );
  OAI211_X1 U16685 ( .C1(n13286), .C2(n16579), .A(n13285), .B(n13284), .ZN(
        n13287) );
  NOR2_X1 U16686 ( .A1(n13290), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13292) );
  NAND2_X1 U16687 ( .A1(n14761), .A2(n13293), .ZN(n13294) );
  NAND2_X1 U16688 ( .A1(n10400), .A2(n13295), .ZN(n13301) );
  INV_X1 U16689 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20548) );
  AOI22_X1 U16690 ( .A1(n10624), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13296) );
  OAI21_X1 U16691 ( .B1(n13297), .B2(n20548), .A(n13296), .ZN(n13298) );
  AOI21_X1 U16692 ( .B1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n9548), .A(
        n13298), .ZN(n13300) );
  NOR2_X1 U16693 ( .A1(n16810), .A2(n20548), .ZN(n13741) );
  AOI21_X1 U16694 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13741), .ZN(n13302) );
  OAI21_X1 U16695 ( .B1(n16856), .B2(n13303), .A(n13302), .ZN(n13304) );
  INV_X1 U16696 ( .A(n13304), .ZN(n13305) );
  NAND2_X1 U16697 ( .A1(n17946), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17233) );
  INV_X1 U16698 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18864) );
  NAND2_X1 U16699 ( .A1(n17248), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13320) );
  NAND4_X1 U16700 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13321) );
  INV_X1 U16701 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18820) );
  NAND2_X1 U16702 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18774) );
  NAND2_X1 U16703 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18740) );
  NAND2_X1 U16704 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18700) );
  NOR2_X2 U16705 ( .A1(n18696), .A2(n18700), .ZN(n18687) );
  NAND2_X1 U16706 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18647) );
  INV_X1 U16707 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17685) );
  INV_X1 U16708 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17675) );
  XNOR2_X1 U16709 ( .A(n13318), .B(n17675), .ZN(n17672) );
  INV_X1 U16710 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17709) );
  INV_X1 U16711 ( .A(n13312), .ZN(n13328) );
  NOR2_X1 U16712 ( .A1(n17709), .A2(n13328), .ZN(n13327) );
  OAI21_X1 U16713 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n13327), .A(
        n14729), .ZN(n17183) );
  INV_X1 U16714 ( .A(n17183), .ZN(n17696) );
  INV_X1 U16715 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18663) );
  AND2_X1 U16716 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18687), .ZN(
        n18645) );
  NAND2_X1 U16717 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18645), .ZN(
        n13316) );
  NOR2_X1 U16718 ( .A1(n18663), .A2(n13316), .ZN(n13314) );
  NAND2_X1 U16719 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n13313), .ZN(
        n17175) );
  OAI21_X1 U16720 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13314), .A(
        n17175), .ZN(n18649) );
  INV_X1 U16721 ( .A(n18649), .ZN(n17731) );
  INV_X1 U16722 ( .A(n13316), .ZN(n13315) );
  AOI22_X1 U16723 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n13316), .B1(
        n13315), .B2(n18663), .ZN(n18676) );
  INV_X1 U16724 ( .A(n18676), .ZN(n17746) );
  OAI21_X1 U16725 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18645), .A(
        n13316), .ZN(n18682) );
  INV_X1 U16726 ( .A(n18682), .ZN(n17754) );
  INV_X1 U16727 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18727) );
  INV_X1 U16728 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18020) );
  INV_X1 U16729 ( .A(n13317), .ZN(n18728) );
  NOR2_X1 U16730 ( .A1(n18020), .A2(n18728), .ZN(n18697) );
  INV_X1 U16731 ( .A(n18697), .ZN(n17795) );
  NOR2_X1 U16732 ( .A1(n18727), .A2(n17795), .ZN(n13322) );
  XNOR2_X1 U16733 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n13322), .ZN(
        n18706) );
  INV_X1 U16734 ( .A(n18706), .ZN(n17778) );
  NAND2_X1 U16735 ( .A1(n13318), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13319) );
  INV_X1 U16736 ( .A(n13320), .ZN(n17250) );
  NAND2_X1 U16737 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17250), .ZN(
        n17947) );
  NOR2_X1 U16738 ( .A1(n13321), .A2(n17947), .ZN(n17886) );
  NAND3_X1 U16739 ( .A1(n18805), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17886), .ZN(n17858) );
  INV_X1 U16740 ( .A(n17858), .ZN(n17213) );
  NAND2_X1 U16741 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17213), .ZN(
        n17832) );
  NOR2_X1 U16742 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17832), .ZN(
        n17833) );
  AOI21_X1 U16743 ( .B1(n18727), .B2(n17795), .A(n13322), .ZN(n18731) );
  NOR2_X1 U16744 ( .A1(n17778), .A2(n17777), .ZN(n17776) );
  NOR2_X1 U16745 ( .A1(n17776), .A2(n18000), .ZN(n17765) );
  INV_X1 U16746 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21596) );
  INV_X1 U16747 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21558) );
  INV_X1 U16748 ( .A(n13322), .ZN(n13323) );
  AOI221_X1 U16749 ( .B1(n21596), .B2(n21558), .C1(n13323), .C2(n21558), .A(
        n18645), .ZN(n18699) );
  INV_X1 U16750 ( .A(n18699), .ZN(n13324) );
  NOR2_X1 U16751 ( .A1(n17752), .A2(n18000), .ZN(n17745) );
  NOR2_X2 U16752 ( .A1(n17746), .A2(n17745), .ZN(n17744) );
  NOR2_X1 U16753 ( .A1(n17744), .A2(n18000), .ZN(n17730) );
  NOR2_X1 U16754 ( .A1(n17731), .A2(n17730), .ZN(n17729) );
  NOR2_X1 U16755 ( .A1(n17729), .A2(n18000), .ZN(n17720) );
  INV_X1 U16756 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13325) );
  AOI21_X1 U16757 ( .B1(n13325), .B2(n17175), .A(n13312), .ZN(n17721) );
  NOR2_X2 U16758 ( .A1(n17720), .A2(n17721), .ZN(n17719) );
  INV_X1 U16759 ( .A(n17719), .ZN(n13326) );
  AOI21_X1 U16760 ( .B1(n13328), .B2(n17709), .A(n13327), .ZN(n17708) );
  NAND2_X1 U16761 ( .A1(n17704), .A2(n13329), .ZN(n17705) );
  INV_X1 U16762 ( .A(n18000), .ZN(n13330) );
  AND2_X2 U16763 ( .A1(n17705), .A2(n13330), .ZN(n17695) );
  NOR2_X2 U16764 ( .A1(n17696), .A2(n17695), .ZN(n17694) );
  NOR2_X1 U16765 ( .A1(n17694), .A2(n18000), .ZN(n17683) );
  AOI21_X1 U16766 ( .B1(n17685), .B2(n14729), .A(n13318), .ZN(n17682) );
  AND2_X2 U16767 ( .A1(n17684), .A2(n13330), .ZN(n17674) );
  INV_X1 U16768 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19737) );
  NAND3_X1 U16769 ( .A1(n19740), .A2(n19737), .A3(n17653), .ZN(n19633) );
  NAND2_X1 U16770 ( .A1(n13330), .A2(n18025), .ZN(n17959) );
  NOR3_X1 U16771 ( .A1(n17672), .A2(n17674), .A3(n17959), .ZN(n13346) );
  NAND2_X1 U16772 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19736), .ZN(n13333) );
  AOI211_X4 U16773 ( .C1(n17653), .C2(n19617), .A(n19754), .B(n13333), .ZN(
        n18011) );
  NAND2_X1 U16774 ( .A1(n18017), .A2(n18012), .ZN(n18010) );
  NAND2_X1 U16775 ( .A1(n17984), .A2(n17979), .ZN(n17978) );
  INV_X1 U16776 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17923) );
  INV_X1 U16777 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17905) );
  NAND2_X1 U16778 ( .A1(n17910), .A2(n17905), .ZN(n17897) );
  INV_X1 U16779 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17874) );
  NAND2_X1 U16780 ( .A1(n17882), .A2(n17874), .ZN(n17873) );
  INV_X1 U16781 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17857) );
  INV_X1 U16782 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17827) );
  NAND2_X1 U16783 ( .A1(n17835), .A2(n17827), .ZN(n17826) );
  INV_X1 U16784 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17801) );
  NAND2_X1 U16785 ( .A1(n17812), .A2(n17801), .ZN(n17800) );
  INV_X1 U16786 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18049) );
  NAND2_X1 U16787 ( .A1(n17787), .A2(n18049), .ZN(n17779) );
  INV_X1 U16788 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n18106) );
  INV_X1 U16789 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17740) );
  NAND2_X1 U16790 ( .A1(n17728), .A2(n17740), .ZN(n17718) );
  INV_X1 U16791 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17713) );
  NAND2_X1 U16792 ( .A1(n17717), .A2(n17713), .ZN(n17712) );
  NOR2_X2 U16793 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17712), .ZN(n17693) );
  INV_X1 U16794 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21602) );
  NAND2_X1 U16795 ( .A1(n17693), .A2(n21602), .ZN(n17671) );
  NOR2_X1 U16796 ( .A1(n18038), .A2(n17671), .ZN(n17679) );
  INV_X1 U16797 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n18085) );
  NAND2_X1 U16798 ( .A1(n17679), .A2(n18085), .ZN(n13344) );
  INV_X1 U16799 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19697) );
  INV_X1 U16800 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19694) );
  INV_X1 U16801 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19690) );
  INV_X1 U16802 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19686) );
  INV_X1 U16803 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19681) );
  INV_X1 U16804 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19675) );
  INV_X1 U16805 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19673) );
  INV_X1 U16806 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19670) );
  INV_X1 U16807 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19666) );
  NAND3_X1 U16808 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17994) );
  NOR2_X1 U16809 ( .A1(n19656), .A2(n17994), .ZN(n17971) );
  NAND2_X1 U16810 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17971), .ZN(n17954) );
  NOR2_X1 U16811 ( .A1(n19660), .A2(n17954), .ZN(n17935) );
  NAND3_X1 U16812 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(n17935), .ZN(n17912) );
  NOR2_X1 U16813 ( .A1(n19666), .A2(n17912), .ZN(n17913) );
  NAND2_X1 U16814 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n17913), .ZN(n17892) );
  NAND2_X1 U16815 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17885), .ZN(n17869) );
  NOR3_X1 U16816 ( .A1(n19675), .A2(n19673), .A3(n17869), .ZN(n17838) );
  NAND3_X1 U16817 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n17838), .ZN(n17819) );
  NAND2_X1 U16818 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17794), .ZN(n17804) );
  NOR2_X1 U16819 ( .A1(n19686), .A2(n17804), .ZN(n17791) );
  NAND2_X1 U16820 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17791), .ZN(n17768) );
  NOR2_X1 U16821 ( .A1(n19690), .A2(n17768), .ZN(n17771) );
  NAND2_X1 U16822 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17771), .ZN(n17751) );
  NOR2_X1 U16823 ( .A1(n19694), .A2(n17751), .ZN(n17742) );
  NAND2_X1 U16824 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17742), .ZN(n17732) );
  NOR2_X1 U16825 ( .A1(n19697), .A2(n17732), .ZN(n13335) );
  INV_X1 U16826 ( .A(n19756), .ZN(n19751) );
  NOR2_X2 U16827 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19723), .ZN(n19509) );
  NAND2_X1 U16828 ( .A1(n19628), .A2(n19509), .ZN(n19621) );
  NAND3_X1 U16829 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n13335), .A3(n18042), 
        .ZN(n17692) );
  NAND3_X1 U16830 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n13334) );
  OAI211_X1 U16831 ( .C1(n19735), .C2(n19736), .A(n19617), .B(n17653), .ZN(
        n19615) );
  NAND2_X1 U16832 ( .A1(n18042), .A2(n18004), .ZN(n18040) );
  OAI21_X1 U16833 ( .B1(n17692), .B2(n13334), .A(n18040), .ZN(n17691) );
  INV_X1 U16834 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19699) );
  NAND2_X1 U16835 ( .A1(n18034), .A2(n13335), .ZN(n17727) );
  NAND4_X1 U16836 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17703), .ZN(n13338) );
  NOR2_X1 U16837 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n13338), .ZN(n17677) );
  INV_X1 U16838 ( .A(n17677), .ZN(n13336) );
  INV_X1 U16839 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19707) );
  AOI21_X1 U16840 ( .B1(n17691), .B2(n13336), .A(n19707), .ZN(n13342) );
  AOI21_X1 U16841 ( .B1(n19736), .B2(P3_EBX_REG_31__SCAN_IN), .A(n19754), .ZN(
        n13337) );
  NOR3_X1 U16842 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n11958), .A3(n13338), 
        .ZN(n13339) );
  AOI21_X1 U16843 ( .B1(n17997), .B2(P3_EBX_REG_31__SCAN_IN), .A(n13339), .ZN(
        n13340) );
  INV_X1 U16844 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14734) );
  NAND2_X1 U16845 ( .A1(n13347), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U16846 ( .A1(n13374), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20606), .B2(n20291), .ZN(n13349) );
  INV_X1 U16847 ( .A(n13353), .ZN(n13354) );
  NAND2_X1 U16848 ( .A1(n13351), .A2(n13354), .ZN(n13355) );
  NAND2_X1 U16849 ( .A1(n13374), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13356) );
  NAND2_X1 U16850 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20235) );
  NAND2_X1 U16851 ( .A1(n20591), .A2(n20291), .ZN(n20137) );
  NAND2_X1 U16852 ( .A1(n20235), .A2(n20137), .ZN(n20012) );
  INV_X1 U16853 ( .A(n20012), .ZN(n20083) );
  NAND2_X1 U16854 ( .A1(n20083), .A2(n20606), .ZN(n20211) );
  NAND2_X1 U16855 ( .A1(n13356), .A2(n20211), .ZN(n13357) );
  NAND2_X1 U16856 ( .A1(n13361), .A2(n13360), .ZN(n13365) );
  NAND2_X1 U16857 ( .A1(n20235), .A2(n20582), .ZN(n13363) );
  NAND2_X1 U16858 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20413) );
  INV_X1 U16859 ( .A(n20413), .ZN(n13362) );
  NAND2_X1 U16860 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13362), .ZN(
        n19844) );
  AND2_X1 U16861 ( .A1(n13363), .A2(n19844), .ZN(n20011) );
  AOI22_X1 U16862 ( .A1(n13374), .A2(n17154), .B1(n20606), .B2(n20011), .ZN(
        n13364) );
  NAND2_X1 U16863 ( .A1(n14099), .A2(n14098), .ZN(n13370) );
  INV_X1 U16864 ( .A(n13366), .ZN(n13367) );
  NAND2_X1 U16865 ( .A1(n13368), .A2(n13367), .ZN(n13369) );
  INV_X1 U16866 ( .A(n20235), .ZN(n13372) );
  NAND2_X1 U16867 ( .A1(n20574), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20079) );
  INV_X1 U16868 ( .A(n20079), .ZN(n20082) );
  NAND2_X1 U16869 ( .A1(n13372), .A2(n20082), .ZN(n20142) );
  NAND2_X1 U16870 ( .A1(n19844), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13373) );
  NAND2_X1 U16871 ( .A1(n20142), .A2(n13373), .ZN(n20292) );
  AOI22_X1 U16872 ( .A1(n13374), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20606), .B2(n20292), .ZN(n13375) );
  INV_X1 U16873 ( .A(n13377), .ZN(n13378) );
  AOI22_X1 U16874 ( .A1(n13379), .A2(n13378), .B1(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13347), .ZN(n13380) );
  AND4_X1 U16875 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__5__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13381) );
  AND2_X1 U16876 ( .A1(n14399), .A2(n13381), .ZN(n13382) );
  NAND2_X1 U16877 ( .A1(n14186), .A2(n13382), .ZN(n14264) );
  NAND3_X1 U16878 ( .A1(n14266), .A2(n14410), .A3(n14329), .ZN(n13383) );
  NOR2_X1 U16879 ( .A1(n14264), .A2(n13383), .ZN(n13384) );
  AOI22_X1 U16880 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13389) );
  AOI22_X1 U16881 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13388) );
  AOI22_X1 U16882 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13387) );
  AOI22_X1 U16883 ( .A1(n11346), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13386) );
  NAND4_X1 U16884 ( .A1(n13389), .A2(n13388), .A3(n13387), .A4(n13386), .ZN(
        n13399) );
  AOI22_X1 U16885 ( .A1(n13534), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13397) );
  INV_X1 U16886 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13392) );
  NAND2_X1 U16887 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13391) );
  NAND2_X1 U16888 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13390) );
  OAI211_X1 U16889 ( .C1(n10727), .C2(n13392), .A(n13391), .B(n13390), .ZN(
        n13393) );
  INV_X1 U16890 ( .A(n13393), .ZN(n13396) );
  AOI22_X1 U16891 ( .A1(n13541), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U16892 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13394) );
  NAND4_X1 U16893 ( .A1(n13397), .A2(n13396), .A3(n13395), .A4(n13394), .ZN(
        n13398) );
  NOR2_X1 U16894 ( .A1(n13399), .A2(n13398), .ZN(n14675) );
  AOI22_X1 U16895 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10780), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U16896 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11327), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U16897 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13527), .ZN(n13401) );
  AOI22_X1 U16898 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11346), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13400) );
  NAND4_X1 U16899 ( .A1(n13403), .A2(n13402), .A3(n13401), .A4(n13400), .ZN(
        n13413) );
  AOI22_X1 U16900 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n13533), .B1(
        n13534), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U16901 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13405) );
  NAND2_X1 U16902 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13404) );
  OAI211_X1 U16903 ( .C1(n10727), .C2(n13406), .A(n13405), .B(n13404), .ZN(
        n13407) );
  INV_X1 U16904 ( .A(n13407), .ZN(n13410) );
  AOI22_X1 U16905 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13540), .B1(
        n13541), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13409) );
  NAND2_X1 U16906 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13408) );
  NAND4_X1 U16907 ( .A1(n13411), .A2(n13410), .A3(n13409), .A4(n13408), .ZN(
        n13412) );
  NOR2_X1 U16908 ( .A1(n13413), .A2(n13412), .ZN(n14681) );
  AOI22_X1 U16909 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10780), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U16910 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n13526), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U16911 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U16912 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n11346), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13414) );
  NAND4_X1 U16913 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13428) );
  INV_X1 U16914 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13423) );
  INV_X1 U16915 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13419) );
  INV_X1 U16916 ( .A(n13540), .ZN(n13495) );
  INV_X1 U16917 ( .A(n13541), .ZN(n13497) );
  INV_X1 U16918 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13418) );
  OAI22_X1 U16919 ( .A1(n13419), .A2(n13495), .B1(n13497), .B2(n13418), .ZN(
        n13420) );
  AOI21_X1 U16920 ( .B1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n13542), .A(
        n13420), .ZN(n13422) );
  AOI22_X1 U16921 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13535), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13421) );
  OAI211_X1 U16922 ( .C1(n13423), .C2(n10727), .A(n13422), .B(n13421), .ZN(
        n13427) );
  INV_X1 U16923 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13424) );
  OAI22_X1 U16924 ( .A1(n13425), .A2(n10733), .B1(n13465), .B2(n13424), .ZN(
        n13426) );
  AOI22_X1 U16925 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10780), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13432) );
  AOI22_X1 U16926 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11327), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U16927 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U16928 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n11346), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13429) );
  NAND4_X1 U16929 ( .A1(n13432), .A2(n13431), .A3(n13430), .A4(n13429), .ZN(
        n13443) );
  OAI22_X1 U16930 ( .A1(n13434), .A2(n10733), .B1(n13465), .B2(n13433), .ZN(
        n13442) );
  AOI22_X1 U16931 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13540), .B1(
        n13541), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13435) );
  OAI21_X1 U16932 ( .B1(n13437), .B2(n13436), .A(n13435), .ZN(n13441) );
  AOI22_X1 U16933 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13535), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13438) );
  OAI21_X1 U16934 ( .B1(n13439), .B2(n10727), .A(n13438), .ZN(n13440) );
  NOR4_X1 U16935 ( .A1(n13443), .A2(n13442), .A3(n13441), .A4(n13440), .ZN(
        n16434) );
  AOI22_X1 U16936 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10780), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13447) );
  AOI22_X1 U16937 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13526), .B1(
        n11327), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U16938 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13445) );
  AOI22_X1 U16939 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11346), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13444) );
  NAND4_X1 U16940 ( .A1(n13447), .A2(n13446), .A3(n13445), .A4(n13444), .ZN(
        n13458) );
  INV_X1 U16941 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13453) );
  INV_X1 U16942 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13449) );
  INV_X1 U16943 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13448) );
  OAI22_X1 U16944 ( .A1(n13449), .A2(n13495), .B1(n13497), .B2(n13448), .ZN(
        n13450) );
  AOI21_X1 U16945 ( .B1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n13542), .A(
        n13450), .ZN(n13452) );
  AOI22_X1 U16946 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13535), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13451) );
  OAI211_X1 U16947 ( .C1(n13453), .C2(n10727), .A(n13452), .B(n13451), .ZN(
        n13457) );
  INV_X1 U16948 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13454) );
  OAI22_X1 U16949 ( .A1(n13455), .A2(n10733), .B1(n13465), .B2(n13454), .ZN(
        n13456) );
  OR3_X1 U16950 ( .A1(n13458), .A2(n13457), .A3(n13456), .ZN(n16429) );
  INV_X1 U16951 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13464) );
  INV_X1 U16952 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13460) );
  INV_X1 U16953 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13459) );
  OAI22_X1 U16954 ( .A1(n13497), .A2(n13460), .B1(n13495), .B2(n13459), .ZN(
        n13461) );
  AOI21_X1 U16955 ( .B1(n13542), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n13461), .ZN(n13463) );
  AOI22_X1 U16956 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13462) );
  OAI211_X1 U16957 ( .C1(n10727), .C2(n13464), .A(n13463), .B(n13462), .ZN(
        n13473) );
  INV_X1 U16958 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13635) );
  OAI22_X1 U16959 ( .A1(n10733), .A2(n13466), .B1(n13465), .B2(n13635), .ZN(
        n13472) );
  AOI22_X1 U16960 ( .A1(n10780), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13470) );
  AOI22_X1 U16961 ( .A1(n11327), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13469) );
  AOI22_X1 U16962 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13527), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U16963 ( .A1(n11346), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13467) );
  NAND4_X1 U16964 ( .A1(n13470), .A2(n13469), .A3(n13468), .A4(n13467), .ZN(
        n13471) );
  NOR3_X1 U16965 ( .A1(n13473), .A2(n13472), .A3(n13471), .ZN(n16424) );
  OAI22_X1 U16966 ( .A1(n13477), .A2(n13476), .B1(n13475), .B2(n13474), .ZN(
        n13493) );
  INV_X1 U16967 ( .A(n13526), .ZN(n13479) );
  OAI22_X1 U16968 ( .A1(n13481), .A2(n13480), .B1(n13479), .B2(n13478), .ZN(
        n13492) );
  INV_X1 U16969 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13484) );
  OAI22_X1 U16970 ( .A1(n13485), .A2(n13484), .B1(n13483), .B2(n13482), .ZN(
        n13491) );
  OAI22_X1 U16971 ( .A1(n13489), .A2(n13488), .B1(n13487), .B2(n13486), .ZN(
        n13490) );
  NOR4_X1 U16972 ( .A1(n13493), .A2(n13492), .A3(n13491), .A4(n13490), .ZN(
        n13504) );
  AOI22_X1 U16973 ( .A1(n13534), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13503) );
  INV_X1 U16974 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13496) );
  INV_X1 U16975 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13494) );
  OAI22_X1 U16976 ( .A1(n13497), .A2(n13496), .B1(n13495), .B2(n13494), .ZN(
        n13501) );
  AOI22_X1 U16977 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13498) );
  OAI21_X1 U16978 ( .B1(n10727), .B2(n13499), .A(n13498), .ZN(n13500) );
  AOI211_X1 U16979 ( .C1(n13542), .C2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n13501), .B(n13500), .ZN(n13502) );
  NAND3_X1 U16980 ( .A1(n13504), .A2(n13503), .A3(n13502), .ZN(n16419) );
  AOI22_X1 U16981 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U16982 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U16983 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9579), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13515) );
  INV_X1 U16984 ( .A(n13507), .ZN(n13510) );
  INV_X1 U16985 ( .A(n13508), .ZN(n13509) );
  NAND2_X1 U16986 ( .A1(n13510), .A2(n13509), .ZN(n13687) );
  NAND2_X1 U16987 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13513) );
  NAND2_X1 U16988 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13512) );
  AND3_X1 U16989 ( .A1(n13687), .A2(n13513), .A3(n13512), .ZN(n13514) );
  NAND4_X1 U16990 ( .A1(n13517), .A2(n13516), .A3(n13515), .A4(n13514), .ZN(
        n13525) );
  AOI22_X1 U16991 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13523) );
  AOI22_X1 U16992 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U16993 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n9578), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13521) );
  INV_X1 U16994 ( .A(n13687), .ZN(n13676) );
  NAND2_X1 U16995 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13519) );
  NAND2_X1 U16996 ( .A1(n13684), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13518) );
  AND3_X1 U16997 ( .A1(n13676), .A2(n13519), .A3(n13518), .ZN(n13520) );
  NAND4_X1 U16998 ( .A1(n13523), .A2(n13522), .A3(n13521), .A4(n13520), .ZN(
        n13524) );
  NAND2_X1 U16999 ( .A1(n13525), .A2(n13524), .ZN(n13573) );
  AOI22_X1 U17000 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10780), .B1(
        n10757), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13532) );
  AOI22_X1 U17001 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11327), .B1(
        n13526), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13531) );
  AOI22_X1 U17002 ( .A1(n13528), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n13527), .ZN(n13530) );
  AOI22_X1 U17003 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n11346), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13529) );
  NAND4_X1 U17004 ( .A1(n13532), .A2(n13531), .A3(n13530), .A4(n13529), .ZN(
        n13548) );
  AOI22_X1 U17005 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n13534), .B1(
        n13533), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13546) );
  INV_X1 U17006 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U17007 ( .A1(n13535), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13537) );
  NAND2_X1 U17008 ( .A1(n10686), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n13536) );
  OAI211_X1 U17009 ( .C1(n10727), .C2(n13538), .A(n13537), .B(n13536), .ZN(
        n13539) );
  INV_X1 U17010 ( .A(n13539), .ZN(n13545) );
  AOI22_X1 U17011 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13541), .B1(
        n13540), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13544) );
  NAND2_X1 U17012 ( .A1(n13542), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13543) );
  NAND4_X1 U17013 ( .A1(n13546), .A2(n13545), .A3(n13544), .A4(n13543), .ZN(
        n13547) );
  OR2_X1 U17014 ( .A1(n13548), .A2(n13547), .ZN(n13566) );
  AOI22_X1 U17015 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13555) );
  AOI22_X1 U17016 ( .A1(n9575), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13678), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13554) );
  AOI22_X1 U17017 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13682), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13553) );
  NAND2_X1 U17018 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13551) );
  NAND2_X1 U17019 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13550) );
  AND3_X1 U17020 ( .A1(n13687), .A2(n13551), .A3(n13550), .ZN(n13552) );
  NAND4_X1 U17021 ( .A1(n13555), .A2(n13554), .A3(n13553), .A4(n13552), .ZN(
        n13563) );
  AOI22_X1 U17022 ( .A1(n13506), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13561) );
  AOI22_X1 U17023 ( .A1(n13505), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9589), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13560) );
  AOI22_X1 U17024 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13682), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13559) );
  NAND2_X1 U17025 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13557) );
  NAND2_X1 U17026 ( .A1(n13684), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13556) );
  AND3_X1 U17027 ( .A1(n13676), .A2(n13557), .A3(n13556), .ZN(n13558) );
  NAND4_X1 U17028 ( .A1(n13561), .A2(n13560), .A3(n13559), .A4(n13558), .ZN(
        n13562) );
  NAND2_X1 U17029 ( .A1(n13566), .A2(n13571), .ZN(n13564) );
  INV_X1 U17030 ( .A(n14186), .ZN(n13628) );
  NOR2_X1 U17031 ( .A1(n13564), .A2(n13573), .ZN(n13592) );
  AOI211_X1 U17032 ( .C1(n13573), .C2(n13564), .A(n13628), .B(n13592), .ZN(
        n16403) );
  INV_X1 U17033 ( .A(n13564), .ZN(n13565) );
  NAND2_X1 U17034 ( .A1(n13565), .A2(n17491), .ZN(n13570) );
  INV_X1 U17035 ( .A(n13566), .ZN(n13568) );
  NAND2_X1 U17036 ( .A1(n20620), .A2(n13571), .ZN(n13567) );
  NAND2_X1 U17037 ( .A1(n13568), .A2(n13567), .ZN(n13569) );
  NAND2_X1 U17038 ( .A1(n16403), .A2(n16407), .ZN(n13576) );
  INV_X1 U17039 ( .A(n13571), .ZN(n13572) );
  NOR2_X1 U17040 ( .A1(n17491), .A2(n13572), .ZN(n16414) );
  INV_X1 U17041 ( .A(n13573), .ZN(n16404) );
  NAND2_X1 U17042 ( .A1(n16414), .A2(n16404), .ZN(n13574) );
  AOI22_X1 U17043 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13577), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13583) );
  AOI22_X1 U17044 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13582) );
  AOI22_X1 U17045 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13682), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13581) );
  NAND2_X1 U17046 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n13579) );
  NAND2_X1 U17047 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13578) );
  AND3_X1 U17048 ( .A1(n13687), .A2(n13579), .A3(n13578), .ZN(n13580) );
  NAND4_X1 U17049 ( .A1(n13583), .A2(n13582), .A3(n13581), .A4(n13580), .ZN(
        n13591) );
  AOI22_X1 U17050 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13589) );
  AOI22_X1 U17051 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U17052 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9578), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13587) );
  NAND2_X1 U17053 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13585) );
  NAND2_X1 U17054 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13584) );
  AND3_X1 U17055 ( .A1(n13676), .A2(n13585), .A3(n13584), .ZN(n13586) );
  NAND4_X1 U17056 ( .A1(n13589), .A2(n13588), .A3(n13587), .A4(n13586), .ZN(
        n13590) );
  AND2_X1 U17057 ( .A1(n13591), .A2(n13590), .ZN(n13608) );
  NAND2_X1 U17058 ( .A1(n13592), .A2(n13608), .ZN(n13611) );
  OAI211_X1 U17059 ( .C1(n13592), .C2(n13608), .A(n14186), .B(n13611), .ZN(
        n13610) );
  AOI22_X1 U17060 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9595), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13599) );
  AOI22_X1 U17061 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U17062 ( .A1(n13683), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13511), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13597) );
  NAND2_X1 U17063 ( .A1(n9578), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13595) );
  NAND2_X1 U17064 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n13594) );
  AND3_X1 U17065 ( .A1(n13687), .A2(n13595), .A3(n13594), .ZN(n13596) );
  NAND4_X1 U17066 ( .A1(n13599), .A2(n13598), .A3(n13597), .A4(n13596), .ZN(
        n13607) );
  AOI22_X1 U17067 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13605) );
  AOI22_X1 U17068 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13604) );
  AOI22_X1 U17069 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13682), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13603) );
  NAND2_X1 U17070 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13601) );
  NAND2_X1 U17071 ( .A1(n13684), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13600) );
  AND3_X1 U17072 ( .A1(n13676), .A2(n13601), .A3(n13600), .ZN(n13602) );
  NAND4_X1 U17073 ( .A1(n13605), .A2(n13604), .A3(n13603), .A4(n13602), .ZN(
        n13606) );
  NAND2_X1 U17074 ( .A1(n13607), .A2(n13606), .ZN(n16389) );
  NAND2_X1 U17075 ( .A1(n9593), .A2(n13608), .ZN(n16399) );
  NOR3_X2 U17076 ( .A1(n16400), .A2(n16389), .A3(n16399), .ZN(n16376) );
  INV_X1 U17077 ( .A(n13611), .ZN(n13613) );
  INV_X1 U17078 ( .A(n16389), .ZN(n13612) );
  OAI211_X1 U17079 ( .C1(n13613), .C2(n13612), .A(n14186), .B(n13629), .ZN(
        n16391) );
  AOI22_X1 U17080 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13619) );
  AOI22_X1 U17081 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U17082 ( .A1(n10564), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13682), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U17083 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n13615) );
  NAND2_X1 U17084 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n13614) );
  AND3_X1 U17085 ( .A1(n13687), .A2(n13615), .A3(n13614), .ZN(n13616) );
  NAND4_X1 U17086 ( .A1(n13619), .A2(n13618), .A3(n13617), .A4(n13616), .ZN(
        n13627) );
  AOI22_X1 U17087 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13625) );
  AOI22_X1 U17088 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13624) );
  AOI22_X1 U17089 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9578), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U17090 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13621) );
  NAND2_X1 U17091 ( .A1(n13684), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13620) );
  AND3_X1 U17092 ( .A1(n13676), .A2(n13621), .A3(n13620), .ZN(n13622) );
  NAND4_X1 U17093 ( .A1(n13625), .A2(n13624), .A3(n13623), .A4(n13622), .ZN(
        n13626) );
  NAND2_X1 U17094 ( .A1(n13627), .A2(n13626), .ZN(n13631) );
  AOI21_X1 U17095 ( .B1(n13629), .B2(n13631), .A(n13628), .ZN(n13630) );
  NAND2_X1 U17096 ( .A1(n13630), .A2(n16377), .ZN(n16383) );
  INV_X1 U17097 ( .A(n13631), .ZN(n13632) );
  NAND2_X1 U17098 ( .A1(n9593), .A2(n13632), .ZN(n16382) );
  NAND2_X1 U17099 ( .A1(n16383), .A2(n16382), .ZN(n13652) );
  NAND2_X1 U17100 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13633) );
  NAND2_X1 U17101 ( .A1(n13676), .A2(n13633), .ZN(n13638) );
  OAI22_X1 U17102 ( .A1(n9588), .A2(n13635), .B1(n9562), .B2(n13634), .ZN(
        n13637) );
  AOI22_X1 U17103 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U17104 ( .A1(n10564), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13639) );
  NAND3_X1 U17105 ( .A1(n13641), .A2(n13640), .A3(n13639), .ZN(n13651) );
  NAND2_X1 U17106 ( .A1(n13684), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13642) );
  NAND2_X1 U17107 ( .A1(n13687), .A2(n13642), .ZN(n13646) );
  INV_X1 U17108 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13643) );
  OAI22_X1 U17109 ( .A1(n10496), .A2(n13644), .B1(n13549), .B2(n13643), .ZN(
        n13645) );
  AOI211_X1 U17110 ( .C1(n13511), .C2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n13646), .B(n13645), .ZN(n13649) );
  AOI22_X1 U17111 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13648) );
  AOI22_X1 U17112 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13647) );
  NAND3_X1 U17113 ( .A1(n13649), .A2(n13648), .A3(n13647), .ZN(n13650) );
  AND2_X1 U17114 ( .A1(n13651), .A2(n13650), .ZN(n16378) );
  OAI21_X2 U17115 ( .B1(n16376), .B2(n16375), .A(n10485), .ZN(n16372) );
  AOI22_X1 U17116 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U17117 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13653) );
  NAND2_X1 U17118 ( .A1(n13654), .A2(n13653), .ZN(n13667) );
  AOI22_X1 U17119 ( .A1(n10564), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9578), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13657) );
  NAND2_X1 U17120 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13656) );
  NAND2_X1 U17121 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13655) );
  NAND4_X1 U17122 ( .A1(n13657), .A2(n13687), .A3(n13656), .A4(n13655), .ZN(
        n13666) );
  AOI22_X1 U17123 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13683), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13660) );
  AOI22_X1 U17124 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13659) );
  NAND2_X1 U17125 ( .A1(n13660), .A2(n13659), .ZN(n13665) );
  AOI22_X1 U17126 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13682), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13663) );
  NAND2_X1 U17127 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13662) );
  NAND2_X1 U17128 ( .A1(n13684), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13661) );
  NAND4_X1 U17129 ( .A1(n13663), .A2(n13676), .A3(n13662), .A4(n13661), .ZN(
        n13664) );
  OAI22_X1 U17130 ( .A1(n13667), .A2(n13666), .B1(n13665), .B2(n13664), .ZN(
        n13670) );
  INV_X1 U17131 ( .A(n16378), .ZN(n13668) );
  NOR3_X1 U17132 ( .A1(n16377), .A2(n9593), .A3(n13668), .ZN(n13669) );
  XOR2_X1 U17133 ( .A(n13670), .B(n13669), .Z(n16371) );
  INV_X1 U17134 ( .A(n13669), .ZN(n13671) );
  OAI21_X2 U17135 ( .B1(n16372), .B2(n16371), .A(n10466), .ZN(n13695) );
  AOI22_X1 U17136 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10564), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U17137 ( .A1(n13683), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13672) );
  NAND2_X1 U17138 ( .A1(n13673), .A2(n13672), .ZN(n13692) );
  AOI22_X1 U17139 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9578), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13677) );
  NAND2_X1 U17140 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13675) );
  NAND2_X1 U17141 ( .A1(n9576), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13674) );
  NAND4_X1 U17142 ( .A1(n13677), .A2(n13676), .A3(n13675), .A4(n13674), .ZN(
        n13691) );
  AOI22_X1 U17143 ( .A1(n13636), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10564), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13681) );
  AOI22_X1 U17144 ( .A1(n13679), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13658), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13680) );
  NAND2_X1 U17145 ( .A1(n13681), .A2(n13680), .ZN(n13690) );
  AOI22_X1 U17146 ( .A1(n13683), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13682), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13688) );
  NAND2_X1 U17147 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n13686) );
  NAND2_X1 U17148 ( .A1(n13684), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13685) );
  NAND4_X1 U17149 ( .A1(n13688), .A2(n13687), .A3(n13686), .A4(n13685), .ZN(
        n13689) );
  OAI22_X1 U17150 ( .A1(n13692), .A2(n13691), .B1(n13690), .B2(n13689), .ZN(
        n13693) );
  XNOR2_X1 U17151 ( .A(n13695), .B(n13694), .ZN(n14809) );
  NAND2_X1 U17152 ( .A1(n14570), .A2(n14206), .ZN(n13698) );
  AND3_X1 U17153 ( .A1(n11247), .A2(n14574), .A3(n20613), .ZN(n13696) );
  NAND2_X1 U17154 ( .A1(n11494), .A2(n13696), .ZN(n13697) );
  NAND2_X1 U17155 ( .A1(n13698), .A2(n13697), .ZN(n14215) );
  NAND2_X1 U17156 ( .A1(n13701), .A2(n13700), .ZN(n13702) );
  NOR2_X1 U17157 ( .A1(n13699), .A2(n13702), .ZN(n13703) );
  INV_X1 U17158 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n13724) );
  AND2_X1 U17159 ( .A1(n19795), .A2(n13708), .ZN(n13985) );
  NOR4_X1 U17160 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13712) );
  NOR4_X1 U17161 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13711) );
  NOR4_X1 U17162 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13710) );
  NOR4_X1 U17163 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13709) );
  AND4_X1 U17164 ( .A1(n13712), .A2(n13711), .A3(n13710), .A4(n13709), .ZN(
        n13717) );
  NOR4_X1 U17165 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13715) );
  NOR4_X1 U17166 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13714) );
  NOR4_X1 U17167 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13713) );
  AND4_X1 U17168 ( .A1(n13715), .A2(n13714), .A3(n13713), .A4(n20499), .ZN(
        n13716) );
  NAND2_X1 U17169 ( .A1(n13717), .A2(n13716), .ZN(n13718) );
  NAND2_X1 U17170 ( .A1(n13985), .A2(n19839), .ZN(n16546) );
  AND2_X1 U17171 ( .A1(n9590), .A2(n19895), .ZN(n13720) );
  INV_X1 U17172 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n13722) );
  NAND2_X1 U17173 ( .A1(n19839), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13721) );
  OAI21_X1 U17174 ( .B1(n19839), .B2(n13722), .A(n13721), .ZN(n16553) );
  AOI22_X1 U17175 ( .A1(n16543), .A2(n16553), .B1(n19796), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n13723) );
  OAI21_X1 U17176 ( .B1(n13724), .B2(n16546), .A(n13723), .ZN(n13725) );
  INV_X1 U17177 ( .A(n13725), .ZN(n13727) );
  NAND2_X1 U17178 ( .A1(n16541), .A2(BUF2_REG_30__SCAN_IN), .ZN(n13726) );
  NAND2_X1 U17179 ( .A1(n13727), .A2(n13726), .ZN(n13728) );
  OAI21_X1 U17180 ( .B1(n14809), .B2(n16562), .A(n13730), .ZN(P2_U2889) );
  AOI22_X1 U17181 ( .A1(n11298), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n13732), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13733) );
  OAI21_X1 U17182 ( .B1(n13734), .B2(n20548), .A(n13733), .ZN(n13735) );
  XNOR2_X2 U17183 ( .A(n13736), .B(n13735), .ZN(n16440) );
  OAI21_X1 U17184 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17098), .A(
        n13737), .ZN(n13742) );
  NOR4_X1 U17185 ( .A1(n16865), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13739), .A4(n13738), .ZN(n13740) );
  AOI211_X1 U17186 ( .C1(n13742), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n13741), .B(n13740), .ZN(n13743) );
  OAI21_X1 U17187 ( .B1(n16369), .B2(n17116), .A(n13743), .ZN(n13744) );
  INV_X1 U17188 ( .A(n13744), .ZN(n13746) );
  INV_X1 U17189 ( .A(n13748), .ZN(n13749) );
  OR2_X1 U17190 ( .A1(n13750), .A2(n13749), .ZN(n13751) );
  INV_X1 U17191 ( .A(n15459), .ZN(n15450) );
  OAI21_X1 U17192 ( .B1(n15450), .B2(n15661), .A(n9581), .ZN(n13753) );
  INV_X1 U17193 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U17194 ( .A1(n20666), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15660) );
  OAI21_X1 U17195 ( .B1(n15530), .B2(n14907), .A(n15660), .ZN(n13754) );
  INV_X1 U17196 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21520) );
  NOR3_X1 U17197 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21520), .ZN(n13758) );
  NOR4_X1 U17198 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13757) );
  NAND4_X1 U17199 ( .A1(n20838), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13758), .A4(
        n13757), .ZN(U214) );
  INV_X1 U17200 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20594) );
  NOR2_X1 U17201 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n20594), .ZN(n13760) );
  NOR4_X1 U17202 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13759) );
  NAND4_X1 U17203 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13760), .A3(n13759), .A4(
        n21590), .ZN(n13761) );
  NOR2_X1 U17204 ( .A1(n19837), .A2(n13761), .ZN(n17564) );
  NAND2_X1 U17205 ( .A1(n17564), .A2(U214), .ZN(U212) );
  AND2_X1 U17206 ( .A1(n15070), .A2(n13763), .ZN(n15041) );
  INV_X1 U17207 ( .A(n13945), .ZN(n13766) );
  NOR2_X1 U17208 ( .A1(n13946), .A2(n13766), .ZN(n13869) );
  NAND2_X1 U17209 ( .A1(n13869), .A2(n13767), .ZN(n13866) );
  NOR2_X1 U17210 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21526) );
  NAND2_X1 U17211 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21526), .ZN(n15933) );
  NAND2_X1 U17212 ( .A1(n12451), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13768) );
  MUX2_X1 U17213 ( .A(n15933), .B(n13768), .S(n14376), .Z(n13769) );
  NAND2_X1 U17214 ( .A1(n20771), .A2(n13769), .ZN(n13770) );
  NOR2_X1 U17215 ( .A1(n15472), .A2(n15255), .ZN(n13802) );
  NAND2_X1 U17216 ( .A1(n15045), .A2(n13772), .ZN(n13773) );
  NAND2_X1 U17217 ( .A1(n15034), .A2(n13773), .ZN(n15701) );
  AND2_X1 U17218 ( .A1(n20854), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13793) );
  INV_X1 U17219 ( .A(n13793), .ZN(n13774) );
  AND2_X1 U17220 ( .A1(n21523), .A2(n21050), .ZN(n15923) );
  NOR2_X1 U17221 ( .A1(n13774), .A2(n15923), .ZN(n13775) );
  NOR2_X1 U17222 ( .A1(n15701), .A2(n20678), .ZN(n13801) );
  AND2_X1 U17223 ( .A1(n13776), .A2(n15923), .ZN(n13794) );
  INV_X1 U17224 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21623) );
  NAND4_X1 U17225 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n15256)
         );
  NAND3_X1 U17226 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n15248) );
  NOR3_X1 U17227 ( .A1(n21623), .A2(n15256), .A3(n15248), .ZN(n15235) );
  NAND2_X1 U17228 ( .A1(n15270), .A2(n15235), .ZN(n13777) );
  NAND2_X1 U17229 ( .A1(n20673), .A2(n13777), .ZN(n15242) );
  AND2_X1 U17230 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n15169) );
  AND2_X1 U17231 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n13778) );
  NAND2_X1 U17232 ( .A1(n15169), .A2(n13778), .ZN(n15117) );
  AND4_X1 U17233 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(P1_REIP_REG_17__SCAN_IN), .A4(P1_REIP_REG_16__SCAN_IN), .ZN(n13779) );
  NAND2_X1 U17234 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n13779), .ZN(n13780) );
  NOR2_X1 U17235 ( .A1(n15117), .A2(n13780), .ZN(n13784) );
  INV_X1 U17236 ( .A(n13784), .ZN(n13781) );
  NAND2_X1 U17237 ( .A1(n20673), .A2(n13781), .ZN(n13782) );
  NAND2_X1 U17238 ( .A1(n15242), .A2(n13782), .ZN(n15107) );
  AND3_X1 U17239 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14867) );
  NOR2_X1 U17240 ( .A1(n15287), .A2(n14867), .ZN(n13783) );
  NOR2_X1 U17241 ( .A1(n15107), .A2(n13783), .ZN(n15064) );
  NAND2_X1 U17242 ( .A1(n15235), .A2(n13784), .ZN(n15077) );
  NAND2_X1 U17243 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n13785) );
  OR2_X1 U17244 ( .A1(n15077), .A2(n13785), .ZN(n13786) );
  NOR2_X1 U17245 ( .A1(n15287), .A2(n13786), .ZN(n15058) );
  INV_X1 U17246 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21484) );
  AND2_X1 U17247 ( .A1(n21484), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n13787) );
  NAND2_X1 U17248 ( .A1(n15058), .A2(n13787), .ZN(n15048) );
  INV_X1 U17249 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21486) );
  AOI21_X1 U17250 ( .B1(n15064), .B2(n15048), .A(n21486), .ZN(n13800) );
  AND2_X1 U17251 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n13788) );
  NAND2_X1 U17252 ( .A1(n15058), .A2(n13788), .ZN(n15027) );
  AND2_X2 U17253 ( .A1(n13790), .A2(n13789), .ZN(n15294) );
  INV_X1 U17254 ( .A(n15475), .ZN(n13791) );
  OAI22_X1 U17255 ( .A1(n9558), .A2(n13791), .B1(n15471), .B2(n20694), .ZN(
        n13792) );
  INV_X1 U17256 ( .A(n13792), .ZN(n13798) );
  NOR2_X1 U17257 ( .A1(n13794), .A2(n13793), .ZN(n13795) );
  NAND2_X1 U17258 ( .A1(n20691), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n13797) );
  OAI211_X1 U17259 ( .C1(n15027), .C2(P1_REIP_REG_22__SCAN_IN), .A(n13798), 
        .B(n13797), .ZN(n13799) );
  OR4_X1 U17260 ( .A1(n13802), .A2(n13801), .A3(n13800), .A4(n13799), .ZN(
        P1_U2818) );
  INV_X1 U17261 ( .A(n13803), .ZN(n13805) );
  INV_X1 U17262 ( .A(n18998), .ZN(n19073) );
  NAND2_X1 U17263 ( .A1(n19073), .A2(n17314), .ZN(n18978) );
  INV_X1 U17264 ( .A(n18978), .ZN(n17336) );
  NAND2_X1 U17265 ( .A1(n18998), .A2(n19020), .ZN(n17306) );
  OAI211_X1 U17266 ( .C1(n13805), .C2(n17336), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n17306), .ZN(n13804) );
  AOI21_X1 U17267 ( .B1(n19586), .B2(n14082), .A(n13804), .ZN(n14122) );
  AOI221_X1 U17268 ( .B1(n14122), .B2(n19114), .C1(n17276), .C2(n19114), .A(
        n14157), .ZN(n13814) );
  INV_X1 U17269 ( .A(n14082), .ZN(n13806) );
  OAI21_X1 U17270 ( .B1(n19073), .B2(n19020), .A(n17314), .ZN(n14087) );
  AOI22_X1 U17271 ( .A1(n19586), .A2(n13806), .B1(n13805), .B2(n14087), .ZN(
        n18981) );
  NOR4_X1 U17272 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18981), .A3(
        n9934), .A4(n19121), .ZN(n13813) );
  AOI21_X1 U17273 ( .B1(n14157), .B2(n13808), .A(n13807), .ZN(n18879) );
  AND2_X1 U17274 ( .A1(n19119), .A2(n18879), .ZN(n13812) );
  INV_X1 U17275 ( .A(n17301), .ZN(n19115) );
  XNOR2_X1 U17276 ( .A(n13809), .B(n13810), .ZN(n18881) );
  OAI22_X1 U17277 ( .A1(n19115), .A2(n18881), .B1(n19120), .B2(n19656), .ZN(
        n13811) );
  OR4_X1 U17278 ( .A1(n13814), .A2(n13813), .A3(n13812), .A4(n13811), .ZN(
        P3_U2858) );
  INV_X1 U17279 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n13815) );
  NOR2_X1 U17280 ( .A1(n21442), .A2(n13815), .ZN(n21443) );
  INV_X1 U17281 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21452) );
  INV_X1 U17282 ( .A(HOLD), .ZN(n21441) );
  OAI222_X1 U17283 ( .A1(n21443), .A2(P1_STATE_REG_1__SCAN_IN), .B1(n21443), 
        .B2(HOLD), .C1(n21452), .C2(n21441), .ZN(n13816) );
  OAI211_X1 U17284 ( .C1(n21523), .C2(n20628), .A(n13816), .B(n15925), .ZN(
        P1_U3195) );
  MUX2_X1 U17285 ( .A(P2_STATEBS16_REG_SCAN_IN), .B(n20613), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n13818) );
  INV_X1 U17286 ( .A(n14591), .ZN(n20614) );
  NAND2_X1 U17287 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13817), .ZN(n14595) );
  OAI211_X1 U17288 ( .C1(n13818), .C2(P2_STATE2_REG_2__SCAN_IN), .A(n20614), 
        .B(n14595), .ZN(n13819) );
  INV_X1 U17289 ( .A(n13819), .ZN(P2_U3178) );
  INV_X1 U17290 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n13821) );
  NAND2_X1 U17291 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20607), .ZN(n13820) );
  OAI22_X1 U17292 ( .A1(n13823), .A2(n13821), .B1(n13820), .B2(n20614), .ZN(
        P2_U2816) );
  AND2_X1 U17293 ( .A1(n20606), .A2(n17141), .ZN(n13824) );
  INV_X1 U17294 ( .A(n13831), .ZN(n13829) );
  AOI211_X1 U17295 ( .C1(P2_MEMORYFETCH_REG_SCAN_IN), .C2(n16368), .A(n13824), 
        .B(n13829), .ZN(n13822) );
  INV_X1 U17296 ( .A(n13822), .ZN(P2_U2814) );
  INV_X1 U17297 ( .A(n13823), .ZN(n20610) );
  OAI21_X1 U17298 ( .B1(n13824), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n20610), 
        .ZN(n13825) );
  OAI21_X1 U17299 ( .B1(n20619), .B2(n20610), .A(n13825), .ZN(P2_U3612) );
  NAND2_X1 U17300 ( .A1(n20619), .A2(n20618), .ZN(n13827) );
  INV_X1 U17301 ( .A(n14574), .ZN(n13826) );
  AOI211_X1 U17302 ( .C1(n20613), .C2(n13827), .A(n13826), .B(n9805), .ZN(
        n14575) );
  INV_X1 U17303 ( .A(n14601), .ZN(n14226) );
  NOR2_X1 U17304 ( .A1(n14575), .A2(n14226), .ZN(n20604) );
  OAI21_X1 U17305 ( .B1(n20604), .B2(n17498), .A(n13828), .ZN(P2_U2819) );
  INV_X1 U17306 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13835) );
  INV_X1 U17307 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13834) );
  OAI21_X2 U17308 ( .B1(n9593), .B2(n20613), .A(n13829), .ZN(n13863) );
  INV_X1 U17309 ( .A(n13863), .ZN(n13877) );
  NAND2_X1 U17310 ( .A1(n20620), .A2(n20613), .ZN(n13830) );
  INV_X1 U17311 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n13833) );
  INV_X1 U17312 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13832) );
  MUX2_X1 U17313 ( .A(n13833), .B(n13832), .S(n19839), .Z(n16551) );
  OAI222_X1 U17314 ( .A1(n13929), .A2(n13835), .B1(n13834), .B2(n13877), .C1(
        n13836), .C2(n16551), .ZN(P2_U2982) );
  INV_X1 U17315 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13964) );
  INV_X1 U17316 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n13838) );
  NAND2_X1 U17317 ( .A1(n19839), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13837) );
  OAI21_X1 U17318 ( .B1(n19839), .B2(n13838), .A(n13837), .ZN(n19898) );
  NAND2_X1 U17319 ( .A1(n13897), .A2(n19898), .ZN(n13899) );
  NAND2_X1 U17320 ( .A1(n13863), .A2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13839) );
  OAI211_X1 U17321 ( .C1(n13929), .C2(n13964), .A(n13899), .B(n13839), .ZN(
        P2_U2959) );
  INV_X1 U17322 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n21593) );
  NAND2_X1 U17323 ( .A1(n19837), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13841) );
  NAND2_X1 U17324 ( .A1(n19839), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13840) );
  AND2_X1 U17325 ( .A1(n13841), .A2(n13840), .ZN(n19849) );
  INV_X1 U17326 ( .A(n19849), .ZN(n16542) );
  NAND2_X1 U17327 ( .A1(n13897), .A2(n16542), .ZN(n13906) );
  NAND2_X1 U17328 ( .A1(n13863), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13842) );
  OAI211_X1 U17329 ( .C1(n13929), .C2(n21593), .A(n13906), .B(n13842), .ZN(
        P2_U2952) );
  INV_X1 U17330 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13934) );
  INV_X1 U17331 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n13844) );
  NAND2_X1 U17332 ( .A1(n19839), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13843) );
  OAI21_X1 U17333 ( .B1(n19839), .B2(n13844), .A(n13843), .ZN(n16456) );
  NAND2_X1 U17334 ( .A1(n13897), .A2(n16456), .ZN(n13901) );
  NAND2_X1 U17335 ( .A1(n13863), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13845) );
  OAI211_X1 U17336 ( .C1(n13929), .C2(n13934), .A(n13901), .B(n13845), .ZN(
        P2_U2963) );
  INV_X1 U17337 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13968) );
  MUX2_X1 U17338 ( .A(BUF2_REG_10__SCAN_IN), .B(BUF1_REG_10__SCAN_IN), .S(
        n19839), .Z(n16464) );
  NAND2_X1 U17339 ( .A1(n13897), .A2(n16464), .ZN(n13891) );
  NAND2_X1 U17340 ( .A1(n13863), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13846) );
  OAI211_X1 U17341 ( .C1(n13929), .C2(n13968), .A(n13891), .B(n13846), .ZN(
        P2_U2962) );
  INV_X1 U17342 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13936) );
  INV_X1 U17343 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n13848) );
  NAND2_X1 U17344 ( .A1(n19839), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13847) );
  OAI21_X1 U17345 ( .B1(n19839), .B2(n13848), .A(n13847), .ZN(n16443) );
  NAND2_X1 U17346 ( .A1(n13897), .A2(n16443), .ZN(n13878) );
  NAND2_X1 U17347 ( .A1(n13863), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13849) );
  OAI211_X1 U17348 ( .C1(n13929), .C2(n13936), .A(n13878), .B(n13849), .ZN(
        P2_U2965) );
  INV_X1 U17349 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13981) );
  INV_X1 U17350 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n13851) );
  NAND2_X1 U17351 ( .A1(n19839), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13850) );
  OAI21_X1 U17352 ( .B1(n19839), .B2(n13851), .A(n13850), .ZN(n16473) );
  NAND2_X1 U17353 ( .A1(n13897), .A2(n16473), .ZN(n13903) );
  NAND2_X1 U17354 ( .A1(n13863), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13852) );
  OAI211_X1 U17355 ( .C1(n13929), .C2(n13981), .A(n13903), .B(n13852), .ZN(
        P2_U2961) );
  INV_X1 U17356 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19806) );
  NAND2_X1 U17357 ( .A1(n13897), .A2(n16553), .ZN(n13862) );
  NAND2_X1 U17358 ( .A1(n13863), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13853) );
  OAI211_X1 U17359 ( .C1(n19806), .C2(n13929), .A(n13862), .B(n13853), .ZN(
        P2_U2981) );
  INV_X1 U17360 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13966) );
  INV_X1 U17361 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n13855) );
  NAND2_X1 U17362 ( .A1(n19839), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13854) );
  OAI21_X1 U17363 ( .B1(n19839), .B2(n13855), .A(n13854), .ZN(n16480) );
  NAND2_X1 U17364 ( .A1(n13897), .A2(n16480), .ZN(n13865) );
  NAND2_X1 U17365 ( .A1(n13863), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13856) );
  OAI211_X1 U17366 ( .C1(n13966), .C2(n13929), .A(n13865), .B(n13856), .ZN(
        P2_U2960) );
  INV_X1 U17367 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19810) );
  INV_X1 U17368 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18494) );
  NAND2_X1 U17369 ( .A1(n19839), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13857) );
  OAI21_X1 U17370 ( .B1(n19839), .B2(n18494), .A(n13857), .ZN(n16449) );
  NAND2_X1 U17371 ( .A1(n13897), .A2(n16449), .ZN(n13860) );
  NAND2_X1 U17372 ( .A1(n13863), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13858) );
  OAI211_X1 U17373 ( .C1(n19810), .C2(n13929), .A(n13860), .B(n13858), .ZN(
        P2_U2979) );
  INV_X1 U17374 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13932) );
  NAND2_X1 U17375 ( .A1(n13863), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13859) );
  OAI211_X1 U17376 ( .C1(n13932), .C2(n13929), .A(n13860), .B(n13859), .ZN(
        P2_U2964) );
  INV_X1 U17377 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13938) );
  NAND2_X1 U17378 ( .A1(n13863), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13861) );
  OAI211_X1 U17379 ( .C1(n13938), .C2(n13929), .A(n13862), .B(n13861), .ZN(
        P2_U2966) );
  INV_X1 U17380 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19818) );
  NAND2_X1 U17381 ( .A1(n13863), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13864) );
  OAI211_X1 U17382 ( .C1(n19818), .C2(n13929), .A(n13865), .B(n13864), .ZN(
        P2_U2975) );
  INV_X1 U17383 ( .A(n13866), .ZN(n13923) );
  INV_X1 U17384 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n13867) );
  AND2_X1 U17385 ( .A1(n14448), .A2(n10478), .ZN(n13922) );
  OAI21_X1 U17386 ( .B1(n13923), .B2(n13867), .A(n13922), .ZN(P1_U2801) );
  OAI22_X1 U17387 ( .A1(n14374), .A2(n15253), .B1(n10102), .B2(n13869), .ZN(
        n13940) );
  OAI21_X1 U17388 ( .B1(n13940), .B2(n15940), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n13870) );
  OAI21_X1 U17389 ( .B1(n10478), .B2(n14376), .A(n13870), .ZN(P1_U2803) );
  OAI21_X1 U17390 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16356), .A(
        n13953), .ZN(n13990) );
  OAI21_X1 U17391 ( .B1(n13872), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13871), .ZN(n13989) );
  NAND2_X1 U17392 ( .A1(n16837), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13995) );
  OAI21_X1 U17393 ( .B1(n16846), .B2(n13989), .A(n13995), .ZN(n13873) );
  AOI21_X1 U17394 ( .B1(n16366), .B2(n16827), .A(n13873), .ZN(n13876) );
  OAI21_X1 U17395 ( .B1(n16858), .B2(n13874), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13875) );
  OAI211_X1 U17396 ( .C1(n13990), .C2(n16863), .A(n13876), .B(n13875), .ZN(
        P2_U3014) );
  AOI22_X1 U17397 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13879) );
  NAND2_X1 U17398 ( .A1(n13879), .A2(n13878), .ZN(P2_U2980) );
  AOI22_X1 U17399 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13882) );
  INV_X1 U17400 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n13881) );
  NAND2_X1 U17401 ( .A1(n19839), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13880) );
  OAI21_X1 U17402 ( .B1(n19839), .B2(n13881), .A(n13880), .ZN(n19886) );
  NAND2_X1 U17403 ( .A1(n13897), .A2(n19886), .ZN(n13915) );
  NAND2_X1 U17404 ( .A1(n13882), .A2(n13915), .ZN(P2_U2973) );
  AOI22_X1 U17405 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13884) );
  NAND2_X1 U17406 ( .A1(n19839), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13883) );
  OAI21_X1 U17407 ( .B1(n19839), .B2(n19149), .A(n13883), .ZN(n19864) );
  NAND2_X1 U17408 ( .A1(n13897), .A2(n19864), .ZN(n13917) );
  NAND2_X1 U17409 ( .A1(n13884), .A2(n13917), .ZN(P2_U2969) );
  AOI22_X1 U17410 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13887) );
  NAND2_X1 U17411 ( .A1(n19837), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13886) );
  NAND2_X1 U17412 ( .A1(n19839), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13885) );
  AND2_X1 U17413 ( .A1(n13886), .A2(n13885), .ZN(n19877) );
  INV_X1 U17414 ( .A(n19877), .ZN(n16510) );
  NAND2_X1 U17415 ( .A1(n13897), .A2(n16510), .ZN(n13913) );
  NAND2_X1 U17416 ( .A1(n13887), .A2(n13913), .ZN(P2_U2971) );
  AOI22_X1 U17417 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13890) );
  NAND2_X1 U17418 ( .A1(n19837), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13889) );
  NAND2_X1 U17419 ( .A1(n19839), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13888) );
  AND2_X1 U17420 ( .A1(n13889), .A2(n13888), .ZN(n19871) );
  INV_X1 U17421 ( .A(n19871), .ZN(n16519) );
  NAND2_X1 U17422 ( .A1(n13897), .A2(n16519), .ZN(n13911) );
  NAND2_X1 U17423 ( .A1(n13890), .A2(n13911), .ZN(P2_U2970) );
  AOI22_X1 U17424 ( .A1(P2_LWORD_REG_10__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n13892) );
  NAND2_X1 U17425 ( .A1(n13892), .A2(n13891), .ZN(P2_U2977) );
  AOI22_X1 U17426 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13894) );
  INV_X1 U17427 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n19143) );
  NAND2_X1 U17428 ( .A1(n19839), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13893) );
  OAI21_X1 U17429 ( .B1(n19839), .B2(n19143), .A(n13893), .ZN(n19859) );
  NAND2_X1 U17430 ( .A1(n13897), .A2(n19859), .ZN(n13909) );
  NAND2_X1 U17431 ( .A1(n13894), .A2(n13909), .ZN(P2_U2968) );
  AOI22_X1 U17432 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13898) );
  INV_X1 U17433 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n13896) );
  NAND2_X1 U17434 ( .A1(n19839), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13895) );
  OAI21_X1 U17435 ( .B1(n19839), .B2(n13896), .A(n13895), .ZN(n19881) );
  NAND2_X1 U17436 ( .A1(n13897), .A2(n19881), .ZN(n13920) );
  NAND2_X1 U17437 ( .A1(n13898), .A2(n13920), .ZN(P2_U2972) );
  AOI22_X1 U17438 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13900) );
  NAND2_X1 U17439 ( .A1(n13900), .A2(n13899), .ZN(P2_U2974) );
  AOI22_X1 U17440 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13902) );
  NAND2_X1 U17441 ( .A1(n13902), .A2(n13901), .ZN(P2_U2978) );
  AOI22_X1 U17442 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13904) );
  NAND2_X1 U17443 ( .A1(n13904), .A2(n13903), .ZN(P2_U2976) );
  AOI22_X1 U17444 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n13918), .B1(n13905), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13907) );
  NAND2_X1 U17445 ( .A1(n13907), .A2(n13906), .ZN(P2_U2967) );
  INV_X1 U17446 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13975) );
  NAND2_X1 U17447 ( .A1(n13918), .A2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13908) );
  OAI211_X1 U17448 ( .C1(n13929), .C2(n13975), .A(n13909), .B(n13908), .ZN(
        P2_U2953) );
  INV_X1 U17449 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13972) );
  NAND2_X1 U17450 ( .A1(n13918), .A2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13910) );
  OAI211_X1 U17451 ( .C1(n13929), .C2(n13972), .A(n13911), .B(n13910), .ZN(
        P2_U2955) );
  INV_X1 U17452 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13962) );
  NAND2_X1 U17453 ( .A1(n13918), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13912) );
  OAI211_X1 U17454 ( .C1(n13929), .C2(n13962), .A(n13913), .B(n13912), .ZN(
        P2_U2956) );
  INV_X1 U17455 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13978) );
  NAND2_X1 U17456 ( .A1(n13918), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13914) );
  OAI211_X1 U17457 ( .C1(n13929), .C2(n13978), .A(n13915), .B(n13914), .ZN(
        P2_U2958) );
  INV_X1 U17458 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n21571) );
  NAND2_X1 U17459 ( .A1(n13918), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13916) );
  OAI211_X1 U17460 ( .C1(n13929), .C2(n21571), .A(n13917), .B(n13916), .ZN(
        P2_U2954) );
  INV_X1 U17461 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13970) );
  NAND2_X1 U17462 ( .A1(n13918), .A2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13919) );
  OAI211_X1 U17463 ( .C1(n13929), .C2(n13970), .A(n13920), .B(n13919), .ZN(
        P2_U2957) );
  INV_X1 U17464 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n13921) );
  NAND2_X1 U17465 ( .A1(n13922), .A2(n13921), .ZN(n13924) );
  INV_X1 U17466 ( .A(n13924), .ZN(n13926) );
  OAI22_X1 U17467 ( .A1(n13924), .A2(n13923), .B1(n15253), .B2(n10191), .ZN(
        n13925) );
  OAI21_X1 U17468 ( .B1(n13926), .B2(n21521), .A(n13925), .ZN(P1_U3487) );
  NAND2_X1 U17469 ( .A1(n14577), .A2(n14601), .ZN(n13927) );
  OR2_X1 U17470 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n21689), .ZN(n20611) );
  INV_X2 U17471 ( .A(n19828), .ZN(n19832) );
  AOI22_X1 U17472 ( .A1(n19833), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13931) );
  OAI21_X1 U17473 ( .B1(n13932), .B2(n13980), .A(n13931), .ZN(P2_U2923) );
  AOI22_X1 U17474 ( .A1(n19833), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13933) );
  OAI21_X1 U17475 ( .B1(n13934), .B2(n13980), .A(n13933), .ZN(P2_U2924) );
  AOI22_X1 U17476 ( .A1(n19833), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13935) );
  OAI21_X1 U17477 ( .B1(n13936), .B2(n13980), .A(n13935), .ZN(P2_U2922) );
  AOI22_X1 U17478 ( .A1(n19833), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13937) );
  OAI21_X1 U17479 ( .B1(n13938), .B2(n13980), .A(n13937), .ZN(P2_U2921) );
  NAND2_X1 U17480 ( .A1(n10084), .A2(n15260), .ZN(n13939) );
  INV_X1 U17481 ( .A(n21523), .ZN(n21447) );
  AOI21_X1 U17482 ( .B1(n13939), .B2(n15925), .A(n21447), .ZN(n21525) );
  NOR2_X1 U17483 ( .A1(n13940), .A2(n21525), .ZN(n15915) );
  NOR2_X1 U17484 ( .A1(n15915), .A2(n15940), .ZN(n20635) );
  INV_X1 U17485 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13951) );
  MUX2_X1 U17486 ( .A(n13944), .B(n13943), .S(n14013), .Z(n13948) );
  NOR2_X1 U17487 ( .A1(n13946), .A2(n13945), .ZN(n13947) );
  OAI21_X1 U17488 ( .B1(n13948), .B2(n13947), .A(n20885), .ZN(n15917) );
  INV_X1 U17489 ( .A(n15917), .ZN(n13949) );
  NAND2_X1 U17490 ( .A1(n20635), .A2(n13949), .ZN(n13950) );
  OAI21_X1 U17491 ( .B1(n20635), .B2(n13951), .A(n13950), .ZN(P1_U3484) );
  NAND2_X1 U17492 ( .A1(n16837), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n14054) );
  OAI21_X1 U17493 ( .B1(n16839), .B2(n16338), .A(n14054), .ZN(n13959) );
  XNOR2_X1 U17494 ( .A(n16334), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13952) );
  XNOR2_X1 U17495 ( .A(n13953), .B(n13952), .ZN(n14053) );
  INV_X1 U17496 ( .A(n14053), .ZN(n13957) );
  OR2_X1 U17497 ( .A1(n13954), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13956) );
  NAND2_X1 U17498 ( .A1(n13956), .A2(n13955), .ZN(n14057) );
  OAI22_X1 U17499 ( .A1(n16863), .A2(n13957), .B1(n16846), .B2(n14057), .ZN(
        n13958) );
  AOI211_X1 U17500 ( .C1(n16842), .C2(n16338), .A(n13959), .B(n13958), .ZN(
        n13960) );
  OAI21_X1 U17501 ( .B1(n10646), .B2(n19838), .A(n13960), .ZN(P2_U3013) );
  INV_X2 U17502 ( .A(n20611), .ZN(n19833) );
  AOI22_X1 U17503 ( .A1(n19833), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13961) );
  OAI21_X1 U17504 ( .B1(n13962), .B2(n13980), .A(n13961), .ZN(P2_U2931) );
  AOI22_X1 U17505 ( .A1(n19833), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13963) );
  OAI21_X1 U17506 ( .B1(n13964), .B2(n13980), .A(n13963), .ZN(P2_U2928) );
  AOI22_X1 U17507 ( .A1(n19833), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13965) );
  OAI21_X1 U17508 ( .B1(n13966), .B2(n13980), .A(n13965), .ZN(P2_U2927) );
  AOI22_X1 U17509 ( .A1(n19833), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13967) );
  OAI21_X1 U17510 ( .B1(n13968), .B2(n13980), .A(n13967), .ZN(P2_U2925) );
  AOI22_X1 U17511 ( .A1(n19833), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13969) );
  OAI21_X1 U17512 ( .B1(n13970), .B2(n13980), .A(n13969), .ZN(P2_U2930) );
  AOI22_X1 U17513 ( .A1(n19833), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13971) );
  OAI21_X1 U17514 ( .B1(n13972), .B2(n13980), .A(n13971), .ZN(P2_U2932) );
  AOI22_X1 U17515 ( .A1(n19833), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13973) );
  OAI21_X1 U17516 ( .B1(n21593), .B2(n13980), .A(n13973), .ZN(P2_U2935) );
  AOI22_X1 U17517 ( .A1(n19833), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13974) );
  OAI21_X1 U17518 ( .B1(n13975), .B2(n13980), .A(n13974), .ZN(P2_U2934) );
  AOI22_X1 U17519 ( .A1(n19833), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13976) );
  OAI21_X1 U17520 ( .B1(n21571), .B2(n13980), .A(n13976), .ZN(P2_U2933) );
  AOI22_X1 U17521 ( .A1(n19833), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13977) );
  OAI21_X1 U17522 ( .B1(n13978), .B2(n13980), .A(n13977), .ZN(P2_U2929) );
  AOI22_X1 U17523 ( .A1(n19833), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13979) );
  OAI21_X1 U17524 ( .B1(n13981), .B2(n13980), .A(n13979), .ZN(P2_U2926) );
  INV_X1 U17525 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19822) );
  INV_X1 U17526 ( .A(n13983), .ZN(n13984) );
  XNOR2_X1 U17527 ( .A(n13982), .B(n13984), .ZN(n17094) );
  INV_X1 U17528 ( .A(n17094), .ZN(n16272) );
  INV_X1 U17529 ( .A(n16543), .ZN(n13987) );
  INV_X1 U17530 ( .A(n13985), .ZN(n13986) );
  INV_X1 U17531 ( .A(n19886), .ZN(n13988) );
  OAI222_X1 U17532 ( .A1(n19822), .A2(n19795), .B1(n16272), .B2(n16565), .C1(
        n19803), .C2(n13988), .ZN(P2_U2913) );
  OAI22_X1 U17533 ( .A1(n17139), .A2(n13990), .B1(n17124), .B2(n13989), .ZN(
        n13997) );
  OR2_X1 U17534 ( .A1(n13992), .A2(n13991), .ZN(n13994) );
  AND2_X1 U17535 ( .A1(n13994), .A2(n13993), .ZN(n19800) );
  INV_X1 U17536 ( .A(n19800), .ZN(n16352) );
  OAI21_X1 U17537 ( .B1(n17134), .B2(n16352), .A(n13995), .ZN(n13996) );
  AOI211_X1 U17538 ( .C1(n16366), .C2(n17127), .A(n13997), .B(n13996), .ZN(
        n13999) );
  MUX2_X1 U17539 ( .A(n17098), .B(n14785), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13998) );
  NAND2_X1 U17540 ( .A1(n13999), .A2(n13998), .ZN(P2_U3046) );
  INV_X1 U17541 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19820) );
  OAI21_X1 U17542 ( .B1(n14002), .B2(n14001), .A(n14000), .ZN(n17086) );
  INV_X1 U17543 ( .A(n19898), .ZN(n14003) );
  OAI222_X1 U17544 ( .A1(n19820), .A2(n19795), .B1(n17086), .B2(n16565), .C1(
        n19803), .C2(n14003), .ZN(P2_U2912) );
  MUX2_X1 U17545 ( .A(n14008), .B(n10646), .S(n16430), .Z(n14009) );
  OAI21_X1 U17546 ( .B1(n20009), .B2(n16433), .A(n14009), .ZN(P2_U2886) );
  OAI21_X1 U17547 ( .B1(n21447), .B2(n15925), .A(n14010), .ZN(n14012) );
  INV_X1 U17548 ( .A(n14925), .ZN(n14339) );
  NAND3_X1 U17549 ( .A1(n14339), .A2(n14336), .A3(n14343), .ZN(n14011) );
  NAND2_X1 U17550 ( .A1(n14012), .A2(n14011), .ZN(n14014) );
  MUX2_X1 U17551 ( .A(n14014), .B(n14344), .S(n14013), .Z(n14019) );
  OAI21_X1 U17552 ( .B1(n15260), .B2(n20859), .A(n14015), .ZN(n14016) );
  NOR2_X1 U17553 ( .A1(n14017), .A2(n14016), .ZN(n14018) );
  NAND2_X1 U17554 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17555) );
  NAND2_X1 U17555 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14378), .ZN(n17560) );
  INV_X1 U17556 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20634) );
  OAI22_X1 U17557 ( .A1(n15906), .A2(n15940), .B1(n17560), .B2(n20634), .ZN(
        n14021) );
  AOI21_X1 U17558 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n14376), .A(n14021), 
        .ZN(n15900) );
  INV_X1 U17559 ( .A(n15900), .ZN(n14929) );
  INV_X1 U17560 ( .A(n20995), .ZN(n21237) );
  XNOR2_X1 U17561 ( .A(n14020), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n15262) );
  INV_X1 U17562 ( .A(n14335), .ZN(n14366) );
  NAND4_X1 U17563 ( .A1(n15262), .A2(n14926), .A3(n14366), .A4(n14021), .ZN(
        n14022) );
  OAI21_X1 U17564 ( .B1(n14929), .B2(n14369), .A(n14022), .ZN(P1_U3468) );
  NAND2_X1 U17565 ( .A1(n19589), .A2(n19617), .ZN(n14026) );
  NOR2_X1 U17566 ( .A1(n19736), .A2(n10217), .ZN(n19614) );
  NAND2_X1 U17567 ( .A1(n19592), .A2(n14024), .ZN(n14504) );
  OAI211_X1 U17568 ( .C1(n14026), .C2(n18537), .A(n14025), .B(n14504), .ZN(
        n14027) );
  NOR2_X1 U17569 ( .A1(n14501), .A2(n14027), .ZN(n19602) );
  OR2_X1 U17570 ( .A1(n19602), .A2(n19623), .ZN(n14029) );
  NAND2_X1 U17571 ( .A1(n19740), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19139) );
  INV_X1 U17572 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19128) );
  NAND3_X1 U17573 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19721)
         );
  OR2_X1 U17574 ( .A1(n19128), .A2(n19721), .ZN(n17480) );
  AND2_X1 U17575 ( .A1(n19139), .A2(n17480), .ZN(n14028) );
  NAND2_X1 U17576 ( .A1(n14029), .A2(n14028), .ZN(n17489) );
  NOR2_X1 U17577 ( .A1(n14508), .A2(n18998), .ZN(n14035) );
  MUX2_X1 U17578 ( .A(n14035), .B(n17314), .S(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n19571) );
  INV_X1 U17579 ( .A(n19571), .ZN(n19572) );
  INV_X1 U17580 ( .A(n18043), .ZN(n17487) );
  INV_X1 U17581 ( .A(n19612), .ZN(n17359) );
  OAI22_X1 U17582 ( .A1(n17359), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18536), .ZN(n14030) );
  AOI21_X1 U17583 ( .B1(n19572), .B2(n17487), .A(n14030), .ZN(n14032) );
  NAND2_X1 U17584 ( .A1(n14076), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14031) );
  OAI21_X1 U17585 ( .B1(n14076), .B2(n14032), .A(n14031), .ZN(P3_U3290) );
  NOR2_X1 U17586 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19122), .ZN(
        n14063) );
  INV_X1 U17587 ( .A(n14033), .ZN(n14034) );
  INV_X1 U17588 ( .A(n17351), .ZN(n14061) );
  NAND2_X1 U17589 ( .A1(n14034), .A2(n14061), .ZN(n14249) );
  OAI22_X1 U17590 ( .A1(n14063), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n14035), .B2(n14249), .ZN(n19574) );
  INV_X1 U17591 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14750) );
  AOI22_X1 U17592 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n11902), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14750), .ZN(n17358) );
  NAND2_X1 U17593 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17357) );
  INV_X1 U17594 ( .A(n17357), .ZN(n14037) );
  INV_X1 U17595 ( .A(n14249), .ZN(n14036) );
  AOI222_X1 U17596 ( .A1(n19574), .A2(n17487), .B1(n17358), .B2(n14037), .C1(
        n14036), .C2(n19612), .ZN(n14039) );
  NAND2_X1 U17597 ( .A1(n14076), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14038) );
  OAI21_X1 U17598 ( .B1(n14039), .B2(n14076), .A(n14038), .ZN(P3_U3289) );
  AOI21_X1 U17599 ( .B1(n14041), .B2(n14000), .A(n11364), .ZN(n17072) );
  INV_X1 U17600 ( .A(n17072), .ZN(n14043) );
  AOI22_X1 U17601 ( .A1(n19793), .A2(n16480), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19796), .ZN(n14042) );
  OAI21_X1 U17602 ( .B1(n14043), .B2(n16565), .A(n14042), .ZN(P2_U2911) );
  NAND2_X1 U17603 ( .A1(n17491), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14045) );
  NAND4_X1 U17604 ( .A1(n14046), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14045), 
        .A4(n20607), .ZN(n14047) );
  MUX2_X1 U17605 ( .A(n13350), .B(n16349), .S(n16438), .Z(n14048) );
  OAI21_X1 U17606 ( .B1(n21692), .B2(n16433), .A(n14048), .ZN(P2_U2887) );
  INV_X1 U17607 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14692) );
  AOI211_X1 U17608 ( .C1(n14056), .C2(n14692), .A(n14788), .B(n17098), .ZN(
        n14060) );
  OR2_X1 U17609 ( .A1(n14051), .A2(n14050), .ZN(n14052) );
  NAND2_X1 U17610 ( .A1(n14049), .A2(n14052), .ZN(n20589) );
  INV_X1 U17611 ( .A(n20589), .ZN(n16557) );
  AOI22_X1 U17612 ( .A1(n9574), .A2(n17127), .B1(n14053), .B2(n9563), .ZN(
        n14055) );
  OAI211_X1 U17613 ( .C1(n16557), .C2(n17134), .A(n14055), .B(n14054), .ZN(
        n14059) );
  OAI22_X1 U17614 ( .A1(n17124), .A2(n14057), .B1(n14785), .B2(n14056), .ZN(
        n14058) );
  OR3_X1 U17615 ( .A1(n14060), .A2(n14059), .A3(n14058), .ZN(P2_U3045) );
  NAND2_X1 U17616 ( .A1(n14061), .A2(n17346), .ZN(n17343) );
  INV_X1 U17617 ( .A(n17343), .ZN(n14062) );
  OAI22_X1 U17618 ( .A1(n14063), .A2(n14065), .B1(n14062), .B2(n18971), .ZN(
        n19599) );
  NOR2_X1 U17619 ( .A1(n18043), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14067) );
  NOR2_X1 U17620 ( .A1(n14065), .A2(n14064), .ZN(n14071) );
  NOR2_X1 U17621 ( .A1(n14071), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14066) );
  NOR2_X1 U17622 ( .A1(n9560), .A2(n14066), .ZN(n18005) );
  AOI22_X1 U17623 ( .A1(n19599), .A2(n14067), .B1(n19612), .B2(n18005), .ZN(
        n14077) );
  OAI21_X1 U17624 ( .B1(n14070), .B2(n14069), .A(n14068), .ZN(n17349) );
  INV_X1 U17625 ( .A(n14071), .ZN(n17344) );
  OAI21_X1 U17626 ( .B1(n17314), .B2(n11564), .A(n17343), .ZN(n14072) );
  AOI21_X1 U17627 ( .B1(n17349), .B2(n17344), .A(n14072), .ZN(n19600) );
  NOR2_X1 U17628 ( .A1(n19600), .A2(n18043), .ZN(n14073) );
  NOR2_X1 U17629 ( .A1(n14073), .A2(n14076), .ZN(n14075) );
  OAI22_X1 U17630 ( .A1(n14077), .A2(n14076), .B1(n14075), .B2(n14074), .ZN(
        P3_U3285) );
  NAND2_X1 U17631 ( .A1(n14040), .A2(n14079), .ZN(n14080) );
  AND2_X1 U17632 ( .A1(n14078), .A2(n14080), .ZN(n17061) );
  INV_X1 U17633 ( .A(n17061), .ZN(n16234) );
  INV_X1 U17634 ( .A(n16473), .ZN(n14081) );
  INV_X1 U17635 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19816) );
  OAI222_X1 U17636 ( .A1(n16234), .A2(n16565), .B1(n14081), .B2(n19803), .C1(
        n19816), .C2(n19795), .ZN(P2_U2910) );
  INV_X1 U17637 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14097) );
  NOR2_X1 U17638 ( .A1(n19020), .A2(n11902), .ZN(n14083) );
  AOI21_X1 U17639 ( .B1(n14083), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n14082), .ZN(n14090) );
  XNOR2_X1 U17640 ( .A(n14085), .B(n14084), .ZN(n18903) );
  OAI21_X1 U17641 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17336), .A(
        n17306), .ZN(n14086) );
  AOI22_X1 U17642 ( .A1(n19585), .A2(n18903), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14086), .ZN(n14089) );
  NAND3_X1 U17643 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14087), .A3(
        n14097), .ZN(n14088) );
  OAI211_X1 U17644 ( .C1(n14090), .C2(n18971), .A(n14089), .B(n14088), .ZN(
        n14091) );
  NAND2_X1 U17645 ( .A1(n14091), .A2(n19053), .ZN(n14096) );
  XNOR2_X1 U17646 ( .A(n14092), .B(n14093), .ZN(n18898) );
  INV_X1 U17647 ( .A(n18898), .ZN(n14094) );
  INV_X1 U17648 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19653) );
  NOR2_X1 U17649 ( .A1(n19120), .A2(n19653), .ZN(n18902) );
  AOI21_X1 U17650 ( .B1(n17301), .B2(n14094), .A(n18902), .ZN(n14095) );
  OAI211_X1 U17651 ( .C1(n19114), .C2(n14097), .A(n14096), .B(n14095), .ZN(
        P3_U2860) );
  MUX2_X1 U17652 ( .A(n13361), .B(P2_EBX_REG_2__SCAN_IN), .S(n16438), .Z(
        n14101) );
  AOI21_X1 U17653 ( .B1(n20578), .B2(n16435), .A(n14101), .ZN(n14102) );
  INV_X1 U17654 ( .A(n14102), .ZN(P2_U2885) );
  INV_X1 U17655 ( .A(n14103), .ZN(n14106) );
  OAI21_X1 U17656 ( .B1(n14106), .B2(n14105), .A(n14104), .ZN(n15301) );
  OAI21_X1 U17657 ( .B1(n14108), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14107), .ZN(n14184) );
  NAND2_X1 U17658 ( .A1(n20666), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14178) );
  OAI21_X1 U17659 ( .B1(n20772), .B2(n14109), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14110) );
  OAI211_X1 U17660 ( .C1(n14184), .C2(n20633), .A(n14178), .B(n14110), .ZN(
        n14111) );
  INV_X1 U17661 ( .A(n14111), .ZN(n14112) );
  OAI21_X1 U17662 ( .B1(n20837), .B2(n15301), .A(n14112), .ZN(P1_U2999) );
  AOI21_X1 U17663 ( .B1(n14114), .B2(n15883), .A(n14113), .ZN(n15293) );
  INV_X1 U17664 ( .A(n20712), .ZN(n15320) );
  AOI22_X1 U17665 ( .A1(n20707), .A2(n15293), .B1(P1_EBX_REG_0__SCAN_IN), .B2(
        n15320), .ZN(n14115) );
  OAI21_X1 U17666 ( .B1(n15301), .B2(n15330), .A(n14115), .ZN(P1_U2872) );
  AOI21_X1 U17667 ( .B1(n14118), .B2(n14117), .A(n14116), .ZN(n18892) );
  XNOR2_X1 U17668 ( .A(n14119), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18888) );
  NAND2_X1 U17669 ( .A1(n19008), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14121) );
  INV_X1 U17670 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19655) );
  NOR2_X1 U17671 ( .A1(n19055), .A2(n19655), .ZN(n18891) );
  INV_X1 U17672 ( .A(n18891), .ZN(n14120) );
  OAI211_X1 U17673 ( .C1(n19115), .C2(n18888), .A(n14121), .B(n14120), .ZN(
        n14124) );
  AOI211_X1 U17674 ( .C1(n18981), .C2(n9934), .A(n14122), .B(n19121), .ZN(
        n14123) );
  AOI211_X1 U17675 ( .C1(n19119), .C2(n18892), .A(n14124), .B(n14123), .ZN(
        n14125) );
  INV_X1 U17676 ( .A(n14125), .ZN(P3_U2859) );
  OR2_X1 U17677 ( .A1(n12106), .A2(n12036), .ZN(n14127) );
  INV_X1 U17678 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20742) );
  INV_X1 U17679 ( .A(n14127), .ZN(n14128) );
  NAND2_X1 U17680 ( .A1(n20836), .A2(DATAI_0_), .ZN(n14130) );
  NAND2_X1 U17681 ( .A1(n20838), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14129) );
  AND2_X1 U17682 ( .A1(n14130), .A2(n14129), .ZN(n20847) );
  OAI222_X1 U17683 ( .A1(n15301), .A2(n15415), .B1(n15413), .B2(n20742), .C1(
        n15412), .C2(n20847), .ZN(P1_U2904) );
  OAI21_X1 U17684 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(n15292) );
  INV_X1 U17685 ( .A(DATAI_1_), .ZN(n14135) );
  NAND2_X1 U17686 ( .A1(n20838), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14134) );
  OAI21_X1 U17687 ( .B1(n20838), .B2(n14135), .A(n14134), .ZN(n20856) );
  INV_X1 U17688 ( .A(n20856), .ZN(n14136) );
  OAI222_X1 U17689 ( .A1(n15292), .A2(n15415), .B1(n15413), .B2(n12211), .C1(
        n15412), .C2(n14136), .ZN(P1_U2903) );
  INV_X1 U17690 ( .A(n19859), .ZN(n14141) );
  XNOR2_X1 U17691 ( .A(n20009), .B(n20589), .ZN(n14137) );
  NAND2_X1 U17692 ( .A1(n19840), .A2(n19800), .ZN(n19799) );
  NAND2_X1 U17693 ( .A1(n14137), .A2(n19799), .ZN(n16558) );
  OAI21_X1 U17694 ( .B1(n14137), .B2(n19799), .A(n16558), .ZN(n14138) );
  INV_X1 U17695 ( .A(n16562), .ZN(n19798) );
  NAND2_X1 U17696 ( .A1(n14138), .A2(n19798), .ZN(n14140) );
  AOI22_X1 U17697 ( .A1(n19797), .A2(n20589), .B1(n19796), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n14139) );
  OAI211_X1 U17698 ( .C1(n19803), .C2(n14141), .A(n14140), .B(n14139), .ZN(
        P2_U2918) );
  INV_X1 U17699 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14143) );
  XNOR2_X1 U17700 ( .A(n14142), .B(n14934), .ZN(n15282) );
  OAI222_X1 U17701 ( .A1(n15330), .A2(n15292), .B1(n14143), .B2(n20712), .C1(
        n15328), .C2(n15282), .ZN(P1_U2871) );
  XNOR2_X1 U17702 ( .A(n14145), .B(n14278), .ZN(n17264) );
  INV_X1 U17703 ( .A(n17264), .ZN(n14150) );
  AOI211_X1 U17704 ( .C1(n17314), .C2(n19020), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n17276), .ZN(n14148) );
  OR3_X1 U17705 ( .A1(n19121), .A2(n19029), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19124) );
  AOI21_X1 U17706 ( .B1(n19114), .B2(n19124), .A(n11902), .ZN(n14147) );
  XNOR2_X1 U17707 ( .A(n14145), .B(n14144), .ZN(n17262) );
  NAND2_X1 U17708 ( .A1(n19089), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n17260) );
  OAI21_X1 U17709 ( .B1(n19115), .B2(n17262), .A(n17260), .ZN(n14146) );
  NOR3_X1 U17710 ( .A1(n14148), .A2(n14147), .A3(n14146), .ZN(n14149) );
  OAI21_X1 U17711 ( .B1(n19044), .B2(n14150), .A(n14149), .ZN(P3_U2861) );
  AOI21_X1 U17712 ( .B1(n9748), .B2(n14152), .A(n14151), .ZN(n18873) );
  INV_X1 U17713 ( .A(n18873), .ZN(n14162) );
  AND2_X1 U17714 ( .A1(n14153), .A2(n17306), .ZN(n14154) );
  OAI22_X1 U17715 ( .A1(n14155), .A2(n18971), .B1(n17336), .B2(n14154), .ZN(
        n14389) );
  INV_X1 U17716 ( .A(n14389), .ZN(n14156) );
  OAI21_X1 U17717 ( .B1(n14156), .B2(n19121), .A(n19114), .ZN(n14174) );
  OR2_X1 U17718 ( .A1(n19121), .A2(n18981), .ZN(n14388) );
  NOR3_X1 U17719 ( .A1(n9934), .A2(n14157), .A3(n14388), .ZN(n14158) );
  AOI22_X1 U17720 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14174), .B1(
        n14158), .B2(n9939), .ZN(n14161) );
  XOR2_X1 U17721 ( .A(n14159), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18870) );
  AOI22_X1 U17722 ( .A1(n17301), .A2(n18870), .B1(n19089), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n14160) );
  OAI211_X1 U17723 ( .C1(n19044), .C2(n14162), .A(n14161), .B(n14160), .ZN(
        P3_U2857) );
  AOI21_X1 U17724 ( .B1(n14165), .B2(n14078), .A(n14164), .ZN(n17049) );
  INV_X1 U17725 ( .A(n17049), .ZN(n14167) );
  INV_X1 U17726 ( .A(n16464), .ZN(n14166) );
  INV_X1 U17727 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19814) );
  OAI222_X1 U17728 ( .A1(n14167), .A2(n16565), .B1(n14166), .B2(n19803), .C1(
        n19814), .C2(n19795), .ZN(P2_U2909) );
  AOI21_X1 U17729 ( .B1(n14169), .B2(n14390), .A(n14168), .ZN(n18867) );
  INV_X1 U17730 ( .A(n18867), .ZN(n14177) );
  NOR3_X1 U17731 ( .A1(n18981), .A2(n18980), .A3(n19121), .ZN(n14173) );
  XNOR2_X1 U17732 ( .A(n14171), .B(n14170), .ZN(n18862) );
  OAI22_X1 U17733 ( .A1(n19115), .A2(n18862), .B1(n19120), .B2(n19660), .ZN(
        n14172) );
  AOI21_X1 U17734 ( .B1(n14173), .B2(n14390), .A(n14172), .ZN(n14176) );
  NAND2_X1 U17735 ( .A1(n14174), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14175) );
  OAI211_X1 U17736 ( .C1(n14177), .C2(n19044), .A(n14176), .B(n14175), .ZN(
        P3_U2856) );
  INV_X1 U17737 ( .A(n14178), .ZN(n14182) );
  AOI21_X1 U17738 ( .B1(n20811), .B2(n15883), .A(n15817), .ZN(n20833) );
  INV_X1 U17739 ( .A(n20811), .ZN(n14179) );
  AND3_X1 U17740 ( .A1(n14179), .A2(n15883), .A3(n15703), .ZN(n14180) );
  AOI21_X1 U17741 ( .B1(n20833), .B2(n15802), .A(n14180), .ZN(n14181) );
  AOI211_X1 U17742 ( .C1(n20823), .C2(n15293), .A(n14182), .B(n14181), .ZN(
        n14183) );
  OAI21_X1 U17743 ( .B1(n15862), .B2(n14184), .A(n14183), .ZN(P1_U3031) );
  AND2_X1 U17744 ( .A1(n14186), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14187) );
  NAND2_X1 U17745 ( .A1(n14185), .A2(n14187), .ZN(n14237) );
  OR2_X1 U17746 ( .A1(n14185), .A2(n14187), .ZN(n14188) );
  NAND2_X1 U17747 ( .A1(n14237), .A2(n14188), .ZN(n19779) );
  NAND2_X1 U17748 ( .A1(n14191), .A2(n14190), .ZN(n14192) );
  NAND2_X1 U17749 ( .A1(n14189), .A2(n14192), .ZN(n16860) );
  NOR2_X1 U17750 ( .A1(n16860), .A2(n16438), .ZN(n14193) );
  AOI21_X1 U17751 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n16438), .A(n14193), .ZN(
        n14194) );
  OAI21_X1 U17752 ( .B1(n19779), .B2(n16433), .A(n14194), .ZN(P2_U2883) );
  OAI21_X1 U17753 ( .B1(n14164), .B2(n14195), .A(n10348), .ZN(n17036) );
  INV_X1 U17754 ( .A(n16456), .ZN(n14196) );
  INV_X1 U17755 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19812) );
  OAI222_X1 U17756 ( .A1(n17036), .A2(n16565), .B1(n14196), .B2(n19803), .C1(
        n19812), .C2(n19795), .ZN(P2_U2908) );
  INV_X1 U17757 ( .A(n20567), .ZN(n20177) );
  INV_X1 U17758 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n21574) );
  MUX2_X1 U17759 ( .A(n21574), .B(n10648), .S(n16430), .Z(n14200) );
  OAI21_X1 U17760 ( .B1(n20177), .B2(n16433), .A(n14200), .ZN(P2_U2884) );
  AND2_X1 U17761 ( .A1(n14570), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17151) );
  AOI21_X1 U17762 ( .B1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n17154), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14201) );
  NOR2_X1 U17763 ( .A1(n14202), .A2(n14201), .ZN(n14205) );
  NAND2_X1 U17764 ( .A1(n11236), .A2(n14203), .ZN(n14537) );
  OAI21_X1 U17765 ( .B1(n13511), .B2(n10669), .A(n10733), .ZN(n14204) );
  AOI22_X1 U17766 ( .A1(n11235), .A2(n14205), .B1(n14537), .B2(n14204), .ZN(
        n14214) );
  INV_X1 U17767 ( .A(n14206), .ZN(n14572) );
  AND2_X1 U17768 ( .A1(n14572), .A2(n14571), .ZN(n14539) );
  INV_X1 U17769 ( .A(n14556), .ZN(n14207) );
  NAND2_X1 U17770 ( .A1(n14207), .A2(n14541), .ZN(n14536) );
  INV_X1 U17771 ( .A(n14536), .ZN(n14208) );
  NOR2_X1 U17772 ( .A1(n14539), .A2(n14208), .ZN(n14211) );
  INV_X1 U17773 ( .A(n14539), .ZN(n14209) );
  NAND2_X1 U17774 ( .A1(n14209), .A2(n14208), .ZN(n14544) );
  INV_X1 U17775 ( .A(n14544), .ZN(n14210) );
  MUX2_X1 U17776 ( .A(n14211), .B(n14210), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14212) );
  INV_X1 U17777 ( .A(n14212), .ZN(n14213) );
  OAI211_X1 U17778 ( .C1(n10648), .C2(n14535), .A(n14214), .B(n14213), .ZN(
        n14534) );
  AOI22_X1 U17779 ( .A1(n20567), .A2(n17151), .B1(n17490), .B2(n14534), .ZN(
        n14228) );
  INV_X1 U17780 ( .A(n14215), .ZN(n14223) );
  INV_X1 U17781 ( .A(n14216), .ZN(n14217) );
  AND2_X1 U17782 ( .A1(n14218), .A2(n14217), .ZN(n14222) );
  NAND2_X1 U17783 ( .A1(n14577), .A2(n20613), .ZN(n14219) );
  OR2_X1 U17784 ( .A1(n14220), .A2(n14219), .ZN(n14221) );
  INV_X1 U17785 ( .A(n14595), .ZN(n17500) );
  AND2_X1 U17786 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(n17500), .ZN(n14224) );
  AOI21_X1 U17787 ( .B1(n13189), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n14224), 
        .ZN(n14225) );
  OAI21_X1 U17788 ( .B1(n14582), .B2(n14226), .A(n14225), .ZN(n17497) );
  NAND2_X1 U17789 ( .A1(n17156), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14227) );
  OAI21_X1 U17790 ( .B1(n14228), .B2(n17156), .A(n14227), .ZN(P2_U3596) );
  NAND2_X1 U17791 ( .A1(n20804), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20820) );
  OAI21_X1 U17792 ( .B1(n15530), .B2(n14233), .A(n20820), .ZN(n14232) );
  OAI21_X1 U17793 ( .B1(n14230), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n14229), .ZN(n20824) );
  NOR2_X1 U17794 ( .A1(n20824), .A2(n20633), .ZN(n14231) );
  AOI211_X1 U17795 ( .C1(n15533), .C2(n14233), .A(n14232), .B(n14231), .ZN(
        n14234) );
  OAI21_X1 U17796 ( .B1(n20837), .B2(n15292), .A(n14234), .ZN(P1_U2998) );
  INV_X1 U17797 ( .A(n14237), .ZN(n14235) );
  OAI21_X1 U17798 ( .B1(n14235), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n16435), .ZN(n14243) );
  INV_X1 U17799 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14236) );
  AND2_X1 U17800 ( .A1(n14189), .A2(n14238), .ZN(n14240) );
  OR2_X1 U17801 ( .A1(n14240), .A2(n14239), .ZN(n17117) );
  MUX2_X1 U17802 ( .A(n17117), .B(n14241), .S(n16438), .Z(n14242) );
  OAI21_X1 U17803 ( .B1(n14243), .B2(n14414), .A(n14242), .ZN(P2_U2882) );
  NAND2_X1 U17804 ( .A1(n19756), .A2(n19140), .ZN(n18046) );
  INV_X1 U17805 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18001) );
  OAI21_X1 U17806 ( .B1(n18001), .B2(n17959), .A(n18015), .ZN(n14246) );
  OAI21_X1 U17807 ( .B1(n18000), .B2(n18001), .A(n18025), .ZN(n17965) );
  INV_X1 U17808 ( .A(n17965), .ZN(n14245) );
  OAI22_X1 U17809 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18004), .B1(n18388), 
        .B2(n18039), .ZN(n14244) );
  AOI221_X1 U17810 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n14246), .C1(
        n18020), .C2(n14245), .A(n14244), .ZN(n14248) );
  NOR2_X1 U17811 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18016) );
  AOI21_X1 U17812 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n18016), .ZN(n18386) );
  AOI22_X1 U17813 ( .A1(n18011), .A2(n18386), .B1(n17983), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n14247) );
  OAI211_X1 U17814 ( .C1(n14249), .C2(n18046), .A(n14248), .B(n14247), .ZN(
        P3_U2670) );
  INV_X1 U17815 ( .A(n14250), .ZN(n14251) );
  AOI21_X1 U17816 ( .B1(n14252), .B2(n10348), .A(n14251), .ZN(n17020) );
  INV_X1 U17817 ( .A(n17020), .ZN(n16199) );
  AOI22_X1 U17818 ( .A1(n19793), .A2(n16449), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19796), .ZN(n14253) );
  OAI21_X1 U17819 ( .B1(n16199), .B2(n16565), .A(n14253), .ZN(P2_U2907) );
  OAI21_X1 U17820 ( .B1(n14256), .B2(n14255), .A(n14254), .ZN(n20810) );
  INV_X1 U17821 ( .A(n14257), .ZN(n14258) );
  AOI21_X1 U17822 ( .B1(n14259), .B2(n14131), .A(n14258), .ZN(n20703) );
  NOR2_X1 U17823 ( .A1(n20783), .A2(n20696), .ZN(n14262) );
  INV_X1 U17824 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20695) );
  INV_X1 U17825 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n14260) );
  OAI22_X1 U17826 ( .A1(n15530), .A2(n20695), .B1(n20771), .B2(n14260), .ZN(
        n14261) );
  AOI211_X1 U17827 ( .C1(n20703), .C2(n20778), .A(n14262), .B(n14261), .ZN(
        n14263) );
  OAI21_X1 U17828 ( .B1(n20633), .B2(n20810), .A(n14263), .ZN(P1_U2997) );
  INV_X1 U17829 ( .A(n14185), .ZN(n14265) );
  NOR2_X1 U17830 ( .A1(n14265), .A2(n14264), .ZN(n14397) );
  NAND2_X1 U17831 ( .A1(n14397), .A2(n14266), .ZN(n14407) );
  OAI211_X1 U17832 ( .C1(n14397), .C2(n14266), .A(n14407), .B(n16435), .ZN(
        n14271) );
  OAI21_X1 U17833 ( .B1(n14267), .B2(n14269), .A(n14268), .ZN(n17058) );
  INV_X1 U17834 ( .A(n17058), .ZN(n16779) );
  NAND2_X1 U17835 ( .A1(n16779), .A2(n16430), .ZN(n14270) );
  OAI211_X1 U17836 ( .C1(n16430), .C2(n14272), .A(n14271), .B(n14270), .ZN(
        P2_U2878) );
  INV_X1 U17837 ( .A(n20703), .ZN(n14294) );
  NAND2_X1 U17838 ( .A1(n20836), .A2(DATAI_2_), .ZN(n14274) );
  NAND2_X1 U17839 ( .A1(n20838), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14273) );
  AND2_X1 U17840 ( .A1(n14274), .A2(n14273), .ZN(n20861) );
  OAI222_X1 U17841 ( .A1(n15415), .A2(n14294), .B1(n15413), .B2(n12207), .C1(
        n15412), .C2(n20861), .ZN(P1_U2902) );
  INV_X1 U17842 ( .A(n19589), .ZN(n17655) );
  NOR2_X1 U17843 ( .A1(n14275), .A2(n17655), .ZN(n19593) );
  INV_X1 U17844 ( .A(n14728), .ZN(n18897) );
  NAND2_X1 U17845 ( .A1(n14278), .A2(n14277), .ZN(n19118) );
  NOR2_X1 U17846 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19737), .ZN(n18801) );
  NAND2_X1 U17847 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19127) );
  NAND2_X1 U17848 ( .A1(n19723), .A2(n19127), .ZN(n19742) );
  INV_X1 U17849 ( .A(n19742), .ZN(n14279) );
  NAND2_X1 U17850 ( .A1(n14279), .A2(n19740), .ZN(n14280) );
  NAND3_X1 U17851 ( .A1(n18536), .A2(n18737), .A3(n18906), .ZN(n14282) );
  INV_X1 U17852 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n14281) );
  NOR2_X1 U17853 ( .A1(n19120), .A2(n14281), .ZN(n19117) );
  AOI21_X1 U17854 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n14282), .A(
        n19117), .ZN(n14284) );
  NOR2_X4 U17855 ( .A1(n9644), .A2(n19736), .ZN(n18904) );
  NAND2_X1 U17856 ( .A1(n18904), .A2(n19118), .ZN(n14283) );
  OAI211_X1 U17857 ( .C1(n18897), .C2(n19118), .A(n14284), .B(n14283), .ZN(
        P3_U2830) );
  XNOR2_X1 U17858 ( .A(n14414), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14290) );
  OR2_X1 U17859 ( .A1(n14239), .A2(n14286), .ZN(n14287) );
  AND2_X1 U17860 ( .A1(n14285), .A2(n14287), .ZN(n17093) );
  INV_X1 U17861 ( .A(n17093), .ZN(n14288) );
  MUX2_X1 U17862 ( .A(n14288), .B(n16262), .S(n16438), .Z(n14289) );
  OAI21_X1 U17863 ( .B1(n14290), .B2(n16433), .A(n14289), .ZN(P2_U2881) );
  OR2_X1 U17864 ( .A1(n14292), .A2(n14291), .ZN(n14293) );
  NAND2_X1 U17865 ( .A1(n14430), .A2(n14293), .ZN(n20807) );
  INV_X1 U17866 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14295) );
  OAI222_X1 U17867 ( .A1(n20807), .A2(n15328), .B1(n14295), .B2(n20712), .C1(
        n14294), .C2(n15330), .ZN(P1_U2870) );
  NOR2_X1 U17868 ( .A1(n14298), .A2(n14297), .ZN(n14299) );
  OR2_X1 U17869 ( .A1(n14296), .A2(n14299), .ZN(n15281) );
  XNOR2_X1 U17870 ( .A(n14430), .B(n14426), .ZN(n20798) );
  AOI22_X1 U17871 ( .A1(n20707), .A2(n20798), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n15320), .ZN(n14300) );
  OAI21_X1 U17872 ( .B1(n15281), .B2(n15330), .A(n14300), .ZN(P1_U2869) );
  INV_X1 U17873 ( .A(DATAI_3_), .ZN(n14302) );
  NAND2_X1 U17874 ( .A1(n20838), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14301) );
  OAI21_X1 U17875 ( .B1(n20838), .B2(n14302), .A(n14301), .ZN(n20866) );
  INV_X1 U17876 ( .A(n20866), .ZN(n14303) );
  OAI222_X1 U17877 ( .A1(n15281), .A2(n15415), .B1(n15413), .B2(n12259), .C1(
        n15412), .C2(n14303), .ZN(P1_U2901) );
  INV_X1 U17878 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n21572) );
  OAI21_X1 U17879 ( .B1(n14448), .B2(n20854), .A(n14305), .ZN(n14307) );
  INV_X1 U17880 ( .A(n15925), .ZN(n14306) );
  OR2_X1 U17881 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17555), .ZN(n20735) );
  INV_X2 U17882 ( .A(n20735), .ZN(n21524) );
  NOR2_X4 U17883 ( .A1(n20721), .A2(n21524), .ZN(n20736) );
  AOI22_X1 U17884 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14308) );
  OAI21_X1 U17885 ( .B1(n21572), .B2(n20713), .A(n14308), .ZN(P1_U2909) );
  INV_X1 U17886 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14310) );
  AOI22_X1 U17887 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14309) );
  OAI21_X1 U17888 ( .B1(n14310), .B2(n20713), .A(n14309), .ZN(P1_U2920) );
  INV_X1 U17889 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14312) );
  AOI22_X1 U17890 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14311) );
  OAI21_X1 U17891 ( .B1(n14312), .B2(n20713), .A(n14311), .ZN(P1_U2908) );
  AOI22_X1 U17892 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14313) );
  OAI21_X1 U17893 ( .B1(n12563), .B2(n20713), .A(n14313), .ZN(P1_U2917) );
  AOI22_X1 U17894 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14314) );
  OAI21_X1 U17895 ( .B1(n15381), .B2(n20713), .A(n14314), .ZN(P1_U2918) );
  AOI22_X1 U17896 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14315) );
  OAI21_X1 U17897 ( .B1(n12729), .B2(n20713), .A(n14315), .ZN(P1_U2907) );
  AOI22_X1 U17898 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14316) );
  OAI21_X1 U17899 ( .B1(n15333), .B2(n20713), .A(n14316), .ZN(P1_U2906) );
  INV_X1 U17900 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15349) );
  AOI22_X1 U17901 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14317) );
  OAI21_X1 U17902 ( .B1(n15349), .B2(n20713), .A(n14317), .ZN(P1_U2911) );
  AOI22_X1 U17903 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14318) );
  OAI21_X1 U17904 ( .B1(n15361), .B2(n20713), .A(n14318), .ZN(P1_U2913) );
  INV_X1 U17905 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U17906 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14319) );
  OAI21_X1 U17907 ( .B1(n14320), .B2(n20713), .A(n14319), .ZN(P1_U2916) );
  INV_X1 U17908 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14322) );
  AOI22_X1 U17909 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14321) );
  OAI21_X1 U17910 ( .B1(n14322), .B2(n20713), .A(n14321), .ZN(P1_U2910) );
  AOI22_X1 U17911 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14323) );
  OAI21_X1 U17912 ( .B1(n15369), .B2(n20713), .A(n14323), .ZN(P1_U2915) );
  AOI21_X1 U17913 ( .B1(n14326), .B2(n10395), .A(n14325), .ZN(n17027) );
  INV_X1 U17914 ( .A(n17027), .ZN(n16751) );
  INV_X1 U17915 ( .A(n14410), .ZN(n14327) );
  NOR2_X1 U17916 ( .A1(n14407), .A2(n14327), .ZN(n14408) );
  OAI211_X1 U17917 ( .C1(n14408), .C2(n14329), .A(n16435), .B(n14328), .ZN(
        n14331) );
  NAND2_X1 U17918 ( .A1(n16438), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14330) );
  OAI211_X1 U17919 ( .C1(n16751), .C2(n16438), .A(n14331), .B(n14330), .ZN(
        P2_U2876) );
  NOR2_X1 U17920 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15884), .ZN(n14370) );
  INV_X1 U17921 ( .A(n14332), .ZN(n20844) );
  NAND4_X1 U17922 ( .A1(n14336), .A2(n14335), .A3(n14334), .A4(n14333), .ZN(
        n14337) );
  OR2_X1 U17923 ( .A1(n14338), .A2(n14337), .ZN(n15882) );
  AND2_X1 U17924 ( .A1(n10077), .A2(n14925), .ZN(n15881) );
  NOR2_X1 U17925 ( .A1(n14339), .A2(n10077), .ZN(n14340) );
  MUX2_X1 U17926 ( .A(n15881), .B(n14340), .S(n14342), .Z(n14348) );
  XNOR2_X1 U17927 ( .A(n14341), .B(n14342), .ZN(n15891) );
  NAND2_X1 U17928 ( .A1(n9580), .A2(n15891), .ZN(n14346) );
  NAND2_X1 U17929 ( .A1(n14344), .A2(n14343), .ZN(n14356) );
  INV_X1 U17930 ( .A(n14356), .ZN(n14345) );
  OAI22_X1 U17931 ( .A1(n15882), .A2(n14346), .B1(n14345), .B2(n15891), .ZN(
        n14347) );
  AOI211_X1 U17932 ( .C1(n20844), .C2(n15882), .A(n14348), .B(n14347), .ZN(
        n15894) );
  INV_X1 U17933 ( .A(n15894), .ZN(n14349) );
  MUX2_X1 U17934 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14349), .S(
        n14367), .Z(n15912) );
  AOI22_X1 U17935 ( .A1(n14370), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15912), .B2(n15884), .ZN(n14364) );
  AOI21_X1 U17936 ( .B1(n14341), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14351) );
  NOR2_X1 U17937 ( .A1(n12746), .A2(n14351), .ZN(n15896) );
  NAND2_X1 U17938 ( .A1(n9580), .A2(n15896), .ZN(n14360) );
  INV_X1 U17939 ( .A(n14355), .ZN(n14353) );
  NAND2_X1 U17940 ( .A1(n14353), .A2(n14352), .ZN(n14354) );
  AOI22_X1 U17941 ( .A1(n15881), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n14925), .B2(n14354), .ZN(n14359) );
  MUX2_X1 U17942 ( .A(n14355), .B(n11964), .S(n14341), .Z(n14357) );
  OAI211_X1 U17943 ( .C1(n15882), .C2(n14360), .A(n14359), .B(n14358), .ZN(
        n14361) );
  AOI21_X1 U17944 ( .B1(n21119), .B2(n15882), .A(n14361), .ZN(n15899) );
  MUX2_X1 U17945 ( .A(n11964), .B(n15899), .S(n14367), .Z(n15914) );
  INV_X1 U17946 ( .A(n15914), .ZN(n14362) );
  AOI22_X1 U17947 ( .A1(n14370), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n15884), .B2(n14362), .ZN(n14363) );
  NOR2_X1 U17948 ( .A1(n14364), .A2(n14363), .ZN(n15920) );
  INV_X1 U17949 ( .A(n14365), .ZN(n15879) );
  NAND2_X1 U17950 ( .A1(n15920), .A2(n15879), .ZN(n14379) );
  NAND2_X1 U17951 ( .A1(n15262), .A2(n14366), .ZN(n14368) );
  NAND2_X1 U17952 ( .A1(n14368), .A2(n14367), .ZN(n14373) );
  AOI21_X1 U17953 ( .B1(n15906), .B2(n14369), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n14372) );
  AND2_X1 U17954 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n14370), .ZN(
        n14371) );
  AOI21_X1 U17955 ( .B1(n14373), .B2(n14372), .A(n14371), .ZN(n15919) );
  AND3_X1 U17956 ( .A1(n14379), .A2(n15919), .A3(n20634), .ZN(n14377) );
  AND3_X1 U17957 ( .A1(n14379), .A2(n15919), .A3(n14378), .ZN(n15935) );
  INV_X1 U17958 ( .A(n12223), .ZN(n15297) );
  AND2_X1 U17959 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21248), .ZN(n15875) );
  OAI22_X1 U17960 ( .A1(n12880), .A2(n21382), .B1(n15297), .B2(n15875), .ZN(
        n14380) );
  OAI21_X1 U17961 ( .B1(n15935), .B2(n14380), .A(n20834), .ZN(n14381) );
  OAI21_X1 U17962 ( .B1(n20834), .B2(n21294), .A(n14381), .ZN(P1_U3478) );
  AOI21_X1 U17963 ( .B1(n14383), .B2(n14250), .A(n14382), .ZN(n17007) );
  INV_X1 U17964 ( .A(n17007), .ZN(n16185) );
  INV_X1 U17965 ( .A(n16443), .ZN(n14384) );
  INV_X1 U17966 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19808) );
  OAI222_X1 U17967 ( .A1(n16185), .A2(n16565), .B1(n14384), .B2(n19803), .C1(
        n19808), .C2(n19795), .ZN(P2_U2906) );
  XNOR2_X1 U17968 ( .A(n17254), .B(n10316), .ZN(n17259) );
  AOI21_X1 U17969 ( .B1(n14387), .B2(n21579), .A(n14386), .ZN(n17256) );
  NOR4_X1 U17970 ( .A1(n19113), .A2(n14390), .A3(n18980), .A4(n14388), .ZN(
        n14393) );
  AOI211_X1 U17971 ( .C1(n18995), .C2(n14390), .A(n19113), .B(n14389), .ZN(
        n19106) );
  OAI21_X1 U17972 ( .B1(n19106), .B2(n17276), .A(n19114), .ZN(n14392) );
  NAND2_X1 U17973 ( .A1(n19089), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17251) );
  INV_X1 U17974 ( .A(n17251), .ZN(n14391) );
  AOI221_X1 U17975 ( .B1(n14393), .B2(n21579), .C1(n14392), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n14391), .ZN(n14394) );
  OAI21_X1 U17976 ( .B1(n17254), .B2(n19037), .A(n14394), .ZN(n14395) );
  AOI21_X1 U17977 ( .B1(n19119), .B2(n17256), .A(n14395), .ZN(n14396) );
  OAI21_X1 U17978 ( .B1(n17259), .B2(n19058), .A(n14396), .ZN(P3_U2854) );
  INV_X1 U17979 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n16235) );
  AND3_X1 U17980 ( .A1(n14414), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14416) );
  INV_X1 U17981 ( .A(n14397), .ZN(n14398) );
  OAI211_X1 U17982 ( .C1(n14416), .C2(n14399), .A(n16435), .B(n14398), .ZN(
        n14405) );
  AND2_X1 U17983 ( .A1(n14400), .A2(n14401), .ZN(n14402) );
  OR2_X1 U17984 ( .A1(n14402), .A2(n14267), .ZN(n17069) );
  INV_X1 U17985 ( .A(n17069), .ZN(n14403) );
  NAND2_X1 U17986 ( .A1(n14403), .A2(n16430), .ZN(n14404) );
  OAI211_X1 U17987 ( .C1(n16430), .C2(n16235), .A(n14405), .B(n14404), .ZN(
        P2_U2879) );
  AOI21_X1 U17988 ( .B1(n14406), .B2(n14268), .A(n14324), .ZN(n16760) );
  INV_X1 U17989 ( .A(n16760), .ZN(n17046) );
  INV_X1 U17990 ( .A(n14407), .ZN(n14411) );
  INV_X1 U17991 ( .A(n14408), .ZN(n14409) );
  OAI211_X1 U17992 ( .C1(n14411), .C2(n14410), .A(n14409), .B(n16435), .ZN(
        n14413) );
  NAND2_X1 U17993 ( .A1(n16438), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14412) );
  OAI211_X1 U17994 ( .C1(n17046), .C2(n16438), .A(n14413), .B(n14412), .ZN(
        P2_U2877) );
  AOI21_X1 U17995 ( .B1(n14414), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14415) );
  OR3_X1 U17996 ( .A1(n14416), .A2(n14415), .A3(n16433), .ZN(n14421) );
  NAND2_X1 U17997 ( .A1(n14285), .A2(n14417), .ZN(n14418) );
  NAND2_X1 U17998 ( .A1(n14400), .A2(n14418), .ZN(n16815) );
  MUX2_X1 U17999 ( .A(n16815), .B(n14419), .S(n16438), .Z(n14420) );
  NAND2_X1 U18000 ( .A1(n14421), .A2(n14420), .ZN(P2_U2880) );
  NAND2_X1 U18001 ( .A1(n20836), .A2(DATAI_4_), .ZN(n14423) );
  NAND2_X1 U18002 ( .A1(n20838), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14422) );
  AND2_X1 U18003 ( .A1(n14423), .A2(n14422), .ZN(n20871) );
  INV_X1 U18004 ( .A(n14424), .ZN(n14425) );
  XNOR2_X1 U18005 ( .A(n14296), .B(n14425), .ZN(n20777) );
  INV_X1 U18006 ( .A(n20777), .ZN(n15269) );
  INV_X1 U18007 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20733) );
  OAI222_X1 U18008 ( .A1(n15412), .A2(n20871), .B1(n15415), .B2(n15269), .C1(
        n20733), .C2(n15413), .ZN(P1_U2900) );
  INV_X1 U18009 ( .A(n14426), .ZN(n14429) );
  INV_X1 U18010 ( .A(n14427), .ZN(n14428) );
  OAI21_X1 U18011 ( .B1(n14430), .B2(n14429), .A(n14428), .ZN(n14431) );
  NAND2_X1 U18012 ( .A1(n14431), .A2(n14531), .ZN(n20787) );
  OAI222_X1 U18013 ( .A1(n20787), .A2(n15328), .B1(n14432), .B2(n20712), .C1(
        n15330), .C2(n15269), .ZN(P1_U2868) );
  NOR2_X1 U18014 ( .A1(n14325), .A2(n14433), .ZN(n14434) );
  OR2_X1 U18015 ( .A1(n14440), .A2(n14434), .ZN(n17018) );
  NAND2_X1 U18016 ( .A1(n16735), .A2(n16430), .ZN(n14438) );
  OAI211_X1 U18017 ( .C1(n10412), .C2(n14436), .A(n16435), .B(n14435), .ZN(
        n14437) );
  OAI211_X1 U18018 ( .C1(n16430), .C2(n16191), .A(n14438), .B(n14437), .ZN(
        P2_U2875) );
  NAND2_X1 U18019 ( .A1(n14440), .A2(n14439), .ZN(n14654) );
  OAI21_X1 U18020 ( .B1(n14440), .B2(n14439), .A(n14654), .ZN(n17004) );
  INV_X1 U18021 ( .A(n14435), .ZN(n14443) );
  OAI211_X1 U18022 ( .C1(n14443), .C2(n14442), .A(n16435), .B(n14441), .ZN(
        n14445) );
  NAND2_X1 U18023 ( .A1(n16438), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n14444) );
  OAI211_X1 U18024 ( .C1(n17004), .C2(n16438), .A(n14445), .B(n14444), .ZN(
        P2_U2874) );
  NOR2_X1 U18025 ( .A1(n14446), .A2(n21523), .ZN(n14447) );
  NAND2_X1 U18026 ( .A1(n20836), .A2(DATAI_9_), .ZN(n14450) );
  NAND2_X1 U18027 ( .A1(n20838), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14449) );
  AND2_X1 U18028 ( .A1(n14450), .A2(n14449), .ZN(n15408) );
  INV_X1 U18029 ( .A(n15408), .ZN(n14451) );
  NAND2_X1 U18030 ( .A1(n20756), .A2(n14451), .ZN(n20760) );
  AOI22_X1 U18031 ( .A1(n14493), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14452) );
  NAND2_X1 U18032 ( .A1(n20760), .A2(n14452), .ZN(P1_U2946) );
  NAND2_X1 U18033 ( .A1(n20836), .A2(DATAI_7_), .ZN(n14454) );
  NAND2_X1 U18034 ( .A1(n20838), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14453) );
  AND2_X1 U18035 ( .A1(n14454), .A2(n14453), .ZN(n20888) );
  INV_X1 U18036 ( .A(n20888), .ZN(n14455) );
  NAND2_X1 U18037 ( .A1(n20756), .A2(n14455), .ZN(n14478) );
  AOI22_X1 U18038 ( .A1(n14493), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n14456) );
  NAND2_X1 U18039 ( .A1(n14478), .A2(n14456), .ZN(P1_U2959) );
  NAND2_X1 U18040 ( .A1(n20836), .A2(DATAI_5_), .ZN(n14458) );
  NAND2_X1 U18041 ( .A1(n20838), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14457) );
  AND2_X1 U18042 ( .A1(n14458), .A2(n14457), .ZN(n20875) );
  INV_X1 U18043 ( .A(n20875), .ZN(n14459) );
  NAND2_X1 U18044 ( .A1(n20756), .A2(n14459), .ZN(n14490) );
  AOI22_X1 U18045 ( .A1(n14493), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n14460) );
  NAND2_X1 U18046 ( .A1(n14490), .A2(n14460), .ZN(P1_U2957) );
  INV_X1 U18047 ( .A(n20861), .ZN(n14461) );
  NAND2_X1 U18048 ( .A1(n20756), .A2(n14461), .ZN(n14482) );
  AOI22_X1 U18049 ( .A1(n14493), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U18050 ( .A1(n14482), .A2(n14462), .ZN(P1_U2939) );
  NAND2_X1 U18051 ( .A1(n20836), .A2(DATAI_6_), .ZN(n14464) );
  NAND2_X1 U18052 ( .A1(n20838), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14463) );
  AND2_X1 U18053 ( .A1(n14464), .A2(n14463), .ZN(n20880) );
  INV_X1 U18054 ( .A(n20880), .ZN(n14465) );
  NAND2_X1 U18055 ( .A1(n20756), .A2(n14465), .ZN(n14480) );
  AOI22_X1 U18056 ( .A1(n14493), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n14466) );
  NAND2_X1 U18057 ( .A1(n14480), .A2(n14466), .ZN(P1_U2958) );
  INV_X1 U18058 ( .A(n20871), .ZN(n14467) );
  NAND2_X1 U18059 ( .A1(n20756), .A2(n14467), .ZN(n14492) );
  AOI22_X1 U18060 ( .A1(n14493), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n14468) );
  NAND2_X1 U18061 ( .A1(n14492), .A2(n14468), .ZN(P1_U2956) );
  NAND2_X1 U18062 ( .A1(n20756), .A2(n20866), .ZN(n14486) );
  AOI22_X1 U18063 ( .A1(n14493), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n14469) );
  NAND2_X1 U18064 ( .A1(n14486), .A2(n14469), .ZN(P1_U2955) );
  INV_X1 U18065 ( .A(n20847), .ZN(n14470) );
  NAND2_X1 U18066 ( .A1(n20756), .A2(n14470), .ZN(n14488) );
  AOI22_X1 U18067 ( .A1(n14493), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14471) );
  NAND2_X1 U18068 ( .A1(n14488), .A2(n14471), .ZN(P1_U2937) );
  NAND2_X1 U18069 ( .A1(n20756), .A2(n20856), .ZN(n14484) );
  AOI22_X1 U18070 ( .A1(n14493), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n14472) );
  NAND2_X1 U18071 ( .A1(n14484), .A2(n14472), .ZN(P1_U2953) );
  NAND2_X1 U18072 ( .A1(n20836), .A2(DATAI_11_), .ZN(n14474) );
  NAND2_X1 U18073 ( .A1(n20838), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14473) );
  AND2_X1 U18074 ( .A1(n14474), .A2(n14473), .ZN(n15405) );
  INV_X1 U18075 ( .A(n15405), .ZN(n14475) );
  NAND2_X1 U18076 ( .A1(n20756), .A2(n14475), .ZN(n14495) );
  AOI22_X1 U18077 ( .A1(n14493), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20768), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n14476) );
  NAND2_X1 U18078 ( .A1(n14495), .A2(n14476), .ZN(P1_U2963) );
  AOI22_X1 U18079 ( .A1(n14493), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14477) );
  NAND2_X1 U18080 ( .A1(n14478), .A2(n14477), .ZN(P1_U2944) );
  AOI22_X1 U18081 ( .A1(n14493), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14479) );
  NAND2_X1 U18082 ( .A1(n14480), .A2(n14479), .ZN(P1_U2943) );
  AOI22_X1 U18083 ( .A1(n14493), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n14481) );
  NAND2_X1 U18084 ( .A1(n14482), .A2(n14481), .ZN(P1_U2954) );
  AOI22_X1 U18085 ( .A1(n14493), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14483) );
  NAND2_X1 U18086 ( .A1(n14484), .A2(n14483), .ZN(P1_U2938) );
  AOI22_X1 U18087 ( .A1(n14493), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14485) );
  NAND2_X1 U18088 ( .A1(n14486), .A2(n14485), .ZN(P1_U2940) );
  AOI22_X1 U18089 ( .A1(n14493), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n14487) );
  NAND2_X1 U18090 ( .A1(n14488), .A2(n14487), .ZN(P1_U2952) );
  AOI22_X1 U18091 ( .A1(n14493), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14489) );
  NAND2_X1 U18092 ( .A1(n14490), .A2(n14489), .ZN(P1_U2942) );
  AOI22_X1 U18093 ( .A1(n14493), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14491) );
  NAND2_X1 U18094 ( .A1(n14492), .A2(n14491), .ZN(P1_U2941) );
  AOI22_X1 U18095 ( .A1(n14493), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14494) );
  NAND2_X1 U18096 ( .A1(n14495), .A2(n14494), .ZN(P1_U2948) );
  INV_X1 U18097 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14499) );
  INV_X1 U18098 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20719) );
  INV_X1 U18099 ( .A(n20756), .ZN(n14497) );
  MUX2_X1 U18100 ( .A(DATAI_15_), .B(BUF1_REG_15__SCAN_IN), .S(n20838), .Z(
        n15396) );
  INV_X1 U18101 ( .A(n15396), .ZN(n14496) );
  OAI222_X1 U18102 ( .A1(n14500), .A2(n14499), .B1(n14498), .B2(n20719), .C1(
        n14497), .C2(n14496), .ZN(P1_U2967) );
  INV_X1 U18103 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18608) );
  INV_X1 U18104 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18606) );
  NAND2_X1 U18105 ( .A1(n14501), .A2(n19743), .ZN(n14507) );
  NAND3_X1 U18106 ( .A1(n19157), .A2(n11836), .A3(n14502), .ZN(n14503) );
  NAND2_X1 U18107 ( .A1(n14711), .A2(n14505), .ZN(n14506) );
  NOR3_X1 U18108 ( .A1(n18608), .A2(n18606), .A3(n18438), .ZN(n14515) );
  NAND2_X1 U18109 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n14518), .ZN(n18535) );
  INV_X1 U18110 ( .A(n18535), .ZN(n18523) );
  NOR2_X1 U18111 ( .A1(n11836), .A2(n14663), .ZN(n18533) );
  AOI21_X1 U18112 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18522), .A(n14518), .ZN(
        n14511) );
  AOI22_X1 U18113 ( .A1(n14509), .A2(n18530), .B1(n18531), .B2(
        BUF2_REG_3__SCAN_IN), .ZN(n14510) );
  OAI21_X1 U18114 ( .B1(n18523), .B2(n14511), .A(n14510), .ZN(P3_U2732) );
  AOI22_X1 U18115 ( .A1(n14512), .A2(n18530), .B1(n18531), .B2(
        BUF2_REG_0__SCAN_IN), .ZN(n14514) );
  NAND2_X1 U18116 ( .A1(n14663), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n14513) );
  OAI211_X1 U18117 ( .C1(n18438), .C2(P3_EAX_REG_0__SCAN_IN), .A(n14514), .B(
        n14513), .ZN(P3_U2735) );
  AOI21_X1 U18118 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18522), .A(n14515), .ZN(
        n14519) );
  AOI22_X1 U18119 ( .A1(n14516), .A2(n18530), .B1(n18531), .B2(
        BUF2_REG_2__SCAN_IN), .ZN(n14517) );
  OAI21_X1 U18120 ( .B1(n14519), .B2(n14518), .A(n14517), .ZN(P3_U2733) );
  XNOR2_X1 U18121 ( .A(n14520), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14524) );
  AND2_X1 U18122 ( .A1(n14522), .A2(n14521), .ZN(n14523) );
  NOR2_X1 U18123 ( .A1(n14524), .A2(n14523), .ZN(n20773) );
  AOI21_X1 U18124 ( .B1(n14524), .B2(n14523), .A(n20773), .ZN(n20800) );
  NAND2_X1 U18125 ( .A1(n20800), .A2(n20779), .ZN(n14527) );
  AND2_X1 U18126 ( .A1(n20804), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20797) );
  NOR2_X1 U18127 ( .A1(n20783), .A2(n15274), .ZN(n14525) );
  AOI211_X1 U18128 ( .C1(n20772), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20797), .B(n14525), .ZN(n14526) );
  OAI211_X1 U18129 ( .C1(n20837), .C2(n15281), .A(n14527), .B(n14526), .ZN(
        P1_U2996) );
  AOI21_X1 U18130 ( .B1(n14530), .B2(n14529), .A(n14528), .ZN(n20686) );
  INV_X1 U18131 ( .A(n20686), .ZN(n14533) );
  INV_X1 U18132 ( .A(n14531), .ZN(n17538) );
  XNOR2_X1 U18133 ( .A(n17538), .B(n17537), .ZN(n20677) );
  OAI222_X1 U18134 ( .A1(n15330), .A2(n14533), .B1(n14532), .B2(n20712), .C1(
        n15328), .C2(n20677), .ZN(P1_U2867) );
  OAI222_X1 U18135 ( .A1(n15415), .A2(n14533), .B1(n15413), .B2(n12303), .C1(
        n15412), .C2(n20875), .ZN(P1_U2899) );
  AOI22_X1 U18136 ( .A1(n14582), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n14534), .B2(n14565), .ZN(n14586) );
  INV_X1 U18137 ( .A(n14535), .ZN(n14555) );
  NAND2_X1 U18138 ( .A1(n14537), .A2(n14536), .ZN(n14538) );
  MUX2_X1 U18139 ( .A(n14539), .B(n14538), .S(n9562), .Z(n14545) );
  AND2_X1 U18140 ( .A1(n14541), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14542) );
  OAI21_X1 U18141 ( .B1(n14540), .B2(n14542), .A(n11235), .ZN(n14543) );
  NAND3_X1 U18142 ( .A1(n14545), .A2(n14544), .A3(n14543), .ZN(n14546) );
  AOI21_X1 U18143 ( .B1(n13361), .B2(n14555), .A(n14546), .ZN(n17149) );
  NOR2_X1 U18144 ( .A1(n14565), .A2(n17154), .ZN(n14547) );
  AOI21_X1 U18145 ( .B1(n17149), .B2(n14565), .A(n14547), .ZN(n14568) );
  INV_X1 U18146 ( .A(n14568), .ZN(n14585) );
  NAND2_X1 U18147 ( .A1(n16366), .A2(n14555), .ZN(n14554) );
  INV_X1 U18148 ( .A(n11235), .ZN(n14552) );
  INV_X1 U18149 ( .A(n14548), .ZN(n14549) );
  OR2_X1 U18150 ( .A1(n11496), .A2(n14549), .ZN(n14557) );
  INV_X1 U18151 ( .A(n14557), .ZN(n14551) );
  MUX2_X1 U18152 ( .A(n14552), .B(n14551), .S(n14550), .Z(n14553) );
  NAND2_X1 U18153 ( .A1(n14554), .A2(n14553), .ZN(n14693) );
  NAND2_X1 U18154 ( .A1(n9574), .A2(n14555), .ZN(n14561) );
  AOI22_X1 U18155 ( .A1(n11235), .A2(n14559), .B1(n14558), .B2(n14557), .ZN(
        n14560) );
  NAND2_X1 U18156 ( .A1(n14561), .A2(n14560), .ZN(n17146) );
  INV_X1 U18157 ( .A(n17146), .ZN(n14564) );
  INV_X1 U18158 ( .A(n20137), .ZN(n14562) );
  AOI21_X1 U18159 ( .B1(n14693), .B2(n20591), .A(n14562), .ZN(n14563) );
  AOI22_X1 U18160 ( .A1(n17149), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n14564), .B2(n14563), .ZN(n14566) );
  OAI211_X1 U18161 ( .C1(n20235), .C2(n14693), .A(n14566), .B(n14565), .ZN(
        n14567) );
  AOI222_X1 U18162 ( .A1(n14586), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .B1(n14586), .B2(n14567), .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .C2(n14567), .ZN(n14569) );
  NAND2_X1 U18163 ( .A1(n20574), .A2(n20582), .ZN(n19970) );
  INV_X1 U18164 ( .A(n19970), .ZN(n19941) );
  OAI221_X1 U18165 ( .B1(n14569), .B2(n19941), .C1(n14569), .C2(n14568), .A(
        n10865), .ZN(n14584) );
  MUX2_X1 U18166 ( .A(n14572), .B(n14571), .S(n14570), .Z(n14573) );
  OAI21_X1 U18167 ( .B1(n9805), .B2(n14574), .A(n14573), .ZN(n20599) );
  OAI21_X1 U18168 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n14575), .ZN(n14579) );
  INV_X1 U18169 ( .A(n17492), .ZN(n14576) );
  NAND3_X1 U18170 ( .A1(n14577), .A2(n9593), .A3(n14576), .ZN(n14578) );
  OAI211_X1 U18171 ( .C1(n14580), .C2(n10858), .A(n14579), .B(n14578), .ZN(
        n14581) );
  AOI211_X1 U18172 ( .C1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n14582), .A(
        n20599), .B(n14581), .ZN(n14583) );
  OAI211_X1 U18173 ( .C1(n14586), .C2(n14585), .A(n14584), .B(n14583), .ZN(
        n14597) );
  OAI21_X1 U18174 ( .B1(n14597), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14588) );
  AOI211_X1 U18175 ( .C1(n10050), .C2(n14587), .A(n20608), .B(n20326), .ZN(
        n14590) );
  NAND2_X1 U18176 ( .A1(n14588), .A2(n14590), .ZN(n14602) );
  NAND2_X1 U18177 ( .A1(n14602), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14606) );
  INV_X1 U18178 ( .A(n14606), .ZN(n14589) );
  OAI21_X1 U18179 ( .B1(n14589), .B2(n20607), .A(n14595), .ZN(P2_U3593) );
  INV_X1 U18180 ( .A(n20613), .ZN(n20612) );
  AOI22_X1 U18181 ( .A1(n17151), .A2(n14591), .B1(n14590), .B2(n20612), .ZN(
        n14592) );
  OAI21_X1 U18182 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n14592), .A(n14606), 
        .ZN(n14599) );
  INV_X1 U18183 ( .A(n17499), .ZN(n20601) );
  NAND3_X1 U18184 ( .A1(n20326), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20612), 
        .ZN(n14594) );
  OAI211_X1 U18185 ( .C1(n20601), .C2(n14595), .A(n14594), .B(n14593), .ZN(
        n14596) );
  AOI21_X1 U18186 ( .B1(n14597), .B2(n14601), .A(n14596), .ZN(n14598) );
  NAND2_X1 U18187 ( .A1(n14599), .A2(n14598), .ZN(P2_U3176) );
  NAND2_X1 U18188 ( .A1(n20613), .A2(n17490), .ZN(n14605) );
  OAI21_X1 U18189 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n13189), .A(n14602), 
        .ZN(n14600) );
  NAND3_X1 U18190 ( .A1(n14600), .A2(n20612), .A3(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n14604) );
  AOI21_X1 U18191 ( .B1(n14602), .B2(n14601), .A(n16292), .ZN(n14603) );
  OAI211_X1 U18192 ( .C1(n14606), .C2(n14605), .A(n14604), .B(n14603), .ZN(
        P2_U3177) );
  OR2_X1 U18193 ( .A1(n14654), .A2(n14608), .ZN(n14656) );
  INV_X1 U18194 ( .A(n14656), .ZN(n14607) );
  AOI21_X1 U18195 ( .B1(n14608), .B2(n14654), .A(n14607), .ZN(n16983) );
  NAND2_X1 U18196 ( .A1(n16983), .A2(n16430), .ZN(n14613) );
  INV_X1 U18197 ( .A(n14441), .ZN(n14611) );
  INV_X1 U18198 ( .A(n14660), .ZN(n14609) );
  OAI211_X1 U18199 ( .C1(n14611), .C2(n14610), .A(n14609), .B(n16435), .ZN(
        n14612) );
  OAI211_X1 U18200 ( .C1(n16430), .C2(n10995), .A(n14613), .B(n14612), .ZN(
        P2_U2873) );
  XNOR2_X1 U18201 ( .A(n14615), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14616) );
  XNOR2_X1 U18202 ( .A(n14614), .B(n14616), .ZN(n15620) );
  INV_X1 U18203 ( .A(n14618), .ZN(n15327) );
  INV_X1 U18204 ( .A(n14619), .ZN(n14620) );
  AOI21_X1 U18205 ( .B1(n14617), .B2(n15327), .A(n14620), .ZN(n14621) );
  OR2_X1 U18206 ( .A1(n15224), .A2(n14621), .ZN(n15323) );
  NAND2_X1 U18207 ( .A1(n14622), .A2(n20784), .ZN(n17552) );
  INV_X1 U18208 ( .A(n17552), .ZN(n14627) );
  INV_X1 U18209 ( .A(n15816), .ZN(n20814) );
  NAND2_X1 U18210 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14623) );
  AND2_X1 U18211 ( .A1(n15816), .A2(n14623), .ZN(n14624) );
  OR2_X1 U18212 ( .A1(n14624), .A2(n15817), .ZN(n15846) );
  INV_X1 U18213 ( .A(n15846), .ZN(n20792) );
  NAND2_X1 U18214 ( .A1(n20811), .A2(n14625), .ZN(n14626) );
  OAI211_X1 U18215 ( .C1(n20814), .C2(n20784), .A(n20792), .B(n14626), .ZN(
        n17548) );
  AOI211_X1 U18216 ( .C1(n14628), .C2(n14627), .A(n17514), .B(n17548), .ZN(
        n17544) );
  INV_X1 U18217 ( .A(n17544), .ZN(n17529) );
  NAND3_X1 U18218 ( .A1(n17529), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n17528), .ZN(n14629) );
  NAND2_X1 U18219 ( .A1(n20804), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15615) );
  OAI211_X1 U18220 ( .C1(n20808), .C2(n15323), .A(n14629), .B(n15615), .ZN(
        n14630) );
  INV_X1 U18221 ( .A(n14630), .ZN(n14633) );
  NAND2_X1 U18222 ( .A1(n17535), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17534) );
  INV_X1 U18223 ( .A(n17534), .ZN(n14631) );
  OAI211_X1 U18224 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n14631), .B(n15841), .ZN(n14632) );
  OAI211_X1 U18225 ( .C1(n15620), .C2(n15862), .A(n14633), .B(n14632), .ZN(
        P1_U3023) );
  XNOR2_X1 U18226 ( .A(n16847), .B(n14634), .ZN(n16849) );
  XNOR2_X1 U18227 ( .A(n16849), .B(n16848), .ZN(n14652) );
  XOR2_X1 U18228 ( .A(n14635), .B(n14636), .Z(n14650) );
  NAND2_X1 U18229 ( .A1(n16837), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n14644) );
  OAI21_X1 U18230 ( .B1(n16839), .B2(n14637), .A(n14644), .ZN(n14638) );
  AOI21_X1 U18231 ( .B1(n16842), .B2(n16308), .A(n14638), .ZN(n14639) );
  OAI21_X1 U18232 ( .B1(n10648), .B2(n19838), .A(n14639), .ZN(n14640) );
  AOI21_X1 U18233 ( .B1(n14650), .B2(n13307), .A(n14640), .ZN(n14641) );
  OAI21_X1 U18234 ( .B1(n14652), .B2(n16863), .A(n14641), .ZN(P2_U3011) );
  XNOR2_X1 U18235 ( .A(n14642), .B(n14643), .ZN(n20565) );
  INV_X1 U18236 ( .A(n14644), .ZN(n14645) );
  MUX2_X1 U18237 ( .A(n14646), .B(n17095), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n14647) );
  OAI211_X1 U18238 ( .C1(n20565), .C2(n17134), .A(n14648), .B(n14647), .ZN(
        n14649) );
  AOI21_X1 U18239 ( .B1(n14650), .B2(n17136), .A(n14649), .ZN(n14651) );
  OAI21_X1 U18240 ( .B1(n14652), .B2(n17139), .A(n14651), .ZN(P2_U3043) );
  OR2_X1 U18241 ( .A1(n14654), .A2(n14653), .ZN(n14670) );
  INV_X1 U18242 ( .A(n14670), .ZN(n14655) );
  AOI21_X1 U18243 ( .B1(n14657), .B2(n14656), .A(n14655), .ZN(n16696) );
  INV_X1 U18244 ( .A(n16696), .ZN(n16977) );
  OAI211_X1 U18245 ( .C1(n14660), .C2(n14659), .A(n14658), .B(n16435), .ZN(
        n14662) );
  NAND2_X1 U18246 ( .A1(n16438), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14661) );
  OAI211_X1 U18247 ( .C1(n16977), .C2(n16438), .A(n14662), .B(n14661), .ZN(
        P2_U2872) );
  AOI21_X1 U18248 ( .B1(n11836), .B2(n18606), .A(n14663), .ZN(n14668) );
  NAND2_X1 U18249 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18512), .ZN(n14664) );
  OAI22_X1 U18250 ( .A1(n19143), .A2(n18528), .B1(P3_EAX_REG_1__SCAN_IN), .B2(
        n14664), .ZN(n14665) );
  AOI21_X1 U18251 ( .B1(n14666), .B2(n18530), .A(n14665), .ZN(n14667) );
  OAI21_X1 U18252 ( .B1(n14668), .B2(n18608), .A(n14667), .ZN(P3_U2734) );
  AND2_X1 U18253 ( .A1(n14670), .A2(n14669), .ZN(n14672) );
  INV_X1 U18254 ( .A(n14673), .ZN(n14674) );
  AOI21_X1 U18255 ( .B1(n14675), .B2(n14658), .A(n14674), .ZN(n16540) );
  NAND2_X1 U18256 ( .A1(n16540), .A2(n16435), .ZN(n14677) );
  NAND2_X1 U18257 ( .A1(n16438), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n14676) );
  OAI211_X1 U18258 ( .C1(n16963), .C2(n16438), .A(n14677), .B(n14676), .ZN(
        P2_U2871) );
  XOR2_X1 U18259 ( .A(n14679), .B(n14678), .Z(n20709) );
  INV_X1 U18260 ( .A(n20709), .ZN(n14680) );
  OAI222_X1 U18261 ( .A1(n15412), .A2(n20880), .B1(n15415), .B2(n14680), .C1(
        n21595), .C2(n15413), .ZN(P1_U2898) );
  AND2_X1 U18262 ( .A1(n14673), .A2(n14681), .ZN(n14683) );
  OR2_X1 U18263 ( .A1(n14683), .A2(n14682), .ZN(n16539) );
  NAND2_X1 U18264 ( .A1(n16676), .A2(n16430), .ZN(n14685) );
  NAND2_X1 U18265 ( .A1(n16438), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14684) );
  OAI211_X1 U18266 ( .C1(n16539), .C2(n16433), .A(n14685), .B(n14684), .ZN(
        P2_U2870) );
  OAI21_X1 U18267 ( .B1(n14682), .B2(n14687), .A(n14686), .ZN(n16532) );
  INV_X1 U18268 ( .A(n16089), .ZN(n14688) );
  AOI21_X1 U18269 ( .B1(n14689), .B2(n13149), .A(n14688), .ZN(n16956) );
  NAND2_X1 U18270 ( .A1(n16956), .A2(n16430), .ZN(n14691) );
  NAND2_X1 U18271 ( .A1(n16438), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14690) );
  OAI211_X1 U18272 ( .C1(n16532), .C2(n16433), .A(n14691), .B(n14690), .ZN(
        P2_U2869) );
  INV_X1 U18273 ( .A(n16331), .ZN(n16363) );
  MUX2_X1 U18274 ( .A(n16363), .B(n14692), .S(n13243), .Z(n17142) );
  AOI222_X1 U18275 ( .A1(n17142), .A2(P2_STATE2_REG_1__SCAN_IN), .B1(n14044), 
        .B2(n17151), .C1(n14693), .C2(n17490), .ZN(n14695) );
  NAND2_X1 U18276 ( .A1(n17156), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14694) );
  OAI21_X1 U18277 ( .B1(n14695), .B2(n17156), .A(n14694), .ZN(P2_U3601) );
  INV_X1 U18278 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14698) );
  AOI22_X1 U18279 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14697) );
  NAND2_X1 U18280 ( .A1(n18170), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14696) );
  OAI211_X1 U18281 ( .C1(n14698), .C2(n18218), .A(n14697), .B(n14696), .ZN(
        n14699) );
  INV_X1 U18282 ( .A(n14699), .ZN(n14702) );
  AOI22_X1 U18283 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14701) );
  AOI22_X1 U18284 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14700) );
  NAND3_X1 U18285 ( .A1(n14702), .A2(n14701), .A3(n14700), .ZN(n14709) );
  INV_X1 U18286 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18229) );
  AOI22_X1 U18287 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14703) );
  OAI21_X1 U18288 ( .B1(n18352), .B2(n18229), .A(n14703), .ZN(n14704) );
  AOI21_X1 U18289 ( .B1(n9560), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(n14704), .ZN(n14707) );
  AOI22_X1 U18290 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14706) );
  AOI22_X1 U18291 ( .A1(n9556), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11628), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14705) );
  NAND3_X1 U18292 ( .A1(n14707), .A2(n14706), .A3(n14705), .ZN(n14708) );
  NOR2_X1 U18293 ( .A1(n14709), .A2(n14708), .ZN(n18511) );
  INV_X1 U18294 ( .A(n18511), .ZN(n14716) );
  INV_X1 U18295 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17944) );
  INV_X1 U18296 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n18373) );
  NAND2_X1 U18297 ( .A1(n11836), .A2(n14713), .ZN(n18372) );
  NOR2_X1 U18298 ( .A1(n18373), .A2(n18372), .ZN(n18369) );
  AOI21_X1 U18299 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18369), .A(
        P3_EBX_REG_8__SCAN_IN), .ZN(n14714) );
  NOR2_X1 U18300 ( .A1(n18366), .A2(n14714), .ZN(n14715) );
  MUX2_X1 U18301 ( .A(n14716), .B(n14715), .S(n9564), .Z(P3_U2695) );
  AOI21_X1 U18302 ( .B1(n11722), .B2(n11723), .A(n18712), .ZN(n14721) );
  AOI21_X1 U18303 ( .B1(n14717), .B2(n17300), .A(n14721), .ZN(n14718) );
  AND2_X1 U18304 ( .A1(n14750), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14743) );
  NOR2_X1 U18305 ( .A1(n14718), .A2(n14743), .ZN(n14725) );
  NAND2_X1 U18306 ( .A1(n10316), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14719) );
  MUX2_X1 U18307 ( .A(n10316), .B(n14719), .S(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(n14724) );
  AND2_X1 U18308 ( .A1(n14720), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14723) );
  OAI22_X1 U18309 ( .A1(n14721), .A2(n14741), .B1(n10316), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14722) );
  OAI22_X2 U18310 ( .A1(n14725), .A2(n14724), .B1(n14723), .B2(n14722), .ZN(
        n14755) );
  NAND2_X1 U18311 ( .A1(n17160), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14726) );
  XNOR2_X1 U18312 ( .A(n14726), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14753) );
  NAND2_X1 U18313 ( .A1(n17159), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14727) );
  AOI22_X1 U18314 ( .A1(n14727), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n17159), .B2(n14743), .ZN(n14745) );
  NAND2_X1 U18315 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18799) );
  INV_X1 U18316 ( .A(n14729), .ZN(n14731) );
  NAND2_X1 U18317 ( .A1(n18536), .A2(n19737), .ZN(n19739) );
  NAND3_X1 U18318 ( .A1(n14730), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17166) );
  NOR2_X1 U18319 ( .A1(n17685), .A2(n17166), .ZN(n14733) );
  OR2_X1 U18320 ( .A1(n19479), .A2(n14733), .ZN(n17167) );
  OAI211_X1 U18321 ( .C1(n18737), .C2(n14731), .A(n18906), .B(n17167), .ZN(
        n17164) );
  NOR2_X1 U18322 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18725), .ZN(
        n17161) );
  NOR2_X1 U18323 ( .A1(n17164), .A2(n17161), .ZN(n14882) );
  NOR2_X1 U18324 ( .A1(n14882), .A2(n14734), .ZN(n14736) );
  NAND2_X1 U18325 ( .A1(n19479), .A2(n14732), .ZN(n18818) );
  XOR2_X1 U18326 ( .A(n14734), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n14735) );
  NAND2_X1 U18327 ( .A1(n19089), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n14748) );
  OAI21_X1 U18328 ( .B1(n14745), .B2(n18810), .A(n14737), .ZN(n14738) );
  AOI21_X1 U18329 ( .B1(n14753), .B2(n18904), .A(n14738), .ZN(n14739) );
  OAI21_X1 U18330 ( .B1(n14755), .B2(n18829), .A(n14739), .ZN(P3_U2799) );
  INV_X1 U18331 ( .A(n17276), .ZN(n14742) );
  AOI21_X1 U18332 ( .B1(n14742), .B2(n14741), .A(n14740), .ZN(n14751) );
  INV_X1 U18333 ( .A(n14743), .ZN(n14744) );
  NOR4_X1 U18334 ( .A1(n18909), .A2(n17315), .A3(n14877), .A4(n14744), .ZN(
        n14747) );
  NOR2_X1 U18335 ( .A1(n14745), .A2(n19048), .ZN(n14746) );
  OAI21_X1 U18336 ( .B1(n14747), .B2(n14746), .A(n19053), .ZN(n14749) );
  OAI211_X1 U18337 ( .C1(n14751), .C2(n14750), .A(n14749), .B(n14748), .ZN(
        n14752) );
  AOI21_X1 U18338 ( .B1(n14753), .B2(n19119), .A(n14752), .ZN(n14754) );
  OAI21_X1 U18339 ( .B1(n14755), .B2(n19058), .A(n14754), .ZN(P3_U2831) );
  NOR3_X1 U18340 ( .A1(n14756), .A2(n14766), .A3(n16362), .ZN(n14760) );
  AOI22_X1 U18341 ( .A1(P2_REIP_REG_31__SCAN_IN), .A2(n16288), .B1(n16337), 
        .B2(P2_EBX_REG_31__SCAN_IN), .ZN(n14757) );
  OAI21_X1 U18342 ( .B1(n14758), .B2(n16340), .A(n14757), .ZN(n14759) );
  NAND2_X1 U18343 ( .A1(n16440), .A2(n16342), .ZN(n14762) );
  OAI211_X1 U18344 ( .C1(n16369), .C2(n16304), .A(n14763), .B(n14762), .ZN(
        P2_U2824) );
  AOI21_X1 U18345 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14765), .ZN(n14768) );
  NAND2_X1 U18346 ( .A1(n16842), .A2(n14766), .ZN(n14767) );
  OAI211_X1 U18347 ( .C1(n14806), .C2(n19838), .A(n14768), .B(n14767), .ZN(
        n14769) );
  AOI21_X1 U18348 ( .B1(n13307), .B2(n14770), .A(n14769), .ZN(n14771) );
  OAI21_X1 U18349 ( .B1(n14772), .B2(n16863), .A(n14771), .ZN(P2_U2984) );
  XNOR2_X1 U18350 ( .A(n14774), .B(n14773), .ZN(n14801) );
  INV_X1 U18351 ( .A(n14801), .ZN(n14782) );
  XNOR2_X1 U18352 ( .A(n14776), .B(n14775), .ZN(n14793) );
  INV_X1 U18353 ( .A(n16320), .ZN(n14779) );
  INV_X1 U18354 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20496) );
  NOR2_X1 U18355 ( .A1(n16810), .A2(n20496), .ZN(n14803) );
  INV_X1 U18356 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14777) );
  NOR2_X1 U18357 ( .A1(n16839), .A2(n14777), .ZN(n14778) );
  AOI211_X1 U18358 ( .C1(n16842), .C2(n14779), .A(n14803), .B(n14778), .ZN(
        n14780) );
  OAI21_X1 U18359 ( .B1(n14793), .B2(n16846), .A(n14780), .ZN(n14781) );
  AOI21_X1 U18360 ( .B1(n16836), .B2(n14782), .A(n14781), .ZN(n14783) );
  OAI21_X1 U18361 ( .B1(n14784), .B2(n19838), .A(n14783), .ZN(P2_U3012) );
  INV_X1 U18362 ( .A(n14785), .ZN(n14796) );
  AOI21_X1 U18363 ( .B1(n14789), .B2(n14787), .A(n14786), .ZN(n14795) );
  AOI22_X1 U18364 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14790), .B1(
        n14789), .B2(n14788), .ZN(n14792) );
  OAI22_X1 U18365 ( .A1(n14793), .A2(n17124), .B1(n14792), .B2(n14791), .ZN(
        n14794) );
  AOI211_X1 U18366 ( .C1(n14796), .C2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n14795), .B(n14794), .ZN(n14805) );
  OR2_X1 U18367 ( .A1(n14798), .A2(n14797), .ZN(n14799) );
  NAND2_X1 U18368 ( .A1(n14800), .A2(n14799), .ZN(n20576) );
  NOR2_X1 U18369 ( .A1(n17139), .A2(n14801), .ZN(n14802) );
  AOI211_X1 U18370 ( .C1(n17121), .C2(n20576), .A(n14803), .B(n14802), .ZN(
        n14804) );
  NOR2_X1 U18371 ( .A1(n14806), .A2(n16438), .ZN(n14807) );
  AOI21_X1 U18372 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16438), .A(n14807), .ZN(
        n14808) );
  OAI21_X1 U18373 ( .B1(n14809), .B2(n16433), .A(n14808), .ZN(P2_U2857) );
  NAND2_X1 U18374 ( .A1(n14836), .A2(n9698), .ZN(n14814) );
  NAND2_X1 U18375 ( .A1(n14837), .A2(n14832), .ZN(n14813) );
  XNOR2_X1 U18376 ( .A(n14814), .B(n14813), .ZN(n16647) );
  XNOR2_X1 U18377 ( .A(n16654), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16645) );
  AND2_X1 U18378 ( .A1(n16088), .A2(n14817), .ZN(n14845) );
  INV_X1 U18379 ( .A(n14845), .ZN(n14816) );
  OAI21_X1 U18380 ( .B1(n16088), .B2(n14817), .A(n14816), .ZN(n16643) );
  NAND3_X1 U18381 ( .A1(n17031), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14818), .ZN(n14894) );
  INV_X1 U18382 ( .A(n14894), .ZN(n14823) );
  NOR2_X1 U18383 ( .A1(n16810), .A2(n20525), .ZN(n16641) );
  NOR2_X1 U18384 ( .A1(n17098), .A2(n14818), .ZN(n14819) );
  NOR2_X1 U18385 ( .A1(n17028), .A2(n14819), .ZN(n16953) );
  NOR2_X1 U18386 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n14820), .ZN(
        n14821) );
  NAND2_X1 U18387 ( .A1(n17031), .A2(n14821), .ZN(n16938) );
  AOI21_X1 U18388 ( .B1(n16953), .B2(n16938), .A(n14893), .ZN(n14822) );
  AOI211_X1 U18389 ( .C1(n14823), .C2(n14893), .A(n16641), .B(n14822), .ZN(
        n14829) );
  NAND2_X1 U18390 ( .A1(n16103), .A2(n14824), .ZN(n16086) );
  NAND2_X1 U18391 ( .A1(n16103), .A2(n14825), .ZN(n14889) );
  INV_X1 U18392 ( .A(n14889), .ZN(n14826) );
  AOI21_X1 U18393 ( .B1(n14827), .B2(n16086), .A(n14826), .ZN(n16515) );
  NAND2_X1 U18394 ( .A1(n16515), .A2(n17121), .ZN(n14828) );
  OAI211_X1 U18395 ( .C1(n16643), .C2(n17116), .A(n14829), .B(n14828), .ZN(
        n14830) );
  AOI21_X1 U18396 ( .B1(n16645), .B2(n17136), .A(n14830), .ZN(n14831) );
  OAI21_X1 U18397 ( .B1(n16647), .B2(n17139), .A(n14831), .ZN(P2_U3026) );
  INV_X1 U18398 ( .A(n14832), .ZN(n14834) );
  INV_X1 U18399 ( .A(n9698), .ZN(n14833) );
  NOR2_X1 U18400 ( .A1(n14834), .A2(n14833), .ZN(n14835) );
  XNOR2_X1 U18401 ( .A(n14840), .B(n10454), .ZN(n14902) );
  NAND2_X1 U18402 ( .A1(n16088), .A2(n14843), .ZN(n16052) );
  OAI21_X1 U18403 ( .B1(n14845), .B2(n14844), .A(n16052), .ZN(n16427) );
  NOR2_X1 U18404 ( .A1(n16810), .A2(n20527), .ZN(n14895) );
  AOI21_X1 U18405 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14895), .ZN(n14847) );
  NAND2_X1 U18406 ( .A1(n16842), .A2(n16066), .ZN(n14846) );
  OAI211_X1 U18407 ( .C1(n16427), .C2(n19838), .A(n14847), .B(n14846), .ZN(
        n14848) );
  OAI21_X1 U18408 ( .B1(n14902), .B2(n16863), .A(n14849), .ZN(P2_U2993) );
  NAND2_X1 U18409 ( .A1(n15533), .A2(n14951), .ZN(n14851) );
  OAI211_X1 U18410 ( .C1(n15530), .C2(n14952), .A(n14851), .B(n14850), .ZN(
        n14852) );
  AOI21_X1 U18411 ( .B1(n14950), .B2(n20778), .A(n14852), .ZN(n14853) );
  OAI21_X1 U18412 ( .B1(n20633), .B2(n14854), .A(n14853), .ZN(P1_U2969) );
  INV_X1 U18413 ( .A(n14856), .ZN(n14858) );
  NAND2_X1 U18414 ( .A1(n13750), .A2(n14857), .ZN(n14974) );
  NAND2_X1 U18415 ( .A1(n14905), .A2(n14859), .ZN(n14860) );
  NAND2_X1 U18416 ( .A1(n14977), .A2(n14860), .ZN(n14865) );
  OAI222_X1 U18417 ( .A1(n15437), .A2(n15330), .B1(n21565), .B2(n20712), .C1(
        n14865), .C2(n15328), .ZN(P1_U2845) );
  NAND3_X1 U18418 ( .A1(n15413), .A2(n14861), .A3(n20885), .ZN(n15390) );
  OAI22_X1 U18419 ( .A1(n15390), .A2(n15405), .B1(n15413), .B2(n21572), .ZN(
        n14862) );
  AOI21_X1 U18420 ( .B1(n15392), .B2(BUF1_REG_27__SCAN_IN), .A(n14862), .ZN(
        n14864) );
  NAND2_X1 U18421 ( .A1(n15393), .A2(DATAI_27_), .ZN(n14863) );
  OAI211_X1 U18422 ( .C1(n15437), .C2(n15415), .A(n14864), .B(n14863), .ZN(
        P1_U2877) );
  INV_X1 U18423 ( .A(n14865), .ZN(n15657) );
  INV_X1 U18424 ( .A(n15287), .ZN(n20690) );
  AND3_X1 U18425 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .ZN(n14866) );
  NAND2_X1 U18426 ( .A1(n14867), .A2(n14866), .ZN(n15000) );
  NOR2_X1 U18427 ( .A1(n15077), .A2(n15000), .ZN(n15014) );
  AND3_X1 U18428 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_26__SCAN_IN), .ZN(n14868) );
  NAND2_X1 U18429 ( .A1(n15014), .A2(n14868), .ZN(n14938) );
  INV_X1 U18430 ( .A(n15270), .ZN(n20689) );
  AOI21_X1 U18431 ( .B1(n20690), .B2(n14938), .A(n20689), .ZN(n14913) );
  INV_X1 U18432 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21495) );
  OAI22_X1 U18433 ( .A1(n9558), .A2(n15439), .B1(n14869), .B2(n20694), .ZN(
        n14871) );
  NOR3_X1 U18434 ( .A1(n15287), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14938), 
        .ZN(n14870) );
  AOI211_X1 U18435 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n20681), .A(n14871), .B(
        n14870), .ZN(n14872) );
  OAI21_X1 U18436 ( .B1(n14913), .B2(n21495), .A(n14872), .ZN(n14873) );
  AOI21_X1 U18437 ( .B1(n15657), .B2(n20693), .A(n14873), .ZN(n14874) );
  OAI21_X1 U18438 ( .B1(n15437), .B2(n15255), .A(n14874), .ZN(P1_U2813) );
  OAI22_X1 U18439 ( .A1(n17160), .A2(n18811), .B1(n17159), .B2(n18810), .ZN(
        n17171) );
  INV_X1 U18440 ( .A(n18795), .ZN(n14875) );
  INV_X1 U18441 ( .A(n18809), .ZN(n19078) );
  NAND2_X1 U18442 ( .A1(n18904), .A2(n19078), .ZN(n14876) );
  NAND2_X1 U18443 ( .A1(n17216), .A2(n14876), .ZN(n17226) );
  INV_X1 U18444 ( .A(n18985), .ZN(n17294) );
  NAND2_X1 U18445 ( .A1(n18780), .A2(n17176), .ZN(n17195) );
  NOR3_X1 U18446 ( .A1(n17195), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14877), .ZN(n14884) );
  NAND2_X1 U18447 ( .A1(n18824), .A2(n17672), .ZN(n14881) );
  AOI21_X1 U18448 ( .B1(n14879), .B2(n17675), .A(n14878), .ZN(n14880) );
  OAI211_X1 U18449 ( .C1(n14882), .C2(n17675), .A(n14881), .B(n14880), .ZN(
        n14883) );
  AOI211_X1 U18450 ( .C1(n17171), .C2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14884), .B(n14883), .ZN(n14885) );
  OAI21_X1 U18451 ( .B1(n14886), .B2(n18829), .A(n14885), .ZN(P3_U2800) );
  NAND2_X1 U18452 ( .A1(n16103), .A2(n14887), .ZN(n16061) );
  INV_X1 U18453 ( .A(n16061), .ZN(n14888) );
  AOI21_X1 U18454 ( .B1(n14890), .B2(n14889), .A(n14888), .ZN(n16507) );
  NAND2_X1 U18455 ( .A1(n16507), .A2(n17121), .ZN(n14899) );
  OR2_X1 U18456 ( .A1(n14891), .A2(n17032), .ZN(n16929) );
  INV_X1 U18457 ( .A(n16929), .ZN(n14897) );
  OAI21_X1 U18458 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(n14896) );
  AOI21_X1 U18459 ( .B1(n14897), .B2(n14896), .A(n14895), .ZN(n14898) );
  OAI211_X1 U18460 ( .C1(n16427), .C2(n17116), .A(n14899), .B(n14898), .ZN(
        n14900) );
  OAI21_X1 U18461 ( .B1(n14902), .B2(n17139), .A(n14901), .ZN(P2_U3025) );
  NAND2_X1 U18462 ( .A1(n14995), .A2(n14903), .ZN(n14904) );
  NAND2_X1 U18463 ( .A1(n14905), .A2(n14904), .ZN(n14916) );
  INV_X1 U18464 ( .A(n14916), .ZN(n15665) );
  INV_X1 U18465 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21493) );
  INV_X1 U18466 ( .A(n14906), .ZN(n14908) );
  OAI22_X1 U18467 ( .A1(n9558), .A2(n14908), .B1(n14907), .B2(n20694), .ZN(
        n14909) );
  AOI21_X1 U18468 ( .B1(n20691), .B2(P1_EBX_REG_26__SCAN_IN), .A(n14909), .ZN(
        n14912) );
  NAND2_X1 U18469 ( .A1(n15014), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14910) );
  NOR2_X1 U18470 ( .A1(n15287), .A2(n14910), .ZN(n14999) );
  NAND3_X1 U18471 ( .A1(n14999), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14938), 
        .ZN(n14911) );
  OAI211_X1 U18472 ( .C1(n14913), .C2(n21493), .A(n14912), .B(n14911), .ZN(
        n14914) );
  AOI21_X1 U18473 ( .B1(n15665), .B2(n20693), .A(n14914), .ZN(n14915) );
  OAI21_X1 U18474 ( .B1(n14922), .B2(n15255), .A(n14915), .ZN(P1_U2814) );
  OAI222_X1 U18475 ( .A1(n14922), .A2(n15330), .B1(n21666), .B2(n20712), .C1(
        n14916), .C2(n15328), .ZN(P1_U2846) );
  NAND2_X1 U18476 ( .A1(n20836), .A2(DATAI_10_), .ZN(n14918) );
  NAND2_X1 U18477 ( .A1(n20838), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14917) );
  AND2_X1 U18478 ( .A1(n14918), .A2(n14917), .ZN(n20746) );
  OAI22_X1 U18479 ( .A1(n15390), .A2(n20746), .B1(n15413), .B2(n14322), .ZN(
        n14919) );
  AOI21_X1 U18480 ( .B1(n15392), .B2(BUF1_REG_26__SCAN_IN), .A(n14919), .ZN(
        n14921) );
  NAND2_X1 U18481 ( .A1(n15393), .A2(DATAI_26_), .ZN(n14920) );
  OAI211_X1 U18482 ( .C1(n14922), .C2(n15415), .A(n14921), .B(n14920), .ZN(
        P1_U2878) );
  AOI21_X1 U18483 ( .B1(n12223), .B2(n15882), .A(n14923), .ZN(n15904) );
  INV_X1 U18484 ( .A(n14926), .ZN(n15898) );
  INV_X1 U18485 ( .A(n15931), .ZN(n15892) );
  AOI22_X1 U18486 ( .A1(n15892), .A2(n14930), .B1(n15883), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n14924) );
  OAI21_X1 U18487 ( .B1(n15904), .B2(n15898), .A(n14924), .ZN(n14927) );
  AND2_X1 U18488 ( .A1(n14925), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15902) );
  AOI22_X1 U18489 ( .A1(n14929), .A2(n14927), .B1(n14926), .B2(n15902), .ZN(
        n14928) );
  OAI21_X1 U18490 ( .B1(n14930), .B2(n14929), .A(n14928), .ZN(P1_U3474) );
  INV_X1 U18491 ( .A(n14931), .ZN(n14949) );
  MUX2_X1 U18492 ( .A(n14933), .B(n9577), .S(n14932), .Z(n14937) );
  INV_X1 U18493 ( .A(n14935), .ZN(n14936) );
  NAND2_X1 U18494 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14942) );
  NOR2_X1 U18495 ( .A1(n21495), .A2(n14938), .ZN(n14980) );
  AND2_X1 U18496 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n14980), .ZN(n14940) );
  NAND2_X1 U18497 ( .A1(n15270), .A2(n14940), .ZN(n14939) );
  AND2_X1 U18498 ( .A1(n20673), .A2(n14939), .ZN(n14979) );
  AOI21_X1 U18499 ( .B1(n20673), .B2(n14942), .A(n14979), .ZN(n14955) );
  AOI22_X1 U18500 ( .A1(n20681), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20674), .ZN(n14945) );
  INV_X1 U18501 ( .A(n14940), .ZN(n14941) );
  NOR2_X1 U18502 ( .A1(n15287), .A2(n14941), .ZN(n14968) );
  INV_X1 U18503 ( .A(n14942), .ZN(n14943) );
  NAND3_X1 U18504 ( .A1(n14968), .A2(n14943), .A3(n14946), .ZN(n14944) );
  OAI211_X1 U18505 ( .C1(n14955), .C2(n14946), .A(n14945), .B(n14944), .ZN(
        n14947) );
  OAI21_X1 U18506 ( .B1(n14949), .B2(n15255), .A(n14948), .ZN(P1_U2809) );
  NAND2_X1 U18507 ( .A1(n14950), .A2(n20668), .ZN(n14959) );
  INV_X1 U18508 ( .A(n14951), .ZN(n14953) );
  OAI22_X1 U18509 ( .A1(n9558), .A2(n14953), .B1(n14952), .B2(n20694), .ZN(
        n14957) );
  AOI21_X1 U18510 ( .B1(n14968), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14954) );
  NOR2_X1 U18511 ( .A1(n14955), .A2(n14954), .ZN(n14956) );
  AOI211_X1 U18512 ( .C1(n20681), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14957), .B(
        n14956), .ZN(n14958) );
  OAI211_X1 U18513 ( .C1(n14960), .C2(n20678), .A(n14959), .B(n14958), .ZN(
        P1_U2810) );
  XNOR2_X1 U18514 ( .A(n14976), .B(n14964), .ZN(n15635) );
  INV_X1 U18515 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21498) );
  NAND2_X1 U18516 ( .A1(n20691), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14966) );
  NAND2_X1 U18517 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14965) );
  OAI211_X1 U18518 ( .C1(n9558), .C2(n15418), .A(n14966), .B(n14965), .ZN(
        n14967) );
  AOI21_X1 U18519 ( .B1(n14968), .B2(n21498), .A(n14967), .ZN(n14970) );
  NAND2_X1 U18520 ( .A1(n14979), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14969) );
  OAI211_X1 U18521 ( .C1(n15635), .C2(n20678), .A(n14970), .B(n14969), .ZN(
        n14971) );
  AOI21_X1 U18522 ( .B1(n15420), .B2(n20668), .A(n14971), .ZN(n14972) );
  INV_X1 U18523 ( .A(n14972), .ZN(P1_U2811) );
  INV_X1 U18524 ( .A(n15430), .ZN(n15348) );
  AOI21_X1 U18525 ( .B1(n14978), .B2(n14977), .A(n14976), .ZN(n15644) );
  INV_X1 U18526 ( .A(n14979), .ZN(n14985) );
  AOI21_X1 U18527 ( .B1(n20690), .B2(n14980), .A(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14984) );
  OAI22_X1 U18528 ( .A1(n9558), .A2(n15428), .B1(n14981), .B2(n20694), .ZN(
        n14982) );
  AOI21_X1 U18529 ( .B1(n20691), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14982), .ZN(
        n14983) );
  OAI21_X1 U18530 ( .B1(n14985), .B2(n14984), .A(n14983), .ZN(n14986) );
  AOI21_X1 U18531 ( .B1(n15644), .B2(n20693), .A(n14986), .ZN(n14987) );
  OAI21_X1 U18532 ( .B1(n15348), .B2(n15255), .A(n14987), .ZN(P1_U2812) );
  INV_X1 U18533 ( .A(n14988), .ZN(n14992) );
  INV_X1 U18534 ( .A(n14989), .ZN(n14991) );
  INV_X1 U18535 ( .A(n13750), .ZN(n14990) );
  INV_X1 U18536 ( .A(n15353), .ZN(n15448) );
  OR2_X1 U18537 ( .A1(n15009), .A2(n14993), .ZN(n14994) );
  NAND2_X1 U18538 ( .A1(n14995), .A2(n14994), .ZN(n15678) );
  INV_X1 U18539 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21491) );
  NAND2_X1 U18540 ( .A1(n20691), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n14997) );
  NAND2_X1 U18541 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14996) );
  OAI211_X1 U18542 ( .C1(n9558), .C2(n15446), .A(n14997), .B(n14996), .ZN(
        n14998) );
  AOI21_X1 U18543 ( .B1(n14999), .B2(n21491), .A(n14998), .ZN(n15004) );
  AND2_X1 U18544 ( .A1(n20673), .A2(n15000), .ZN(n15001) );
  OR2_X1 U18545 ( .A1(n15107), .A2(n15001), .ZN(n15031) );
  NOR2_X1 U18546 ( .A1(n15287), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15002) );
  OAI21_X1 U18547 ( .B1(n15031), .B2(n15002), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15003) );
  OAI211_X1 U18548 ( .C1(n15678), .C2(n20678), .A(n15004), .B(n15003), .ZN(
        n15005) );
  AOI21_X1 U18549 ( .B1(n15448), .B2(n20668), .A(n15005), .ZN(n15006) );
  INV_X1 U18550 ( .A(n15006), .ZN(P1_U2815) );
  NOR2_X1 U18551 ( .A1(n15036), .A2(n15007), .ZN(n15008) );
  OR2_X1 U18552 ( .A1(n15009), .A2(n15008), .ZN(n15682) );
  OAI21_X1 U18553 ( .B1(n15011), .B2(n15012), .A(n14988), .ZN(n15360) );
  INV_X1 U18554 ( .A(n15360), .ZN(n15457) );
  NAND2_X1 U18555 ( .A1(n15457), .A2(n20668), .ZN(n15022) );
  INV_X1 U18556 ( .A(n15455), .ZN(n15013) );
  NAND2_X1 U18557 ( .A1(n15294), .A2(n15013), .ZN(n15019) );
  INV_X1 U18558 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21489) );
  NAND2_X1 U18559 ( .A1(n15014), .A2(n21489), .ZN(n15015) );
  OR2_X1 U18560 ( .A1(n15287), .A2(n15015), .ZN(n15018) );
  NAND2_X1 U18561 ( .A1(n20681), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n15017) );
  NAND2_X1 U18562 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15016) );
  NAND4_X1 U18563 ( .A1(n15019), .A2(n15018), .A3(n15017), .A4(n15016), .ZN(
        n15020) );
  AOI21_X1 U18564 ( .B1(n15031), .B2(P1_REIP_REG_24__SCAN_IN), .A(n15020), 
        .ZN(n15021) );
  OAI211_X1 U18565 ( .C1(n15682), .C2(n20678), .A(n15022), .B(n15021), .ZN(
        P1_U2816) );
  INV_X1 U18566 ( .A(n13764), .ZN(n15025) );
  INV_X1 U18567 ( .A(n15011), .ZN(n15023) );
  INV_X1 U18568 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15026) );
  OAI21_X1 U18569 ( .B1(n15027), .B2(n21486), .A(n15026), .ZN(n15032) );
  NAND2_X1 U18570 ( .A1(n20681), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n15029) );
  NAND2_X1 U18571 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15028) );
  OAI211_X1 U18572 ( .C1(n9558), .C2(n15463), .A(n15029), .B(n15028), .ZN(
        n15030) );
  AOI21_X1 U18573 ( .B1(n15032), .B2(n15031), .A(n15030), .ZN(n15038) );
  AND2_X1 U18574 ( .A1(n15034), .A2(n15033), .ZN(n15035) );
  NOR2_X1 U18575 ( .A1(n15036), .A2(n15035), .ZN(n15693) );
  NAND2_X1 U18576 ( .A1(n15693), .A2(n20693), .ZN(n15037) );
  OAI211_X1 U18577 ( .C1(n15461), .C2(n15255), .A(n15038), .B(n15037), .ZN(
        P1_U2817) );
  AOI21_X1 U18578 ( .B1(n15042), .B2(n15040), .A(n15041), .ZN(n15485) );
  INV_X1 U18579 ( .A(n15485), .ZN(n15373) );
  OR2_X1 U18580 ( .A1(n15056), .A2(n15043), .ZN(n15044) );
  NAND2_X1 U18581 ( .A1(n15045), .A2(n15044), .ZN(n15310) );
  INV_X1 U18582 ( .A(n15310), .ZN(n15726) );
  OAI22_X1 U18583 ( .A1(n9558), .A2(n15483), .B1(n15046), .B2(n20694), .ZN(
        n15047) );
  AOI21_X1 U18584 ( .B1(n20691), .B2(P1_EBX_REG_21__SCAN_IN), .A(n15047), .ZN(
        n15049) );
  OAI211_X1 U18585 ( .C1(n15064), .C2(n21484), .A(n15049), .B(n15048), .ZN(
        n15050) );
  AOI21_X1 U18586 ( .B1(n20693), .B2(n15726), .A(n15050), .ZN(n15051) );
  OAI21_X1 U18587 ( .B1(n15373), .B2(n15255), .A(n15051), .ZN(P1_U2819) );
  INV_X1 U18588 ( .A(n15052), .ZN(n15054) );
  INV_X1 U18589 ( .A(n15491), .ZN(n15067) );
  AOI21_X1 U18590 ( .B1(n10124), .B2(n15069), .A(n15055), .ZN(n15057) );
  OR2_X1 U18591 ( .A1(n15057), .A2(n15056), .ZN(n15730) );
  NOR2_X1 U18592 ( .A1(n15730), .A2(n20678), .ZN(n15066) );
  NOR2_X1 U18593 ( .A1(n15058), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15063) );
  INV_X1 U18594 ( .A(n15494), .ZN(n15059) );
  OAI22_X1 U18595 ( .A1(n9558), .A2(n15059), .B1(n15490), .B2(n20694), .ZN(
        n15060) );
  INV_X1 U18596 ( .A(n15060), .ZN(n15062) );
  NAND2_X1 U18597 ( .A1(n20691), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n15061) );
  OAI211_X1 U18598 ( .C1(n15064), .C2(n15063), .A(n15062), .B(n15061), .ZN(
        n15065) );
  AOI211_X1 U18599 ( .C1(n15067), .C2(n20668), .A(n15066), .B(n15065), .ZN(
        n15068) );
  INV_X1 U18600 ( .A(n15068), .ZN(P1_U2820) );
  XNOR2_X1 U18601 ( .A(n10124), .B(n15069), .ZN(n15743) );
  AOI21_X1 U18602 ( .B1(n15070), .B2(n15087), .A(n15071), .ZN(n15072) );
  NAND2_X1 U18603 ( .A1(n15503), .A2(n20668), .ZN(n15083) );
  INV_X1 U18604 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21479) );
  NOR3_X1 U18605 ( .A1(n15287), .A2(n15077), .A3(n21479), .ZN(n15075) );
  INV_X1 U18606 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21480) );
  NOR2_X1 U18607 ( .A1(n20694), .A2(n15073), .ZN(n15074) );
  AOI211_X1 U18608 ( .C1(n15075), .C2(n21480), .A(n20666), .B(n15074), .ZN(
        n15076) );
  OAI21_X1 U18609 ( .B1(n15501), .B2(n9558), .A(n15076), .ZN(n15081) );
  INV_X1 U18610 ( .A(n15107), .ZN(n15079) );
  OR2_X1 U18611 ( .A1(n15077), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15078) );
  OR2_X1 U18612 ( .A1(n15287), .A2(n15078), .ZN(n15092) );
  AOI21_X1 U18613 ( .B1(n15079), .B2(n15092), .A(n21480), .ZN(n15080) );
  AOI211_X1 U18614 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n20681), .A(n15081), .B(
        n15080), .ZN(n15082) );
  OAI211_X1 U18615 ( .C1(n15743), .C2(n20678), .A(n15083), .B(n15082), .ZN(
        P1_U2821) );
  OAI21_X1 U18616 ( .B1(n15121), .B2(n15104), .A(n15084), .ZN(n15086) );
  NAND2_X1 U18617 ( .A1(n15086), .A2(n15085), .ZN(n15757) );
  XNOR2_X1 U18618 ( .A(n15070), .B(n15087), .ZN(n15511) );
  INV_X1 U18619 ( .A(n15511), .ZN(n15088) );
  NAND2_X1 U18620 ( .A1(n15088), .A2(n20668), .ZN(n15097) );
  INV_X1 U18621 ( .A(n15089), .ZN(n15509) );
  NAND2_X1 U18622 ( .A1(n15294), .A2(n15509), .ZN(n15094) );
  NAND2_X1 U18623 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15090) );
  AND2_X1 U18624 ( .A1(n15090), .A2(n20771), .ZN(n15093) );
  NAND2_X1 U18625 ( .A1(n20681), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n15091) );
  NAND4_X1 U18626 ( .A1(n15094), .A2(n15093), .A3(n15092), .A4(n15091), .ZN(
        n15095) );
  AOI21_X1 U18627 ( .B1(n15107), .B2(P1_REIP_REG_18__SCAN_IN), .A(n15095), 
        .ZN(n15096) );
  OAI211_X1 U18628 ( .C1(n15757), .C2(n20678), .A(n15097), .B(n15096), .ZN(
        P1_U2822) );
  OAI21_X1 U18629 ( .B1(n13762), .B2(n15099), .A(n15098), .ZN(n15519) );
  INV_X1 U18630 ( .A(n15235), .ZN(n15100) );
  OR2_X1 U18631 ( .A1(n15287), .A2(n15100), .ZN(n15212) );
  NAND2_X1 U18632 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15113) );
  NOR2_X1 U18633 ( .A1(n15212), .A2(n15113), .ZN(n15170) );
  INV_X1 U18634 ( .A(n15117), .ZN(n15115) );
  NAND3_X1 U18635 ( .A1(n15170), .A2(n15115), .A3(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15125) );
  INV_X1 U18636 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21476) );
  INV_X1 U18637 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15101) );
  OAI21_X1 U18638 ( .B1(n15125), .B2(n21476), .A(n15101), .ZN(n15108) );
  OAI21_X1 U18639 ( .B1(n20694), .B2(n15518), .A(n20771), .ZN(n15102) );
  AOI21_X1 U18640 ( .B1(n15294), .B2(n15522), .A(n15102), .ZN(n15103) );
  OAI21_X1 U18641 ( .B1(n15228), .B2(n15315), .A(n15103), .ZN(n15106) );
  XNOR2_X1 U18642 ( .A(n15121), .B(n15104), .ZN(n15767) );
  NOR2_X1 U18643 ( .A1(n15767), .A2(n20678), .ZN(n15105) );
  AOI211_X1 U18644 ( .C1(n15108), .C2(n15107), .A(n15106), .B(n15105), .ZN(
        n15109) );
  OAI21_X1 U18645 ( .B1(n15519), .B2(n15255), .A(n15109), .ZN(P1_U2823) );
  INV_X1 U18646 ( .A(n13762), .ZN(n15111) );
  OAI21_X1 U18647 ( .B1(n15112), .B2(n15110), .A(n15111), .ZN(n15536) );
  NAND2_X1 U18648 ( .A1(n20673), .A2(n15113), .ZN(n15114) );
  OR2_X1 U18649 ( .A1(n15287), .A2(n15115), .ZN(n15116) );
  NAND2_X1 U18650 ( .A1(n15217), .A2(n15116), .ZN(n15159) );
  INV_X1 U18651 ( .A(n15159), .ZN(n15119) );
  NOR2_X1 U18652 ( .A1(n15117), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15118) );
  NAND2_X1 U18653 ( .A1(n15170), .A2(n15118), .ZN(n15143) );
  NAND2_X1 U18654 ( .A1(n15119), .A2(n15143), .ZN(n15130) );
  INV_X1 U18655 ( .A(n15139), .ZN(n15154) );
  OAI21_X1 U18656 ( .B1(n15154), .B2(n15137), .A(n15120), .ZN(n15122) );
  NAND2_X1 U18657 ( .A1(n15122), .A2(n15121), .ZN(n15777) );
  INV_X1 U18658 ( .A(n15532), .ZN(n15124) );
  NAND2_X1 U18659 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15123) );
  OAI211_X1 U18660 ( .C1(n9558), .C2(n15124), .A(n20771), .B(n15123), .ZN(
        n15127) );
  NOR2_X1 U18661 ( .A1(n15125), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15126) );
  AOI211_X1 U18662 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n20681), .A(n15127), .B(
        n15126), .ZN(n15128) );
  OAI21_X1 U18663 ( .B1(n20678), .B2(n15777), .A(n15128), .ZN(n15129) );
  AOI21_X1 U18664 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n15130), .A(n15129), 
        .ZN(n15131) );
  OAI21_X1 U18665 ( .B1(n15536), .B2(n15255), .A(n15131), .ZN(P1_U2824) );
  INV_X1 U18666 ( .A(n15132), .ZN(n15133) );
  NAND2_X1 U18667 ( .A1(n15132), .A2(n15163), .ZN(n15164) );
  OAI21_X1 U18668 ( .B1(n15193), .B2(n15133), .A(n15164), .ZN(n15134) );
  INV_X1 U18669 ( .A(n15110), .ZN(n15135) );
  INV_X1 U18670 ( .A(n15137), .ZN(n15138) );
  XNOR2_X1 U18671 ( .A(n15139), .B(n15138), .ZN(n15782) );
  NOR2_X1 U18672 ( .A1(n15782), .A2(n20678), .ZN(n15145) );
  NAND2_X1 U18673 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15140) );
  OAI211_X1 U18674 ( .C1(n9558), .C2(n15545), .A(n20771), .B(n15140), .ZN(
        n15141) );
  INV_X1 U18675 ( .A(n15141), .ZN(n15142) );
  OAI211_X1 U18676 ( .C1(n21557), .C2(n15228), .A(n15143), .B(n15142), .ZN(
        n15144) );
  AOI211_X1 U18677 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15159), .A(n15145), 
        .B(n15144), .ZN(n15146) );
  OAI21_X1 U18678 ( .B1(n15543), .B2(n15255), .A(n15146), .ZN(P1_U2825) );
  INV_X1 U18679 ( .A(n15147), .ZN(n15150) );
  INV_X1 U18680 ( .A(n15166), .ZN(n15149) );
  AOI21_X1 U18681 ( .B1(n15150), .B2(n15149), .A(n15148), .ZN(n15558) );
  INV_X1 U18682 ( .A(n15558), .ZN(n15399) );
  AOI21_X1 U18683 ( .B1(n20674), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20666), .ZN(n15151) );
  OAI21_X1 U18684 ( .B1(n9558), .B2(n15556), .A(n15151), .ZN(n15157) );
  INV_X1 U18685 ( .A(n15184), .ZN(n15153) );
  OAI21_X1 U18686 ( .B1(n15153), .B2(n15168), .A(n15152), .ZN(n15155) );
  NAND2_X1 U18687 ( .A1(n15155), .A2(n15154), .ZN(n15794) );
  NOR2_X1 U18688 ( .A1(n15794), .A2(n20678), .ZN(n15156) );
  AOI211_X1 U18689 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n20681), .A(n15157), .B(
        n15156), .ZN(n15162) );
  INV_X1 U18690 ( .A(n15170), .ZN(n15198) );
  NAND3_X1 U18691 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n15158) );
  NOR2_X1 U18692 ( .A1(n15198), .A2(n15158), .ZN(n15160) );
  OAI21_X1 U18693 ( .B1(n15160), .B2(P1_REIP_REG_14__SCAN_IN), .A(n15159), 
        .ZN(n15161) );
  OAI211_X1 U18694 ( .C1(n15399), .C2(n15255), .A(n15162), .B(n15161), .ZN(
        P1_U2826) );
  OAI21_X1 U18695 ( .B1(n15132), .B2(n15163), .A(n15164), .ZN(n15192) );
  OAI21_X1 U18696 ( .B1(n15192), .B2(n15193), .A(n15164), .ZN(n15180) );
  NAND2_X1 U18697 ( .A1(n15180), .A2(n15179), .ZN(n15178) );
  INV_X1 U18698 ( .A(n15165), .ZN(n15167) );
  AOI21_X1 U18699 ( .B1(n15178), .B2(n15167), .A(n15166), .ZN(n15570) );
  INV_X1 U18700 ( .A(n15570), .ZN(n15403) );
  INV_X1 U18701 ( .A(n20673), .ZN(n15257) );
  OAI21_X1 U18702 ( .B1(n15257), .B2(n15169), .A(n15217), .ZN(n15188) );
  XNOR2_X1 U18703 ( .A(n15184), .B(n15168), .ZN(n15806) );
  INV_X1 U18704 ( .A(n15806), .ZN(n15175) );
  INV_X1 U18705 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21470) );
  NAND3_X1 U18706 ( .A1(n15170), .A2(n15169), .A3(n21470), .ZN(n15174) );
  NAND2_X1 U18707 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15171) );
  OAI211_X1 U18708 ( .C1(n9558), .C2(n15568), .A(n20771), .B(n15171), .ZN(
        n15172) );
  AOI21_X1 U18709 ( .B1(n20691), .B2(P1_EBX_REG_13__SCAN_IN), .A(n15172), .ZN(
        n15173) );
  OAI211_X1 U18710 ( .C1(n15175), .C2(n20678), .A(n15174), .B(n15173), .ZN(
        n15176) );
  AOI21_X1 U18711 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15188), .A(n15176), 
        .ZN(n15177) );
  OAI21_X1 U18712 ( .B1(n15403), .B2(n15255), .A(n15177), .ZN(P1_U2827) );
  OAI21_X1 U18713 ( .B1(n15180), .B2(n15179), .A(n15178), .ZN(n15576) );
  AOI21_X1 U18714 ( .B1(n20674), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20666), .ZN(n15181) );
  OAI21_X1 U18715 ( .B1(n9558), .B2(n15578), .A(n15181), .ZN(n15187) );
  INV_X1 U18716 ( .A(n15207), .ZN(n15183) );
  AOI21_X1 U18717 ( .B1(n15183), .B2(n15194), .A(n15182), .ZN(n15185) );
  OR2_X1 U18718 ( .A1(n15185), .A2(n15184), .ZN(n15820) );
  NOR2_X1 U18719 ( .A1(n20678), .A2(n15820), .ZN(n15186) );
  AOI211_X1 U18720 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n20681), .A(n15187), .B(
        n15186), .ZN(n15191) );
  INV_X1 U18721 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21466) );
  NOR2_X1 U18722 ( .A1(n15198), .A2(n21466), .ZN(n15189) );
  OAI21_X1 U18723 ( .B1(n15189), .B2(P1_REIP_REG_12__SCAN_IN), .A(n15188), 
        .ZN(n15190) );
  OAI211_X1 U18724 ( .C1(n15576), .C2(n15255), .A(n15191), .B(n15190), .ZN(
        P1_U2828) );
  XOR2_X1 U18725 ( .A(n15193), .B(n15192), .Z(n15591) );
  NAND2_X1 U18726 ( .A1(n15591), .A2(n20668), .ZN(n15201) );
  XNOR2_X1 U18727 ( .A(n15207), .B(n15194), .ZN(n15830) );
  AOI21_X1 U18728 ( .B1(n20674), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20666), .ZN(n15195) );
  OAI21_X1 U18729 ( .B1(n9558), .B2(n15589), .A(n15195), .ZN(n15196) );
  AOI21_X1 U18730 ( .B1(n20691), .B2(P1_EBX_REG_11__SCAN_IN), .A(n15196), .ZN(
        n15197) );
  OAI21_X1 U18731 ( .B1(n15198), .B2(P1_REIP_REG_11__SCAN_IN), .A(n15197), 
        .ZN(n15199) );
  AOI21_X1 U18732 ( .B1(n20693), .B2(n15830), .A(n15199), .ZN(n15200) );
  OAI211_X1 U18733 ( .C1(n15217), .C2(n21466), .A(n15201), .B(n15200), .ZN(
        P1_U2829) );
  NAND2_X1 U18734 ( .A1(n15202), .A2(n15203), .ZN(n15204) );
  AND2_X1 U18735 ( .A1(n15133), .A2(n15204), .ZN(n15604) );
  INV_X1 U18736 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15216) );
  NAND2_X1 U18737 ( .A1(n15226), .A2(n15205), .ZN(n15206) );
  NAND2_X1 U18738 ( .A1(n15207), .A2(n15206), .ZN(n15850) );
  INV_X1 U18739 ( .A(n15850), .ZN(n15208) );
  AOI22_X1 U18740 ( .A1(n20693), .A2(n15208), .B1(n20691), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n15209) );
  OAI211_X1 U18741 ( .C1(n20694), .C2(n15210), .A(n15209), .B(n20771), .ZN(
        n15211) );
  AOI21_X1 U18742 ( .B1(n15294), .B2(n15600), .A(n15211), .ZN(n15215) );
  INV_X1 U18743 ( .A(n15212), .ZN(n15213) );
  NAND3_X1 U18744 ( .A1(n15213), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n15216), 
        .ZN(n15214) );
  OAI211_X1 U18745 ( .C1(n15217), .C2(n15216), .A(n15215), .B(n15214), .ZN(
        n15218) );
  AOI21_X1 U18746 ( .B1(n15604), .B2(n20668), .A(n15218), .ZN(n15219) );
  INV_X1 U18747 ( .A(n15219), .ZN(P1_U2830) );
  OAI21_X1 U18748 ( .B1(n15221), .B2(n15222), .A(n15202), .ZN(n15608) );
  OR2_X1 U18749 ( .A1(n15224), .A2(n15223), .ZN(n15225) );
  NAND2_X1 U18750 ( .A1(n15226), .A2(n15225), .ZN(n15857) );
  INV_X1 U18751 ( .A(n15857), .ZN(n15234) );
  INV_X1 U18752 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21464) );
  OAI22_X1 U18753 ( .A1(n15242), .A2(n21464), .B1(n15228), .B2(n15227), .ZN(
        n15229) );
  INV_X1 U18754 ( .A(n15229), .ZN(n15230) );
  OAI211_X1 U18755 ( .C1(n20694), .C2(n15231), .A(n15230), .B(n20771), .ZN(
        n15233) );
  NOR2_X1 U18756 ( .A1(n9558), .A2(n15610), .ZN(n15232) );
  AOI211_X1 U18757 ( .C1(n15234), .C2(n20693), .A(n15233), .B(n15232), .ZN(
        n15237) );
  NAND3_X1 U18758 ( .A1(n20690), .A2(n15235), .A3(n21464), .ZN(n15236) );
  OAI211_X1 U18759 ( .C1(n15608), .C2(n15255), .A(n15237), .B(n15236), .ZN(
        P1_U2831) );
  INV_X1 U18760 ( .A(n15238), .ZN(n15241) );
  INV_X1 U18761 ( .A(n15239), .ZN(n15240) );
  AOI21_X1 U18762 ( .B1(n15241), .B2(n15240), .A(n15221), .ZN(n15618) );
  INV_X1 U18763 ( .A(n15618), .ZN(n15411) );
  INV_X1 U18764 ( .A(n15242), .ZN(n15251) );
  AOI21_X1 U18765 ( .B1(n20674), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20666), .ZN(n15243) );
  OAI21_X1 U18766 ( .B1(n9558), .B2(n15616), .A(n15243), .ZN(n15244) );
  AOI21_X1 U18767 ( .B1(n20691), .B2(P1_EBX_REG_8__SCAN_IN), .A(n15244), .ZN(
        n15245) );
  OAI21_X1 U18768 ( .B1(n20678), .B2(n15323), .A(n15245), .ZN(n15250) );
  NAND2_X1 U18769 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n15247) );
  INV_X1 U18770 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n15246) );
  NOR2_X1 U18771 ( .A1(n15247), .A2(n20700), .ZN(n15267) );
  NAND2_X1 U18772 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n15267), .ZN(n20688) );
  NOR3_X1 U18773 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n15248), .A3(n20688), .ZN(
        n15249) );
  AOI211_X1 U18774 ( .C1(P1_REIP_REG_8__SCAN_IN), .C2(n15251), .A(n15250), .B(
        n15249), .ZN(n15252) );
  OAI21_X1 U18775 ( .B1(n15411), .B2(n15255), .A(n15252), .ZN(P1_U2832) );
  NAND2_X1 U18776 ( .A1(n21521), .A2(n15253), .ZN(n15254) );
  INV_X1 U18777 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21457) );
  NOR2_X1 U18778 ( .A1(n20689), .A2(n15256), .ZN(n20684) );
  NOR3_X1 U18779 ( .A1(n20684), .A2(n15257), .A3(n21457), .ZN(n15266) );
  NAND2_X1 U18780 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15258) );
  OAI211_X1 U18781 ( .C1(n9558), .C2(n20782), .A(n20771), .B(n15258), .ZN(
        n15259) );
  AOI21_X1 U18782 ( .B1(n20681), .B2(P1_EBX_REG_4__SCAN_IN), .A(n15259), .ZN(
        n15264) );
  NOR2_X1 U18783 ( .A1(n15261), .A2(n15260), .ZN(n20698) );
  NAND2_X1 U18784 ( .A1(n15262), .A2(n20698), .ZN(n15263) );
  OAI211_X1 U18785 ( .C1(n20787), .C2(n20678), .A(n15264), .B(n15263), .ZN(
        n15265) );
  AOI211_X1 U18786 ( .C1(n15267), .C2(n21457), .A(n15266), .B(n15265), .ZN(
        n15268) );
  OAI21_X1 U18787 ( .B1(n15269), .B2(n20672), .A(n15268), .ZN(P1_U2836) );
  OR2_X1 U18788 ( .A1(n14260), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n15278) );
  NAND2_X1 U18789 ( .A1(n20681), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n15273) );
  OAI221_X1 U18790 ( .B1(n15287), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n15287), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n15270), .ZN(n15271) );
  AOI22_X1 U18791 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n15271), .ZN(n15272) );
  OAI211_X1 U18792 ( .C1(n9558), .C2(n15274), .A(n15273), .B(n15272), .ZN(
        n15275) );
  INV_X1 U18793 ( .A(n15275), .ZN(n15277) );
  NAND2_X1 U18794 ( .A1(n20693), .A2(n20798), .ZN(n15276) );
  OAI211_X1 U18795 ( .C1(n15278), .C2(n20700), .A(n15277), .B(n15276), .ZN(
        n15279) );
  AOI21_X1 U18796 ( .B1(n20698), .B2(n21119), .A(n15279), .ZN(n15280) );
  OAI21_X1 U18797 ( .B1(n15281), .B2(n20672), .A(n15280), .ZN(P1_U2837) );
  INV_X1 U18798 ( .A(n15282), .ZN(n20822) );
  AOI22_X1 U18799 ( .A1(n20693), .A2(n20822), .B1(n20691), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n15291) );
  AOI22_X1 U18800 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20689), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n15286) );
  NAND2_X1 U18801 ( .A1(n20698), .A2(n21329), .ZN(n15285) );
  OAI211_X1 U18802 ( .C1(n9558), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15286), .B(n15285), .ZN(n15289) );
  NOR2_X1 U18803 ( .A1(n15287), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n15288) );
  NOR2_X1 U18804 ( .A1(n15289), .A2(n15288), .ZN(n15290) );
  OAI211_X1 U18805 ( .C1(n15292), .C2(n20672), .A(n15291), .B(n15290), .ZN(
        P1_U2839) );
  INV_X1 U18806 ( .A(n20698), .ZN(n15298) );
  AOI22_X1 U18807 ( .A1(n20693), .A2(n15293), .B1(n20691), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n15296) );
  OAI21_X1 U18808 ( .B1(n15294), .B2(n20674), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15295) );
  OAI211_X1 U18809 ( .C1(n15298), .C2(n15297), .A(n15296), .B(n15295), .ZN(
        n15299) );
  AOI21_X1 U18810 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n20673), .A(n15299), .ZN(
        n15300) );
  OAI21_X1 U18811 ( .B1(n20672), .B2(n15301), .A(n15300), .ZN(P1_U2840) );
  INV_X1 U18812 ( .A(n15627), .ZN(n15303) );
  INV_X1 U18813 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15302) );
  OAI22_X1 U18814 ( .A1(n15303), .A2(n15328), .B1(n20712), .B2(n15302), .ZN(
        P1_U2841) );
  OAI222_X1 U18815 ( .A1(n15343), .A2(n15330), .B1(n15304), .B2(n20712), .C1(
        n15328), .C2(n15635), .ZN(P1_U2843) );
  AOI22_X1 U18816 ( .A1(n15644), .A2(n20707), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n15320), .ZN(n15305) );
  OAI21_X1 U18817 ( .B1(n15348), .B2(n15330), .A(n15305), .ZN(P1_U2844) );
  OAI222_X1 U18818 ( .A1(n15353), .A2(n15330), .B1(n15306), .B2(n20712), .C1(
        n15678), .C2(n15328), .ZN(P1_U2847) );
  INV_X1 U18819 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15307) );
  OAI222_X1 U18820 ( .A1(n15360), .A2(n15330), .B1(n15307), .B2(n20712), .C1(
        n15682), .C2(n15328), .ZN(P1_U2848) );
  AOI22_X1 U18821 ( .A1(n15693), .A2(n20707), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n15320), .ZN(n15308) );
  OAI21_X1 U18822 ( .B1(n15461), .B2(n15330), .A(n15308), .ZN(P1_U2849) );
  INV_X1 U18823 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15309) );
  OAI222_X1 U18824 ( .A1(n15472), .A2(n15330), .B1(n15309), .B2(n20712), .C1(
        n15701), .C2(n15328), .ZN(P1_U2850) );
  OAI222_X1 U18825 ( .A1(n15373), .A2(n15330), .B1(n15311), .B2(n20712), .C1(
        n15310), .C2(n15328), .ZN(P1_U2851) );
  OAI222_X1 U18826 ( .A1(n15491), .A2(n15330), .B1(n15312), .B2(n20712), .C1(
        n15730), .C2(n15328), .ZN(P1_U2852) );
  INV_X1 U18827 ( .A(n15503), .ZN(n15380) );
  OAI222_X1 U18828 ( .A1(n15380), .A2(n15330), .B1(n15313), .B2(n20712), .C1(
        n15328), .C2(n15743), .ZN(P1_U2853) );
  INV_X1 U18829 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15314) );
  OAI222_X1 U18830 ( .A1(n15757), .A2(n15328), .B1(n15314), .B2(n20712), .C1(
        n15330), .C2(n15511), .ZN(P1_U2854) );
  OAI222_X1 U18831 ( .A1(n15519), .A2(n15330), .B1(n15315), .B2(n20712), .C1(
        n15328), .C2(n15767), .ZN(P1_U2855) );
  INV_X1 U18832 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15316) );
  OAI222_X1 U18833 ( .A1(n15536), .A2(n15330), .B1(n15316), .B2(n20712), .C1(
        n15777), .C2(n15328), .ZN(P1_U2856) );
  OAI222_X1 U18834 ( .A1(n15543), .A2(n15330), .B1(n21557), .B2(n20712), .C1(
        n15328), .C2(n15782), .ZN(P1_U2857) );
  INV_X1 U18835 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15317) );
  OAI222_X1 U18836 ( .A1(n15399), .A2(n15330), .B1(n15317), .B2(n20712), .C1(
        n15794), .C2(n15328), .ZN(P1_U2858) );
  AOI22_X1 U18837 ( .A1(n15806), .A2(n20707), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n15320), .ZN(n15318) );
  OAI21_X1 U18838 ( .B1(n15403), .B2(n15330), .A(n15318), .ZN(P1_U2859) );
  OAI222_X1 U18839 ( .A1(n15820), .A2(n15328), .B1(n15319), .B2(n20712), .C1(
        n15576), .C2(n15330), .ZN(P1_U2860) );
  INV_X1 U18840 ( .A(n15591), .ZN(n15406) );
  AOI22_X1 U18841 ( .A1(n15830), .A2(n20707), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n15320), .ZN(n15321) );
  OAI21_X1 U18842 ( .B1(n15406), .B2(n15330), .A(n15321), .ZN(P1_U2861) );
  INV_X1 U18843 ( .A(n15604), .ZN(n15407) );
  INV_X1 U18844 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15322) );
  OAI222_X1 U18845 ( .A1(n15407), .A2(n15330), .B1(n15322), .B2(n20712), .C1(
        n15850), .C2(n15328), .ZN(P1_U2862) );
  OAI222_X1 U18846 ( .A1(n15608), .A2(n15330), .B1(n20712), .B2(n15227), .C1(
        n15857), .C2(n15328), .ZN(P1_U2863) );
  OAI222_X1 U18847 ( .A1(n15411), .A2(n15330), .B1(n15324), .B2(n20712), .C1(
        n15323), .C2(n15328), .ZN(P1_U2864) );
  AOI21_X1 U18848 ( .B1(n15326), .B2(n15325), .A(n15239), .ZN(n20658) );
  INV_X1 U18849 ( .A(n20658), .ZN(n15414) );
  XNOR2_X1 U18850 ( .A(n14617), .B(n15327), .ZN(n20655) );
  OAI222_X1 U18851 ( .A1(n15330), .A2(n15414), .B1(n15329), .B2(n20712), .C1(
        n15328), .C2(n20655), .ZN(P1_U2865) );
  NAND2_X1 U18852 ( .A1(n20836), .A2(DATAI_14_), .ZN(n15332) );
  NAND2_X1 U18853 ( .A1(n20838), .A2(BUF1_REG_14__SCAN_IN), .ZN(n15331) );
  AND2_X1 U18854 ( .A1(n15332), .A2(n15331), .ZN(n20754) );
  OAI22_X1 U18855 ( .A1(n15390), .A2(n20754), .B1(n15413), .B2(n15333), .ZN(
        n15334) );
  AOI21_X1 U18856 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n15392), .A(n15334), .ZN(
        n15336) );
  NAND2_X1 U18857 ( .A1(n15393), .A2(DATAI_30_), .ZN(n15335) );
  OAI211_X1 U18858 ( .C1(n15337), .C2(n15415), .A(n15336), .B(n15335), .ZN(
        P1_U2874) );
  INV_X1 U18859 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n17568) );
  INV_X1 U18860 ( .A(n15390), .ZN(n15385) );
  INV_X1 U18861 ( .A(DATAI_13_), .ZN(n15339) );
  NAND2_X1 U18862 ( .A1(n20838), .A2(BUF1_REG_13__SCAN_IN), .ZN(n15338) );
  OAI21_X1 U18863 ( .B1(n20838), .B2(n15339), .A(n15338), .ZN(n20752) );
  AOI22_X1 U18864 ( .A1(n15385), .A2(n20752), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15400), .ZN(n15340) );
  OAI21_X1 U18865 ( .B1(n15387), .B2(n17568), .A(n15340), .ZN(n15341) );
  AOI21_X1 U18866 ( .B1(n15393), .B2(DATAI_29_), .A(n15341), .ZN(n15342) );
  OAI21_X1 U18867 ( .B1(n15343), .B2(n15415), .A(n15342), .ZN(P1_U2875) );
  INV_X1 U18868 ( .A(DATAI_12_), .ZN(n15344) );
  INV_X1 U18869 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17588) );
  MUX2_X1 U18870 ( .A(n15344), .B(n17588), .S(n20838), .Z(n20749) );
  OAI22_X1 U18871 ( .A1(n15390), .A2(n20749), .B1(n15413), .B2(n14312), .ZN(
        n15345) );
  AOI21_X1 U18872 ( .B1(n15392), .B2(BUF1_REG_28__SCAN_IN), .A(n15345), .ZN(
        n15347) );
  NAND2_X1 U18873 ( .A1(n15393), .A2(DATAI_28_), .ZN(n15346) );
  OAI211_X1 U18874 ( .C1(n15348), .C2(n15415), .A(n15347), .B(n15346), .ZN(
        P1_U2876) );
  OAI22_X1 U18875 ( .A1(n15390), .A2(n15408), .B1(n15413), .B2(n15349), .ZN(
        n15350) );
  AOI21_X1 U18876 ( .B1(n15392), .B2(BUF1_REG_25__SCAN_IN), .A(n15350), .ZN(
        n15352) );
  NAND2_X1 U18877 ( .A1(n15393), .A2(DATAI_25_), .ZN(n15351) );
  OAI211_X1 U18878 ( .C1(n15353), .C2(n15415), .A(n15352), .B(n15351), .ZN(
        P1_U2879) );
  NAND2_X1 U18879 ( .A1(n20836), .A2(DATAI_8_), .ZN(n15355) );
  NAND2_X1 U18880 ( .A1(n20838), .A2(BUF1_REG_8__SCAN_IN), .ZN(n15354) );
  AND2_X1 U18881 ( .A1(n15355), .A2(n15354), .ZN(n20743) );
  OAI22_X1 U18882 ( .A1(n15390), .A2(n20743), .B1(n15413), .B2(n15356), .ZN(
        n15357) );
  AOI21_X1 U18883 ( .B1(n15392), .B2(BUF1_REG_24__SCAN_IN), .A(n15357), .ZN(
        n15359) );
  NAND2_X1 U18884 ( .A1(n15393), .A2(DATAI_24_), .ZN(n15358) );
  OAI211_X1 U18885 ( .C1(n15360), .C2(n15415), .A(n15359), .B(n15358), .ZN(
        P1_U2880) );
  OAI22_X1 U18886 ( .A1(n15390), .A2(n20888), .B1(n15413), .B2(n15361), .ZN(
        n15362) );
  AOI21_X1 U18887 ( .B1(n15392), .B2(BUF1_REG_23__SCAN_IN), .A(n15362), .ZN(
        n15364) );
  NAND2_X1 U18888 ( .A1(n15393), .A2(DATAI_23_), .ZN(n15363) );
  OAI211_X1 U18889 ( .C1(n15461), .C2(n15415), .A(n15364), .B(n15363), .ZN(
        P1_U2881) );
  INV_X1 U18890 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15365) );
  OAI22_X1 U18891 ( .A1(n15390), .A2(n20880), .B1(n15413), .B2(n15365), .ZN(
        n15366) );
  AOI21_X1 U18892 ( .B1(n15392), .B2(BUF1_REG_22__SCAN_IN), .A(n15366), .ZN(
        n15368) );
  NAND2_X1 U18893 ( .A1(n15393), .A2(DATAI_22_), .ZN(n15367) );
  OAI211_X1 U18894 ( .C1(n15472), .C2(n15415), .A(n15368), .B(n15367), .ZN(
        P1_U2882) );
  OAI22_X1 U18895 ( .A1(n15390), .A2(n20875), .B1(n15413), .B2(n15369), .ZN(
        n15370) );
  AOI21_X1 U18896 ( .B1(n15392), .B2(BUF1_REG_21__SCAN_IN), .A(n15370), .ZN(
        n15372) );
  NAND2_X1 U18897 ( .A1(n15393), .A2(DATAI_21_), .ZN(n15371) );
  OAI211_X1 U18898 ( .C1(n15373), .C2(n15415), .A(n15372), .B(n15371), .ZN(
        P1_U2883) );
  OAI22_X1 U18899 ( .A1(n15390), .A2(n20871), .B1(n15413), .B2(n14320), .ZN(
        n15374) );
  AOI21_X1 U18900 ( .B1(n15392), .B2(BUF1_REG_20__SCAN_IN), .A(n15374), .ZN(
        n15376) );
  NAND2_X1 U18901 ( .A1(n15393), .A2(DATAI_20_), .ZN(n15375) );
  OAI211_X1 U18902 ( .C1(n15491), .C2(n15415), .A(n15376), .B(n15375), .ZN(
        P1_U2884) );
  INV_X1 U18903 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U18904 ( .A1(n15385), .A2(n20866), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15400), .ZN(n15377) );
  OAI21_X1 U18905 ( .B1(n15387), .B2(n19868), .A(n15377), .ZN(n15378) );
  AOI21_X1 U18906 ( .B1(n15393), .B2(DATAI_19_), .A(n15378), .ZN(n15379) );
  OAI21_X1 U18907 ( .B1(n15380), .B2(n15415), .A(n15379), .ZN(P1_U2885) );
  OAI22_X1 U18908 ( .A1(n15390), .A2(n20861), .B1(n15413), .B2(n15381), .ZN(
        n15382) );
  AOI21_X1 U18909 ( .B1(n15392), .B2(BUF1_REG_18__SCAN_IN), .A(n15382), .ZN(
        n15384) );
  NAND2_X1 U18910 ( .A1(n15393), .A2(DATAI_18_), .ZN(n15383) );
  OAI211_X1 U18911 ( .C1(n15511), .C2(n15415), .A(n15384), .B(n15383), .ZN(
        P1_U2886) );
  INV_X1 U18912 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n17580) );
  AOI22_X1 U18913 ( .A1(n15385), .A2(n20856), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n15400), .ZN(n15386) );
  OAI21_X1 U18914 ( .B1(n15387), .B2(n17580), .A(n15386), .ZN(n15388) );
  AOI21_X1 U18915 ( .B1(n15393), .B2(DATAI_17_), .A(n15388), .ZN(n15389) );
  OAI21_X1 U18916 ( .B1(n15519), .B2(n15415), .A(n15389), .ZN(P1_U2887) );
  OAI22_X1 U18917 ( .A1(n15390), .A2(n20847), .B1(n15413), .B2(n14310), .ZN(
        n15391) );
  AOI21_X1 U18918 ( .B1(n15392), .B2(BUF1_REG_16__SCAN_IN), .A(n15391), .ZN(
        n15395) );
  NAND2_X1 U18919 ( .A1(n15393), .A2(DATAI_16_), .ZN(n15394) );
  OAI211_X1 U18920 ( .C1(n15536), .C2(n15415), .A(n15395), .B(n15394), .ZN(
        P1_U2888) );
  AOI22_X1 U18921 ( .A1(n15401), .A2(n15396), .B1(n15400), .B2(
        P1_EAX_REG_15__SCAN_IN), .ZN(n15397) );
  OAI21_X1 U18922 ( .B1(n15543), .B2(n15415), .A(n15397), .ZN(P1_U2889) );
  INV_X1 U18923 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15398) );
  OAI222_X1 U18924 ( .A1(n15399), .A2(n15415), .B1(n15398), .B2(n15413), .C1(
        n15412), .C2(n20754), .ZN(P1_U2890) );
  AOI22_X1 U18925 ( .A1(n15401), .A2(n20752), .B1(n15400), .B2(
        P1_EAX_REG_13__SCAN_IN), .ZN(n15402) );
  OAI21_X1 U18926 ( .B1(n15403), .B2(n15415), .A(n15402), .ZN(P1_U2891) );
  INV_X1 U18927 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15404) );
  OAI222_X1 U18928 ( .A1(n15576), .A2(n15415), .B1(n15404), .B2(n15413), .C1(
        n15412), .C2(n20749), .ZN(P1_U2892) );
  OAI222_X1 U18929 ( .A1(n15406), .A2(n15415), .B1(n21575), .B2(n15413), .C1(
        n15412), .C2(n15405), .ZN(P1_U2893) );
  OAI222_X1 U18930 ( .A1(n15407), .A2(n15415), .B1(n20726), .B2(n15413), .C1(
        n15412), .C2(n20746), .ZN(P1_U2894) );
  INV_X1 U18931 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15409) );
  OAI222_X1 U18932 ( .A1(n15608), .A2(n15415), .B1(n15409), .B2(n15413), .C1(
        n15412), .C2(n15408), .ZN(P1_U2895) );
  INV_X1 U18933 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n15410) );
  OAI222_X1 U18934 ( .A1(n15411), .A2(n15415), .B1(n15410), .B2(n15413), .C1(
        n15412), .C2(n20743), .ZN(P1_U2896) );
  OAI222_X1 U18935 ( .A1(n15415), .A2(n15414), .B1(n15413), .B2(n12333), .C1(
        n15412), .C2(n20888), .ZN(P1_U2897) );
  NAND2_X1 U18936 ( .A1(n20804), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15634) );
  NAND2_X1 U18937 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15417) );
  OAI211_X1 U18938 ( .C1(n20783), .C2(n15418), .A(n15634), .B(n15417), .ZN(
        n15419) );
  AOI21_X1 U18939 ( .B1(n15420), .B2(n20778), .A(n15419), .ZN(n15421) );
  OAI21_X1 U18940 ( .B1(n15640), .B2(n20633), .A(n15421), .ZN(P1_U2970) );
  INV_X1 U18941 ( .A(n15425), .ZN(n15424) );
  NOR4_X1 U18942 ( .A1(n15422), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15423) );
  NAND2_X1 U18943 ( .A1(n15424), .A2(n15423), .ZN(n15426) );
  NAND2_X1 U18944 ( .A1(n20804), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15641) );
  NAND2_X1 U18945 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15427) );
  OAI211_X1 U18946 ( .C1(n20783), .C2(n15428), .A(n15641), .B(n15427), .ZN(
        n15429) );
  AOI21_X1 U18947 ( .B1(n15430), .B2(n20778), .A(n15429), .ZN(n15431) );
  NAND2_X1 U18948 ( .A1(n15433), .A2(n15432), .ZN(n15434) );
  MUX2_X1 U18949 ( .A(n15435), .B(n15434), .S(n15583), .Z(n15436) );
  NAND2_X1 U18950 ( .A1(n20666), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15651) );
  NAND2_X1 U18951 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15438) );
  OAI211_X1 U18952 ( .C1(n20783), .C2(n15439), .A(n15651), .B(n15438), .ZN(
        n15440) );
  NAND2_X1 U18953 ( .A1(n15441), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15451) );
  MUX2_X1 U18954 ( .A(n15689), .B(n15442), .S(n10434), .Z(n15443) );
  XNOR2_X1 U18955 ( .A(n15444), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15681) );
  NAND2_X1 U18956 ( .A1(n20666), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15673) );
  NAND2_X1 U18957 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15445) );
  OAI211_X1 U18958 ( .C1(n20783), .C2(n15446), .A(n15673), .B(n15445), .ZN(
        n15447) );
  AOI21_X1 U18959 ( .B1(n15448), .B2(n20778), .A(n15447), .ZN(n15449) );
  OAI21_X1 U18960 ( .B1(n20633), .B2(n15681), .A(n15449), .ZN(P1_U2974) );
  NAND2_X1 U18961 ( .A1(n15450), .A2(n15451), .ZN(n15452) );
  MUX2_X1 U18962 ( .A(n15452), .B(n15451), .S(n15583), .Z(n15453) );
  XNOR2_X1 U18963 ( .A(n15453), .B(n15689), .ZN(n15692) );
  NAND2_X1 U18964 ( .A1(n20666), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15683) );
  NAND2_X1 U18965 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15454) );
  OAI211_X1 U18966 ( .C1(n20783), .C2(n15455), .A(n15683), .B(n15454), .ZN(
        n15456) );
  AOI21_X1 U18967 ( .B1(n15457), .B2(n20778), .A(n15456), .ZN(n15458) );
  OAI21_X1 U18968 ( .B1(n20633), .B2(n15692), .A(n15458), .ZN(P1_U2975) );
  XNOR2_X1 U18969 ( .A(n9581), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15460) );
  XNOR2_X1 U18970 ( .A(n15459), .B(n15460), .ZN(n15700) );
  INV_X1 U18971 ( .A(n15461), .ZN(n15465) );
  NAND2_X1 U18972 ( .A1(n20804), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15694) );
  NAND2_X1 U18973 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15462) );
  OAI211_X1 U18974 ( .C1(n20783), .C2(n15463), .A(n15694), .B(n15462), .ZN(
        n15464) );
  AOI21_X1 U18975 ( .B1(n15465), .B2(n20778), .A(n15464), .ZN(n15466) );
  OAI21_X1 U18976 ( .B1(n15700), .B2(n20633), .A(n15466), .ZN(P1_U2976) );
  NAND3_X1 U18977 ( .A1(n15496), .A2(n15711), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15469) );
  AOI21_X1 U18978 ( .B1(n15583), .B2(n15469), .A(n15468), .ZN(n15470) );
  XNOR2_X1 U18979 ( .A(n15470), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15720) );
  NAND2_X1 U18980 ( .A1(n20666), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15715) );
  OAI21_X1 U18981 ( .B1(n15530), .B2(n15471), .A(n15715), .ZN(n15474) );
  NOR2_X1 U18982 ( .A1(n15472), .A2(n20837), .ZN(n15473) );
  AOI211_X1 U18983 ( .C1(n15533), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        n15476) );
  OAI21_X1 U18984 ( .B1(n20633), .B2(n15720), .A(n15476), .ZN(P1_U2977) );
  NAND2_X1 U18985 ( .A1(n15497), .A2(n10092), .ZN(n15478) );
  NOR2_X1 U18986 ( .A1(n15583), .A2(n15478), .ZN(n15479) );
  NAND2_X1 U18987 ( .A1(n15477), .A2(n15479), .ZN(n15487) );
  MUX2_X1 U18988 ( .A(n15488), .B(n15487), .S(n15733), .Z(n15481) );
  XNOR2_X1 U18989 ( .A(n15481), .B(n15480), .ZN(n15729) );
  NAND2_X1 U18990 ( .A1(n20804), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15722) );
  NAND2_X1 U18991 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15482) );
  OAI211_X1 U18992 ( .C1(n20783), .C2(n15483), .A(n15722), .B(n15482), .ZN(
        n15484) );
  AOI21_X1 U18993 ( .B1(n15485), .B2(n20778), .A(n15484), .ZN(n15486) );
  OAI21_X1 U18994 ( .B1(n15729), .B2(n20633), .A(n15486), .ZN(P1_U2978) );
  NAND2_X1 U18995 ( .A1(n15488), .A2(n15487), .ZN(n15489) );
  NAND2_X1 U18996 ( .A1(n20666), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15735) );
  OAI21_X1 U18997 ( .B1(n15530), .B2(n15490), .A(n15735), .ZN(n15493) );
  NOR2_X1 U18998 ( .A1(n15491), .A2(n20837), .ZN(n15492) );
  AOI211_X1 U18999 ( .C1(n15533), .C2(n15494), .A(n15493), .B(n15492), .ZN(
        n15495) );
  OAI21_X1 U19000 ( .B1(n15737), .B2(n20633), .A(n15495), .ZN(P1_U2979) );
  AOI21_X1 U19001 ( .B1(n15595), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15496), .ZN(n15499) );
  XNOR2_X1 U19002 ( .A(n9581), .B(n15497), .ZN(n15498) );
  XNOR2_X1 U19003 ( .A(n15499), .B(n15498), .ZN(n15748) );
  NAND2_X1 U19004 ( .A1(n20666), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15741) );
  NAND2_X1 U19005 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15500) );
  OAI211_X1 U19006 ( .C1(n20783), .C2(n15501), .A(n15741), .B(n15500), .ZN(
        n15502) );
  AOI21_X1 U19007 ( .B1(n15503), .B2(n20778), .A(n15502), .ZN(n15504) );
  OAI21_X1 U19008 ( .B1(n15748), .B2(n20633), .A(n15504), .ZN(P1_U2980) );
  NAND2_X1 U19009 ( .A1(n20666), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15756) );
  OAI21_X1 U19010 ( .B1(n15530), .B2(n15505), .A(n15756), .ZN(n15508) );
  OAI21_X1 U19011 ( .B1(n10430), .B2(n15506), .A(n15467), .ZN(n15763) );
  NOR2_X1 U19012 ( .A1(n15763), .A2(n20633), .ZN(n15507) );
  AOI211_X1 U19013 ( .C1(n15533), .C2(n15509), .A(n15508), .B(n15507), .ZN(
        n15510) );
  OAI21_X1 U19014 ( .B1(n15511), .B2(n20837), .A(n15510), .ZN(P1_U2981) );
  NAND2_X1 U19015 ( .A1(n15527), .A2(n15516), .ZN(n15515) );
  NAND2_X1 U19016 ( .A1(n15583), .A2(n15842), .ZN(n15513) );
  NAND2_X1 U19017 ( .A1(n15594), .A2(n15513), .ZN(n15593) );
  NAND2_X1 U19018 ( .A1(n10434), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15538) );
  XNOR2_X1 U19019 ( .A(n15517), .B(n15764), .ZN(n15772) );
  NAND2_X1 U19020 ( .A1(n20666), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15766) );
  OAI21_X1 U19021 ( .B1(n15530), .B2(n15518), .A(n15766), .ZN(n15521) );
  NOR2_X1 U19022 ( .A1(n15519), .A2(n20837), .ZN(n15520) );
  AOI211_X1 U19023 ( .C1(n15533), .C2(n15522), .A(n15521), .B(n15520), .ZN(
        n15523) );
  OAI21_X1 U19024 ( .B1(n20633), .B2(n15772), .A(n15523), .ZN(P1_U2982) );
  AOI21_X1 U19025 ( .B1(n15525), .B2(n15537), .A(n15524), .ZN(n15528) );
  INV_X1 U19026 ( .A(n15524), .ZN(n15526) );
  OAI22_X1 U19027 ( .A1(n15528), .A2(n15527), .B1(n15526), .B2(n15525), .ZN(
        n15780) );
  NAND2_X1 U19028 ( .A1(n15780), .A2(n20779), .ZN(n15535) );
  NAND2_X1 U19029 ( .A1(n20666), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15775) );
  OAI21_X1 U19030 ( .B1(n15530), .B2(n15529), .A(n15775), .ZN(n15531) );
  AOI21_X1 U19031 ( .B1(n15533), .B2(n15532), .A(n15531), .ZN(n15534) );
  OAI211_X1 U19032 ( .C1(n20837), .C2(n15536), .A(n15535), .B(n15534), .ZN(
        P1_U2983) );
  NAND2_X1 U19033 ( .A1(n15538), .A2(n15537), .ZN(n15542) );
  NAND2_X1 U19034 ( .A1(n15540), .A2(n15539), .ZN(n15541) );
  XOR2_X1 U19035 ( .A(n15542), .B(n15541), .Z(n15790) );
  INV_X1 U19036 ( .A(n15543), .ZN(n15547) );
  NAND2_X1 U19037 ( .A1(n20804), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15783) );
  NAND2_X1 U19038 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15544) );
  OAI211_X1 U19039 ( .C1(n20783), .C2(n15545), .A(n15783), .B(n15544), .ZN(
        n15546) );
  AOI21_X1 U19040 ( .B1(n15547), .B2(n20778), .A(n15546), .ZN(n15548) );
  OAI21_X1 U19041 ( .B1(n15790), .B2(n20633), .A(n15548), .ZN(P1_U2984) );
  INV_X1 U19042 ( .A(n15549), .ZN(n15550) );
  AOI21_X1 U19043 ( .B1(n15552), .B2(n15551), .A(n15550), .ZN(n15554) );
  XNOR2_X1 U19044 ( .A(n15583), .B(n15797), .ZN(n15553) );
  XNOR2_X1 U19045 ( .A(n15554), .B(n15553), .ZN(n15800) );
  NAND2_X1 U19046 ( .A1(n20666), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15793) );
  NAND2_X1 U19047 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15555) );
  OAI211_X1 U19048 ( .C1(n20783), .C2(n15556), .A(n15793), .B(n15555), .ZN(
        n15557) );
  AOI21_X1 U19049 ( .B1(n15558), .B2(n20778), .A(n15557), .ZN(n15559) );
  OAI21_X1 U19050 ( .B1(n15800), .B2(n20633), .A(n15559), .ZN(P1_U2985) );
  INV_X1 U19051 ( .A(n15593), .ZN(n15582) );
  INV_X1 U19052 ( .A(n15560), .ZN(n15561) );
  AOI21_X1 U19053 ( .B1(n15582), .B2(n15562), .A(n15561), .ZN(n15574) );
  AND2_X1 U19054 ( .A1(n15563), .A2(n15564), .ZN(n15573) );
  NAND2_X1 U19055 ( .A1(n15574), .A2(n15573), .ZN(n15572) );
  NAND2_X1 U19056 ( .A1(n15572), .A2(n15564), .ZN(n15566) );
  XNOR2_X1 U19057 ( .A(n15566), .B(n15565), .ZN(n15813) );
  NAND2_X1 U19058 ( .A1(n20804), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15807) );
  NAND2_X1 U19059 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15567) );
  OAI211_X1 U19060 ( .C1(n20783), .C2(n15568), .A(n15807), .B(n15567), .ZN(
        n15569) );
  AOI21_X1 U19061 ( .B1(n15570), .B2(n20778), .A(n15569), .ZN(n15571) );
  OAI21_X1 U19062 ( .B1(n20633), .B2(n15813), .A(n15571), .ZN(P1_U2986) );
  OAI21_X1 U19063 ( .B1(n15574), .B2(n15573), .A(n15572), .ZN(n15575) );
  INV_X1 U19064 ( .A(n15575), .ZN(n15829) );
  INV_X1 U19065 ( .A(n15576), .ZN(n15580) );
  NAND2_X1 U19066 ( .A1(n20666), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15819) );
  NAND2_X1 U19067 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15577) );
  OAI211_X1 U19068 ( .C1(n20783), .C2(n15578), .A(n15819), .B(n15577), .ZN(
        n15579) );
  AOI21_X1 U19069 ( .B1(n15580), .B2(n20778), .A(n15579), .ZN(n15581) );
  OAI21_X1 U19070 ( .B1(n15829), .B2(n20633), .A(n15581), .ZN(P1_U2987) );
  NAND3_X1 U19071 ( .A1(n15582), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15583), .ZN(n15586) );
  INV_X1 U19072 ( .A(n15594), .ZN(n15585) );
  NOR2_X1 U19073 ( .A1(n15583), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15584) );
  NAND2_X1 U19074 ( .A1(n15585), .A2(n15584), .ZN(n15598) );
  NAND2_X1 U19075 ( .A1(n15586), .A2(n15598), .ZN(n15587) );
  XNOR2_X1 U19076 ( .A(n15587), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15839) );
  NAND2_X1 U19077 ( .A1(n20666), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15831) );
  NAND2_X1 U19078 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15588) );
  OAI211_X1 U19079 ( .C1(n20783), .C2(n15589), .A(n15831), .B(n15588), .ZN(
        n15590) );
  AOI21_X1 U19080 ( .B1(n15591), .B2(n20778), .A(n15590), .ZN(n15592) );
  OAI21_X1 U19081 ( .B1(n15839), .B2(n20633), .A(n15592), .ZN(P1_U2988) );
  XNOR2_X1 U19082 ( .A(n15593), .B(n10090), .ZN(n15597) );
  NAND2_X1 U19083 ( .A1(n15594), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15596) );
  MUX2_X1 U19084 ( .A(n15597), .B(n15596), .S(n15595), .Z(n15599) );
  NAND2_X1 U19085 ( .A1(n15599), .A2(n15598), .ZN(n15840) );
  NAND2_X1 U19086 ( .A1(n15840), .A2(n20779), .ZN(n15606) );
  INV_X1 U19087 ( .A(n15600), .ZN(n15602) );
  NAND2_X1 U19088 ( .A1(n20804), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15848) );
  NAND2_X1 U19089 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15601) );
  OAI211_X1 U19090 ( .C1(n20783), .C2(n15602), .A(n15848), .B(n15601), .ZN(
        n15603) );
  AOI21_X1 U19091 ( .B1(n15604), .B2(n20778), .A(n15603), .ZN(n15605) );
  NAND2_X1 U19092 ( .A1(n15606), .A2(n15605), .ZN(P1_U2989) );
  XNOR2_X1 U19093 ( .A(n15583), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15607) );
  INV_X1 U19094 ( .A(n15608), .ZN(n15612) );
  NAND2_X1 U19095 ( .A1(n20666), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15856) );
  NAND2_X1 U19096 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15609) );
  OAI211_X1 U19097 ( .C1(n20783), .C2(n15610), .A(n15856), .B(n15609), .ZN(
        n15611) );
  AOI21_X1 U19098 ( .B1(n15612), .B2(n20778), .A(n15611), .ZN(n15613) );
  OAI21_X1 U19099 ( .B1(n15863), .B2(n20633), .A(n15613), .ZN(P1_U2990) );
  NAND2_X1 U19100 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15614) );
  OAI211_X1 U19101 ( .C1(n20783), .C2(n15616), .A(n15615), .B(n15614), .ZN(
        n15617) );
  AOI21_X1 U19102 ( .B1(n15618), .B2(n20778), .A(n15617), .ZN(n15619) );
  OAI21_X1 U19103 ( .B1(n15620), .B2(n20633), .A(n15619), .ZN(P1_U2991) );
  NOR4_X1 U19104 ( .A1(n15631), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15621), .A4(n15637), .ZN(n15626) );
  AND3_X1 U19105 ( .A1(n15623), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15622), .ZN(n15624) );
  NOR3_X1 U19106 ( .A1(n15626), .A2(n15625), .A3(n15624), .ZN(n15629) );
  NAND2_X1 U19107 ( .A1(n15627), .A2(n20823), .ZN(n15628) );
  OAI211_X1 U19108 ( .C1(n15630), .C2(n15862), .A(n15629), .B(n15628), .ZN(
        P1_U3000) );
  INV_X1 U19109 ( .A(n15631), .ZN(n15638) );
  NAND2_X1 U19110 ( .A1(n15632), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15633) );
  OAI211_X1 U19111 ( .C1(n15635), .C2(n20808), .A(n15634), .B(n15633), .ZN(
        n15636) );
  AOI21_X1 U19112 ( .B1(n15638), .B2(n15637), .A(n15636), .ZN(n15639) );
  OAI21_X1 U19113 ( .B1(n15640), .B2(n15862), .A(n15639), .ZN(P1_U3002) );
  OAI21_X1 U19114 ( .B1(n15653), .B2(n15642), .A(n15641), .ZN(n15643) );
  AOI21_X1 U19115 ( .B1(n15644), .B2(n20823), .A(n15643), .ZN(n15649) );
  INV_X1 U19116 ( .A(n15654), .ZN(n15647) );
  NAND3_X1 U19117 ( .A1(n15647), .A2(n15646), .A3(n15645), .ZN(n15648) );
  OAI211_X1 U19118 ( .C1(n15650), .C2(n15862), .A(n15649), .B(n15648), .ZN(
        P1_U3003) );
  OAI21_X1 U19119 ( .B1(n15653), .B2(n15652), .A(n15651), .ZN(n15656) );
  NOR2_X1 U19120 ( .A1(n15654), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15655) );
  AOI211_X1 U19121 ( .C1(n20823), .C2(n15657), .A(n15656), .B(n15655), .ZN(
        n15658) );
  OAI21_X1 U19122 ( .B1(n15659), .B2(n15862), .A(n15658), .ZN(P1_U3004) );
  INV_X1 U19123 ( .A(n15660), .ZN(n15664) );
  INV_X1 U19124 ( .A(n15698), .ZN(n15662) );
  NOR3_X1 U19125 ( .A1(n15662), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15661), .ZN(n15663) );
  AOI211_X1 U19126 ( .C1(n20823), .C2(n15665), .A(n15664), .B(n15663), .ZN(
        n15671) );
  AND2_X1 U19127 ( .A1(n15667), .A2(n15666), .ZN(n15668) );
  NAND2_X1 U19128 ( .A1(n15698), .A2(n15668), .ZN(n15677) );
  INV_X1 U19129 ( .A(n15677), .ZN(n15669) );
  OAI21_X1 U19130 ( .B1(n15669), .B2(n15675), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15670) );
  OAI211_X1 U19131 ( .C1(n15672), .C2(n15862), .A(n15671), .B(n15670), .ZN(
        P1_U3005) );
  INV_X1 U19132 ( .A(n15673), .ZN(n15674) );
  AOI21_X1 U19133 ( .B1(n15675), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15674), .ZN(n15676) );
  OAI211_X1 U19134 ( .C1(n20808), .C2(n15678), .A(n15677), .B(n15676), .ZN(
        n15679) );
  INV_X1 U19135 ( .A(n15679), .ZN(n15680) );
  OAI21_X1 U19136 ( .B1(n15681), .B2(n15862), .A(n15680), .ZN(P1_U3006) );
  INV_X1 U19137 ( .A(n15682), .ZN(n15688) );
  INV_X1 U19138 ( .A(n15683), .ZN(n15687) );
  INV_X1 U19139 ( .A(n15684), .ZN(n15696) );
  OAI21_X1 U19140 ( .B1(n15823), .B2(n20811), .A(n10076), .ZN(n15685) );
  AOI21_X1 U19141 ( .B1(n15696), .B2(n15685), .A(n15689), .ZN(n15686) );
  AOI211_X1 U19142 ( .C1(n15688), .C2(n20823), .A(n15687), .B(n15686), .ZN(
        n15691) );
  NAND3_X1 U19143 ( .A1(n15698), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15689), .ZN(n15690) );
  OAI211_X1 U19144 ( .C1(n15692), .C2(n15862), .A(n15691), .B(n15690), .ZN(
        P1_U3007) );
  NAND2_X1 U19145 ( .A1(n15693), .A2(n20823), .ZN(n15695) );
  OAI211_X1 U19146 ( .C1(n15696), .C2(n10076), .A(n15695), .B(n15694), .ZN(
        n15697) );
  AOI21_X1 U19147 ( .B1(n15698), .B2(n10076), .A(n15697), .ZN(n15699) );
  OAI21_X1 U19148 ( .B1(n15700), .B2(n15862), .A(n15699), .ZN(P1_U3008) );
  INV_X1 U19149 ( .A(n15701), .ZN(n15718) );
  NAND2_X1 U19150 ( .A1(n20811), .A2(n15749), .ZN(n15705) );
  INV_X1 U19151 ( .A(n15702), .ZN(n15801) );
  OR3_X1 U19152 ( .A1(n15703), .A2(n15883), .A3(n15801), .ZN(n15704) );
  NAND2_X1 U19153 ( .A1(n15705), .A2(n15704), .ZN(n15805) );
  AND2_X1 U19154 ( .A1(n15707), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15706) );
  NAND2_X1 U19155 ( .A1(n15805), .A2(n15706), .ZN(n15731) );
  INV_X1 U19156 ( .A(n15707), .ZN(n15708) );
  OR3_X1 U19157 ( .A1(n15802), .A2(n15709), .A3(n15708), .ZN(n15710) );
  NAND2_X1 U19158 ( .A1(n15731), .A2(n15710), .ZN(n15740) );
  NAND2_X1 U19159 ( .A1(n15740), .A2(n15711), .ZN(n15723) );
  INV_X1 U19160 ( .A(n15723), .ZN(n15713) );
  OAI211_X1 U19161 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15713), .B(n15712), .ZN(
        n15714) );
  OAI211_X1 U19162 ( .C1(n15721), .C2(n15716), .A(n15715), .B(n15714), .ZN(
        n15717) );
  AOI21_X1 U19163 ( .B1(n20823), .B2(n15718), .A(n15717), .ZN(n15719) );
  OAI21_X1 U19164 ( .B1(n15720), .B2(n15862), .A(n15719), .ZN(P1_U3009) );
  INV_X1 U19165 ( .A(n15721), .ZN(n15725) );
  OAI21_X1 U19166 ( .B1(n15723), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15722), .ZN(n15724) );
  AOI21_X1 U19167 ( .B1(n15725), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15724), .ZN(n15728) );
  NAND2_X1 U19168 ( .A1(n15726), .A2(n20823), .ZN(n15727) );
  OAI211_X1 U19169 ( .C1(n15729), .C2(n15862), .A(n15728), .B(n15727), .ZN(
        P1_U3010) );
  INV_X1 U19170 ( .A(n15730), .ZN(n15739) );
  AOI21_X1 U19171 ( .B1(n15731), .B2(n15802), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15732) );
  OAI21_X1 U19172 ( .B1(n15746), .B2(n15732), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15736) );
  NAND3_X1 U19173 ( .A1(n15740), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15733), .ZN(n15734) );
  NAND3_X1 U19174 ( .A1(n15736), .A2(n15735), .A3(n15734), .ZN(n15738) );
  INV_X1 U19175 ( .A(n15740), .ZN(n15742) );
  OAI21_X1 U19176 ( .B1(n15742), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15741), .ZN(n15745) );
  NOR2_X1 U19177 ( .A1(n15743), .A2(n20808), .ZN(n15744) );
  AOI211_X1 U19178 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15746), .A(
        n15745), .B(n15744), .ZN(n15747) );
  OAI21_X1 U19179 ( .B1(n15748), .B2(n15862), .A(n15747), .ZN(P1_U3012) );
  INV_X1 U19180 ( .A(n15749), .ZN(n15750) );
  NAND2_X1 U19181 ( .A1(n20811), .A2(n15750), .ZN(n15751) );
  AND2_X1 U19182 ( .A1(n15752), .A2(n15751), .ZN(n15791) );
  AOI22_X1 U19183 ( .A1(n20826), .A2(n15797), .B1(n20811), .B2(n15803), .ZN(
        n15753) );
  AND2_X1 U19184 ( .A1(n15791), .A2(n15753), .ZN(n15785) );
  OAI21_X1 U19185 ( .B1(n15755), .B2(n15754), .A(n15785), .ZN(n15769) );
  OAI21_X1 U19186 ( .B1(n15757), .B2(n20808), .A(n15756), .ZN(n15761) );
  INV_X1 U19187 ( .A(n15758), .ZN(n15798) );
  NAND2_X1 U19188 ( .A1(n15798), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15773) );
  NOR3_X1 U19189 ( .A1(n15773), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15759), .ZN(n15760) );
  AOI211_X1 U19190 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15769), .A(
        n15761), .B(n15760), .ZN(n15762) );
  OAI21_X1 U19191 ( .B1(n15862), .B2(n15763), .A(n15762), .ZN(P1_U3013) );
  NAND2_X1 U19192 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15765) );
  OAI21_X1 U19193 ( .B1(n15773), .B2(n15765), .A(n15764), .ZN(n15770) );
  OAI21_X1 U19194 ( .B1(n15767), .B2(n20808), .A(n15766), .ZN(n15768) );
  AOI21_X1 U19195 ( .B1(n15770), .B2(n15769), .A(n15768), .ZN(n15771) );
  OAI21_X1 U19196 ( .B1(n15772), .B2(n15862), .A(n15771), .ZN(P1_U3014) );
  INV_X1 U19197 ( .A(n15773), .ZN(n15774) );
  NAND2_X1 U19198 ( .A1(n15774), .A2(n15784), .ZN(n15788) );
  AOI21_X1 U19199 ( .B1(n15788), .B2(n15785), .A(n10088), .ZN(n15779) );
  NAND3_X1 U19200 ( .A1(n15774), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n10088), .ZN(n15776) );
  OAI211_X1 U19201 ( .C1(n20808), .C2(n15777), .A(n15776), .B(n15775), .ZN(
        n15778) );
  AOI211_X1 U19202 ( .C1(n15780), .C2(n20828), .A(n15779), .B(n15778), .ZN(
        n15781) );
  INV_X1 U19203 ( .A(n15781), .ZN(P1_U3015) );
  INV_X1 U19204 ( .A(n15782), .ZN(n15787) );
  OAI21_X1 U19205 ( .B1(n15785), .B2(n15784), .A(n15783), .ZN(n15786) );
  AOI21_X1 U19206 ( .B1(n20823), .B2(n15787), .A(n15786), .ZN(n15789) );
  OAI211_X1 U19207 ( .C1(n15790), .C2(n15862), .A(n15789), .B(n15788), .ZN(
        P1_U3016) );
  INV_X1 U19208 ( .A(n15791), .ZN(n15811) );
  AOI21_X1 U19209 ( .B1(n15803), .B2(n15805), .A(n15811), .ZN(n15792) );
  NOR2_X1 U19210 ( .A1(n15792), .A2(n15797), .ZN(n15796) );
  OAI21_X1 U19211 ( .B1(n15794), .B2(n20808), .A(n15793), .ZN(n15795) );
  AOI211_X1 U19212 ( .C1(n15798), .C2(n15797), .A(n15796), .B(n15795), .ZN(
        n15799) );
  OAI21_X1 U19213 ( .B1(n15800), .B2(n15862), .A(n15799), .ZN(P1_U3017) );
  NOR2_X1 U19214 ( .A1(n15802), .A2(n15801), .ZN(n15804) );
  OAI21_X1 U19215 ( .B1(n15805), .B2(n15804), .A(n15803), .ZN(n15809) );
  NAND2_X1 U19216 ( .A1(n15806), .A2(n20823), .ZN(n15808) );
  NAND3_X1 U19217 ( .A1(n15809), .A2(n15808), .A3(n15807), .ZN(n15810) );
  AOI21_X1 U19218 ( .B1(n15811), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15810), .ZN(n15812) );
  OAI21_X1 U19219 ( .B1(n15813), .B2(n15862), .A(n15812), .ZN(P1_U3018) );
  AOI22_X1 U19220 ( .A1(n15816), .A2(n15815), .B1(n20811), .B2(n15814), .ZN(
        n15818) );
  INV_X1 U19221 ( .A(n15817), .ZN(n20813) );
  NAND2_X1 U19222 ( .A1(n15818), .A2(n20813), .ZN(n15837) );
  OAI21_X1 U19223 ( .B1(n15820), .B2(n20808), .A(n15819), .ZN(n15827) );
  AOI21_X1 U19224 ( .B1(n17535), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15825) );
  AOI21_X1 U19225 ( .B1(n15823), .B2(n15822), .A(n15821), .ZN(n15824) );
  NOR3_X1 U19226 ( .A1(n15825), .A2(n15824), .A3(n15833), .ZN(n15826) );
  AOI211_X1 U19227 ( .C1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15837), .A(
        n15827), .B(n15826), .ZN(n15828) );
  OAI21_X1 U19228 ( .B1(n15829), .B2(n15862), .A(n15828), .ZN(P1_U3019) );
  INV_X1 U19229 ( .A(n15830), .ZN(n15832) );
  OAI21_X1 U19230 ( .B1(n15832), .B2(n20808), .A(n15831), .ZN(n15836) );
  INV_X1 U19231 ( .A(n17535), .ZN(n15834) );
  NOR3_X1 U19232 ( .A1(n15834), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15833), .ZN(n15835) );
  AOI211_X1 U19233 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15837), .A(
        n15836), .B(n15835), .ZN(n15838) );
  OAI21_X1 U19234 ( .B1(n15839), .B2(n15862), .A(n15838), .ZN(P1_U3020) );
  NAND2_X1 U19235 ( .A1(n15840), .A2(n20828), .ZN(n15854) );
  NOR2_X1 U19236 ( .A1(n17534), .A2(n15841), .ZN(n15847) );
  NAND2_X1 U19237 ( .A1(n15847), .A2(n15842), .ZN(n15860) );
  NAND2_X1 U19238 ( .A1(n15844), .A2(n15843), .ZN(n15845) );
  OAI21_X1 U19239 ( .B1(n15846), .B2(n15845), .A(n17528), .ZN(n15855) );
  AOI21_X1 U19240 ( .B1(n15860), .B2(n15855), .A(n10090), .ZN(n15852) );
  NAND3_X1 U19241 ( .A1(n15847), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n10090), .ZN(n15849) );
  OAI211_X1 U19242 ( .C1(n20808), .C2(n15850), .A(n15849), .B(n15848), .ZN(
        n15851) );
  NOR2_X1 U19243 ( .A1(n15852), .A2(n15851), .ZN(n15853) );
  NAND2_X1 U19244 ( .A1(n15854), .A2(n15853), .ZN(P1_U3021) );
  INV_X1 U19245 ( .A(n15855), .ZN(n15859) );
  OAI21_X1 U19246 ( .B1(n20808), .B2(n15857), .A(n15856), .ZN(n15858) );
  AOI21_X1 U19247 ( .B1(n15859), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15858), .ZN(n15861) );
  OAI211_X1 U19248 ( .C1(n15863), .C2(n15862), .A(n15861), .B(n15860), .ZN(
        P1_U3022) );
  NAND2_X1 U19249 ( .A1(n9599), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21378) );
  OAI211_X1 U19250 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n9599), .A(n21378), 
        .B(n21210), .ZN(n15865) );
  OAI21_X1 U19251 ( .B1(n15284), .B2(n15875), .A(n15865), .ZN(n15866) );
  MUX2_X1 U19252 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15866), .S(
        n20834), .Z(P1_U3477) );
  INV_X1 U19253 ( .A(n15867), .ZN(n15871) );
  XNOR2_X1 U19254 ( .A(n15867), .B(n21378), .ZN(n15868) );
  OAI22_X1 U19255 ( .A1(n15868), .A2(n21382), .B1(n14332), .B2(n15875), .ZN(
        n15869) );
  MUX2_X1 U19256 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15869), .S(
        n20834), .Z(P1_U3476) );
  INV_X1 U19257 ( .A(n21119), .ZN(n15876) );
  AOI21_X1 U19258 ( .B1(n21211), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n15870), 
        .ZN(n15872) );
  NOR2_X1 U19259 ( .A1(n21087), .A2(n21378), .ZN(n21091) );
  OAI21_X1 U19260 ( .B1(n15872), .B2(n21091), .A(n21210), .ZN(n15874) );
  OR2_X1 U19261 ( .A1(n9599), .A2(n21050), .ZN(n21149) );
  OR3_X1 U19262 ( .A1(n21379), .A2(n21382), .A3(n21149), .ZN(n21298) );
  OAI211_X1 U19263 ( .C1(n15876), .C2(n15875), .A(n15874), .B(n21298), .ZN(
        n15877) );
  MUX2_X1 U19264 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15877), .S(
        n20834), .Z(P1_U3475) );
  INV_X1 U19265 ( .A(n14341), .ZN(n15878) );
  AOI211_X1 U19266 ( .C1(n21329), .C2(n15882), .A(n15881), .B(n15880), .ZN(
        n15905) );
  NOR2_X1 U19267 ( .A1(n15884), .A2(n15883), .ZN(n15890) );
  INV_X1 U19268 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15885) );
  AOI22_X1 U19269 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20832), .B2(n15885), .ZN(
        n15889) );
  INV_X1 U19270 ( .A(n15889), .ZN(n15886) );
  AOI22_X1 U19271 ( .A1(n15892), .A2(n9759), .B1(n15890), .B2(n15886), .ZN(
        n15887) );
  OAI21_X1 U19272 ( .B1(n15905), .B2(n15898), .A(n15887), .ZN(n15888) );
  MUX2_X1 U19273 ( .A(n15888), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15900), .Z(P1_U3473) );
  AOI22_X1 U19274 ( .A1(n15892), .A2(n15891), .B1(n15890), .B2(n15889), .ZN(
        n15893) );
  OAI21_X1 U19275 ( .B1(n15894), .B2(n15898), .A(n15893), .ZN(n15895) );
  MUX2_X1 U19276 ( .A(n15895), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15900), .Z(P1_U3472) );
  INV_X1 U19277 ( .A(n15896), .ZN(n15897) );
  OAI22_X1 U19278 ( .A1(n15899), .A2(n15898), .B1(n15897), .B2(n15931), .ZN(
        n15901) );
  MUX2_X1 U19279 ( .A(n15901), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15900), .Z(P1_U3469) );
  NOR2_X1 U19280 ( .A1(n15902), .A2(n21294), .ZN(n15903) );
  AND2_X1 U19281 ( .A1(n15904), .A2(n15903), .ZN(n15908) );
  AOI211_X1 U19282 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n15908), .A(
        n15906), .B(n15905), .ZN(n15907) );
  INV_X1 U19283 ( .A(n15907), .ZN(n15910) );
  OR2_X1 U19284 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15908), .ZN(
        n15909) );
  NAND2_X1 U19285 ( .A1(n15910), .A2(n15909), .ZN(n15911) );
  AOI222_X1 U19286 ( .A1(n15912), .A2(n21120), .B1(n15912), .B2(n15911), .C1(
        n21120), .C2(n15911), .ZN(n15913) );
  AOI222_X1 U19287 ( .A1(n15914), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .B1(n15914), .B2(n15913), .C1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .C2(n15913), .ZN(n15922) );
  OAI21_X1 U19288 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15915), .ZN(n15916) );
  NAND4_X1 U19289 ( .A1(n15919), .A2(n15918), .A3(n15917), .A4(n15916), .ZN(
        n15921) );
  AOI211_X1 U19290 ( .C1(n15922), .C2(n20835), .A(n15921), .B(n15920), .ZN(
        n15941) );
  INV_X1 U19291 ( .A(n15923), .ZN(n15924) );
  NOR3_X1 U19292 ( .A1(n15926), .A2(n15925), .A3(n15924), .ZN(n15930) );
  INV_X1 U19293 ( .A(n15944), .ZN(n15928) );
  AOI21_X1 U19294 ( .B1(n15928), .B2(n21447), .A(n15927), .ZN(n15929) );
  NOR2_X1 U19295 ( .A1(n15930), .A2(n15929), .ZN(n17553) );
  OAI221_X1 U19296 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15941), 
        .A(n17553), .ZN(n17561) );
  INV_X1 U19297 ( .A(n21526), .ZN(n17556) );
  NOR2_X1 U19298 ( .A1(n17556), .A2(n15931), .ZN(n15932) );
  NOR2_X1 U19299 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15932), .ZN(n15938) );
  INV_X1 U19300 ( .A(n15933), .ZN(n15934) );
  AOI211_X1 U19301 ( .C1(n21447), .C2(n21373), .A(n15935), .B(n15934), .ZN(
        n15936) );
  NAND2_X1 U19302 ( .A1(n17561), .A2(n15936), .ZN(n15937) );
  AOI22_X1 U19303 ( .A1(n17561), .A2(n15938), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15937), .ZN(n15939) );
  OAI21_X1 U19304 ( .B1(n15941), .B2(n15940), .A(n15939), .ZN(P1_U3161) );
  NOR2_X1 U19305 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21447), .ZN(n15942) );
  MUX2_X1 U19306 ( .A(P1_STATEBS16_REG_SCAN_IN), .B(n15942), .S(
        P1_STATE2_REG_0__SCAN_IN), .Z(n15943) );
  NAND2_X1 U19307 ( .A1(n15943), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n17554) );
  NAND3_X1 U19308 ( .A1(n17554), .A2(n15945), .A3(n15944), .ZN(P1_U3163) );
  INV_X1 U19309 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n15946) );
  OAI22_X1 U19310 ( .A1(n20541), .A2(n16351), .B1(n16350), .B2(n15946), .ZN(
        n15948) );
  INV_X1 U19311 ( .A(n16567), .ZN(n15947) );
  AOI21_X1 U19312 ( .B1(n15949), .B2(n16292), .A(n16358), .ZN(n15952) );
  OAI21_X1 U19313 ( .B1(n15952), .B2(n16567), .A(n15951), .ZN(n15953) );
  INV_X1 U19314 ( .A(n15953), .ZN(n15954) );
  NAND2_X1 U19315 ( .A1(n15955), .A2(n16342), .ZN(n15956) );
  INV_X1 U19316 ( .A(n11233), .ZN(n15957) );
  OAI21_X1 U19317 ( .B1(n15976), .B2(n15958), .A(n15957), .ZN(n16872) );
  XOR2_X1 U19318 ( .A(n16583), .B(n15959), .Z(n15965) );
  AOI22_X1 U19319 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n16288), .B1(n16337), 
        .B2(P2_EBX_REG_28__SCAN_IN), .ZN(n15960) );
  OAI21_X1 U19320 ( .B1(n15961), .B2(n16340), .A(n15960), .ZN(n15964) );
  NOR2_X1 U19321 ( .A1(n15962), .A2(n16335), .ZN(n15963) );
  AOI211_X1 U19322 ( .C1(n16292), .C2(n15965), .A(n15964), .B(n15963), .ZN(
        n15970) );
  AOI21_X1 U19323 ( .B1(n15968), .B2(n15971), .A(n15967), .ZN(n16869) );
  NAND2_X1 U19324 ( .A1(n16869), .A2(n16342), .ZN(n15969) );
  OAI211_X1 U19325 ( .C1(n16872), .C2(n16304), .A(n15970), .B(n15969), .ZN(
        P2_U2827) );
  OAI21_X1 U19326 ( .B1(n15973), .B2(n15972), .A(n15971), .ZN(n16877) );
  AND2_X1 U19327 ( .A1(n15975), .A2(n15974), .ZN(n15977) );
  OR2_X1 U19328 ( .A1(n15977), .A2(n15976), .ZN(n16882) );
  INV_X1 U19329 ( .A(n16882), .ZN(n15990) );
  NOR2_X1 U19330 ( .A1(n15978), .A2(n16335), .ZN(n15989) );
  AOI21_X1 U19331 ( .B1(n15983), .B2(n16292), .A(n16358), .ZN(n15987) );
  NOR2_X1 U19332 ( .A1(n16340), .A2(n15979), .ZN(n15982) );
  INV_X1 U19333 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15980) );
  OAI22_X1 U19334 ( .A1(n20538), .A2(n16351), .B1(n16350), .B2(n15980), .ZN(
        n15981) );
  NOR2_X1 U19335 ( .A1(n15982), .A2(n15981), .ZN(n15986) );
  INV_X1 U19336 ( .A(n15983), .ZN(n15984) );
  NAND3_X1 U19337 ( .A1(n15984), .A2(n16305), .A3(n16589), .ZN(n15985) );
  OAI211_X1 U19338 ( .C1(n15987), .C2(n16589), .A(n15986), .B(n15985), .ZN(
        n15988) );
  AOI211_X1 U19339 ( .C1(n15990), .C2(n16365), .A(n15989), .B(n15988), .ZN(
        n15991) );
  OAI21_X1 U19340 ( .B1(n16877), .B2(n16353), .A(n15991), .ZN(P2_U2828) );
  XNOR2_X1 U19341 ( .A(n15992), .B(n15993), .ZN(n15996) );
  AOI22_X1 U19342 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n16288), .B1(n16337), 
        .B2(P2_EBX_REG_26__SCAN_IN), .ZN(n15995) );
  NAND2_X1 U19343 ( .A1(n16359), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15994) );
  OAI211_X1 U19344 ( .C1(n15996), .C2(n16345), .A(n15995), .B(n15994), .ZN(
        n15997) );
  AOI21_X1 U19345 ( .B1(n15998), .B2(n16357), .A(n15997), .ZN(n16000) );
  NAND2_X1 U19346 ( .A1(n16469), .A2(n16342), .ZN(n15999) );
  OAI211_X1 U19347 ( .C1(n16394), .C2(n16304), .A(n16000), .B(n15999), .ZN(
        P2_U2829) );
  NAND2_X1 U19348 ( .A1(n16001), .A2(n16002), .ZN(n16003) );
  NAND2_X1 U19349 ( .A1(n11142), .A2(n16003), .ZN(n16894) );
  OAI21_X1 U19350 ( .B1(n16004), .B2(n16345), .A(n16339), .ZN(n16012) );
  INV_X1 U19351 ( .A(n16602), .ZN(n16005) );
  NAND3_X1 U19352 ( .A1(n16004), .A2(n16305), .A3(n16005), .ZN(n16007) );
  AOI22_X1 U19353 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n16288), .B1(n16337), 
        .B2(P2_EBX_REG_25__SCAN_IN), .ZN(n16006) );
  OAI211_X1 U19354 ( .C1(n16340), .C2(n16600), .A(n16007), .B(n16006), .ZN(
        n16011) );
  XNOR2_X1 U19355 ( .A(n16008), .B(P2_EBX_REG_25__SCAN_IN), .ZN(n16009) );
  NOR2_X1 U19356 ( .A1(n16009), .A2(n16335), .ZN(n16010) );
  AOI211_X1 U19357 ( .C1(n16602), .C2(n16012), .A(n16011), .B(n16010), .ZN(
        n16017) );
  AND2_X1 U19358 ( .A1(n16022), .A2(n16013), .ZN(n16014) );
  NOR2_X1 U19359 ( .A1(n16015), .A2(n16014), .ZN(n16891) );
  NAND2_X1 U19360 ( .A1(n16891), .A2(n16342), .ZN(n16016) );
  OAI211_X1 U19361 ( .C1(n16894), .C2(n16304), .A(n16017), .B(n16016), .ZN(
        P2_U2830) );
  OR2_X1 U19362 ( .A1(n16018), .A2(n16019), .ZN(n16020) );
  NAND2_X1 U19363 ( .A1(n16001), .A2(n16020), .ZN(n16903) );
  INV_X1 U19364 ( .A(n16022), .ZN(n16023) );
  AOI21_X1 U19365 ( .B1(n16024), .B2(n16021), .A(n16023), .ZN(n16906) );
  NAND2_X1 U19366 ( .A1(n16906), .A2(n16342), .ZN(n16034) );
  XOR2_X1 U19367 ( .A(n16621), .B(n16025), .Z(n16032) );
  INV_X1 U19368 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16027) );
  AOI22_X1 U19369 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n16288), .B1(n16337), 
        .B2(P2_EBX_REG_24__SCAN_IN), .ZN(n16026) );
  OAI21_X1 U19370 ( .B1(n16027), .B2(n16340), .A(n16026), .ZN(n16031) );
  AOI211_X1 U19371 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n16029), .A(n16335), .B(
        n16028), .ZN(n16030) );
  AOI211_X1 U19372 ( .C1(n16292), .C2(n16032), .A(n16031), .B(n16030), .ZN(
        n16033) );
  OAI211_X1 U19373 ( .C1(n16304), .C2(n16903), .A(n16034), .B(n16033), .ZN(
        P2_U2831) );
  AND2_X1 U19374 ( .A1(n16035), .A2(n16036), .ZN(n16037) );
  NOR2_X1 U19375 ( .A1(n16018), .A2(n16037), .ZN(n16913) );
  INV_X1 U19376 ( .A(n16913), .ZN(n16050) );
  AOI21_X1 U19377 ( .B1(n9663), .B2(n16292), .A(n16358), .ZN(n16043) );
  OAI22_X1 U19378 ( .A1(n20531), .A2(n16351), .B1(n16350), .B2(n16038), .ZN(
        n16041) );
  INV_X1 U19379 ( .A(n16626), .ZN(n16039) );
  NOR3_X1 U19380 ( .A1(n9663), .A2(n16039), .A3(n16362), .ZN(n16040) );
  AOI211_X1 U19381 ( .C1(n16359), .C2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16041), .B(n16040), .ZN(n16042) );
  OAI21_X1 U19382 ( .B1(n16043), .B2(n16626), .A(n16042), .ZN(n16044) );
  AOI21_X1 U19383 ( .B1(n16045), .B2(n16357), .A(n16044), .ZN(n16049) );
  OR2_X1 U19384 ( .A1(n9655), .A2(n16046), .ZN(n16047) );
  AND2_X1 U19385 ( .A1(n16047), .A2(n16021), .ZN(n16921) );
  NAND2_X1 U19386 ( .A1(n16921), .A2(n16342), .ZN(n16048) );
  OAI211_X1 U19387 ( .C1(n16050), .C2(n16304), .A(n16049), .B(n16048), .ZN(
        P2_U2832) );
  INV_X1 U19388 ( .A(n16035), .ZN(n16051) );
  AOI21_X1 U19389 ( .B1(n16053), .B2(n16052), .A(n16051), .ZN(n16923) );
  INV_X1 U19390 ( .A(n16923), .ZN(n16422) );
  XOR2_X1 U19391 ( .A(n16635), .B(n16054), .Z(n16060) );
  INV_X1 U19392 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16056) );
  AOI22_X1 U19393 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n16288), .B1(n16337), 
        .B2(P2_EBX_REG_22__SCAN_IN), .ZN(n16055) );
  OAI21_X1 U19394 ( .B1(n16056), .B2(n16340), .A(n16055), .ZN(n16059) );
  NOR2_X1 U19395 ( .A1(n16057), .A2(n16335), .ZN(n16058) );
  AOI211_X1 U19396 ( .C1(n16292), .C2(n16060), .A(n16059), .B(n16058), .ZN(
        n16064) );
  AOI21_X1 U19397 ( .B1(n16062), .B2(n16061), .A(n9655), .ZN(n16931) );
  NAND2_X1 U19398 ( .A1(n16931), .A2(n16342), .ZN(n16063) );
  OAI211_X1 U19399 ( .C1(n16422), .C2(n16304), .A(n16064), .B(n16063), .ZN(
        P2_U2833) );
  NAND2_X1 U19400 ( .A1(n16507), .A2(n16342), .ZN(n16074) );
  NAND2_X1 U19401 ( .A1(n16065), .A2(n16249), .ZN(n16076) );
  XNOR2_X1 U19402 ( .A(n16076), .B(n16066), .ZN(n16072) );
  INV_X1 U19403 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16068) );
  AOI22_X1 U19404 ( .A1(P2_REIP_REG_21__SCAN_IN), .A2(n16288), .B1(n16337), 
        .B2(P2_EBX_REG_21__SCAN_IN), .ZN(n16067) );
  OAI21_X1 U19405 ( .B1(n16068), .B2(n16340), .A(n16067), .ZN(n16071) );
  NOR2_X1 U19406 ( .A1(n16069), .A2(n16335), .ZN(n16070) );
  AOI211_X1 U19407 ( .C1(n16292), .C2(n16072), .A(n16071), .B(n16070), .ZN(
        n16073) );
  OAI211_X1 U19408 ( .C1(n16304), .C2(n16427), .A(n16074), .B(n16073), .ZN(
        P2_U2834) );
  INV_X1 U19409 ( .A(n16639), .ZN(n16078) );
  INV_X1 U19410 ( .A(n16075), .ZN(n16077) );
  AOI211_X1 U19411 ( .C1(n16078), .C2(n16077), .A(n16345), .B(n16076), .ZN(
        n16082) );
  AOI22_X1 U19412 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n16288), .B1(n16337), 
        .B2(P2_EBX_REG_20__SCAN_IN), .ZN(n16080) );
  NAND2_X1 U19413 ( .A1(n16359), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16079) );
  OAI211_X1 U19414 ( .C1(n16339), .C2(n16639), .A(n16080), .B(n16079), .ZN(
        n16081) );
  AOI211_X1 U19415 ( .C1(n16083), .C2(n16357), .A(n16082), .B(n16081), .ZN(
        n16085) );
  NAND2_X1 U19416 ( .A1(n16515), .A2(n16342), .ZN(n16084) );
  OAI211_X1 U19417 ( .C1(n16643), .C2(n16304), .A(n16085), .B(n16084), .ZN(
        P2_U2835) );
  AND2_X1 U19418 ( .A1(n16103), .A2(n16102), .ZN(n16105) );
  OAI21_X1 U19419 ( .B1(n16105), .B2(n16087), .A(n16086), .ZN(n16943) );
  AOI21_X1 U19420 ( .B1(n16090), .B2(n16089), .A(n16088), .ZN(n16941) );
  NOR2_X1 U19421 ( .A1(n16091), .A2(n13243), .ZN(n16092) );
  XOR2_X1 U19422 ( .A(n16658), .B(n16092), .Z(n16099) );
  NAND2_X1 U19423 ( .A1(n16093), .A2(n16357), .ZN(n16098) );
  AOI21_X1 U19424 ( .B1(n16288), .B2(P2_REIP_REG_19__SCAN_IN), .A(n16837), 
        .ZN(n16094) );
  OAI21_X1 U19425 ( .B1(n16095), .B2(n16350), .A(n16094), .ZN(n16096) );
  AOI21_X1 U19426 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16359), .A(
        n16096), .ZN(n16097) );
  OAI211_X1 U19427 ( .C1(n16345), .C2(n16099), .A(n16098), .B(n16097), .ZN(
        n16100) );
  AOI21_X1 U19428 ( .B1(n16941), .B2(n16365), .A(n16100), .ZN(n16101) );
  OAI21_X1 U19429 ( .B1(n16943), .B2(n16353), .A(n16101), .ZN(P2_U2836) );
  NOR2_X1 U19430 ( .A1(n16103), .A2(n16102), .ZN(n16104) );
  NAND2_X1 U19431 ( .A1(n16956), .A2(n16365), .ZN(n16116) );
  INV_X1 U19432 ( .A(n16109), .ZN(n16106) );
  AOI21_X1 U19433 ( .B1(n16106), .B2(n16292), .A(n16358), .ZN(n16112) );
  AOI21_X1 U19434 ( .B1(n16337), .B2(P2_EBX_REG_18__SCAN_IN), .A(n16837), .ZN(
        n16107) );
  OAI21_X1 U19435 ( .B1(n20521), .B2(n16351), .A(n16107), .ZN(n16108) );
  AOI21_X1 U19436 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16359), .A(
        n16108), .ZN(n16111) );
  NAND3_X1 U19437 ( .A1(n16109), .A2(n16305), .A3(n16666), .ZN(n16110) );
  OAI211_X1 U19438 ( .C1(n16112), .C2(n16666), .A(n16111), .B(n16110), .ZN(
        n16113) );
  AOI21_X1 U19439 ( .B1(n16114), .B2(n16357), .A(n16113), .ZN(n16115) );
  OAI211_X1 U19440 ( .C1(n16353), .C2(n16948), .A(n16116), .B(n16115), .ZN(
        P2_U2837) );
  OAI21_X1 U19441 ( .B1(n16118), .B2(n16345), .A(n16339), .ZN(n16123) );
  NOR2_X1 U19442 ( .A1(n16351), .A2(n20519), .ZN(n16117) );
  AOI211_X1 U19443 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n16337), .A(n16837), .B(
        n16117), .ZN(n16120) );
  NAND3_X1 U19444 ( .A1(n16118), .A2(n16305), .A3(n16672), .ZN(n16119) );
  OAI211_X1 U19445 ( .C1(n16340), .C2(n16121), .A(n16120), .B(n16119), .ZN(
        n16122) );
  AOI21_X1 U19446 ( .B1(n16124), .B2(n16123), .A(n16122), .ZN(n16125) );
  OAI21_X1 U19447 ( .B1(n16126), .B2(n16335), .A(n16125), .ZN(n16127) );
  AOI21_X1 U19448 ( .B1(n16676), .B2(n16365), .A(n16127), .ZN(n16128) );
  OAI21_X1 U19449 ( .B1(n16533), .B2(n16353), .A(n16128), .ZN(P2_U2838) );
  INV_X1 U19450 ( .A(n16129), .ZN(n16130) );
  AOI21_X1 U19451 ( .B1(n16132), .B2(n16131), .A(n16130), .ZN(n16960) );
  INV_X1 U19452 ( .A(n16960), .ZN(n16145) );
  INV_X1 U19453 ( .A(n16963), .ZN(n16686) );
  NOR2_X1 U19454 ( .A1(n16133), .A2(n16335), .ZN(n16143) );
  AOI21_X1 U19455 ( .B1(n16137), .B2(n16292), .A(n16358), .ZN(n16141) );
  NAND2_X1 U19456 ( .A1(n16288), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16134) );
  OAI211_X1 U19457 ( .C1(n16135), .C2(n16350), .A(n16134), .B(n16810), .ZN(
        n16139) );
  INV_X1 U19458 ( .A(n16683), .ZN(n16136) );
  NOR3_X1 U19459 ( .A1(n16137), .A2(n16136), .A3(n16362), .ZN(n16138) );
  AOI211_X1 U19460 ( .C1(n16359), .C2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16139), .B(n16138), .ZN(n16140) );
  OAI21_X1 U19461 ( .B1(n16141), .B2(n16683), .A(n16140), .ZN(n16142) );
  AOI211_X1 U19462 ( .C1(n16686), .C2(n16365), .A(n16143), .B(n16142), .ZN(
        n16144) );
  OAI21_X1 U19463 ( .B1(n16145), .B2(n16353), .A(n16144), .ZN(P2_U2839) );
  NOR2_X1 U19464 ( .A1(n16146), .A2(n13243), .ZN(n16147) );
  XOR2_X1 U19465 ( .A(n16694), .B(n16147), .Z(n16151) );
  NAND2_X1 U19466 ( .A1(n16337), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n16148) );
  OAI211_X1 U19467 ( .C1(n16692), .C2(n16351), .A(n16148), .B(n16810), .ZN(
        n16149) );
  AOI21_X1 U19468 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n16359), .A(
        n16149), .ZN(n16150) );
  OAI21_X1 U19469 ( .B1(n16151), .B2(n16345), .A(n16150), .ZN(n16152) );
  AOI21_X1 U19470 ( .B1(n16153), .B2(n16357), .A(n16152), .ZN(n16156) );
  XNOR2_X1 U19471 ( .A(n9713), .B(n16154), .ZN(n16979) );
  NAND2_X1 U19472 ( .A1(n16979), .A2(n16342), .ZN(n16155) );
  OAI211_X1 U19473 ( .C1(n16977), .C2(n16304), .A(n16156), .B(n16155), .ZN(
        P2_U2840) );
  OAI21_X1 U19474 ( .B1(n14382), .B2(n16157), .A(n9713), .ZN(n16993) );
  AOI21_X1 U19475 ( .B1(n16161), .B2(n16292), .A(n16358), .ZN(n16160) );
  AOI21_X1 U19476 ( .B1(n16337), .B2(P2_EBX_REG_14__SCAN_IN), .A(n16837), .ZN(
        n16159) );
  NAND2_X1 U19477 ( .A1(n16288), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n16158) );
  OAI211_X1 U19478 ( .C1(n16160), .C2(n16709), .A(n16159), .B(n16158), .ZN(
        n16166) );
  INV_X1 U19479 ( .A(n16161), .ZN(n16162) );
  NAND3_X1 U19480 ( .A1(n16162), .A2(n16305), .A3(n16709), .ZN(n16163) );
  OAI21_X1 U19481 ( .B1(n16340), .B2(n16164), .A(n16163), .ZN(n16165) );
  NOR2_X1 U19482 ( .A1(n16166), .A2(n16165), .ZN(n16167) );
  OAI21_X1 U19483 ( .B1(n16168), .B2(n16335), .A(n16167), .ZN(n16169) );
  AOI21_X1 U19484 ( .B1(n16983), .B2(n16365), .A(n16169), .ZN(n16170) );
  OAI21_X1 U19485 ( .B1(n16993), .B2(n16353), .A(n16170), .ZN(P2_U2841) );
  NOR2_X1 U19486 ( .A1(n17004), .A2(n16304), .ZN(n16183) );
  NOR2_X1 U19487 ( .A1(n16171), .A2(n16335), .ZN(n16182) );
  INV_X1 U19488 ( .A(n16721), .ZN(n16172) );
  NAND3_X1 U19489 ( .A1(n16305), .A2(n16172), .A3(n16174), .ZN(n16173) );
  OAI21_X1 U19490 ( .B1(n16340), .B2(n16719), .A(n16173), .ZN(n16181) );
  NAND2_X1 U19491 ( .A1(n16288), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16179) );
  NOR2_X1 U19492 ( .A1(n16174), .A2(n16345), .ZN(n16175) );
  OAI21_X1 U19493 ( .B1(n16175), .B2(n16358), .A(n16721), .ZN(n16178) );
  INV_X1 U19494 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n16176) );
  OR2_X1 U19495 ( .A1(n16350), .A2(n16176), .ZN(n16177) );
  NAND4_X1 U19496 ( .A1(n16179), .A2(n16810), .A3(n16178), .A4(n16177), .ZN(
        n16180) );
  NOR4_X1 U19497 ( .A1(n16183), .A2(n16182), .A3(n16181), .A4(n16180), .ZN(
        n16184) );
  OAI21_X1 U19498 ( .B1(n16185), .B2(n16353), .A(n16184), .ZN(P2_U2842) );
  INV_X1 U19499 ( .A(n16193), .ZN(n16186) );
  AOI21_X1 U19500 ( .B1(n16292), .B2(n16186), .A(n16358), .ZN(n16196) );
  INV_X1 U19501 ( .A(n16187), .ZN(n16733) );
  INV_X1 U19502 ( .A(n16188), .ZN(n16189) );
  AOI22_X1 U19503 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16359), .B1(
        n16189), .B2(n16357), .ZN(n16190) );
  OAI21_X1 U19504 ( .B1(n16191), .B2(n16350), .A(n16190), .ZN(n16192) );
  AOI211_X1 U19505 ( .C1(n16288), .C2(P2_REIP_REG_12__SCAN_IN), .A(n16837), 
        .B(n16192), .ZN(n16195) );
  NAND3_X1 U19506 ( .A1(n16305), .A2(n16733), .A3(n16193), .ZN(n16194) );
  OAI211_X1 U19507 ( .C1(n16196), .C2(n16733), .A(n16195), .B(n16194), .ZN(
        n16197) );
  AOI21_X1 U19508 ( .B1(n16735), .B2(n16365), .A(n16197), .ZN(n16198) );
  OAI21_X1 U19509 ( .B1(n16353), .B2(n16199), .A(n16198), .ZN(P2_U2843) );
  NAND2_X1 U19510 ( .A1(n16249), .A2(n16200), .ZN(n16201) );
  XOR2_X1 U19511 ( .A(n16749), .B(n16201), .Z(n16207) );
  NAND2_X1 U19512 ( .A1(n16202), .A2(n16357), .ZN(n16206) );
  NOR2_X1 U19513 ( .A1(n16350), .A2(n10964), .ZN(n16204) );
  OAI21_X1 U19514 ( .B1(n16351), .B2(n16746), .A(n16810), .ZN(n16203) );
  AOI211_X1 U19515 ( .C1(n16359), .C2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16204), .B(n16203), .ZN(n16205) );
  OAI211_X1 U19516 ( .C1(n16345), .C2(n16207), .A(n16206), .B(n16205), .ZN(
        n16208) );
  AOI21_X1 U19517 ( .B1(n17027), .B2(n16365), .A(n16208), .ZN(n16209) );
  OAI21_X1 U19518 ( .B1(n16353), .B2(n17036), .A(n16209), .ZN(P2_U2844) );
  INV_X1 U19519 ( .A(n16763), .ZN(n16210) );
  NOR2_X1 U19520 ( .A1(n16216), .A2(n16210), .ZN(n16215) );
  INV_X1 U19521 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20510) );
  OAI22_X1 U19522 ( .A1(n16211), .A2(n16335), .B1(n20510), .B2(n16351), .ZN(
        n16212) );
  INV_X1 U19523 ( .A(n16212), .ZN(n16213) );
  OAI211_X1 U19524 ( .C1(n10962), .C2(n16350), .A(n16213), .B(n16810), .ZN(
        n16214) );
  AOI21_X1 U19525 ( .B1(n16305), .B2(n16215), .A(n16214), .ZN(n16220) );
  NAND2_X1 U19526 ( .A1(n16216), .A2(n16292), .ZN(n16217) );
  AOI21_X1 U19527 ( .B1(n16339), .B2(n16217), .A(n16763), .ZN(n16218) );
  AOI21_X1 U19528 ( .B1(n16359), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16218), .ZN(n16219) );
  OAI211_X1 U19529 ( .C1(n17046), .C2(n16304), .A(n16220), .B(n16219), .ZN(
        n16221) );
  AOI21_X1 U19530 ( .B1(n16342), .B2(n17049), .A(n16221), .ZN(n16222) );
  INV_X1 U19531 ( .A(n16222), .ZN(P2_U2845) );
  AOI21_X1 U19532 ( .B1(n16292), .B2(n16227), .A(n16358), .ZN(n16231) );
  AOI22_X1 U19533 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n16288), .B1(n16357), 
        .B2(n16223), .ZN(n16224) );
  OAI21_X1 U19534 ( .B1(n16225), .B2(n16340), .A(n16224), .ZN(n16226) );
  AOI211_X1 U19535 ( .C1(n16337), .C2(P2_EBX_REG_9__SCAN_IN), .A(n16837), .B(
        n16226), .ZN(n16230) );
  INV_X1 U19536 ( .A(n16227), .ZN(n16228) );
  NAND3_X1 U19537 ( .A1(n16305), .A2(n16777), .A3(n16228), .ZN(n16229) );
  OAI211_X1 U19538 ( .C1(n16231), .C2(n16777), .A(n16230), .B(n16229), .ZN(
        n16232) );
  AOI21_X1 U19539 ( .B1(n16779), .B2(n16365), .A(n16232), .ZN(n16233) );
  OAI21_X1 U19540 ( .B1(n16353), .B2(n16234), .A(n16233), .ZN(P2_U2846) );
  NAND2_X1 U19541 ( .A1(n17072), .A2(n16342), .ZN(n16247) );
  INV_X1 U19542 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16786) );
  OR2_X1 U19543 ( .A1(n16340), .A2(n16786), .ZN(n16243) );
  OAI21_X1 U19544 ( .B1(n16235), .B2(n16350), .A(n16810), .ZN(n16236) );
  AOI21_X1 U19545 ( .B1(n16288), .B2(P2_REIP_REG_8__SCAN_IN), .A(n16236), .ZN(
        n16242) );
  INV_X1 U19546 ( .A(n16789), .ZN(n16237) );
  NAND3_X1 U19547 ( .A1(n16305), .A2(n16237), .A3(n16238), .ZN(n16241) );
  NOR2_X1 U19548 ( .A1(n16238), .A2(n16345), .ZN(n16239) );
  OAI21_X1 U19549 ( .B1(n16358), .B2(n16239), .A(n16789), .ZN(n16240) );
  NAND4_X1 U19550 ( .A1(n16243), .A2(n16242), .A3(n16241), .A4(n16240), .ZN(
        n16244) );
  AOI21_X1 U19551 ( .B1(n16245), .B2(n16357), .A(n16244), .ZN(n16246) );
  OAI211_X1 U19552 ( .C1(n17069), .C2(n16304), .A(n16247), .B(n16246), .ZN(
        P2_U2847) );
  INV_X1 U19553 ( .A(n16815), .ZN(n17084) );
  NAND2_X1 U19554 ( .A1(n16249), .A2(n16248), .ZN(n16250) );
  XOR2_X1 U19555 ( .A(n16813), .B(n16250), .Z(n16255) );
  AOI22_X1 U19556 ( .A1(P2_EBX_REG_7__SCAN_IN), .A2(n16337), .B1(n16251), .B2(
        n16357), .ZN(n16252) );
  OAI211_X1 U19557 ( .C1(n20505), .C2(n16351), .A(n16252), .B(n16810), .ZN(
        n16253) );
  AOI21_X1 U19558 ( .B1(n16359), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16253), .ZN(n16254) );
  OAI21_X1 U19559 ( .B1(n16345), .B2(n16255), .A(n16254), .ZN(n16256) );
  AOI21_X1 U19560 ( .B1(n17084), .B2(n16365), .A(n16256), .ZN(n16257) );
  OAI21_X1 U19561 ( .B1(n16353), .B2(n17086), .A(n16257), .ZN(P2_U2848) );
  NAND2_X1 U19562 ( .A1(n16260), .A2(n16292), .ZN(n16258) );
  AOI21_X1 U19563 ( .B1(n16339), .B2(n16258), .A(n16822), .ZN(n16259) );
  AOI21_X1 U19564 ( .B1(n16359), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16259), .ZN(n16268) );
  INV_X1 U19565 ( .A(n16260), .ZN(n16261) );
  NAND3_X1 U19566 ( .A1(n16305), .A2(n16822), .A3(n16261), .ZN(n16265) );
  OAI21_X1 U19567 ( .B1(n16262), .B2(n16350), .A(n16810), .ZN(n16263) );
  INV_X1 U19568 ( .A(n16263), .ZN(n16264) );
  OAI211_X1 U19569 ( .C1(n16351), .C2(n20503), .A(n16265), .B(n16264), .ZN(
        n16266) );
  INV_X1 U19570 ( .A(n16266), .ZN(n16267) );
  OAI211_X1 U19571 ( .C1(n16269), .C2(n16335), .A(n16268), .B(n16267), .ZN(
        n16270) );
  AOI21_X1 U19572 ( .B1(n17093), .B2(n16365), .A(n16270), .ZN(n16271) );
  OAI21_X1 U19573 ( .B1(n16353), .B2(n16272), .A(n16271), .ZN(P2_U2849) );
  XOR2_X1 U19574 ( .A(n16273), .B(n16274), .Z(n17120) );
  INV_X1 U19575 ( .A(n17120), .ZN(n16566) );
  INV_X1 U19576 ( .A(n17117), .ZN(n16286) );
  OAI21_X1 U19577 ( .B1(n16345), .B2(n16275), .A(n16339), .ZN(n16282) );
  INV_X1 U19578 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16838) );
  INV_X1 U19579 ( .A(n16843), .ZN(n16276) );
  NAND3_X1 U19580 ( .A1(n16305), .A2(n16276), .A3(n16275), .ZN(n16277) );
  OAI21_X1 U19581 ( .B1(n16340), .B2(n16838), .A(n16277), .ZN(n16281) );
  INV_X1 U19582 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n16279) );
  AOI21_X1 U19583 ( .B1(n16337), .B2(P2_EBX_REG_5__SCAN_IN), .A(n16837), .ZN(
        n16278) );
  OAI21_X1 U19584 ( .B1(n16279), .B2(n16351), .A(n16278), .ZN(n16280) );
  AOI211_X1 U19585 ( .C1(n16843), .C2(n16282), .A(n16281), .B(n16280), .ZN(
        n16283) );
  OAI21_X1 U19586 ( .B1(n16284), .B2(n16335), .A(n16283), .ZN(n16285) );
  AOI21_X1 U19587 ( .B1(n16286), .B2(n16365), .A(n16285), .ZN(n16287) );
  OAI21_X1 U19588 ( .B1(n16566), .B2(n16353), .A(n16287), .ZN(P2_U2850) );
  INV_X1 U19589 ( .A(n16860), .ZN(n17128) );
  NAND2_X1 U19590 ( .A1(n16288), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n16289) );
  OAI211_X1 U19591 ( .C1(n16290), .C2(n16350), .A(n16289), .B(n16810), .ZN(
        n16291) );
  AOI21_X1 U19592 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16359), .A(
        n16291), .ZN(n16297) );
  AOI21_X1 U19593 ( .B1(n16292), .B2(n16293), .A(n16358), .ZN(n16295) );
  OR2_X1 U19594 ( .A1(n16362), .A2(n16293), .ZN(n16294) );
  MUX2_X1 U19595 ( .A(n16295), .B(n16294), .S(n16855), .Z(n16296) );
  OAI211_X1 U19596 ( .C1(n16335), .C2(n16850), .A(n16297), .B(n16296), .ZN(
        n16302) );
  NAND2_X1 U19597 ( .A1(n16299), .A2(n16298), .ZN(n16300) );
  NAND2_X1 U19598 ( .A1(n16273), .A2(n16300), .ZN(n17133) );
  NOR2_X1 U19599 ( .A1(n17133), .A2(n16353), .ZN(n16301) );
  AOI211_X1 U19600 ( .C1(n17128), .C2(n16365), .A(n16302), .B(n16301), .ZN(
        n16303) );
  OAI21_X1 U19601 ( .B1(n19779), .B2(n16368), .A(n16303), .ZN(P2_U2851) );
  INV_X1 U19602 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20498) );
  OAI22_X1 U19603 ( .A1(n21574), .A2(n16350), .B1(n20498), .B2(n16351), .ZN(
        n16317) );
  NOR2_X1 U19604 ( .A1(n10648), .A2(n16304), .ZN(n16316) );
  NOR2_X1 U19605 ( .A1(n20565), .A2(n16353), .ZN(n16315) );
  NAND2_X1 U19606 ( .A1(n16305), .A2(n16306), .ZN(n16310) );
  NOR2_X1 U19607 ( .A1(n16306), .A2(n16345), .ZN(n16307) );
  NOR2_X1 U19608 ( .A1(n16358), .A2(n16307), .ZN(n16309) );
  MUX2_X1 U19609 ( .A(n16310), .B(n16309), .S(n16308), .Z(n16312) );
  OR2_X1 U19610 ( .A1(n16340), .A2(n14637), .ZN(n16311) );
  OAI211_X1 U19611 ( .C1(n16335), .C2(n16313), .A(n16312), .B(n16311), .ZN(
        n16314) );
  NOR4_X1 U19612 ( .A1(n16317), .A2(n16316), .A3(n16315), .A4(n16314), .ZN(
        n16318) );
  OAI21_X1 U19613 ( .B1(n20177), .B2(n16368), .A(n16318), .ZN(P2_U2852) );
  INV_X1 U19614 ( .A(n20578), .ZN(n16556) );
  NOR2_X1 U19615 ( .A1(n13243), .A2(n16319), .ZN(n16333) );
  XOR2_X1 U19616 ( .A(n16320), .B(n16333), .Z(n16327) );
  OAI22_X1 U19617 ( .A1(n16321), .A2(n16350), .B1(n20496), .B2(n16351), .ZN(
        n16324) );
  NOR2_X1 U19618 ( .A1(n16335), .A2(n16322), .ZN(n16323) );
  AOI211_X1 U19619 ( .C1(n16359), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16324), .B(n16323), .ZN(n16326) );
  NAND2_X1 U19620 ( .A1(n20576), .A2(n16342), .ZN(n16325) );
  OAI211_X1 U19621 ( .C1(n16327), .C2(n16345), .A(n16326), .B(n16325), .ZN(
        n16328) );
  AOI21_X1 U19622 ( .B1(n13361), .B2(n16365), .A(n16328), .ZN(n16329) );
  OAI21_X1 U19623 ( .B1(n16556), .B2(n16368), .A(n16329), .ZN(P2_U2853) );
  NAND2_X1 U19624 ( .A1(n16331), .A2(n16330), .ZN(n16332) );
  NAND2_X1 U19625 ( .A1(n16333), .A2(n16332), .ZN(n17144) );
  OAI22_X1 U19626 ( .A1(n16335), .A2(n16334), .B1(n20494), .B2(n16351), .ZN(
        n16336) );
  AOI21_X1 U19627 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n16337), .A(n16336), .ZN(
        n16344) );
  OAI22_X1 U19628 ( .A1(n16340), .A2(n16338), .B1(n16339), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16341) );
  AOI21_X1 U19629 ( .B1(n16342), .B2(n20589), .A(n16341), .ZN(n16343) );
  OAI211_X1 U19630 ( .C1(n16345), .C2(n17144), .A(n16344), .B(n16343), .ZN(
        n16346) );
  AOI21_X1 U19631 ( .B1(n16365), .B2(n9574), .A(n16346), .ZN(n16348) );
  OAI21_X1 U19632 ( .B1(n20009), .B2(n16368), .A(n16348), .ZN(P2_U2854) );
  INV_X1 U19633 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19770) );
  OAI22_X1 U19634 ( .A1(n19770), .A2(n16351), .B1(n16350), .B2(n16349), .ZN(
        n16355) );
  NOR2_X1 U19635 ( .A1(n16353), .A2(n16352), .ZN(n16354) );
  AOI211_X1 U19636 ( .C1(n16357), .C2(n16356), .A(n16355), .B(n16354), .ZN(
        n16361) );
  OAI21_X1 U19637 ( .B1(n16359), .B2(n16358), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16360) );
  OAI211_X1 U19638 ( .C1(n16363), .C2(n16362), .A(n16361), .B(n16360), .ZN(
        n16364) );
  AOI21_X1 U19639 ( .B1(n16366), .B2(n16365), .A(n16364), .ZN(n16367) );
  OAI21_X1 U19640 ( .B1(n16368), .B2(n21692), .A(n16367), .ZN(P2_U2855) );
  INV_X1 U19641 ( .A(n16369), .ZN(n16370) );
  MUX2_X1 U19642 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16370), .S(n16430), .Z(
        P2_U2856) );
  XNOR2_X1 U19643 ( .A(n16372), .B(n16371), .ZN(n16448) );
  NOR2_X1 U19644 ( .A1(n16571), .A2(n16438), .ZN(n16373) );
  AOI21_X1 U19645 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n16438), .A(n16373), .ZN(
        n16374) );
  OAI21_X1 U19646 ( .B1(n16433), .B2(n16448), .A(n16374), .ZN(P2_U2858) );
  OAI21_X1 U19647 ( .B1(n16385), .B2(n16383), .A(n16377), .ZN(n16379) );
  XNOR2_X1 U19648 ( .A(n16379), .B(n16378), .ZN(n16455) );
  NOR2_X1 U19649 ( .A1(n16872), .A2(n16438), .ZN(n16380) );
  AOI21_X1 U19650 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16438), .A(n16380), .ZN(
        n16381) );
  OAI21_X1 U19651 ( .B1(n16455), .B2(n16433), .A(n16381), .ZN(P2_U2859) );
  XNOR2_X1 U19652 ( .A(n16383), .B(n16382), .ZN(n16384) );
  XNOR2_X1 U19653 ( .A(n16385), .B(n16384), .ZN(n16463) );
  NOR2_X1 U19654 ( .A1(n16882), .A2(n16438), .ZN(n16386) );
  AOI21_X1 U19655 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16438), .A(n16386), .ZN(
        n16387) );
  OAI21_X1 U19656 ( .B1(n16463), .B2(n16433), .A(n16387), .ZN(P2_U2860) );
  NAND2_X1 U19657 ( .A1(n16397), .A2(n16388), .ZN(n16393) );
  NOR2_X1 U19658 ( .A1(n17491), .A2(n16389), .ZN(n16390) );
  XNOR2_X1 U19659 ( .A(n16391), .B(n16390), .ZN(n16392) );
  XNOR2_X1 U19660 ( .A(n16393), .B(n16392), .ZN(n16471) );
  NOR2_X1 U19661 ( .A1(n16394), .A2(n16438), .ZN(n16395) );
  AOI21_X1 U19662 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16438), .A(n16395), .ZN(
        n16396) );
  OAI21_X1 U19663 ( .B1(n16471), .B2(n16433), .A(n16396), .ZN(P2_U2861) );
  INV_X1 U19664 ( .A(n16397), .ZN(n16398) );
  AOI21_X1 U19665 ( .B1(n16400), .B2(n16399), .A(n16398), .ZN(n16472) );
  NAND2_X1 U19666 ( .A1(n16472), .A2(n16435), .ZN(n16402) );
  NAND2_X1 U19667 ( .A1(n16438), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16401) );
  OAI211_X1 U19668 ( .C1(n16438), .C2(n16894), .A(n16402), .B(n16401), .ZN(
        P2_U2862) );
  AOI21_X1 U19669 ( .B1(n9593), .B2(n16404), .A(n16403), .ZN(n16410) );
  OAI21_X1 U19670 ( .B1(n16406), .B2(n16408), .A(n16413), .ZN(n16409) );
  XOR2_X1 U19671 ( .A(n16410), .B(n16409), .Z(n16486) );
  NOR2_X1 U19672 ( .A1(n16903), .A2(n16438), .ZN(n16411) );
  AOI21_X1 U19673 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16438), .A(n16411), .ZN(
        n16412) );
  OAI21_X1 U19674 ( .B1(n16486), .B2(n16433), .A(n16412), .ZN(P2_U2863) );
  OAI21_X1 U19675 ( .B1(n16415), .B2(n16414), .A(n16413), .ZN(n16494) );
  NAND2_X1 U19676 ( .A1(n16913), .A2(n16430), .ZN(n16417) );
  NAND2_X1 U19677 ( .A1(n16438), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16416) );
  OAI211_X1 U19678 ( .C1(n16494), .C2(n16433), .A(n16417), .B(n16416), .ZN(
        P2_U2864) );
  OR2_X1 U19679 ( .A1(n16418), .A2(n16419), .ZN(n16495) );
  NAND3_X1 U19680 ( .A1(n16406), .A2(n16495), .A3(n16435), .ZN(n16421) );
  NAND2_X1 U19681 ( .A1(n16438), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16420) );
  OAI211_X1 U19682 ( .C1(n16422), .C2(n16438), .A(n16421), .B(n16420), .ZN(
        P2_U2865) );
  AOI21_X1 U19683 ( .B1(n16424), .B2(n16423), .A(n16418), .ZN(n16502) );
  NAND2_X1 U19684 ( .A1(n16502), .A2(n16435), .ZN(n16426) );
  NAND2_X1 U19685 ( .A1(n16438), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16425) );
  OAI211_X1 U19686 ( .C1(n16427), .C2(n16438), .A(n16426), .B(n16425), .ZN(
        P2_U2866) );
  OAI21_X1 U19687 ( .B1(n16428), .B2(n16429), .A(n16423), .ZN(n16517) );
  MUX2_X1 U19688 ( .A(n16431), .B(n16643), .S(n16430), .Z(n16432) );
  OAI21_X1 U19689 ( .B1(n16433), .B2(n16517), .A(n16432), .ZN(P2_U2867) );
  INV_X1 U19690 ( .A(n16941), .ZN(n16439) );
  AOI21_X1 U19691 ( .B1(n16434), .B2(n14686), .A(n16428), .ZN(n16518) );
  NAND2_X1 U19692 ( .A1(n16518), .A2(n16435), .ZN(n16437) );
  NAND2_X1 U19693 ( .A1(n16438), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n16436) );
  OAI211_X1 U19694 ( .C1(n16439), .C2(n16438), .A(n16437), .B(n16436), .ZN(
        P2_U2868) );
  NAND2_X1 U19695 ( .A1(n16440), .A2(n19797), .ZN(n16442) );
  AOI22_X1 U19696 ( .A1(n16541), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19796), .ZN(n16441) );
  OAI211_X1 U19697 ( .C1(n17565), .C2(n16546), .A(n16442), .B(n16441), .ZN(
        P2_U2888) );
  NAND2_X1 U19698 ( .A1(n16541), .A2(BUF2_REG_29__SCAN_IN), .ZN(n16445) );
  AOI22_X1 U19699 ( .A1(n16543), .A2(n16443), .B1(n19796), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16444) );
  OAI211_X1 U19700 ( .C1(n16546), .C2(n17568), .A(n16445), .B(n16444), .ZN(
        n16446) );
  AOI21_X1 U19701 ( .B1(n15955), .B2(n19797), .A(n16446), .ZN(n16447) );
  OAI21_X1 U19702 ( .B1(n16448), .B2(n16562), .A(n16447), .ZN(P2_U2890) );
  INV_X1 U19703 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16452) );
  NAND2_X1 U19704 ( .A1(n16541), .A2(BUF2_REG_28__SCAN_IN), .ZN(n16451) );
  AOI22_X1 U19705 ( .A1(n16543), .A2(n16449), .B1(n19796), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16450) );
  OAI211_X1 U19706 ( .C1(n16546), .C2(n16452), .A(n16451), .B(n16450), .ZN(
        n16453) );
  AOI21_X1 U19707 ( .B1(n16869), .B2(n19797), .A(n16453), .ZN(n16454) );
  OAI21_X1 U19708 ( .B1(n16455), .B2(n16562), .A(n16454), .ZN(P2_U2891) );
  INV_X1 U19709 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16458) );
  AOI22_X1 U19710 ( .A1(n16543), .A2(n16456), .B1(n19796), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16457) );
  OAI21_X1 U19711 ( .B1(n16546), .B2(n16458), .A(n16457), .ZN(n16461) );
  NOR2_X1 U19712 ( .A1(n16877), .A2(n16459), .ZN(n16460) );
  AOI211_X1 U19713 ( .C1(n16541), .C2(BUF2_REG_27__SCAN_IN), .A(n16461), .B(
        n16460), .ZN(n16462) );
  OAI21_X1 U19714 ( .B1(n16463), .B2(n16562), .A(n16462), .ZN(P2_U2892) );
  INV_X1 U19715 ( .A(n16541), .ZN(n16491) );
  INV_X1 U19716 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16467) );
  AOI22_X1 U19717 ( .A1(n16543), .A2(n16464), .B1(n19796), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16466) );
  INV_X1 U19718 ( .A(n16546), .ZN(n16487) );
  NAND2_X1 U19719 ( .A1(n16487), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16465) );
  OAI211_X1 U19720 ( .C1(n16491), .C2(n16467), .A(n16466), .B(n16465), .ZN(
        n16468) );
  AOI21_X1 U19721 ( .B1(n16469), .B2(n19797), .A(n16468), .ZN(n16470) );
  OAI21_X1 U19722 ( .B1(n16471), .B2(n16562), .A(n16470), .ZN(P2_U2893) );
  INV_X1 U19723 ( .A(n16472), .ZN(n16479) );
  INV_X1 U19724 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16476) );
  NAND2_X1 U19725 ( .A1(n16541), .A2(BUF2_REG_25__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19726 ( .A1(n16543), .A2(n16473), .B1(n19796), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16474) );
  OAI211_X1 U19727 ( .C1(n16546), .C2(n16476), .A(n16475), .B(n16474), .ZN(
        n16477) );
  AOI21_X1 U19728 ( .B1(n16891), .B2(n19797), .A(n16477), .ZN(n16478) );
  OAI21_X1 U19729 ( .B1(n16479), .B2(n16562), .A(n16478), .ZN(P2_U2894) );
  INV_X1 U19730 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16483) );
  AOI22_X1 U19731 ( .A1(n16543), .A2(n16480), .B1(n19796), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16482) );
  NAND2_X1 U19732 ( .A1(n16487), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16481) );
  OAI211_X1 U19733 ( .C1(n16491), .C2(n16483), .A(n16482), .B(n16481), .ZN(
        n16484) );
  AOI21_X1 U19734 ( .B1(n16906), .B2(n19797), .A(n16484), .ZN(n16485) );
  OAI21_X1 U19735 ( .B1(n16486), .B2(n16562), .A(n16485), .ZN(P2_U2895) );
  INV_X1 U19736 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16490) );
  AOI22_X1 U19737 ( .A1(n16543), .A2(n19898), .B1(n19796), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16489) );
  NAND2_X1 U19738 ( .A1(n16487), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16488) );
  OAI211_X1 U19739 ( .C1(n16491), .C2(n16490), .A(n16489), .B(n16488), .ZN(
        n16492) );
  AOI21_X1 U19740 ( .B1(n16921), .B2(n19797), .A(n16492), .ZN(n16493) );
  OAI21_X1 U19741 ( .B1(n16494), .B2(n16562), .A(n16493), .ZN(P2_U2896) );
  INV_X1 U19742 ( .A(n16495), .ZN(n16501) );
  INV_X1 U19743 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16498) );
  NAND2_X1 U19744 ( .A1(n16541), .A2(BUF2_REG_22__SCAN_IN), .ZN(n16497) );
  AOI22_X1 U19745 ( .A1(n16543), .A2(n19886), .B1(n19796), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16496) );
  OAI211_X1 U19746 ( .C1(n16498), .C2(n16546), .A(n16497), .B(n16496), .ZN(
        n16499) );
  AOI21_X1 U19747 ( .B1(n16931), .B2(n19797), .A(n16499), .ZN(n16500) );
  OAI21_X1 U19748 ( .B1(n16501), .B2(n16562), .A(n16500), .ZN(P2_U2897) );
  INV_X1 U19749 ( .A(n16502), .ZN(n16509) );
  INV_X1 U19750 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16505) );
  NAND2_X1 U19751 ( .A1(n16541), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16504) );
  AOI22_X1 U19752 ( .A1(n16543), .A2(n19881), .B1(n19796), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16503) );
  OAI211_X1 U19753 ( .C1(n16505), .C2(n16546), .A(n16504), .B(n16503), .ZN(
        n16506) );
  AOI21_X1 U19754 ( .B1(n16507), .B2(n19797), .A(n16506), .ZN(n16508) );
  OAI21_X1 U19755 ( .B1(n16509), .B2(n16562), .A(n16508), .ZN(P2_U2898) );
  INV_X1 U19756 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16513) );
  NAND2_X1 U19757 ( .A1(n16541), .A2(BUF2_REG_20__SCAN_IN), .ZN(n16512) );
  AOI22_X1 U19758 ( .A1(n16543), .A2(n16510), .B1(n19796), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16511) );
  OAI211_X1 U19759 ( .C1(n16513), .C2(n16546), .A(n16512), .B(n16511), .ZN(
        n16514) );
  AOI21_X1 U19760 ( .B1(n16515), .B2(n19797), .A(n16514), .ZN(n16516) );
  OAI21_X1 U19761 ( .B1(n16562), .B2(n16517), .A(n16516), .ZN(P2_U2899) );
  INV_X1 U19762 ( .A(n16518), .ZN(n16525) );
  INV_X1 U19763 ( .A(n16943), .ZN(n16523) );
  NAND2_X1 U19764 ( .A1(n16541), .A2(BUF2_REG_19__SCAN_IN), .ZN(n16521) );
  AOI22_X1 U19765 ( .A1(n16543), .A2(n16519), .B1(n19796), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16520) );
  OAI211_X1 U19766 ( .C1(n19868), .C2(n16546), .A(n16521), .B(n16520), .ZN(
        n16522) );
  AOI21_X1 U19767 ( .B1(n16523), .B2(n19797), .A(n16522), .ZN(n16524) );
  OAI21_X1 U19768 ( .B1(n16525), .B2(n16562), .A(n16524), .ZN(P2_U2900) );
  INV_X1 U19769 ( .A(n16948), .ZN(n16530) );
  INV_X1 U19770 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16528) );
  NAND2_X1 U19771 ( .A1(n16541), .A2(BUF2_REG_18__SCAN_IN), .ZN(n16527) );
  AOI22_X1 U19772 ( .A1(n16543), .A2(n19864), .B1(n19796), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16526) );
  OAI211_X1 U19773 ( .C1(n16528), .C2(n16546), .A(n16527), .B(n16526), .ZN(
        n16529) );
  AOI21_X1 U19774 ( .B1(n16530), .B2(n19797), .A(n16529), .ZN(n16531) );
  OAI21_X1 U19775 ( .B1(n16562), .B2(n16532), .A(n16531), .ZN(P2_U2901) );
  INV_X1 U19776 ( .A(n16533), .ZN(n16537) );
  NAND2_X1 U19777 ( .A1(n16541), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16535) );
  AOI22_X1 U19778 ( .A1(n16543), .A2(n19859), .B1(n19796), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16534) );
  OAI211_X1 U19779 ( .C1(n17580), .C2(n16546), .A(n16535), .B(n16534), .ZN(
        n16536) );
  AOI21_X1 U19780 ( .B1(n16537), .B2(n19797), .A(n16536), .ZN(n16538) );
  OAI21_X1 U19781 ( .B1(n16562), .B2(n16539), .A(n16538), .ZN(P2_U2902) );
  INV_X1 U19782 ( .A(n16540), .ZN(n16550) );
  INV_X1 U19783 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16547) );
  NAND2_X1 U19784 ( .A1(n16541), .A2(BUF2_REG_16__SCAN_IN), .ZN(n16545) );
  AOI22_X1 U19785 ( .A1(n16543), .A2(n16542), .B1(n19796), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n16544) );
  OAI211_X1 U19786 ( .C1(n16547), .C2(n16546), .A(n16545), .B(n16544), .ZN(
        n16548) );
  AOI21_X1 U19787 ( .B1(n16960), .B2(n19797), .A(n16548), .ZN(n16549) );
  OAI21_X1 U19788 ( .B1(n16562), .B2(n16550), .A(n16549), .ZN(P2_U2903) );
  INV_X1 U19789 ( .A(n16979), .ZN(n16552) );
  OAI222_X1 U19790 ( .A1(n19795), .A2(n13835), .B1(n16552), .B2(n16565), .C1(
        n19803), .C2(n16551), .ZN(P2_U2904) );
  AOI22_X1 U19791 ( .A1(n19793), .A2(n16553), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19796), .ZN(n16554) );
  OAI21_X1 U19792 ( .B1(n16993), .B2(n16565), .A(n16554), .ZN(P2_U2905) );
  XNOR2_X1 U19793 ( .A(n20567), .B(n20565), .ZN(n19785) );
  INV_X1 U19794 ( .A(n20576), .ZN(n16555) );
  NAND2_X1 U19795 ( .A1(n16556), .A2(n16555), .ZN(n16560) );
  XOR2_X1 U19796 ( .A(n20576), .B(n20578), .Z(n19791) );
  NAND2_X1 U19797 ( .A1(n20009), .A2(n16557), .ZN(n16559) );
  NAND2_X1 U19798 ( .A1(n16559), .A2(n16558), .ZN(n19790) );
  NAND2_X1 U19799 ( .A1(n19791), .A2(n19790), .ZN(n19789) );
  NAND2_X1 U19800 ( .A1(n16560), .A2(n19789), .ZN(n19784) );
  AOI22_X1 U19801 ( .A1(n19785), .A2(n19784), .B1(n20565), .B2(n20177), .ZN(
        n16561) );
  INV_X1 U19802 ( .A(n17133), .ZN(n19777) );
  NOR2_X1 U19803 ( .A1(n16561), .A2(n19777), .ZN(n19778) );
  OR3_X1 U19804 ( .A1(n19778), .A2(n16562), .A3(n19779), .ZN(n16564) );
  AOI22_X1 U19805 ( .A1(n19793), .A2(n19881), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19796), .ZN(n16563) );
  OAI211_X1 U19806 ( .C1(n16566), .C2(n16565), .A(n16564), .B(n16563), .ZN(
        P2_U2914) );
  NOR2_X1 U19807 ( .A1(n16856), .A2(n16567), .ZN(n16568) );
  AOI211_X1 U19808 ( .C1(n16858), .C2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16569), .B(n16568), .ZN(n16570) );
  OAI21_X1 U19809 ( .B1(n16571), .B2(n19838), .A(n16570), .ZN(n16572) );
  INV_X1 U19810 ( .A(n16577), .ZN(n16576) );
  OAI22_X1 U19811 ( .A1(n16588), .A2(n16864), .B1(n16578), .B2(n16576), .ZN(
        n16581) );
  XNOR2_X1 U19812 ( .A(n16579), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16580) );
  XNOR2_X1 U19813 ( .A(n16581), .B(n16580), .ZN(n16876) );
  NOR2_X1 U19814 ( .A1(n16810), .A2(n20539), .ZN(n16867) );
  AOI21_X1 U19815 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16867), .ZN(n16585) );
  NAND2_X1 U19816 ( .A1(n16842), .A2(n16583), .ZN(n16584) );
  OAI211_X1 U19817 ( .C1(n16872), .C2(n19838), .A(n16585), .B(n16584), .ZN(
        n16586) );
  OAI21_X1 U19818 ( .B1(n16876), .B2(n16863), .A(n16587), .ZN(P2_U2986) );
  XOR2_X1 U19819 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n16588), .Z(
        n16886) );
  NOR2_X1 U19820 ( .A1(n16810), .A2(n20538), .ZN(n16879) );
  NOR2_X1 U19821 ( .A1(n16856), .A2(n16589), .ZN(n16590) );
  AOI211_X1 U19822 ( .C1(n16858), .C2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16879), .B(n16590), .ZN(n16591) );
  OAI21_X1 U19823 ( .B1(n16882), .B2(n19838), .A(n16591), .ZN(n16592) );
  OAI21_X1 U19824 ( .B1(n16886), .B2(n16863), .A(n16593), .ZN(P2_U2987) );
  OAI21_X1 U19825 ( .B1(n16617), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16594), .ZN(n16898) );
  INV_X1 U19826 ( .A(n16595), .ZN(n16596) );
  NOR2_X1 U19827 ( .A1(n16597), .A2(n16596), .ZN(n16598) );
  XNOR2_X1 U19828 ( .A(n16599), .B(n16598), .ZN(n16896) );
  INV_X1 U19829 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20534) );
  NOR2_X1 U19830 ( .A1(n16810), .A2(n20534), .ZN(n16889) );
  NOR2_X1 U19831 ( .A1(n16839), .A2(n16600), .ZN(n16601) );
  AOI211_X1 U19832 ( .C1(n16602), .C2(n16842), .A(n16889), .B(n16601), .ZN(
        n16603) );
  OAI21_X1 U19833 ( .B1(n16894), .B2(n19838), .A(n16603), .ZN(n16604) );
  AOI21_X1 U19834 ( .B1(n16836), .B2(n16896), .A(n16604), .ZN(n16605) );
  OAI21_X1 U19835 ( .B1(n16846), .B2(n16898), .A(n16605), .ZN(P2_U2989) );
  INV_X1 U19836 ( .A(n16631), .ZN(n16609) );
  XNOR2_X1 U19837 ( .A(n16610), .B(n16919), .ZN(n16627) );
  AOI21_X1 U19838 ( .B1(n16611), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16912), .ZN(n16616) );
  INV_X1 U19839 ( .A(n16612), .ZN(n16614) );
  NAND2_X1 U19840 ( .A1(n16614), .A2(n16613), .ZN(n16615) );
  XNOR2_X1 U19841 ( .A(n16616), .B(n16615), .ZN(n16910) );
  INV_X1 U19842 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n16619) );
  OR2_X1 U19843 ( .A1(n16810), .A2(n16619), .ZN(n16900) );
  NAND2_X1 U19844 ( .A1(n16858), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16620) );
  OAI211_X1 U19845 ( .C1(n16856), .C2(n16621), .A(n16900), .B(n16620), .ZN(
        n16622) );
  OAI21_X1 U19846 ( .B1(n16910), .B2(n16863), .A(n16623), .ZN(P2_U2990) );
  NOR2_X1 U19847 ( .A1(n16810), .A2(n20531), .ZN(n16915) );
  AOI21_X1 U19848 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16915), .ZN(n16625) );
  OAI21_X1 U19849 ( .B1(n16856), .B2(n16626), .A(n16625), .ZN(n16628) );
  NAND2_X1 U19850 ( .A1(n16631), .A2(n16630), .ZN(n16633) );
  XOR2_X1 U19851 ( .A(n16633), .B(n16632), .Z(n16935) );
  INV_X1 U19852 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20529) );
  NOR2_X1 U19853 ( .A1(n16810), .A2(n20529), .ZN(n16924) );
  AOI21_X1 U19854 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16924), .ZN(n16634) );
  OAI21_X1 U19855 ( .B1(n16856), .B2(n16635), .A(n16634), .ZN(n16636) );
  AOI21_X1 U19856 ( .B1(n16923), .B2(n16827), .A(n16636), .ZN(n16638) );
  NOR2_X1 U19857 ( .A1(n16639), .A2(n16856), .ZN(n16640) );
  AOI211_X1 U19858 ( .C1(n16858), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16641), .B(n16640), .ZN(n16642) );
  OAI21_X1 U19859 ( .B1(n16643), .B2(n19838), .A(n16642), .ZN(n16644) );
  AOI21_X1 U19860 ( .B1(n16645), .B2(n13307), .A(n16644), .ZN(n16646) );
  OAI21_X1 U19861 ( .B1(n16647), .B2(n16863), .A(n16646), .ZN(P2_U2994) );
  INV_X1 U19862 ( .A(n16648), .ZN(n16649) );
  NAND2_X1 U19863 ( .A1(n16651), .A2(n16650), .ZN(n16652) );
  INV_X1 U19864 ( .A(n16654), .ZN(n16655) );
  NAND2_X1 U19865 ( .A1(n16941), .A2(n16827), .ZN(n16657) );
  NOR2_X1 U19866 ( .A1(n16810), .A2(n20523), .ZN(n16936) );
  AOI21_X1 U19867 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16936), .ZN(n16656) );
  OAI211_X1 U19868 ( .C1(n16856), .C2(n16658), .A(n16657), .B(n16656), .ZN(
        n16659) );
  OAI21_X1 U19869 ( .B1(n16946), .B2(n16863), .A(n16660), .ZN(P2_U2995) );
  OAI21_X1 U19870 ( .B1(n16673), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16661), .ZN(n16959) );
  NAND2_X1 U19871 ( .A1(n16947), .A2(n16836), .ZN(n16669) );
  OR2_X1 U19872 ( .A1(n16810), .A2(n20521), .ZN(n16951) );
  NAND2_X1 U19873 ( .A1(n16858), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16665) );
  OAI211_X1 U19874 ( .C1(n16856), .C2(n16666), .A(n16951), .B(n16665), .ZN(
        n16667) );
  AOI21_X1 U19875 ( .B1(n16956), .B2(n16827), .A(n16667), .ZN(n16668) );
  OAI211_X1 U19876 ( .C1(n16846), .C2(n16959), .A(n16669), .B(n16668), .ZN(
        P2_U2996) );
  AOI21_X1 U19877 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16670), .ZN(n16671) );
  OAI21_X1 U19878 ( .B1(n16856), .B2(n16672), .A(n16671), .ZN(n16675) );
  NAND2_X1 U19879 ( .A1(n16679), .A2(n16688), .ZN(n16680) );
  XOR2_X1 U19880 ( .A(n16681), .B(n16680), .Z(n16964) );
  NAND2_X1 U19881 ( .A1(n16837), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16961) );
  NAND2_X1 U19882 ( .A1(n16858), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16682) );
  OAI211_X1 U19883 ( .C1(n16856), .C2(n16683), .A(n16961), .B(n16682), .ZN(
        n16685) );
  NAND2_X1 U19884 ( .A1(n16688), .A2(n16687), .ZN(n16689) );
  XNOR2_X1 U19885 ( .A(n16690), .B(n16689), .ZN(n16982) );
  NOR2_X1 U19886 ( .A1(n16810), .A2(n16692), .ZN(n16972) );
  AOI21_X1 U19887 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16972), .ZN(n16693) );
  OAI21_X1 U19888 ( .B1(n16856), .B2(n16694), .A(n16693), .ZN(n16695) );
  AOI21_X1 U19889 ( .B1(n16696), .B2(n16827), .A(n16695), .ZN(n16697) );
  OAI211_X1 U19890 ( .C1(n16982), .C2(n16863), .A(n16698), .B(n16697), .ZN(
        P2_U2999) );
  NAND2_X1 U19891 ( .A1(n16701), .A2(n16700), .ZN(n16997) );
  NAND2_X1 U19892 ( .A1(n16703), .A2(n16702), .ZN(n16704) );
  XNOR2_X1 U19893 ( .A(n16705), .B(n16704), .ZN(n16995) );
  NAND2_X1 U19894 ( .A1(n16983), .A2(n16827), .ZN(n16708) );
  NOR2_X1 U19895 ( .A1(n16810), .A2(n16706), .ZN(n16988) );
  AOI21_X1 U19896 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16988), .ZN(n16707) );
  OAI211_X1 U19897 ( .C1(n16856), .C2(n16709), .A(n16708), .B(n16707), .ZN(
        n16710) );
  AOI21_X1 U19898 ( .B1(n16995), .B2(n16836), .A(n16710), .ZN(n16711) );
  OAI21_X1 U19899 ( .B1(n16997), .B2(n16846), .A(n16711), .ZN(P2_U3000) );
  XNOR2_X1 U19900 ( .A(n17012), .B(n17002), .ZN(n17011) );
  NAND2_X1 U19901 ( .A1(n16714), .A2(n16757), .ZN(n16741) );
  INV_X1 U19902 ( .A(n16742), .ZN(n16717) );
  INV_X1 U19903 ( .A(n16715), .ZN(n16716) );
  INV_X1 U19904 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16718) );
  NOR2_X1 U19905 ( .A1(n16810), .A2(n16718), .ZN(n16998) );
  NOR2_X1 U19906 ( .A1(n16839), .A2(n16719), .ZN(n16720) );
  AOI211_X1 U19907 ( .C1(n16721), .C2(n16842), .A(n16998), .B(n16720), .ZN(
        n16722) );
  OAI21_X1 U19908 ( .B1(n17004), .B2(n19838), .A(n16722), .ZN(n16723) );
  OAI21_X1 U19909 ( .B1(n17011), .B2(n16846), .A(n16724), .ZN(P2_U3001) );
  INV_X1 U19910 ( .A(n16725), .ZN(n16727) );
  NAND2_X1 U19911 ( .A1(n16727), .A2(n16726), .ZN(n16729) );
  XOR2_X1 U19912 ( .A(n16729), .B(n16728), .Z(n17023) );
  INV_X1 U19913 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n16731) );
  NOR2_X1 U19914 ( .A1(n16810), .A2(n16731), .ZN(n17015) );
  AOI21_X1 U19915 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17015), .ZN(n16732) );
  OAI21_X1 U19916 ( .B1(n16856), .B2(n16733), .A(n16732), .ZN(n16734) );
  AOI21_X1 U19917 ( .B1(n16735), .B2(n16827), .A(n16734), .ZN(n16736) );
  OAI211_X1 U19918 ( .C1(n17023), .C2(n16863), .A(n16737), .B(n16736), .ZN(
        P2_U3002) );
  INV_X1 U19919 ( .A(n16755), .ZN(n16739) );
  NAND2_X1 U19920 ( .A1(n16741), .A2(n16740), .ZN(n16745) );
  NAND2_X1 U19921 ( .A1(n16743), .A2(n16742), .ZN(n16744) );
  XNOR2_X1 U19922 ( .A(n16745), .B(n16744), .ZN(n17038) );
  NOR2_X1 U19923 ( .A1(n16810), .A2(n16746), .ZN(n17026) );
  NOR2_X1 U19924 ( .A1(n16839), .A2(n16747), .ZN(n16748) );
  AOI211_X1 U19925 ( .C1(n16749), .C2(n16842), .A(n17026), .B(n16748), .ZN(
        n16750) );
  OAI21_X1 U19926 ( .B1(n16751), .B2(n19838), .A(n16750), .ZN(n16752) );
  AOI21_X1 U19927 ( .B1(n17038), .B2(n16836), .A(n16752), .ZN(n16753) );
  OAI21_X1 U19928 ( .B1(n17040), .B2(n16846), .A(n16753), .ZN(P2_U3003) );
  OAI21_X1 U19929 ( .B1(n16754), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16755), .ZN(n17053) );
  NAND2_X1 U19930 ( .A1(n16757), .A2(n16756), .ZN(n16758) );
  XNOR2_X1 U19931 ( .A(n16759), .B(n16758), .ZN(n17050) );
  NAND2_X1 U19932 ( .A1(n16760), .A2(n16827), .ZN(n16762) );
  NOR2_X1 U19933 ( .A1(n16810), .A2(n20510), .ZN(n17041) );
  AOI21_X1 U19934 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17041), .ZN(n16761) );
  OAI211_X1 U19935 ( .C1(n16763), .C2(n16856), .A(n16762), .B(n16761), .ZN(
        n16764) );
  AOI21_X1 U19936 ( .B1(n17050), .B2(n16836), .A(n16764), .ZN(n16765) );
  OAI21_X1 U19937 ( .B1(n17053), .B2(n16846), .A(n16765), .ZN(P2_U3004) );
  NAND2_X1 U19938 ( .A1(n16766), .A2(n16767), .ZN(n16805) );
  INV_X1 U19939 ( .A(n16768), .ZN(n16770) );
  OAI21_X1 U19940 ( .B1(n16805), .B2(n16770), .A(n16769), .ZN(n16774) );
  NAND2_X1 U19941 ( .A1(n16772), .A2(n16771), .ZN(n16773) );
  XNOR2_X1 U19942 ( .A(n16774), .B(n16773), .ZN(n17064) );
  NAND2_X1 U19943 ( .A1(n16837), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n17054) );
  NAND2_X1 U19944 ( .A1(n16858), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16776) );
  OAI211_X1 U19945 ( .C1(n16856), .C2(n16777), .A(n17054), .B(n16776), .ZN(
        n16778) );
  AOI21_X1 U19946 ( .B1(n16779), .B2(n16827), .A(n16778), .ZN(n16780) );
  OAI211_X1 U19947 ( .C1(n16863), .C2(n17064), .A(n16781), .B(n16780), .ZN(
        P2_U3005) );
  NAND2_X1 U19948 ( .A1(n16783), .A2(n16782), .ZN(n16785) );
  NAND2_X1 U19949 ( .A1(n16805), .A2(n16806), .ZN(n16804) );
  NAND2_X1 U19950 ( .A1(n16804), .A2(n16808), .ZN(n16784) );
  XOR2_X1 U19951 ( .A(n16785), .B(n16784), .Z(n17077) );
  NAND2_X1 U19952 ( .A1(n16837), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n17066) );
  OAI21_X1 U19953 ( .B1(n16839), .B2(n16786), .A(n17066), .ZN(n16788) );
  NOR2_X1 U19954 ( .A1(n17069), .A2(n19838), .ZN(n16787) );
  AOI211_X1 U19955 ( .C1(n16789), .C2(n16842), .A(n16788), .B(n16787), .ZN(
        n16801) );
  NAND2_X1 U19956 ( .A1(n16790), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16792) );
  NAND2_X1 U19957 ( .A1(n16795), .A2(n16791), .ZN(n16802) );
  NAND2_X1 U19958 ( .A1(n16792), .A2(n16802), .ZN(n16794) );
  OR2_X1 U19959 ( .A1(n16790), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16793) );
  XNOR2_X1 U19960 ( .A(n16795), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16797) );
  NAND2_X1 U19961 ( .A1(n16796), .A2(n16797), .ZN(n17074) );
  INV_X1 U19962 ( .A(n16796), .ZN(n16799) );
  INV_X1 U19963 ( .A(n16797), .ZN(n16798) );
  NAND2_X1 U19964 ( .A1(n16799), .A2(n16798), .ZN(n17073) );
  NAND3_X1 U19965 ( .A1(n17074), .A2(n13307), .A3(n17073), .ZN(n16800) );
  OAI211_X1 U19966 ( .C1(n17077), .C2(n16863), .A(n16801), .B(n16800), .ZN(
        P2_U3006) );
  XNOR2_X1 U19967 ( .A(n16802), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16803) );
  XNOR2_X1 U19968 ( .A(n16790), .B(n16803), .ZN(n17090) );
  INV_X1 U19969 ( .A(n16804), .ZN(n16809) );
  AOI21_X1 U19970 ( .B1(n16808), .B2(n16806), .A(n16805), .ZN(n16807) );
  AOI21_X1 U19971 ( .B1(n16809), .B2(n16808), .A(n16807), .ZN(n17088) );
  NOR2_X1 U19972 ( .A1(n16810), .A2(n20505), .ZN(n17083) );
  NOR2_X1 U19973 ( .A1(n16839), .A2(n16811), .ZN(n16812) );
  AOI211_X1 U19974 ( .C1(n16813), .C2(n16842), .A(n17083), .B(n16812), .ZN(
        n16814) );
  OAI21_X1 U19975 ( .B1(n16815), .B2(n19838), .A(n16814), .ZN(n16816) );
  AOI21_X1 U19976 ( .B1(n17088), .B2(n16836), .A(n16816), .ZN(n16817) );
  OAI21_X1 U19977 ( .B1(n17090), .B2(n16846), .A(n16817), .ZN(P2_U3007) );
  OAI21_X1 U19978 ( .B1(n16834), .B2(n16835), .A(n16818), .ZN(n16820) );
  XNOR2_X1 U19979 ( .A(n16820), .B(n16819), .ZN(n17108) );
  NOR2_X1 U19980 ( .A1(n16810), .A2(n20503), .ZN(n17092) );
  AOI21_X1 U19981 ( .B1(n16858), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17092), .ZN(n16821) );
  OAI21_X1 U19982 ( .B1(n16856), .B2(n16822), .A(n16821), .ZN(n16826) );
  OAI21_X1 U19983 ( .B1(n16823), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n9569), .ZN(n17091) );
  NOR2_X1 U19984 ( .A1(n17091), .A2(n16846), .ZN(n16825) );
  AOI211_X1 U19985 ( .C1(n16827), .C2(n17093), .A(n16826), .B(n16825), .ZN(
        n16828) );
  OAI21_X1 U19986 ( .B1(n16863), .B2(n17108), .A(n16828), .ZN(P2_U3008) );
  OAI21_X1 U19987 ( .B1(n16832), .B2(n16830), .A(n16829), .ZN(n16831) );
  OAI21_X1 U19988 ( .B1(n16833), .B2(n16832), .A(n16831), .ZN(n17125) );
  XOR2_X1 U19989 ( .A(n16835), .B(n16834), .Z(n17109) );
  NAND2_X1 U19990 ( .A1(n17109), .A2(n16836), .ZN(n16845) );
  NAND2_X1 U19991 ( .A1(n16837), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n17115) );
  OAI21_X1 U19992 ( .B1(n16839), .B2(n16838), .A(n17115), .ZN(n16841) );
  NOR2_X1 U19993 ( .A1(n17117), .A2(n19838), .ZN(n16840) );
  AOI211_X1 U19994 ( .C1(n16843), .C2(n16842), .A(n16841), .B(n16840), .ZN(
        n16844) );
  OAI211_X1 U19995 ( .C1(n16846), .C2(n17125), .A(n16845), .B(n16844), .ZN(
        P2_U3009) );
  AOI22_X1 U19996 ( .A1(n16849), .A2(n16848), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16847), .ZN(n16852) );
  XNOR2_X1 U19997 ( .A(n16850), .B(n16853), .ZN(n16851) );
  XNOR2_X1 U19998 ( .A(n16852), .B(n16851), .ZN(n17140) );
  INV_X1 U19999 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20500) );
  NOR2_X1 U20000 ( .A1(n16810), .A2(n20500), .ZN(n17126) );
  NOR2_X1 U20001 ( .A1(n16856), .A2(n16855), .ZN(n16857) );
  AOI211_X1 U20002 ( .C1(n16858), .C2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n17126), .B(n16857), .ZN(n16859) );
  OAI21_X1 U20003 ( .B1(n16860), .B2(n19838), .A(n16859), .ZN(n16861) );
  AOI21_X1 U20004 ( .B1(n17137), .B2(n13307), .A(n16861), .ZN(n16862) );
  OAI21_X1 U20005 ( .B1(n17140), .B2(n16863), .A(n16862), .ZN(P2_U3010) );
  NOR3_X1 U20006 ( .A1(n16865), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16864), .ZN(n16866) );
  AOI211_X1 U20007 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16868), .A(
        n16867), .B(n16866), .ZN(n16871) );
  NAND2_X1 U20008 ( .A1(n16869), .A2(n17121), .ZN(n16870) );
  OAI211_X1 U20009 ( .C1(n16872), .C2(n17116), .A(n16871), .B(n16870), .ZN(
        n16873) );
  AOI21_X1 U20010 ( .B1(n16874), .B2(n17136), .A(n16873), .ZN(n16875) );
  OAI21_X1 U20011 ( .B1(n16876), .B2(n17139), .A(n16875), .ZN(P2_U3018) );
  NOR2_X1 U20012 ( .A1(n16877), .A2(n17134), .ZN(n16884) );
  AOI211_X1 U20013 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16880), .A(
        n16879), .B(n16878), .ZN(n16881) );
  OAI21_X1 U20014 ( .B1(n16882), .B2(n17116), .A(n16881), .ZN(n16883) );
  OAI21_X1 U20015 ( .B1(n16886), .B2(n17139), .A(n16885), .ZN(P2_U3019) );
  NOR2_X1 U20016 ( .A1(n16887), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16888) );
  AOI211_X1 U20017 ( .C1(n16890), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16889), .B(n16888), .ZN(n16893) );
  NAND2_X1 U20018 ( .A1(n16891), .A2(n17121), .ZN(n16892) );
  OAI211_X1 U20019 ( .C1(n16894), .C2(n17116), .A(n16893), .B(n16892), .ZN(
        n16895) );
  AOI21_X1 U20020 ( .B1(n9563), .B2(n16896), .A(n16895), .ZN(n16897) );
  OAI21_X1 U20021 ( .B1(n17124), .B2(n16898), .A(n16897), .ZN(P2_U3021) );
  INV_X1 U20022 ( .A(n16899), .ZN(n16925) );
  NOR2_X1 U20023 ( .A1(n16919), .A2(n16928), .ZN(n16914) );
  AOI21_X1 U20024 ( .B1(n16925), .B2(n16914), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16902) );
  OAI21_X1 U20025 ( .B1(n16902), .B2(n16901), .A(n16900), .ZN(n16905) );
  NOR2_X1 U20026 ( .A1(n16903), .A2(n17116), .ZN(n16904) );
  AOI211_X1 U20027 ( .C1(n16906), .C2(n17121), .A(n16905), .B(n16904), .ZN(
        n16909) );
  NAND2_X1 U20028 ( .A1(n16907), .A2(n17136), .ZN(n16908) );
  OAI211_X1 U20029 ( .C1(n16910), .C2(n17139), .A(n16909), .B(n16908), .ZN(
        P2_U3022) );
  NAND2_X1 U20030 ( .A1(n16913), .A2(n17127), .ZN(n16918) );
  AOI21_X1 U20031 ( .B1(n16919), .B2(n16928), .A(n16914), .ZN(n16916) );
  AOI21_X1 U20032 ( .B1(n16925), .B2(n16916), .A(n16915), .ZN(n16917) );
  OAI211_X1 U20033 ( .C1(n16929), .C2(n16919), .A(n16918), .B(n16917), .ZN(
        n16920) );
  NAND2_X1 U20034 ( .A1(n16923), .A2(n17127), .ZN(n16927) );
  AOI21_X1 U20035 ( .B1(n16925), .B2(n16928), .A(n16924), .ZN(n16926) );
  OAI211_X1 U20036 ( .C1(n16929), .C2(n16928), .A(n16927), .B(n16926), .ZN(
        n16930) );
  AOI21_X1 U20037 ( .B1(n17121), .B2(n16931), .A(n16930), .ZN(n16934) );
  NAND2_X1 U20038 ( .A1(n16932), .A2(n17136), .ZN(n16933) );
  OAI211_X1 U20039 ( .C1(n16935), .C2(n17139), .A(n16934), .B(n16933), .ZN(
        P2_U3024) );
  INV_X1 U20040 ( .A(n16936), .ZN(n16937) );
  OAI211_X1 U20041 ( .C1(n16953), .C2(n16939), .A(n16938), .B(n16937), .ZN(
        n16940) );
  AOI21_X1 U20042 ( .B1(n16941), .B2(n17127), .A(n16940), .ZN(n16942) );
  OAI21_X1 U20043 ( .B1(n17134), .B2(n16943), .A(n16942), .ZN(n16944) );
  OAI21_X1 U20044 ( .B1(n16946), .B2(n17139), .A(n16945), .ZN(P2_U3027) );
  NAND2_X1 U20045 ( .A1(n16947), .A2(n9563), .ZN(n16958) );
  NOR2_X1 U20046 ( .A1(n16948), .A2(n17134), .ZN(n16955) );
  NAND3_X1 U20047 ( .A1(n17031), .A2(n16949), .A3(n16952), .ZN(n16950) );
  OAI211_X1 U20048 ( .C1(n16953), .C2(n16952), .A(n16951), .B(n16950), .ZN(
        n16954) );
  AOI211_X1 U20049 ( .C1(n16956), .C2(n17127), .A(n16955), .B(n16954), .ZN(
        n16957) );
  OAI211_X1 U20050 ( .C1(n16959), .C2(n17124), .A(n16958), .B(n16957), .ZN(
        P2_U3028) );
  NAND2_X1 U20051 ( .A1(n16960), .A2(n17121), .ZN(n16962) );
  OAI211_X1 U20052 ( .C1(n17116), .C2(n16963), .A(n16962), .B(n16961), .ZN(
        n16966) );
  NOR2_X1 U20053 ( .A1(n16964), .A2(n17139), .ZN(n16965) );
  OAI21_X1 U20054 ( .B1(n16970), .B2(n16969), .A(n16968), .ZN(P2_U3030) );
  NAND2_X1 U20055 ( .A1(n16971), .A2(n17136), .ZN(n16981) );
  AOI21_X1 U20056 ( .B1(n16973), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16972), .ZN(n16976) );
  NAND3_X1 U20057 ( .A1(n16990), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16974), .ZN(n16975) );
  OAI211_X1 U20058 ( .C1(n16977), .C2(n17116), .A(n16976), .B(n16975), .ZN(
        n16978) );
  AOI21_X1 U20059 ( .B1(n17121), .B2(n16979), .A(n16978), .ZN(n16980) );
  OAI211_X1 U20060 ( .C1(n16982), .C2(n17139), .A(n16981), .B(n16980), .ZN(
        P2_U3031) );
  NAND2_X1 U20061 ( .A1(n16983), .A2(n17127), .ZN(n16992) );
  NOR2_X1 U20062 ( .A1(n16985), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17014) );
  OAI21_X1 U20063 ( .B1(n17098), .B2(n16984), .A(n17057), .ZN(n17016) );
  NOR2_X1 U20064 ( .A1(n17014), .A2(n17016), .ZN(n17003) );
  INV_X1 U20065 ( .A(n16985), .ZN(n16999) );
  NAND2_X1 U20066 ( .A1(n16999), .A2(n17002), .ZN(n16986) );
  AOI21_X1 U20067 ( .B1(n17003), .B2(n16986), .A(n16989), .ZN(n16987) );
  AOI211_X1 U20068 ( .C1(n16990), .C2(n16989), .A(n16988), .B(n16987), .ZN(
        n16991) );
  OAI211_X1 U20069 ( .C1(n16993), .C2(n17134), .A(n16992), .B(n16991), .ZN(
        n16994) );
  AOI21_X1 U20070 ( .B1(n16995), .B2(n9563), .A(n16994), .ZN(n16996) );
  OAI21_X1 U20071 ( .B1(n16997), .B2(n17124), .A(n16996), .ZN(P2_U3032) );
  INV_X1 U20072 ( .A(n16998), .ZN(n17001) );
  NAND3_X1 U20073 ( .A1(n16999), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n17002), .ZN(n17000) );
  OAI211_X1 U20074 ( .C1(n17003), .C2(n17002), .A(n17001), .B(n17000), .ZN(
        n17006) );
  NOR2_X1 U20075 ( .A1(n17004), .A2(n17116), .ZN(n17005) );
  AOI211_X1 U20076 ( .C1(n17007), .C2(n17121), .A(n17006), .B(n17005), .ZN(
        n17010) );
  NAND2_X1 U20077 ( .A1(n17008), .A2(n9563), .ZN(n17009) );
  OAI211_X1 U20078 ( .C1(n17011), .C2(n17124), .A(n17010), .B(n17009), .ZN(
        P2_U3033) );
  NAND3_X1 U20079 ( .A1(n17013), .A2(n17136), .A3(n17012), .ZN(n17022) );
  AOI211_X1 U20080 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17016), .A(
        n17015), .B(n17014), .ZN(n17017) );
  OAI21_X1 U20081 ( .B1(n17018), .B2(n17116), .A(n17017), .ZN(n17019) );
  AOI21_X1 U20082 ( .B1(n17121), .B2(n17020), .A(n17019), .ZN(n17021) );
  OAI211_X1 U20083 ( .C1(n17023), .C2(n17139), .A(n17022), .B(n17021), .ZN(
        P2_U3034) );
  INV_X1 U20084 ( .A(n17031), .ZN(n17055) );
  NOR3_X1 U20085 ( .A1(n17055), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n17024), .ZN(n17025) );
  AOI211_X1 U20086 ( .C1(n17027), .C2(n17127), .A(n17026), .B(n17025), .ZN(
        n17035) );
  NOR2_X1 U20087 ( .A1(n17028), .A2(n17056), .ZN(n17045) );
  AND2_X1 U20088 ( .A1(n17029), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17030) );
  NAND2_X1 U20089 ( .A1(n17031), .A2(n17030), .ZN(n17043) );
  OAI21_X1 U20090 ( .B1(n17045), .B2(n17032), .A(n17043), .ZN(n17033) );
  NAND2_X1 U20091 ( .A1(n17033), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17034) );
  OAI211_X1 U20092 ( .C1(n17036), .C2(n17134), .A(n17035), .B(n17034), .ZN(
        n17037) );
  AOI21_X1 U20093 ( .B1(n17038), .B2(n9563), .A(n17037), .ZN(n17039) );
  OAI21_X1 U20094 ( .B1(n17040), .B2(n17124), .A(n17039), .ZN(P2_U3035) );
  NAND2_X1 U20095 ( .A1(n17097), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17044) );
  INV_X1 U20096 ( .A(n17041), .ZN(n17042) );
  OAI211_X1 U20097 ( .C1(n17045), .C2(n17044), .A(n17043), .B(n17042), .ZN(
        n17048) );
  NOR2_X1 U20098 ( .A1(n17046), .A2(n17116), .ZN(n17047) );
  AOI211_X1 U20099 ( .C1(n17049), .C2(n17121), .A(n17048), .B(n17047), .ZN(
        n17052) );
  NAND2_X1 U20100 ( .A1(n17050), .A2(n9563), .ZN(n17051) );
  OAI211_X1 U20101 ( .C1(n17053), .C2(n17124), .A(n17052), .B(n17051), .ZN(
        P2_U3036) );
  OAI21_X1 U20102 ( .B1(n17055), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17054), .ZN(n17060) );
  OAI22_X1 U20103 ( .A1(n17058), .A2(n17116), .B1(n17057), .B2(n17056), .ZN(
        n17059) );
  AOI211_X1 U20104 ( .C1(n17121), .C2(n17061), .A(n17060), .B(n17059), .ZN(
        n17062) );
  OAI211_X1 U20105 ( .C1(n17064), .C2(n17139), .A(n17063), .B(n17062), .ZN(
        P2_U3037) );
  OAI211_X1 U20106 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n17078), .B(n17065), .ZN(n17067) );
  NAND2_X1 U20107 ( .A1(n17067), .A2(n17066), .ZN(n17071) );
  OAI22_X1 U20108 ( .A1(n17069), .A2(n17116), .B1(n17068), .B2(n17081), .ZN(
        n17070) );
  AOI211_X1 U20109 ( .C1(n17121), .C2(n17072), .A(n17071), .B(n17070), .ZN(
        n17076) );
  NAND3_X1 U20110 ( .A1(n17074), .A2(n17136), .A3(n17073), .ZN(n17075) );
  OAI211_X1 U20111 ( .C1(n17077), .C2(n17139), .A(n17076), .B(n17075), .ZN(
        P2_U3038) );
  NAND2_X1 U20112 ( .A1(n17078), .A2(n17080), .ZN(n17079) );
  OAI21_X1 U20113 ( .B1(n17081), .B2(n17080), .A(n17079), .ZN(n17082) );
  AOI211_X1 U20114 ( .C1(n17084), .C2(n17127), .A(n17083), .B(n17082), .ZN(
        n17085) );
  OAI21_X1 U20115 ( .B1(n17134), .B2(n17086), .A(n17085), .ZN(n17087) );
  AOI21_X1 U20116 ( .B1(n17088), .B2(n9563), .A(n17087), .ZN(n17089) );
  OAI21_X1 U20117 ( .B1(n17090), .B2(n17124), .A(n17089), .ZN(P2_U3039) );
  INV_X1 U20118 ( .A(n17091), .ZN(n17106) );
  AOI21_X1 U20119 ( .B1(n17093), .B2(n17127), .A(n17092), .ZN(n17104) );
  NAND2_X1 U20120 ( .A1(n17094), .A2(n17121), .ZN(n17103) );
  NAND2_X1 U20121 ( .A1(n17095), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17096) );
  NAND2_X1 U20122 ( .A1(n17097), .A2(n17096), .ZN(n17129) );
  OAI21_X1 U20123 ( .B1(n17098), .B2(n17111), .A(n17129), .ZN(n17099) );
  NAND2_X1 U20124 ( .A1(n17099), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17102) );
  INV_X1 U20125 ( .A(n17130), .ZN(n17113) );
  NAND3_X1 U20126 ( .A1(n17113), .A2(n17111), .A3(n17100), .ZN(n17101) );
  NAND4_X1 U20127 ( .A1(n17104), .A2(n17103), .A3(n17102), .A4(n17101), .ZN(
        n17105) );
  AOI21_X1 U20128 ( .B1(n17106), .B2(n17136), .A(n17105), .ZN(n17107) );
  OAI21_X1 U20129 ( .B1(n17139), .B2(n17108), .A(n17107), .ZN(P2_U3040) );
  NAND2_X1 U20130 ( .A1(n17109), .A2(n9563), .ZN(n17123) );
  NOR2_X1 U20131 ( .A1(n17129), .A2(n17110), .ZN(n17119) );
  INV_X1 U20132 ( .A(n17111), .ZN(n17112) );
  OAI211_X1 U20133 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n17113), .B(n17112), .ZN(n17114) );
  OAI211_X1 U20134 ( .C1(n17117), .C2(n17116), .A(n17115), .B(n17114), .ZN(
        n17118) );
  AOI211_X1 U20135 ( .C1(n17121), .C2(n17120), .A(n17119), .B(n17118), .ZN(
        n17122) );
  OAI211_X1 U20136 ( .C1(n17125), .C2(n17124), .A(n17123), .B(n17122), .ZN(
        P2_U3041) );
  AOI21_X1 U20137 ( .B1(n17128), .B2(n17127), .A(n17126), .ZN(n17132) );
  MUX2_X1 U20138 ( .A(n17130), .B(n17129), .S(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n17131) );
  OAI211_X1 U20139 ( .C1(n17134), .C2(n17133), .A(n17132), .B(n17131), .ZN(
        n17135) );
  AOI21_X1 U20140 ( .B1(n17137), .B2(n17136), .A(n17135), .ZN(n17138) );
  OAI21_X1 U20141 ( .B1(n17140), .B2(n17139), .A(n17138), .ZN(P2_U3042) );
  NOR2_X1 U20142 ( .A1(n17142), .A2(n17141), .ZN(n17152) );
  NAND2_X1 U20143 ( .A1(n13243), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17143) );
  NAND2_X1 U20144 ( .A1(n17144), .A2(n17143), .ZN(n17153) );
  INV_X1 U20145 ( .A(n17153), .ZN(n17145) );
  AOI222_X1 U20146 ( .A1(n17146), .A2(n17490), .B1(n17152), .B2(n17145), .C1(
        n20585), .C2(n17151), .ZN(n17148) );
  NAND2_X1 U20147 ( .A1(n17156), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17147) );
  OAI21_X1 U20148 ( .B1(n17148), .B2(n17156), .A(n17147), .ZN(P2_U3600) );
  INV_X1 U20149 ( .A(n17149), .ZN(n17150) );
  AOI222_X1 U20150 ( .A1(n17153), .A2(n17152), .B1(n20578), .B2(n17151), .C1(
        n17150), .C2(n17490), .ZN(n17157) );
  NAND2_X1 U20151 ( .A1(n17156), .A2(n17154), .ZN(n17155) );
  OAI21_X1 U20152 ( .B1(n17157), .B2(n17156), .A(n17155), .ZN(P2_U3599) );
  XNOR2_X1 U20153 ( .A(n18712), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17285) );
  NOR3_X1 U20154 ( .A1(n11722), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17285), .ZN(n17299) );
  AOI22_X1 U20155 ( .A1(n17299), .A2(n18712), .B1(n11724), .B2(n17290), .ZN(
        n17158) );
  XOR2_X1 U20156 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n17158), .Z(
        n17281) );
  INV_X1 U20157 ( .A(n17267), .ZN(n17288) );
  OAI33_X1 U20158 ( .A1(n18811), .A2(n17160), .A3(n17288), .B1(n17287), .B2(
        n17159), .B3(n18810), .ZN(n17170) );
  INV_X1 U20159 ( .A(n17161), .ZN(n17163) );
  INV_X1 U20160 ( .A(n17682), .ZN(n17162) );
  AOI21_X1 U20161 ( .B1(n18749), .B2(n17163), .A(n17162), .ZN(n17169) );
  NAND2_X1 U20162 ( .A1(n17164), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17165) );
  NAND2_X1 U20163 ( .A1(n19089), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17270) );
  OAI211_X1 U20164 ( .C1(n17167), .C2(n17166), .A(n17165), .B(n17270), .ZN(
        n17168) );
  AOI211_X1 U20165 ( .C1(n17170), .C2(n17290), .A(n17169), .B(n17168), .ZN(
        n17173) );
  NAND2_X1 U20166 ( .A1(n17171), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17172) );
  OAI211_X1 U20167 ( .C1(n17281), .C2(n18829), .A(n17173), .B(n17172), .ZN(
        P3_U2801) );
  XNOR2_X1 U20168 ( .A(n17286), .B(n17285), .ZN(n17187) );
  OAI21_X1 U20169 ( .B1(n14730), .B2(n18799), .A(n18906), .ZN(n17174) );
  AOI21_X1 U20170 ( .B1(n18801), .B2(n17175), .A(n17174), .ZN(n17205) );
  OAI21_X1 U20171 ( .B1(n18725), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17205), .ZN(n17198) );
  NAND3_X1 U20172 ( .A1(n17176), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17300), .ZN(n17296) );
  INV_X1 U20173 ( .A(n17296), .ZN(n17181) );
  INV_X1 U20174 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19703) );
  NOR2_X1 U20175 ( .A1(n19120), .A2(n19703), .ZN(n17298) );
  INV_X1 U20176 ( .A(n14730), .ZN(n17179) );
  OAI211_X1 U20177 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n18818), .B(n17177), .ZN(n17178) );
  NOR2_X1 U20178 ( .A1(n17179), .A2(n17178), .ZN(n17180) );
  AOI211_X1 U20179 ( .C1(n18780), .C2(n17181), .A(n17298), .B(n17180), .ZN(
        n17182) );
  OAI21_X1 U20180 ( .B1(n18749), .B2(n17183), .A(n17182), .ZN(n17184) );
  AOI21_X1 U20181 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17198), .A(
        n17184), .ZN(n17186) );
  INV_X1 U20182 ( .A(n18810), .ZN(n18791) );
  AOI22_X1 U20183 ( .A1(n17288), .A2(n18904), .B1(n18791), .B2(n17287), .ZN(
        n17206) );
  NAND2_X1 U20184 ( .A1(n17206), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17193) );
  AND2_X1 U20185 ( .A1(n18811), .A2(n18810), .ZN(n18695) );
  INV_X1 U20186 ( .A(n18695), .ZN(n18721) );
  NAND3_X1 U20187 ( .A1(n17193), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n18721), .ZN(n17185) );
  OAI211_X1 U20188 ( .C1(n17187), .C2(n18829), .A(n17186), .B(n17185), .ZN(
        P3_U2802) );
  AOI21_X1 U20189 ( .B1(n18712), .B2(n17189), .A(n17188), .ZN(n17322) );
  INV_X1 U20190 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n17190) );
  NOR2_X1 U20191 ( .A1(n19120), .A2(n17190), .ZN(n17317) );
  INV_X1 U20192 ( .A(n17317), .ZN(n17192) );
  NAND3_X1 U20193 ( .A1(n14730), .A2(n18818), .A3(n17709), .ZN(n17191) );
  OAI211_X1 U20194 ( .C1(n18749), .C2(n13329), .A(n17192), .B(n17191), .ZN(
        n17197) );
  INV_X1 U20195 ( .A(n17193), .ZN(n17194) );
  AOI21_X1 U20196 ( .B1(n17316), .B2(n17195), .A(n17194), .ZN(n17196) );
  AOI211_X1 U20197 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17198), .A(
        n17197), .B(n17196), .ZN(n17199) );
  OAI21_X1 U20198 ( .B1(n17322), .B2(n18829), .A(n17199), .ZN(P3_U2803) );
  INV_X1 U20199 ( .A(n17200), .ZN(n17201) );
  AOI21_X1 U20200 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17202), .A(
        n17201), .ZN(n17331) );
  NOR2_X1 U20201 ( .A1(n17323), .A2(n18681), .ZN(n17209) );
  AOI21_X1 U20202 ( .B1(n13313), .B2(n19515), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17204) );
  OAI21_X1 U20203 ( .B1(n18824), .B2(n18730), .A(n17721), .ZN(n17203) );
  NAND2_X1 U20204 ( .A1(n19089), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17327) );
  OAI211_X1 U20205 ( .C1(n17205), .C2(n17204), .A(n17203), .B(n17327), .ZN(
        n17208) );
  NOR2_X1 U20206 ( .A1(n17206), .A2(n11721), .ZN(n17207) );
  AOI211_X1 U20207 ( .C1(n17209), .C2(n11721), .A(n17208), .B(n17207), .ZN(
        n17210) );
  OAI21_X1 U20208 ( .B1(n17331), .B2(n18829), .A(n17210), .ZN(P3_U2804) );
  AOI21_X1 U20209 ( .B1(n18782), .B2(n18997), .A(n18665), .ZN(n17211) );
  INV_X1 U20210 ( .A(n17211), .ZN(n19019) );
  INV_X1 U20211 ( .A(n18818), .ZN(n18739) );
  NOR2_X1 U20212 ( .A1(n18739), .A2(n17212), .ZN(n18775) );
  INV_X1 U20213 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n21625) );
  INV_X1 U20214 ( .A(n18799), .ZN(n18893) );
  INV_X1 U20215 ( .A(n18906), .ZN(n18880) );
  AOI21_X1 U20216 ( .B1(n18893), .B2(n17212), .A(n18880), .ZN(n18784) );
  OAI21_X1 U20217 ( .B1(n17213), .B2(n18737), .A(n18784), .ZN(n18773) );
  INV_X1 U20218 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19677) );
  OAI21_X1 U20219 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17213), .A(
        n17832), .ZN(n17848) );
  OAI22_X1 U20220 ( .A1(n19120), .A2(n19677), .B1(n18749), .B2(n17848), .ZN(
        n17214) );
  AOI221_X1 U20221 ( .B1(n18775), .B2(n21625), .C1(n18773), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17214), .ZN(n17223) );
  INV_X1 U20222 ( .A(n19010), .ZN(n17215) );
  OAI22_X1 U20223 ( .A1(n17216), .A2(n17215), .B1(n18997), .B2(n18810), .ZN(
        n17221) );
  INV_X1 U20224 ( .A(n19021), .ZN(n19045) );
  OR3_X1 U20225 ( .A1(n18795), .A2(n19045), .A3(n18712), .ZN(n17217) );
  NOR2_X1 U20226 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11705), .ZN(
        n18813) );
  AOI21_X1 U20227 ( .B1(n17217), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18813), .ZN(n17218) );
  OAI21_X1 U20228 ( .B1(n17219), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17218), .ZN(n17220) );
  XNOR2_X1 U20229 ( .A(n17220), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19015) );
  AOI22_X1 U20230 ( .A1(n17221), .A2(n18713), .B1(n19015), .B2(n18846), .ZN(
        n17222) );
  OAI211_X1 U20231 ( .C1(n19019), .C2(n18811), .A(n17223), .B(n17222), .ZN(
        P3_U2815) );
  INV_X1 U20232 ( .A(n17227), .ZN(n19080) );
  OR2_X1 U20233 ( .A1(n18835), .A2(n17224), .ZN(n18794) );
  OAI21_X1 U20234 ( .B1(n19080), .B2(n18833), .A(n18794), .ZN(n17225) );
  INV_X1 U20235 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n19081) );
  XNOR2_X1 U20236 ( .A(n17225), .B(n19081), .ZN(n19085) );
  INV_X1 U20237 ( .A(n17226), .ZN(n18812) );
  NAND2_X1 U20238 ( .A1(n17227), .A2(n19081), .ZN(n19087) );
  NOR2_X1 U20239 ( .A1(n18812), .A2(n17227), .ZN(n18840) );
  OR2_X1 U20240 ( .A1(n18810), .A2(n14875), .ZN(n17229) );
  INV_X1 U20241 ( .A(n19078), .ZN(n17293) );
  NAND2_X1 U20242 ( .A1(n18904), .A2(n17293), .ZN(n17228) );
  NAND2_X1 U20243 ( .A1(n17229), .A2(n17228), .ZN(n18841) );
  OAI21_X1 U20244 ( .B1(n18840), .B2(n18841), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17231) );
  NOR2_X1 U20245 ( .A1(n19055), .A2(n19670), .ZN(n19084) );
  INV_X1 U20246 ( .A(n19084), .ZN(n17230) );
  OAI211_X1 U20247 ( .C1(n18812), .C2(n19087), .A(n17231), .B(n17230), .ZN(
        n17236) );
  AND2_X1 U20248 ( .A1(n19515), .A2(n17232), .ZN(n18783) );
  INV_X1 U20249 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17914) );
  NOR2_X1 U20250 ( .A1(n19479), .A2(n17233), .ZN(n18865) );
  NAND2_X1 U20251 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18865), .ZN(
        n18859) );
  NAND2_X1 U20252 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17924) );
  NOR2_X1 U20253 ( .A1(n18859), .A2(n17924), .ZN(n17242) );
  NAND2_X1 U20254 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17242), .ZN(
        n17241) );
  NOR2_X1 U20255 ( .A1(n17914), .A2(n17241), .ZN(n18849) );
  AOI21_X1 U20256 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18860), .A(
        n18849), .ZN(n17234) );
  INV_X1 U20257 ( .A(n17947), .ZN(n17249) );
  NAND3_X1 U20258 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(n17249), .ZN(n17907) );
  NOR2_X1 U20259 ( .A1(n17914), .A2(n17907), .ZN(n17906) );
  INV_X1 U20260 ( .A(n17886), .ZN(n18802) );
  OAI21_X1 U20261 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17906), .A(
        n18802), .ZN(n17896) );
  OAI22_X1 U20262 ( .A1(n18783), .A2(n17234), .B1(n18900), .B2(n17896), .ZN(
        n17235) );
  AOI211_X1 U20263 ( .C1(n18846), .C2(n19085), .A(n17236), .B(n17235), .ZN(
        n17237) );
  INV_X1 U20264 ( .A(n17237), .ZN(P3_U2819) );
  NAND2_X1 U20265 ( .A1(n18835), .A2(n18833), .ZN(n17238) );
  XOR2_X1 U20266 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n17238), .Z(
        n19098) );
  NOR2_X1 U20267 ( .A1(n19120), .A2(n19666), .ZN(n17239) );
  AOI21_X1 U20268 ( .B1(n18841), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17239), .ZN(n17240) );
  OAI21_X1 U20269 ( .B1(n18812), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17240), .ZN(n17246) );
  INV_X1 U20270 ( .A(n17241), .ZN(n18831) );
  AOI21_X1 U20271 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18860), .A(
        n17242), .ZN(n17244) );
  INV_X1 U20272 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21622) );
  NOR2_X1 U20273 ( .A1(n21622), .A2(n17947), .ZN(n17243) );
  OAI21_X1 U20274 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17243), .A(
        n17907), .ZN(n17933) );
  OAI22_X1 U20275 ( .A1(n18831), .A2(n17244), .B1(n18900), .B2(n17933), .ZN(
        n17245) );
  AOI211_X1 U20276 ( .C1(n18846), .C2(n19098), .A(n17246), .B(n17245), .ZN(
        n17247) );
  INV_X1 U20277 ( .A(n17247), .ZN(P3_U2821) );
  OAI21_X1 U20278 ( .B1(n17248), .B2(n18799), .A(n18906), .ZN(n18850) );
  AOI22_X1 U20279 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17947), .B1(
        n17249), .B2(n21622), .ZN(n17937) );
  OAI211_X1 U20280 ( .C1(n17250), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19515), .B(n17924), .ZN(n17252) );
  OAI211_X1 U20281 ( .C1(n18900), .C2(n17937), .A(n17252), .B(n17251), .ZN(
        n17253) );
  AOI21_X1 U20282 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18850), .A(
        n17253), .ZN(n17258) );
  INV_X1 U20283 ( .A(n17254), .ZN(n17255) );
  AOI22_X1 U20284 ( .A1(n17256), .A2(n18904), .B1(n17255), .B2(n18791), .ZN(
        n17257) );
  OAI211_X1 U20285 ( .C1(n17259), .C2(n18829), .A(n17258), .B(n17257), .ZN(
        P3_U2822) );
  AOI22_X1 U20286 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18860), .B1(
        n18884), .B2(n18020), .ZN(n17261) );
  OAI211_X1 U20287 ( .C1(n18897), .C2(n17262), .A(n17261), .B(n17260), .ZN(
        n17263) );
  AOI21_X1 U20288 ( .B1(n18904), .B2(n17264), .A(n17263), .ZN(n17265) );
  INV_X1 U20289 ( .A(n17265), .ZN(P3_U2829) );
  AOI22_X1 U20290 ( .A1(n17267), .A2(n19119), .B1(n19053), .B2(n17266), .ZN(
        n17269) );
  INV_X1 U20291 ( .A(n17290), .ZN(n17268) );
  NOR3_X1 U20292 ( .A1(n17269), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n17268), .ZN(n17272) );
  INV_X1 U20293 ( .A(n17270), .ZN(n17271) );
  NOR2_X1 U20294 ( .A1(n17272), .A2(n17271), .ZN(n17280) );
  AND2_X1 U20295 ( .A1(n17314), .A2(n18971), .ZN(n19090) );
  INV_X1 U20296 ( .A(n19090), .ZN(n17275) );
  INV_X1 U20297 ( .A(n17273), .ZN(n17274) );
  AOI211_X1 U20298 ( .C1(n17316), .C2(n17275), .A(n19121), .B(n17274), .ZN(
        n17289) );
  OAI22_X1 U20299 ( .A1(n17289), .A2(n19089), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17276), .ZN(n17277) );
  OAI21_X1 U20300 ( .B1(n17278), .B2(n17277), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17279) );
  OAI211_X1 U20301 ( .C1(n17281), .C2(n19058), .A(n17280), .B(n17279), .ZN(
        P3_U2833) );
  OAI211_X1 U20302 ( .C1(n17283), .C2(n17316), .A(n19584), .B(n17282), .ZN(
        n17284) );
  AOI21_X1 U20303 ( .B1(n17286), .B2(n17285), .A(n17284), .ZN(n17292) );
  NAND2_X1 U20304 ( .A1(n19077), .A2(n19048), .ZN(n18975) );
  INV_X1 U20305 ( .A(n18975), .ZN(n19070) );
  INV_X1 U20306 ( .A(n19048), .ZN(n19075) );
  AOI22_X1 U20307 ( .A1(n17288), .A2(n19585), .B1(n19075), .B2(n17287), .ZN(
        n17313) );
  OAI211_X1 U20308 ( .C1(n17290), .C2(n19070), .A(n17313), .B(n17289), .ZN(
        n17291) );
  OAI211_X1 U20309 ( .C1(n17292), .C2(n17291), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n19120), .ZN(n17305) );
  NOR2_X1 U20310 ( .A1(n19077), .A2(n17293), .ZN(n18983) );
  NAND2_X1 U20311 ( .A1(n18983), .A2(n17294), .ZN(n17295) );
  OAI211_X1 U20312 ( .C1(n19048), .C2(n18713), .A(n18909), .B(n17295), .ZN(
        n18936) );
  NAND2_X1 U20313 ( .A1(n18936), .A2(n19053), .ZN(n18945) );
  NOR2_X1 U20314 ( .A1(n18945), .A2(n17296), .ZN(n17297) );
  AOI211_X1 U20315 ( .C1(n17299), .C2(n19099), .A(n17298), .B(n17297), .ZN(
        n17304) );
  NAND4_X1 U20316 ( .A1(n17302), .A2(n10316), .A3(n17301), .A4(n17300), .ZN(
        n17303) );
  NAND3_X1 U20317 ( .A1(n17305), .A2(n17304), .A3(n17303), .ZN(P3_U2834) );
  NAND2_X1 U20318 ( .A1(n18928), .A2(n17306), .ZN(n18970) );
  INV_X1 U20319 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17307) );
  NOR2_X1 U20320 ( .A1(n18669), .A2(n17307), .ZN(n18911) );
  INV_X1 U20321 ( .A(n18911), .ZN(n17308) );
  OAI21_X1 U20322 ( .B1(n18970), .B2(n17308), .A(n18978), .ZN(n18908) );
  AOI22_X1 U20323 ( .A1(n18998), .A2(n17309), .B1(n19122), .B2(n11720), .ZN(
        n17312) );
  INV_X1 U20324 ( .A(n17310), .ZN(n17311) );
  AND4_X1 U20325 ( .A1(n17313), .A2(n18908), .A3(n17312), .A4(n17311), .ZN(
        n17324) );
  OAI211_X1 U20326 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17314), .A(
        n17324), .B(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17320) );
  OAI22_X1 U20327 ( .A1(n18945), .A2(n17315), .B1(n19121), .B2(n17316), .ZN(
        n17319) );
  NOR2_X1 U20328 ( .A1(n19114), .A2(n17316), .ZN(n17318) );
  AOI211_X1 U20329 ( .C1(n17320), .C2(n17319), .A(n17318), .B(n17317), .ZN(
        n17321) );
  OAI21_X1 U20330 ( .B1(n17322), .B2(n19058), .A(n17321), .ZN(P3_U2835) );
  NAND3_X1 U20331 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18937), .A3(
        n18936), .ZN(n18922) );
  NOR2_X1 U20332 ( .A1(n17323), .A2(n18922), .ZN(n17326) );
  INV_X1 U20333 ( .A(n17324), .ZN(n17325) );
  MUX2_X1 U20334 ( .A(n17326), .B(n17325), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17329) );
  OAI21_X1 U20335 ( .B1(n19114), .B2(n11721), .A(n17327), .ZN(n17328) );
  AOI21_X1 U20336 ( .B1(n17329), .B2(n19053), .A(n17328), .ZN(n17330) );
  OAI21_X1 U20337 ( .B1(n17331), .B2(n19058), .A(n17330), .ZN(P3_U2836) );
  NAND2_X1 U20338 ( .A1(n17333), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17334) );
  AND2_X1 U20339 ( .A1(n18653), .A2(n17334), .ZN(n18670) );
  NOR2_X1 U20340 ( .A1(n17339), .A2(n18970), .ZN(n18927) );
  NAND2_X1 U20341 ( .A1(n18713), .A2(n19075), .ZN(n19011) );
  AOI211_X1 U20342 ( .C1(n18669), .C2(n18975), .A(n19008), .B(n18947), .ZN(
        n17335) );
  INV_X1 U20343 ( .A(n18972), .ZN(n17337) );
  OAI211_X1 U20344 ( .C1(n18995), .C2(n17338), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18924), .ZN(n17342) );
  NOR2_X1 U20345 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18921), .ZN(
        n18672) );
  NOR2_X1 U20346 ( .A1(n17339), .A2(n18945), .ZN(n17340) );
  INV_X1 U20347 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19695) );
  NOR2_X1 U20348 ( .A1(n19120), .A2(n19695), .ZN(n18661) );
  AOI21_X1 U20349 ( .B1(n18672), .B2(n17340), .A(n18661), .ZN(n17341) );
  OAI211_X1 U20350 ( .C1(n18670), .C2(n19058), .A(n17342), .B(n17341), .ZN(
        P3_U2838) );
  NAND2_X1 U20351 ( .A1(n17344), .A2(n17343), .ZN(n18022) );
  AOI211_X1 U20352 ( .C1(n17345), .C2(n17346), .A(n19588), .B(n11564), .ZN(
        n17356) );
  NAND2_X1 U20353 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18998), .ZN(
        n17347) );
  AOI21_X1 U20354 ( .B1(n17348), .B2(n17347), .A(n17345), .ZN(n17354) );
  AOI21_X1 U20355 ( .B1(n17345), .B2(n17350), .A(n17349), .ZN(n17352) );
  NOR2_X1 U20356 ( .A1(n17352), .A2(n17351), .ZN(n17353) );
  MUX2_X1 U20357 ( .A(n17354), .B(n17353), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n17355) );
  AOI211_X1 U20358 ( .C1(n19586), .C2(n18022), .A(n17356), .B(n17355), .ZN(
        n19570) );
  OAI222_X1 U20359 ( .A1(n18022), .A2(n17359), .B1(n17358), .B2(n17357), .C1(
        n18043), .C2(n19570), .ZN(n17360) );
  MUX2_X1 U20360 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17360), .S(
        n17489), .Z(P3_U3288) );
  AND2_X2 U20361 ( .A1(n18316), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n18317) );
  INV_X1 U20362 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18284) );
  INV_X1 U20363 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17836) );
  INV_X1 U20364 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n18204) );
  NAND2_X1 U20365 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .ZN(n18048) );
  NAND3_X1 U20366 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_26__SCAN_IN), .ZN(n18047) );
  INV_X1 U20367 ( .A(n18047), .ZN(n17361) );
  INV_X1 U20368 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17364) );
  AOI22_X1 U20369 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17363) );
  NAND2_X1 U20370 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n17362) );
  OAI211_X1 U20371 ( .C1(n17364), .C2(n11727), .A(n17363), .B(n17362), .ZN(
        n17365) );
  INV_X1 U20372 ( .A(n17365), .ZN(n17368) );
  AOI22_X1 U20373 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U20374 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9559), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17366) );
  NAND3_X1 U20375 ( .A1(n17368), .A2(n17367), .A3(n17366), .ZN(n17375) );
  INV_X1 U20376 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18157) );
  AOI22_X1 U20377 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17369) );
  OAI21_X1 U20378 ( .B1(n17408), .B2(n18157), .A(n17369), .ZN(n17370) );
  AOI21_X1 U20379 ( .B1(n18345), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17370), .ZN(n17373) );
  AOI22_X1 U20380 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17372) );
  AOI22_X1 U20381 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17371) );
  NAND3_X1 U20382 ( .A1(n17373), .A2(n17372), .A3(n17371), .ZN(n17374) );
  NOR2_X1 U20383 ( .A1(n17375), .A2(n17374), .ZN(n18094) );
  INV_X1 U20384 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17384) );
  INV_X1 U20385 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17378) );
  INV_X1 U20386 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17377) );
  OAI22_X1 U20387 ( .A1(n18325), .A2(n17378), .B1(n11799), .B2(n17377), .ZN(
        n17381) );
  INV_X1 U20388 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18324) );
  OAI22_X1 U20389 ( .A1(n11735), .A2(n18324), .B1(n9567), .B2(n17379), .ZN(
        n17380) );
  AOI211_X1 U20390 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17381), .B(n17380), .ZN(n17383) );
  AOI22_X1 U20391 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17382) );
  OAI211_X1 U20392 ( .C1(n18218), .C2(n17384), .A(n17383), .B(n17382), .ZN(
        n17390) );
  AOI22_X1 U20393 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U20394 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U20395 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9559), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U20396 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17385) );
  NAND4_X1 U20397 ( .A1(n17388), .A2(n17387), .A3(n17386), .A4(n17385), .ZN(
        n17389) );
  NOR2_X1 U20398 ( .A1(n17390), .A2(n17389), .ZN(n18103) );
  INV_X1 U20399 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20400 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U20401 ( .B1(n17408), .B2(n17392), .A(n17391), .ZN(n17393) );
  AOI21_X1 U20402 ( .B1(n18345), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17393), .ZN(n17396) );
  AOI22_X1 U20403 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20404 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17394) );
  NAND3_X1 U20405 ( .A1(n17396), .A2(n17395), .A3(n17394), .ZN(n17406) );
  AOI22_X1 U20406 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17398) );
  NAND2_X1 U20407 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n17397) );
  OAI211_X1 U20408 ( .C1(n17399), .C2(n18352), .A(n17398), .B(n17397), .ZN(
        n17404) );
  INV_X1 U20409 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18235) );
  INV_X1 U20410 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n21672) );
  OAI22_X1 U20411 ( .A1(n18256), .A2(n18235), .B1(n18323), .B2(n21672), .ZN(
        n17403) );
  INV_X1 U20412 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17401) );
  INV_X1 U20413 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17400) );
  OAI22_X1 U20414 ( .A1(n18358), .A2(n17401), .B1(n11727), .B2(n17400), .ZN(
        n17402) );
  OR3_X1 U20415 ( .A1(n17404), .A2(n17403), .A3(n17402), .ZN(n17405) );
  NOR2_X1 U20416 ( .A1(n17406), .A2(n17405), .ZN(n18112) );
  INV_X1 U20417 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18251) );
  AOI22_X1 U20418 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18054), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17407) );
  OAI21_X1 U20419 ( .B1(n17408), .B2(n18251), .A(n17407), .ZN(n17409) );
  AOI21_X1 U20420 ( .B1(n18345), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n17409), .ZN(n17412) );
  AOI22_X1 U20421 ( .A1(n9582), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9559), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U20422 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18334), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17410) );
  NAND3_X1 U20423 ( .A1(n17412), .A2(n17411), .A3(n17410), .ZN(n17421) );
  INV_X1 U20424 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18075) );
  AOI22_X1 U20425 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17414) );
  NAND2_X1 U20426 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n17413) );
  OAI211_X1 U20427 ( .C1(n11623), .C2(n18075), .A(n17414), .B(n17413), .ZN(
        n17415) );
  INV_X1 U20428 ( .A(n17415), .ZN(n17419) );
  AOI22_X1 U20429 ( .A1(n11784), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20430 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9555), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17417) );
  NAND3_X1 U20431 ( .A1(n17419), .A2(n17418), .A3(n17417), .ZN(n17420) );
  NOR2_X1 U20432 ( .A1(n17421), .A2(n17420), .ZN(n18111) );
  NOR2_X1 U20433 ( .A1(n18112), .A2(n18111), .ZN(n18109) );
  INV_X1 U20434 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18206) );
  INV_X1 U20435 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18213) );
  INV_X1 U20436 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18355) );
  OAI22_X1 U20437 ( .A1(n11735), .A2(n18213), .B1(n11799), .B2(n18355), .ZN(
        n17423) );
  INV_X1 U20438 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18343) );
  OAI22_X1 U20439 ( .A1(n18327), .A2(n18343), .B1(n9567), .B2(n18354), .ZN(
        n17422) );
  AOI211_X1 U20440 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n17423), .B(n17422), .ZN(n17425) );
  AOI22_X1 U20441 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17424) );
  OAI211_X1 U20442 ( .C1(n18218), .C2(n18206), .A(n17425), .B(n17424), .ZN(
        n17431) );
  AOI22_X1 U20443 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17429) );
  AOI22_X1 U20444 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20445 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U20446 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17426) );
  NAND4_X1 U20447 ( .A1(n17429), .A2(n17428), .A3(n17427), .A4(n17426), .ZN(
        n17430) );
  OR2_X1 U20448 ( .A1(n17431), .A2(n17430), .ZN(n18108) );
  NAND2_X1 U20449 ( .A1(n18109), .A2(n18108), .ZN(n18107) );
  NOR2_X1 U20450 ( .A1(n18103), .A2(n18107), .ZN(n18099) );
  INV_X1 U20451 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18302) );
  INV_X1 U20452 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18303) );
  INV_X1 U20453 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18168) );
  OAI22_X1 U20454 ( .A1(n11735), .A2(n18303), .B1(n11799), .B2(n18168), .ZN(
        n17434) );
  INV_X1 U20455 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18177) );
  OAI22_X1 U20456 ( .A1(n18327), .A2(n18177), .B1(n9567), .B2(n17432), .ZN(
        n17433) );
  AOI211_X1 U20457 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17434), .B(n17433), .ZN(n17436) );
  AOI22_X1 U20458 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17435) );
  OAI211_X1 U20459 ( .C1(n18218), .C2(n18302), .A(n17436), .B(n17435), .ZN(
        n17442) );
  AOI22_X1 U20460 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20461 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U20462 ( .A1(n9582), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U20463 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17437) );
  NAND4_X1 U20464 ( .A1(n17440), .A2(n17439), .A3(n17438), .A4(n17437), .ZN(
        n17441) );
  OR2_X1 U20465 ( .A1(n17442), .A2(n17441), .ZN(n18098) );
  NAND2_X1 U20466 ( .A1(n18099), .A2(n18098), .ZN(n18097) );
  NOR2_X1 U20467 ( .A1(n18094), .A2(n18097), .ZN(n18088) );
  INV_X1 U20468 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17448) );
  INV_X1 U20469 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17443) );
  OAI22_X1 U20470 ( .A1(n11735), .A2(n17443), .B1(n11799), .B2(n21563), .ZN(
        n17445) );
  INV_X1 U20471 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17470) );
  OAI22_X1 U20472 ( .A1(n18327), .A2(n17470), .B1(n9567), .B2(n17471), .ZN(
        n17444) );
  AOI211_X1 U20473 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n17445), .B(n17444), .ZN(n17447) );
  AOI22_X1 U20474 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17446) );
  OAI211_X1 U20475 ( .C1(n18218), .C2(n17448), .A(n17447), .B(n17446), .ZN(
        n17456) );
  AOI22_X1 U20476 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20477 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U20478 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20479 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17451) );
  NAND4_X1 U20480 ( .A1(n17454), .A2(n17453), .A3(n17452), .A4(n17451), .ZN(
        n17455) );
  OR2_X1 U20481 ( .A1(n17456), .A2(n17455), .ZN(n18089) );
  XNOR2_X1 U20482 ( .A(n18088), .B(n18089), .ZN(n18412) );
  NAND3_X1 U20483 ( .A1(n17458), .A2(P3_EBX_REG_28__SCAN_IN), .A3(n9564), .ZN(
        n17457) );
  OAI221_X1 U20484 ( .B1(n17458), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n9564), 
        .C2(n18412), .A(n17457), .ZN(P3_U2675) );
  AOI22_X1 U20485 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20486 ( .B1(n17408), .B2(n21563), .A(n17459), .ZN(n17460) );
  AOI21_X1 U20487 ( .B1(n9560), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(n17460), .ZN(n17464) );
  AOI22_X1 U20488 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9582), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17463) );
  AOI22_X1 U20489 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17462) );
  NAND3_X1 U20490 ( .A1(n17464), .A2(n17463), .A3(n17462), .ZN(n17476) );
  INV_X1 U20491 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20492 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17467) );
  NAND2_X1 U20493 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n17466) );
  OAI211_X1 U20494 ( .C1(n17468), .C2(n18352), .A(n17467), .B(n17466), .ZN(
        n17474) );
  INV_X1 U20495 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18133) );
  INV_X1 U20496 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17469) );
  OAI22_X1 U20497 ( .A1(n9557), .A2(n18133), .B1(n18323), .B2(n17469), .ZN(
        n17473) );
  OAI22_X1 U20498 ( .A1(n18256), .A2(n17471), .B1(n18321), .B2(n17470), .ZN(
        n17472) );
  OR3_X1 U20499 ( .A1(n17474), .A2(n17473), .A3(n17472), .ZN(n17475) );
  NOR2_X1 U20500 ( .A1(n17476), .A2(n17475), .ZN(n18485) );
  OAI211_X1 U20501 ( .C1(n18301), .C2(P3_EBX_REG_13__SCAN_IN), .A(n9564), .B(
        n18280), .ZN(n17477) );
  OAI21_X1 U20502 ( .B1(n18485), .B2(n9564), .A(n17477), .ZN(P3_U2690) );
  NOR2_X1 U20503 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19723), .ZN(
        n19130) );
  INV_X1 U20504 ( .A(n19130), .ZN(n19180) );
  NOR2_X1 U20505 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17478), .ZN(
        n17486) );
  INV_X1 U20506 ( .A(n17486), .ZN(n17479) );
  NOR2_X1 U20507 ( .A1(n17479), .A2(n11784), .ZN(n19126) );
  OAI211_X1 U20508 ( .C1(n19721), .C2(n19126), .A(n19428), .B(n17480), .ZN(
        n19135) );
  NAND2_X1 U20509 ( .A1(n19180), .A2(n19135), .ZN(n17483) );
  INV_X1 U20510 ( .A(n17483), .ZN(n17482) );
  INV_X1 U20511 ( .A(n19291), .ZN(n19381) );
  OAI22_X1 U20512 ( .A1(n18893), .A2(n19742), .B1(n11865), .B2(n19723), .ZN(
        n17485) );
  NAND3_X1 U20513 ( .A1(n11853), .A2(n19135), .A3(n17485), .ZN(n17481) );
  OAI221_X1 U20514 ( .B1(n11853), .B2(n17482), .C1(n11853), .C2(n19381), .A(
        n17481), .ZN(P3_U2864) );
  NAND2_X1 U20515 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19288) );
  NOR2_X1 U20516 ( .A1(n18893), .A2(n19742), .ZN(n17484) );
  AOI221_X1 U20517 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19288), .C1(n17484), 
        .C2(n19288), .A(n17483), .ZN(n19134) );
  OAI221_X1 U20518 ( .B1(n19291), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19291), .C2(n17485), .A(n19135), .ZN(n19132) );
  AOI22_X1 U20519 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19134), .B1(
        n19132), .B2(n11856), .ZN(P3_U2865) );
  NOR2_X1 U20520 ( .A1(n17486), .A2(n19588), .ZN(n19595) );
  NAND3_X1 U20521 ( .A1(n17489), .A2(n19595), .A3(n17487), .ZN(n17488) );
  OAI21_X1 U20522 ( .B1(n17489), .B2(n19583), .A(n17488), .ZN(P3_U3284) );
  INV_X1 U20523 ( .A(n17490), .ZN(n20563) );
  NOR4_X1 U20524 ( .A1(n17493), .A2(n17492), .A3(n20620), .A4(n20563), .ZN(
        n17494) );
  NAND2_X1 U20525 ( .A1(n17497), .A2(n17494), .ZN(n17495) );
  OAI21_X1 U20526 ( .B1(n17497), .B2(n17496), .A(n17495), .ZN(P2_U3595) );
  INV_X1 U20527 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17639) );
  NOR2_X1 U20528 ( .A1(n20732), .A2(n17639), .ZN(P1_U2905) );
  NAND2_X1 U20529 ( .A1(n17499), .A2(n17498), .ZN(n17501) );
  NAND2_X1 U20530 ( .A1(n17501), .A2(n17500), .ZN(n17502) );
  AND2_X1 U20531 ( .A1(n17502), .A2(n20328), .ZN(n20592) );
  INV_X1 U20532 ( .A(n20592), .ZN(n21695) );
  NOR2_X1 U20533 ( .A1(n10865), .A2(n21695), .ZN(P2_U3047) );
  AND2_X1 U20534 ( .A1(n20804), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n17526) );
  AOI21_X1 U20535 ( .B1(n20772), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n17526), .ZN(n17513) );
  INV_X1 U20536 ( .A(n17504), .ZN(n17506) );
  NOR2_X1 U20537 ( .A1(n17506), .A2(n17505), .ZN(n17517) );
  INV_X1 U20538 ( .A(n17515), .ZN(n17507) );
  OAI22_X1 U20539 ( .A1(n17517), .A2(n17508), .B1(n17507), .B2(n17514), .ZN(
        n17511) );
  XNOR2_X1 U20540 ( .A(n17509), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17510) );
  XNOR2_X1 U20541 ( .A(n17511), .B(n17510), .ZN(n17531) );
  AOI22_X1 U20542 ( .A1(n17531), .A2(n20779), .B1(n20778), .B2(n20658), .ZN(
        n17512) );
  OAI211_X1 U20543 ( .C1(n20783), .C2(n20661), .A(n17513), .B(n17512), .ZN(
        P1_U2992) );
  AOI22_X1 U20544 ( .A1(n20772), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20804), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17519) );
  XNOR2_X1 U20545 ( .A(n17515), .B(n17514), .ZN(n17516) );
  XNOR2_X1 U20546 ( .A(n17517), .B(n17516), .ZN(n17540) );
  AOI22_X1 U20547 ( .A1(n17540), .A2(n20779), .B1(n20778), .B2(n20709), .ZN(
        n17518) );
  OAI211_X1 U20548 ( .C1(n20783), .C2(n20671), .A(n17519), .B(n17518), .ZN(
        P1_U2993) );
  INV_X1 U20549 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n17520) );
  NOR2_X1 U20550 ( .A1(n20771), .A2(n17520), .ZN(n17546) );
  AOI21_X1 U20551 ( .B1(n20772), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n17546), .ZN(n17525) );
  OAI21_X1 U20552 ( .B1(n17522), .B2(n17521), .A(n17504), .ZN(n17523) );
  INV_X1 U20553 ( .A(n17523), .ZN(n17549) );
  AOI22_X1 U20554 ( .A1(n20686), .A2(n20778), .B1(n17549), .B2(n20779), .ZN(
        n17524) );
  OAI211_X1 U20555 ( .C1(n20783), .C2(n20676), .A(n17525), .B(n17524), .ZN(
        P1_U2994) );
  INV_X1 U20556 ( .A(n20655), .ZN(n17527) );
  AOI21_X1 U20557 ( .B1(n20823), .B2(n17527), .A(n17526), .ZN(n17533) );
  AND3_X1 U20558 ( .A1(n17529), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        n17528), .ZN(n17530) );
  AOI21_X1 U20559 ( .B1(n17531), .B2(n20828), .A(n17530), .ZN(n17532) );
  OAI211_X1 U20560 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17534), .A(
        n17533), .B(n17532), .ZN(P1_U3024) );
  NOR2_X1 U20561 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17535), .ZN(
        n17543) );
  AOI21_X1 U20562 ( .B1(n17538), .B2(n17537), .A(n17536), .ZN(n17539) );
  AOI22_X1 U20563 ( .A1(n17540), .A2(n20828), .B1(n20823), .B2(n10459), .ZN(
        n17542) );
  NAND2_X1 U20564 ( .A1(n20804), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n17541) );
  OAI211_X1 U20565 ( .C1(n17544), .C2(n17543), .A(n17542), .B(n17541), .ZN(
        P1_U3025) );
  NAND2_X1 U20566 ( .A1(n20790), .A2(n17545), .ZN(n20803) );
  INV_X1 U20567 ( .A(n20677), .ZN(n17547) );
  AOI21_X1 U20568 ( .B1(n20823), .B2(n17547), .A(n17546), .ZN(n17551) );
  AOI22_X1 U20569 ( .A1(n17549), .A2(n20828), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17548), .ZN(n17550) );
  OAI211_X1 U20570 ( .C1(n17552), .C2(n20803), .A(n17551), .B(n17550), .ZN(
        P1_U3026) );
  AOI21_X1 U20571 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n17561), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17559) );
  AOI21_X1 U20572 ( .B1(n17555), .B2(n17554), .A(n17553), .ZN(n17558) );
  AOI21_X1 U20573 ( .B1(n21248), .B2(n21523), .A(n17556), .ZN(n17557) );
  NOR3_X1 U20574 ( .A1(n17559), .A2(n17558), .A3(n17557), .ZN(P1_U3162) );
  OAI221_X1 U20575 ( .B1(n21248), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n21248), 
        .C2(n17561), .A(n17560), .ZN(P1_U3466) );
  NOR3_X1 U20576 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17563) );
  NOR4_X1 U20577 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17562) );
  NAND4_X1 U20578 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17563), .A3(n17562), .A4(
        U215), .ZN(U213) );
  INV_X2 U20579 ( .A(U214), .ZN(n17601) );
  NOR2_X2 U20580 ( .A1(n17601), .A2(n17564), .ZN(n17605) );
  INV_X1 U20581 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n21639) );
  OAI222_X1 U20582 ( .A1(U214), .A2(n17639), .B1(n17603), .B2(n17565), .C1(
        U212), .C2(n21639), .ZN(U216) );
  AOI22_X1 U20583 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n17600), .ZN(n17566) );
  OAI21_X1 U20584 ( .B1(n13724), .B2(n17603), .A(n17566), .ZN(U217) );
  AOI22_X1 U20585 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17600), .ZN(n17567) );
  OAI21_X1 U20586 ( .B1(n17568), .B2(n17603), .A(n17567), .ZN(U218) );
  AOI22_X1 U20587 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17600), .ZN(n17569) );
  OAI21_X1 U20588 ( .B1(n16452), .B2(n17603), .A(n17569), .ZN(U219) );
  AOI22_X1 U20589 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17600), .ZN(n17570) );
  OAI21_X1 U20590 ( .B1(n16458), .B2(n17603), .A(n17570), .ZN(U220) );
  INV_X1 U20591 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n21580) );
  AOI22_X1 U20592 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17600), .ZN(n17571) );
  OAI21_X1 U20593 ( .B1(n21580), .B2(n17603), .A(n17571), .ZN(U221) );
  AOI22_X1 U20594 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17600), .ZN(n17572) );
  OAI21_X1 U20595 ( .B1(n16476), .B2(n17603), .A(n17572), .ZN(U222) );
  AOI222_X1 U20596 ( .A1(n17600), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(n17605), 
        .B2(BUF1_REG_24__SCAN_IN), .C1(n17601), .C2(P1_DATAO_REG_24__SCAN_IN), 
        .ZN(n17573) );
  INV_X1 U20597 ( .A(n17573), .ZN(U223) );
  INV_X1 U20598 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U20599 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17600), .ZN(n17574) );
  OAI21_X1 U20600 ( .B1(n19890), .B2(n17603), .A(n17574), .ZN(U224) );
  AOI222_X1 U20601 ( .A1(n17600), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(n17605), 
        .B2(BUF1_REG_22__SCAN_IN), .C1(n17601), .C2(P1_DATAO_REG_22__SCAN_IN), 
        .ZN(n17575) );
  INV_X1 U20602 ( .A(n17575), .ZN(U225) );
  AOI22_X1 U20603 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17600), .ZN(n17576) );
  OAI21_X1 U20604 ( .B1(n16505), .B2(n17603), .A(n17576), .ZN(U226) );
  AOI22_X1 U20605 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17600), .ZN(n17577) );
  OAI21_X1 U20606 ( .B1(n16513), .B2(n17603), .A(n17577), .ZN(U227) );
  AOI22_X1 U20607 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17600), .ZN(n17578) );
  OAI21_X1 U20608 ( .B1(n19868), .B2(n17603), .A(n17578), .ZN(U228) );
  AOI22_X1 U20609 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17600), .ZN(n17579) );
  OAI21_X1 U20610 ( .B1(n16528), .B2(n17603), .A(n17579), .ZN(U229) );
  INV_X1 U20611 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n17623) );
  INV_X1 U20612 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n21560) );
  OAI222_X1 U20613 ( .A1(U212), .A2(n17623), .B1(n17603), .B2(n17580), .C1(
        U214), .C2(n21560), .ZN(U230) );
  AOI22_X1 U20614 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17600), .ZN(n17581) );
  OAI21_X1 U20615 ( .B1(n16547), .B2(n17603), .A(n17581), .ZN(U231) );
  AOI22_X1 U20616 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17600), .ZN(n17582) );
  OAI21_X1 U20617 ( .B1(n13832), .B2(n17603), .A(n17582), .ZN(U232) );
  INV_X1 U20618 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n17584) );
  AOI22_X1 U20619 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17600), .ZN(n17583) );
  OAI21_X1 U20620 ( .B1(n17584), .B2(n17603), .A(n17583), .ZN(U233) );
  INV_X1 U20621 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n17586) );
  AOI22_X1 U20622 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17600), .ZN(n17585) );
  OAI21_X1 U20623 ( .B1(n17586), .B2(n17603), .A(n17585), .ZN(U234) );
  AOI22_X1 U20624 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17600), .ZN(n17587) );
  OAI21_X1 U20625 ( .B1(n17588), .B2(n17603), .A(n17587), .ZN(U235) );
  INV_X1 U20626 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n21612) );
  AOI22_X1 U20627 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n17605), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17601), .ZN(n17589) );
  OAI21_X1 U20628 ( .B1(n21612), .B2(U212), .A(n17589), .ZN(U236) );
  INV_X1 U20629 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17616) );
  AOI22_X1 U20630 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n17605), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n17601), .ZN(n17590) );
  OAI21_X1 U20631 ( .B1(n17616), .B2(U212), .A(n17590), .ZN(U237) );
  INV_X1 U20632 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17615) );
  AOI22_X1 U20633 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n17605), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n17601), .ZN(n17591) );
  OAI21_X1 U20634 ( .B1(n17615), .B2(U212), .A(n17591), .ZN(U238) );
  INV_X1 U20635 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17593) );
  AOI22_X1 U20636 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17600), .ZN(n17592) );
  OAI21_X1 U20637 ( .B1(n17593), .B2(n17603), .A(n17592), .ZN(U239) );
  INV_X1 U20638 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17613) );
  AOI22_X1 U20639 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17605), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17601), .ZN(n17594) );
  OAI21_X1 U20640 ( .B1(n17613), .B2(U212), .A(n17594), .ZN(U240) );
  INV_X1 U20641 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17612) );
  AOI22_X1 U20642 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n17605), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n17601), .ZN(n17595) );
  OAI21_X1 U20643 ( .B1(n17612), .B2(U212), .A(n17595), .ZN(U241) );
  INV_X1 U20644 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n20731) );
  AOI22_X1 U20645 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n17605), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17600), .ZN(n17596) );
  OAI21_X1 U20646 ( .B1(n20731), .B2(U214), .A(n17596), .ZN(U242) );
  INV_X1 U20647 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n21587) );
  AOI22_X1 U20648 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n17605), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17600), .ZN(n17597) );
  OAI21_X1 U20649 ( .B1(n21587), .B2(U214), .A(n17597), .ZN(U243) );
  INV_X1 U20650 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n21655) );
  AOI22_X1 U20651 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17605), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17601), .ZN(n17598) );
  OAI21_X1 U20652 ( .B1(n21655), .B2(U212), .A(n17598), .ZN(U244) );
  INV_X1 U20653 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17609) );
  AOI22_X1 U20654 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n17605), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n17601), .ZN(n17599) );
  OAI21_X1 U20655 ( .B1(n17609), .B2(U212), .A(n17599), .ZN(U245) );
  INV_X1 U20656 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n17604) );
  AOI22_X1 U20657 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17601), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17600), .ZN(n17602) );
  OAI21_X1 U20658 ( .B1(n17604), .B2(n17603), .A(n17602), .ZN(U246) );
  INV_X1 U20659 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17607) );
  AOI22_X1 U20660 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n17605), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n17601), .ZN(n17606) );
  OAI21_X1 U20661 ( .B1(n17607), .B2(U212), .A(n17606), .ZN(U247) );
  INV_X1 U20662 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19137) );
  AOI22_X1 U20663 ( .A1(n17638), .A2(n17607), .B1(n19137), .B2(U215), .ZN(U251) );
  INV_X1 U20664 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n17608) );
  AOI22_X1 U20665 ( .A1(n17632), .A2(n17608), .B1(n19143), .B2(U215), .ZN(U252) );
  INV_X1 U20666 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19149) );
  AOI22_X1 U20667 ( .A1(n17632), .A2(n17609), .B1(n19149), .B2(U215), .ZN(U253) );
  INV_X1 U20668 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19152) );
  AOI22_X1 U20669 ( .A1(n17638), .A2(n21655), .B1(n19152), .B2(U215), .ZN(U254) );
  OAI22_X1 U20670 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17638), .ZN(n17610) );
  INV_X1 U20671 ( .A(n17610), .ZN(U255) );
  INV_X1 U20672 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17611) );
  AOI22_X1 U20673 ( .A1(n17632), .A2(n17611), .B1(n13896), .B2(U215), .ZN(U256) );
  AOI22_X1 U20674 ( .A1(n17638), .A2(n17612), .B1(n13881), .B2(U215), .ZN(U257) );
  AOI22_X1 U20675 ( .A1(n17632), .A2(n17613), .B1(n13838), .B2(U215), .ZN(U258) );
  OAI22_X1 U20676 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17638), .ZN(n17614) );
  INV_X1 U20677 ( .A(n17614), .ZN(U259) );
  AOI22_X1 U20678 ( .A1(n17638), .A2(n17615), .B1(n13851), .B2(U215), .ZN(U260) );
  INV_X1 U20679 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18502) );
  AOI22_X1 U20680 ( .A1(n17632), .A2(n17616), .B1(n18502), .B2(U215), .ZN(U261) );
  OAI22_X1 U20681 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n17638), .ZN(n17617) );
  INV_X1 U20682 ( .A(n17617), .ZN(U262) );
  INV_X1 U20683 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17618) );
  AOI22_X1 U20684 ( .A1(n17638), .A2(n17618), .B1(n18494), .B2(U215), .ZN(U263) );
  OAI22_X1 U20685 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17638), .ZN(n17619) );
  INV_X1 U20686 ( .A(n17619), .ZN(U264) );
  OAI22_X1 U20687 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17632), .ZN(n17620) );
  INV_X1 U20688 ( .A(n17620), .ZN(U265) );
  OAI22_X1 U20689 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17638), .ZN(n17621) );
  INV_X1 U20690 ( .A(n17621), .ZN(U266) );
  OAI22_X1 U20691 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17632), .ZN(n17622) );
  INV_X1 U20692 ( .A(n17622), .ZN(U267) );
  INV_X1 U20693 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19144) );
  AOI22_X1 U20694 ( .A1(n17632), .A2(n17623), .B1(n19144), .B2(U215), .ZN(U268) );
  OAI22_X1 U20695 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17638), .ZN(n17624) );
  INV_X1 U20696 ( .A(n17624), .ZN(U269) );
  INV_X1 U20697 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n17625) );
  INV_X1 U20698 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19867) );
  AOI22_X1 U20699 ( .A1(n17638), .A2(n17625), .B1(n19867), .B2(U215), .ZN(U270) );
  OAI22_X1 U20700 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17632), .ZN(n17626) );
  INV_X1 U20701 ( .A(n17626), .ZN(U271) );
  OAI22_X1 U20702 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17638), .ZN(n17627) );
  INV_X1 U20703 ( .A(n17627), .ZN(U272) );
  OAI22_X1 U20704 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17638), .ZN(n17628) );
  INV_X1 U20705 ( .A(n17628), .ZN(U273) );
  INV_X1 U20706 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n17629) );
  AOI22_X1 U20707 ( .A1(n17638), .A2(n17629), .B1(n16490), .B2(U215), .ZN(U274) );
  OAI22_X1 U20708 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17638), .ZN(n17630) );
  INV_X1 U20709 ( .A(n17630), .ZN(U275) );
  INV_X1 U20710 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n17631) );
  INV_X1 U20711 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n19857) );
  AOI22_X1 U20712 ( .A1(n17632), .A2(n17631), .B1(n19857), .B2(U215), .ZN(U276) );
  INV_X1 U20713 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n17633) );
  AOI22_X1 U20714 ( .A1(n17638), .A2(n17633), .B1(n16467), .B2(U215), .ZN(U277) );
  OAI22_X1 U20715 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17638), .ZN(n17634) );
  INV_X1 U20716 ( .A(n17634), .ZN(U278) );
  INV_X1 U20717 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n17635) );
  INV_X1 U20718 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U20719 ( .A1(n17638), .A2(n17635), .B1(n19874), .B2(U215), .ZN(U279) );
  OAI22_X1 U20720 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17638), .ZN(n17636) );
  INV_X1 U20721 ( .A(n17636), .ZN(U280) );
  INV_X1 U20722 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n17637) );
  INV_X1 U20723 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U20724 ( .A1(n17638), .A2(n17637), .B1(n19884), .B2(U215), .ZN(U281) );
  INV_X1 U20725 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19173) );
  AOI22_X1 U20726 ( .A1(n17638), .A2(n21639), .B1(n19173), .B2(U215), .ZN(U282) );
  INV_X1 U20727 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17640) );
  AOI222_X1 U20728 ( .A1(n17640), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(n17639), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n21639), .C2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n17641) );
  INV_X2 U20729 ( .A(n17643), .ZN(n17642) );
  INV_X1 U20730 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19669) );
  INV_X1 U20731 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20511) );
  AOI22_X1 U20732 ( .A1(n17642), .A2(n19669), .B1(n20511), .B2(n17643), .ZN(
        U347) );
  INV_X1 U20733 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19667) );
  INV_X1 U20734 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20509) );
  AOI22_X1 U20735 ( .A1(n17642), .A2(n19667), .B1(n20509), .B2(n17643), .ZN(
        U348) );
  INV_X1 U20736 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19665) );
  INV_X1 U20737 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20507) );
  AOI22_X1 U20738 ( .A1(n17642), .A2(n19665), .B1(n20507), .B2(n17643), .ZN(
        U349) );
  INV_X1 U20739 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19663) );
  INV_X1 U20740 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20506) );
  AOI22_X1 U20741 ( .A1(n17642), .A2(n19663), .B1(n20506), .B2(n17643), .ZN(
        U350) );
  INV_X1 U20742 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19661) );
  INV_X1 U20743 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20504) );
  AOI22_X1 U20744 ( .A1(n17642), .A2(n19661), .B1(n20504), .B2(n17643), .ZN(
        U351) );
  INV_X1 U20745 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19659) );
  INV_X1 U20746 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20502) );
  AOI22_X1 U20747 ( .A1(n17642), .A2(n19659), .B1(n20502), .B2(n17643), .ZN(
        U352) );
  INV_X1 U20748 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19657) );
  INV_X1 U20749 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20501) );
  AOI22_X1 U20750 ( .A1(n17642), .A2(n19657), .B1(n20501), .B2(n17643), .ZN(
        U353) );
  INV_X1 U20751 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n21637) );
  AOI22_X1 U20752 ( .A1(n17642), .A2(n21637), .B1(n20499), .B2(n17643), .ZN(
        U354) );
  INV_X1 U20753 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n21675) );
  INV_X1 U20754 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20547) );
  AOI22_X1 U20755 ( .A1(n17642), .A2(n21675), .B1(n20547), .B2(n17643), .ZN(
        U355) );
  INV_X1 U20756 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19705) );
  INV_X1 U20757 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20543) );
  AOI22_X1 U20758 ( .A1(n17642), .A2(n19705), .B1(n20543), .B2(n17643), .ZN(
        U356) );
  INV_X1 U20759 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19702) );
  INV_X1 U20760 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20540) );
  AOI22_X1 U20761 ( .A1(n17642), .A2(n19702), .B1(n20540), .B2(n17643), .ZN(
        U357) );
  INV_X1 U20762 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19701) );
  INV_X1 U20763 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n21636) );
  AOI22_X1 U20764 ( .A1(n17642), .A2(n19701), .B1(n21636), .B2(n17643), .ZN(
        U358) );
  INV_X1 U20765 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19700) );
  INV_X1 U20766 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20537) );
  AOI22_X1 U20767 ( .A1(n17642), .A2(n19700), .B1(n20537), .B2(n17643), .ZN(
        U359) );
  INV_X1 U20768 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19698) );
  INV_X1 U20769 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20535) );
  AOI22_X1 U20770 ( .A1(n17642), .A2(n19698), .B1(n20535), .B2(n17643), .ZN(
        U360) );
  INV_X1 U20771 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19696) );
  INV_X1 U20772 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20533) );
  AOI22_X1 U20773 ( .A1(n17642), .A2(n19696), .B1(n20533), .B2(n17643), .ZN(
        U361) );
  INV_X1 U20774 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19693) );
  INV_X1 U20775 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20532) );
  AOI22_X1 U20776 ( .A1(n17642), .A2(n19693), .B1(n20532), .B2(n17643), .ZN(
        U362) );
  INV_X1 U20777 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19692) );
  INV_X1 U20778 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20530) );
  AOI22_X1 U20779 ( .A1(n17642), .A2(n19692), .B1(n20530), .B2(n17643), .ZN(
        U363) );
  INV_X1 U20780 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19689) );
  INV_X1 U20781 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20528) );
  AOI22_X1 U20782 ( .A1(n17642), .A2(n19689), .B1(n20528), .B2(n17643), .ZN(
        U364) );
  INV_X1 U20783 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19654) );
  INV_X1 U20784 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20497) );
  AOI22_X1 U20785 ( .A1(n17642), .A2(n19654), .B1(n20497), .B2(n17643), .ZN(
        U365) );
  INV_X1 U20786 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19688) );
  INV_X1 U20787 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20526) );
  AOI22_X1 U20788 ( .A1(n17642), .A2(n19688), .B1(n20526), .B2(n17643), .ZN(
        U366) );
  INV_X1 U20789 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19685) );
  INV_X1 U20790 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20524) );
  AOI22_X1 U20791 ( .A1(n17642), .A2(n19685), .B1(n20524), .B2(n17643), .ZN(
        U367) );
  INV_X1 U20792 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19684) );
  INV_X1 U20793 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20522) );
  AOI22_X1 U20794 ( .A1(n17642), .A2(n19684), .B1(n20522), .B2(n17643), .ZN(
        U368) );
  INV_X1 U20795 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19682) );
  INV_X1 U20796 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20520) );
  AOI22_X1 U20797 ( .A1(n17642), .A2(n19682), .B1(n20520), .B2(n17643), .ZN(
        U369) );
  INV_X1 U20798 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19680) );
  INV_X1 U20799 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20518) );
  AOI22_X1 U20800 ( .A1(n17642), .A2(n19680), .B1(n20518), .B2(n17643), .ZN(
        U370) );
  INV_X1 U20801 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19678) );
  INV_X1 U20802 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20516) );
  AOI22_X1 U20803 ( .A1(n17642), .A2(n19678), .B1(n20516), .B2(n17643), .ZN(
        U371) );
  INV_X1 U20804 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19676) );
  INV_X1 U20805 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20515) );
  AOI22_X1 U20806 ( .A1(n17642), .A2(n19676), .B1(n20515), .B2(n17643), .ZN(
        U372) );
  INV_X1 U20807 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19674) );
  INV_X1 U20808 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20514) );
  AOI22_X1 U20809 ( .A1(n17642), .A2(n19674), .B1(n20514), .B2(n17643), .ZN(
        U373) );
  INV_X1 U20810 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n21658) );
  INV_X1 U20811 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20513) );
  AOI22_X1 U20812 ( .A1(n17642), .A2(n21658), .B1(n20513), .B2(n17643), .ZN(
        U374) );
  INV_X1 U20813 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19671) );
  INV_X1 U20814 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20512) );
  AOI22_X1 U20815 ( .A1(n17642), .A2(n19671), .B1(n20512), .B2(n17643), .ZN(
        U375) );
  INV_X1 U20816 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19651) );
  INV_X1 U20817 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20495) );
  AOI22_X1 U20818 ( .A1(n17642), .A2(n19651), .B1(n20495), .B2(n17643), .ZN(
        U376) );
  INV_X1 U20819 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17645) );
  INV_X1 U20820 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19650) );
  NAND3_X1 U20821 ( .A1(n19650), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n17644) );
  NAND2_X1 U20822 ( .A1(n19647), .A2(n19638), .ZN(n19634) );
  NAND2_X1 U20823 ( .A1(n17644), .A2(n19634), .ZN(n19720) );
  OAI21_X1 U20824 ( .B1(n19647), .B2(n17645), .A(n19717), .ZN(P3_U2633) );
  INV_X1 U20825 ( .A(n19753), .ZN(n17650) );
  INV_X1 U20826 ( .A(n17657), .ZN(n17646) );
  NOR2_X1 U20827 ( .A1(n17647), .A2(n17646), .ZN(n17648) );
  OAI21_X1 U20828 ( .B1(n17648), .B2(n18576), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17649) );
  OAI21_X1 U20829 ( .B1(n17650), .B2(n19740), .A(n17649), .ZN(P3_U2634) );
  AOI21_X1 U20830 ( .B1(n19647), .B2(n19650), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17651) );
  AOI22_X1 U20831 ( .A1(n19749), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17651), 
        .B2(n19731), .ZN(P3_U2635) );
  NOR2_X1 U20832 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n17652) );
  OAI21_X1 U20833 ( .B1(n17652), .B2(BS16), .A(n19720), .ZN(n19718) );
  OAI21_X1 U20834 ( .B1(n19720), .B2(n17653), .A(n19718), .ZN(P3_U2636) );
  INV_X1 U20835 ( .A(n17654), .ZN(n17656) );
  AOI211_X1 U20836 ( .C1(n10217), .C2(n17657), .A(n17656), .B(n17655), .ZN(
        n19580) );
  NOR2_X1 U20837 ( .A1(n19580), .A2(n19623), .ZN(n19733) );
  OAI21_X1 U20838 ( .B1(n19733), .B2(n19128), .A(n9644), .ZN(P3_U2637) );
  NOR4_X1 U20839 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n17661) );
  NOR4_X1 U20840 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17660) );
  NOR4_X1 U20841 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17659) );
  NOR4_X1 U20842 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17658) );
  NAND4_X1 U20843 ( .A1(n17661), .A2(n17660), .A3(n17659), .A4(n17658), .ZN(
        n17667) );
  NOR4_X1 U20844 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17665) );
  AOI211_X1 U20845 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_12__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17664) );
  NOR4_X1 U20846 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n17663) );
  NOR4_X1 U20847 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17662) );
  NAND4_X1 U20848 ( .A1(n17665), .A2(n17664), .A3(n17663), .A4(n17662), .ZN(
        n17666) );
  NOR2_X1 U20849 ( .A1(n17667), .A2(n17666), .ZN(n19730) );
  INV_X1 U20850 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19713) );
  NOR3_X1 U20851 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17669) );
  OAI21_X1 U20852 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17669), .A(n19730), .ZN(
        n17668) );
  OAI21_X1 U20853 ( .B1(n19730), .B2(n19713), .A(n17668), .ZN(P3_U2638) );
  INV_X1 U20854 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19652) );
  INV_X1 U20855 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19719) );
  AOI21_X1 U20856 ( .B1(n19652), .B2(n19719), .A(n17669), .ZN(n17670) );
  INV_X1 U20857 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19710) );
  INV_X1 U20858 ( .A(n19730), .ZN(n19727) );
  AOI22_X1 U20859 ( .A1(n19730), .A2(n17670), .B1(n19710), .B2(n19727), .ZN(
        P3_U2639) );
  NAND2_X1 U20860 ( .A1(n18011), .A2(n17671), .ZN(n17688) );
  INV_X1 U20861 ( .A(n17672), .ZN(n17673) );
  OAI22_X1 U20862 ( .A1(n17675), .A2(n18015), .B1(n11958), .B2(n17691), .ZN(
        n17676) );
  OAI21_X1 U20863 ( .B1(n17997), .B2(n17679), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17680) );
  OAI211_X1 U20864 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17688), .A(n17681), .B(
        n17680), .ZN(P3_U2641) );
  INV_X1 U20865 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19704) );
  NAND3_X1 U20866 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17703), .ZN(n17686) );
  OAI22_X1 U20867 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17686), .B1(n17685), 
        .B2(n18015), .ZN(n17687) );
  INV_X1 U20868 ( .A(n17688), .ZN(n17689) );
  OAI21_X1 U20869 ( .B1(n17693), .B2(n21602), .A(n17689), .ZN(n17690) );
  AOI22_X1 U20870 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18032), .B1(
        P3_EBX_REG_28__SCAN_IN), .B2(n17997), .ZN(n17702) );
  AND2_X1 U20871 ( .A1(n18040), .A2(n17692), .ZN(n17724) );
  AOI211_X1 U20872 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17712), .A(n17693), .B(
        n18038), .ZN(n17698) );
  AOI211_X1 U20873 ( .C1(n17696), .C2(n17695), .A(n17694), .B(n19631), .ZN(
        n17697) );
  NAND2_X1 U20874 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n17699) );
  OAI211_X1 U20875 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17703), .B(n17699), .ZN(n17700) );
  NAND3_X1 U20876 ( .A1(n17702), .A2(n17701), .A3(n17700), .ZN(P3_U2643) );
  INV_X1 U20877 ( .A(n17703), .ZN(n17716) );
  INV_X1 U20878 ( .A(n17704), .ZN(n17707) );
  INV_X1 U20879 ( .A(n17705), .ZN(n17706) );
  AOI211_X1 U20880 ( .C1(n17708), .C2(n17707), .A(n17706), .B(n19631), .ZN(
        n17711) );
  OAI22_X1 U20881 ( .A1(n17709), .A2(n18015), .B1(n17713), .B2(n18039), .ZN(
        n17710) );
  AOI211_X1 U20882 ( .C1(n17724), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17711), 
        .B(n17710), .ZN(n17715) );
  OAI211_X1 U20883 ( .C1(n17717), .C2(n17713), .A(n18011), .B(n17712), .ZN(
        n17714) );
  OAI211_X1 U20884 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17716), .A(n17715), 
        .B(n17714), .ZN(P3_U2644) );
  AOI22_X1 U20885 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18032), .B1(
        P3_EBX_REG_26__SCAN_IN), .B2(n17997), .ZN(n17726) );
  AOI211_X1 U20886 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17718), .A(n17717), .B(
        n18038), .ZN(n17723) );
  AOI211_X1 U20887 ( .C1(n17721), .C2(n17720), .A(n17719), .B(n19631), .ZN(
        n17722) );
  AOI211_X1 U20888 ( .C1(n17724), .C2(P3_REIP_REG_26__SCAN_IN), .A(n17723), 
        .B(n17722), .ZN(n17725) );
  OAI211_X1 U20889 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n17727), .A(n17726), 
        .B(n17725), .ZN(P3_U2645) );
  OR2_X1 U20890 ( .A1(n18038), .A2(n17728), .ZN(n17743) );
  AOI21_X1 U20891 ( .B1(n18011), .B2(n17728), .A(n17997), .ZN(n17739) );
  AOI211_X1 U20892 ( .C1(n17731), .C2(n17730), .A(n17729), .B(n19631), .ZN(
        n17737) );
  NOR2_X1 U20893 ( .A1(n18004), .A2(n17732), .ZN(n17735) );
  OAI21_X1 U20894 ( .B1(n17742), .B2(n18004), .A(n18042), .ZN(n17758) );
  AOI21_X1 U20895 ( .B1(n18034), .B2(n19695), .A(n17758), .ZN(n17733) );
  INV_X1 U20896 ( .A(n17733), .ZN(n17734) );
  MUX2_X1 U20897 ( .A(n17735), .B(n17734), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n17736) );
  AOI211_X1 U20898 ( .C1(n18032), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17737), .B(n17736), .ZN(n17738) );
  OAI221_X1 U20899 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17743), .C1(n17740), 
        .C2(n17739), .A(n17738), .ZN(P3_U2646) );
  NOR2_X1 U20900 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18004), .ZN(n17741) );
  AOI22_X1 U20901 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17997), .B1(n17742), 
        .B2(n17741), .ZN(n17750) );
  AOI21_X1 U20902 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17759), .A(n17743), .ZN(
        n17748) );
  AOI211_X1 U20903 ( .C1(n17746), .C2(n17745), .A(n17744), .B(n19631), .ZN(
        n17747) );
  AOI211_X1 U20904 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n17758), .A(n17748), 
        .B(n17747), .ZN(n17749) );
  OAI211_X1 U20905 ( .C1(n18663), .C2(n18015), .A(n17750), .B(n17749), .ZN(
        P3_U2647) );
  OAI21_X1 U20906 ( .B1(n18004), .B2(n17751), .A(n19694), .ZN(n17757) );
  AOI211_X1 U20907 ( .C1(n17754), .C2(n17753), .A(n17752), .B(n19631), .ZN(
        n17756) );
  INV_X1 U20908 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18686) );
  OAI22_X1 U20909 ( .A1(n18686), .A2(n18015), .B1(n18106), .B2(n18039), .ZN(
        n17755) );
  AOI211_X1 U20910 ( .C1(n17758), .C2(n17757), .A(n17756), .B(n17755), .ZN(
        n17761) );
  OAI211_X1 U20911 ( .C1(n17762), .C2(n18106), .A(n18011), .B(n17759), .ZN(
        n17760) );
  NAND2_X1 U20912 ( .A1(n17761), .A2(n17760), .ZN(P3_U2648) );
  AOI22_X1 U20913 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18032), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n17997), .ZN(n17775) );
  AOI211_X1 U20914 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17779), .A(n17762), .B(
        n18038), .ZN(n17767) );
  INV_X1 U20915 ( .A(n17763), .ZN(n17764) );
  AOI211_X1 U20916 ( .C1(n18699), .C2(n17765), .A(n17764), .B(n19631), .ZN(
        n17766) );
  NOR2_X1 U20917 ( .A1(n17767), .A2(n17766), .ZN(n17774) );
  INV_X1 U20918 ( .A(n17768), .ZN(n17769) );
  OAI21_X1 U20919 ( .B1(n17769), .B2(n18004), .A(n18042), .ZN(n17790) );
  NAND3_X1 U20920 ( .A1(n19690), .A2(n18034), .A3(n17769), .ZN(n17783) );
  INV_X1 U20921 ( .A(n17783), .ZN(n17770) );
  OAI21_X1 U20922 ( .B1(n17790), .B2(n17770), .A(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n17773) );
  INV_X1 U20923 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19691) );
  NAND3_X1 U20924 ( .A1(n18034), .A2(n17771), .A3(n19691), .ZN(n17772) );
  NAND4_X1 U20925 ( .A1(n17775), .A2(n17774), .A3(n17773), .A4(n17772), .ZN(
        P3_U2649) );
  AOI211_X1 U20926 ( .C1(n17778), .C2(n17777), .A(n17776), .B(n19631), .ZN(
        n17782) );
  OAI211_X1 U20927 ( .C1(n17787), .C2(n18049), .A(n18011), .B(n17779), .ZN(
        n17780) );
  OAI21_X1 U20928 ( .B1(n18015), .B2(n21596), .A(n17780), .ZN(n17781) );
  AOI211_X1 U20929 ( .C1(n17790), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17782), 
        .B(n17781), .ZN(n17784) );
  OAI211_X1 U20930 ( .C1(n18039), .C2(n18049), .A(n17784), .B(n17783), .ZN(
        P3_U2650) );
  AOI211_X1 U20931 ( .C1(n18731), .C2(n17786), .A(n17785), .B(n19631), .ZN(
        n17789) );
  AOI211_X1 U20932 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17800), .A(n17787), .B(
        n18038), .ZN(n17788) );
  AOI211_X1 U20933 ( .C1(n17997), .C2(P3_EBX_REG_20__SCAN_IN), .A(n17789), .B(
        n17788), .ZN(n17793) );
  OAI221_X1 U20934 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n18034), .C1(
        P3_REIP_REG_20__SCAN_IN), .C2(n17791), .A(n17790), .ZN(n17792) );
  OAI211_X1 U20935 ( .C1(n18015), .C2(n18727), .A(n17793), .B(n17792), .ZN(
        P3_U2651) );
  NAND2_X1 U20936 ( .A1(n18034), .A2(n19686), .ZN(n17805) );
  INV_X1 U20937 ( .A(n17794), .ZN(n17817) );
  NOR3_X1 U20938 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n18004), .A3(n17817), 
        .ZN(n17807) );
  OAI21_X1 U20939 ( .B1(n17794), .B2(n18004), .A(n18042), .ZN(n17806) );
  INV_X1 U20940 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18752) );
  NOR2_X1 U20941 ( .A1(n18020), .A2(n9741), .ZN(n18738) );
  INV_X1 U20942 ( .A(n18738), .ZN(n17820) );
  NOR2_X1 U20943 ( .A1(n18752), .A2(n17820), .ZN(n17808) );
  AOI21_X1 U20944 ( .B1(n17808), .B2(n17833), .A(n18000), .ZN(n17796) );
  OAI21_X1 U20945 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17808), .A(
        n17795), .ZN(n18743) );
  XOR2_X1 U20946 ( .A(n17796), .B(n18743), .Z(n17798) );
  AOI22_X1 U20947 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18032), .B1(
        P3_EBX_REG_19__SCAN_IN), .B2(n17997), .ZN(n17797) );
  OAI211_X1 U20948 ( .C1(n19631), .C2(n17798), .A(n17797), .B(n19120), .ZN(
        n17799) );
  AOI221_X1 U20949 ( .B1(n17807), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n17806), 
        .C2(P3_REIP_REG_19__SCAN_IN), .A(n17799), .ZN(n17803) );
  OAI211_X1 U20950 ( .C1(n17812), .C2(n17801), .A(n18011), .B(n17800), .ZN(
        n17802) );
  OAI211_X1 U20951 ( .C1(n17805), .C2(n17804), .A(n17803), .B(n17802), .ZN(
        P3_U2652) );
  INV_X1 U20952 ( .A(n17806), .ZN(n17823) );
  INV_X1 U20953 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19683) );
  AOI211_X1 U20954 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17997), .A(n19089), .B(
        n17807), .ZN(n17816) );
  AOI21_X1 U20955 ( .B1(n18752), .B2(n17820), .A(n17808), .ZN(n17809) );
  INV_X1 U20956 ( .A(n17809), .ZN(n18748) );
  INV_X1 U20957 ( .A(n17833), .ZN(n17849) );
  OAI21_X1 U20958 ( .B1(n17820), .B2(n17849), .A(n13330), .ZN(n17811) );
  OAI21_X1 U20959 ( .B1(n18748), .B2(n17811), .A(n18025), .ZN(n17810) );
  AOI21_X1 U20960 ( .B1(n18748), .B2(n17811), .A(n17810), .ZN(n17814) );
  AOI211_X1 U20961 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17826), .A(n17812), .B(
        n18038), .ZN(n17813) );
  AOI211_X1 U20962 ( .C1(n18032), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17814), .B(n17813), .ZN(n17815) );
  OAI211_X1 U20963 ( .C1(n17823), .C2(n19683), .A(n17816), .B(n17815), .ZN(
        P3_U2653) );
  INV_X1 U20964 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17830) );
  NAND2_X1 U20965 ( .A1(n18034), .A2(n17817), .ZN(n17818) );
  OAI22_X1 U20966 ( .A1(n17827), .A2(n18039), .B1(n17819), .B2(n17818), .ZN(
        n17825) );
  AND2_X1 U20967 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18761), .ZN(
        n17831) );
  AOI21_X1 U20968 ( .B1(n17833), .B2(n17831), .A(n18000), .ZN(n17821) );
  OAI21_X1 U20969 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17831), .A(
        n17820), .ZN(n18764) );
  XOR2_X1 U20970 ( .A(n17821), .B(n18764), .Z(n17822) );
  OAI22_X1 U20971 ( .A1(n17823), .A2(n19681), .B1(n19631), .B2(n17822), .ZN(
        n17824) );
  NOR3_X1 U20972 ( .A1(n19089), .A2(n17825), .A3(n17824), .ZN(n17829) );
  OAI211_X1 U20973 ( .C1(n17835), .C2(n17827), .A(n18011), .B(n17826), .ZN(
        n17828) );
  OAI211_X1 U20974 ( .C1(n18015), .C2(n17830), .A(n17829), .B(n17828), .ZN(
        P3_U2654) );
  INV_X1 U20975 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17837) );
  AOI21_X1 U20976 ( .B1(n17837), .B2(n17832), .A(n17831), .ZN(n18772) );
  NOR2_X1 U20977 ( .A1(n17833), .A2(n18000), .ZN(n17834) );
  XNOR2_X1 U20978 ( .A(n18772), .B(n17834), .ZN(n17845) );
  AOI211_X1 U20979 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17854), .A(n17835), .B(
        n18038), .ZN(n17843) );
  OAI22_X1 U20980 ( .A1(n17837), .A2(n18015), .B1(n17836), .B2(n18039), .ZN(
        n17842) );
  NOR3_X1 U20981 ( .A1(n18004), .A2(n19673), .A3(n17869), .ZN(n17863) );
  NAND2_X1 U20982 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17863), .ZN(n17847) );
  NOR2_X1 U20983 ( .A1(n19677), .A2(n17847), .ZN(n17840) );
  NAND2_X1 U20984 ( .A1(n17838), .A2(n18042), .ZN(n17862) );
  OAI21_X1 U20985 ( .B1(n19677), .B2(n17862), .A(n18040), .ZN(n17846) );
  INV_X1 U20986 ( .A(n17846), .ZN(n17839) );
  MUX2_X1 U20987 ( .A(n17840), .B(n17839), .S(P3_REIP_REG_16__SCAN_IN), .Z(
        n17841) );
  NOR3_X1 U20988 ( .A1(n17843), .A2(n17842), .A3(n17841), .ZN(n17844) );
  OAI211_X1 U20989 ( .C1(n17845), .C2(n19631), .A(n17844), .B(n19120), .ZN(
        P3_U2655) );
  AOI21_X1 U20990 ( .B1(n19677), .B2(n17847), .A(n17846), .ZN(n17853) );
  AOI211_X1 U20991 ( .C1(n13330), .C2(n17858), .A(n17965), .B(n17848), .ZN(
        n17852) );
  NAND2_X1 U20992 ( .A1(n17849), .A2(n17848), .ZN(n17850) );
  OAI22_X1 U20993 ( .A1(n21625), .A2(n18015), .B1(n17959), .B2(n17850), .ZN(
        n17851) );
  NOR4_X1 U20994 ( .A1(n19089), .A2(n17853), .A3(n17852), .A4(n17851), .ZN(
        n17856) );
  OAI211_X1 U20995 ( .C1(n17861), .C2(n17857), .A(n18011), .B(n17854), .ZN(
        n17855) );
  OAI211_X1 U20996 ( .C1(n18039), .C2(n17857), .A(n17856), .B(n17855), .ZN(
        P3_U2656) );
  INV_X1 U20997 ( .A(n18805), .ZN(n17860) );
  NOR2_X1 U20998 ( .A1(n17860), .A2(n18802), .ZN(n17859) );
  OAI21_X1 U20999 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17859), .A(
        n17858), .ZN(n18786) );
  NOR2_X1 U21000 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18020), .ZN(
        n18026) );
  AOI21_X1 U21001 ( .B1(n17232), .B2(n18026), .A(n18000), .ZN(n17887) );
  AOI21_X1 U21002 ( .B1(n13330), .B2(n17860), .A(n17887), .ZN(n17872) );
  XNOR2_X1 U21003 ( .A(n18786), .B(n17872), .ZN(n17868) );
  AOI211_X1 U21004 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17873), .A(n17861), .B(
        n18038), .ZN(n17866) );
  OAI211_X1 U21005 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n17863), .A(n18040), 
        .B(n17862), .ZN(n17864) );
  OAI211_X1 U21006 ( .C1(n18284), .C2(n18039), .A(n19055), .B(n17864), .ZN(
        n17865) );
  AOI211_X1 U21007 ( .C1(n18032), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17866), .B(n17865), .ZN(n17867) );
  OAI21_X1 U21008 ( .B1(n17868), .B2(n19631), .A(n17867), .ZN(P3_U2657) );
  NOR2_X1 U21009 ( .A1(n18004), .A2(n17869), .ZN(n17870) );
  AOI22_X1 U21010 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17997), .B1(n17870), 
        .B2(n19673), .ZN(n17881) );
  NAND2_X1 U21011 ( .A1(n18025), .A2(n18000), .ZN(n18029) );
  AOI21_X1 U21012 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18029), .A(
        n17965), .ZN(n17878) );
  NAND2_X1 U21013 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17886), .ZN(
        n17871) );
  AOI22_X1 U21014 ( .A1(n17886), .A2(n18805), .B1(n18803), .B2(n17871), .ZN(
        n18808) );
  NOR3_X1 U21015 ( .A1(n18808), .A2(n17872), .A3(n19631), .ZN(n17877) );
  OAI211_X1 U21016 ( .C1(n17882), .C2(n17874), .A(n18011), .B(n17873), .ZN(
        n17875) );
  OAI21_X1 U21017 ( .B1(n18015), .B2(n18803), .A(n17875), .ZN(n17876) );
  AOI211_X1 U21018 ( .C1(n17878), .C2(n18808), .A(n17877), .B(n17876), .ZN(
        n17880) );
  OAI21_X1 U21019 ( .B1(n17885), .B2(n18004), .A(n18042), .ZN(n17903) );
  NOR2_X1 U21020 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18004), .ZN(n17884) );
  OAI21_X1 U21021 ( .B1(n17903), .B2(n17884), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n17879) );
  NAND4_X1 U21022 ( .A1(n17881), .A2(n17880), .A3(n19055), .A4(n17879), .ZN(
        P3_U2658) );
  AOI211_X1 U21023 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17897), .A(n17882), .B(
        n18038), .ZN(n17883) );
  AOI21_X1 U21024 ( .B1(n18032), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17883), .ZN(n17891) );
  AOI22_X1 U21025 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17997), .B1(n17885), 
        .B2(n17884), .ZN(n17890) );
  AOI22_X1 U21026 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17886), .B1(
        n18802), .B2(n18820), .ZN(n18823) );
  XOR2_X1 U21027 ( .A(n18823), .B(n17887), .Z(n17888) );
  AOI22_X1 U21028 ( .A1(n18025), .A2(n17888), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n17903), .ZN(n17889) );
  NAND4_X1 U21029 ( .A1(n17891), .A2(n17890), .A3(n17889), .A4(n19055), .ZN(
        P3_U2659) );
  OAI21_X1 U21030 ( .B1(n18004), .B2(n17892), .A(n19670), .ZN(n17902) );
  INV_X1 U21031 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17900) );
  AOI21_X1 U21032 ( .B1(n18001), .B2(n17906), .A(n18000), .ZN(n17893) );
  INV_X1 U21033 ( .A(n17893), .ZN(n17895) );
  AOI21_X1 U21034 ( .B1(n17896), .B2(n17895), .A(n19631), .ZN(n17894) );
  OAI21_X1 U21035 ( .B1(n17896), .B2(n17895), .A(n17894), .ZN(n17899) );
  OAI211_X1 U21036 ( .C1(n17910), .C2(n17905), .A(n18011), .B(n17897), .ZN(
        n17898) );
  OAI211_X1 U21037 ( .C1(n18015), .C2(n17900), .A(n17899), .B(n17898), .ZN(
        n17901) );
  AOI21_X1 U21038 ( .B1(n17903), .B2(n17902), .A(n17901), .ZN(n17904) );
  OAI211_X1 U21039 ( .C1(n17905), .C2(n18039), .A(n17904), .B(n19120), .ZN(
        P3_U2660) );
  AOI21_X1 U21040 ( .B1(n17914), .B2(n17907), .A(n17906), .ZN(n18839) );
  NAND2_X1 U21041 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17908) );
  AND2_X1 U21042 ( .A1(n17248), .A2(n18026), .ZN(n17960) );
  NAND2_X1 U21043 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17960), .ZN(
        n17936) );
  OAI21_X1 U21044 ( .B1(n17908), .B2(n17936), .A(n13330), .ZN(n17909) );
  INV_X1 U21045 ( .A(n17909), .ZN(n17925) );
  XNOR2_X1 U21046 ( .A(n18839), .B(n17925), .ZN(n17920) );
  AOI211_X1 U21047 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17921), .A(n17910), .B(
        n18038), .ZN(n17911) );
  AOI211_X1 U21048 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17997), .A(n19089), .B(
        n17911), .ZN(n17919) );
  AOI21_X1 U21049 ( .B1(n17912), .B2(n18034), .A(n17983), .ZN(n17939) );
  INV_X1 U21050 ( .A(n17939), .ZN(n17917) );
  NOR3_X1 U21051 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18004), .A3(n17912), .ZN(
        n17930) );
  NAND2_X1 U21052 ( .A1(n18034), .A2(n17913), .ZN(n17915) );
  OAI22_X1 U21053 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n17915), .B1(n17914), 
        .B2(n18015), .ZN(n17916) );
  AOI221_X1 U21054 ( .B1(n17917), .B2(P3_REIP_REG_10__SCAN_IN), .C1(n17930), 
        .C2(P3_REIP_REG_10__SCAN_IN), .A(n17916), .ZN(n17918) );
  OAI211_X1 U21055 ( .C1(n19631), .C2(n17920), .A(n17919), .B(n17918), .ZN(
        P3_U2661) );
  OAI211_X1 U21056 ( .C1(n17934), .C2(n17923), .A(n18011), .B(n17921), .ZN(
        n17922) );
  OAI211_X1 U21057 ( .C1(n17923), .C2(n18039), .A(n19055), .B(n17922), .ZN(
        n17929) );
  NOR2_X1 U21058 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17924), .ZN(
        n17926) );
  AOI22_X1 U21059 ( .A1(n17926), .A2(n17960), .B1(n17925), .B2(n17933), .ZN(
        n17927) );
  OAI22_X1 U21060 ( .A1(n17927), .A2(n19631), .B1(n19666), .B2(n17939), .ZN(
        n17928) );
  AOI211_X1 U21061 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18032), .A(
        n17929), .B(n17928), .ZN(n17932) );
  INV_X1 U21062 ( .A(n17930), .ZN(n17931) );
  OAI211_X1 U21063 ( .C1(n18029), .C2(n17933), .A(n17932), .B(n17931), .ZN(
        P3_U2662) );
  AOI211_X1 U21064 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17950), .A(n17934), .B(
        n18038), .ZN(n17942) );
  AND2_X1 U21065 ( .A1(n18034), .A2(n17935), .ZN(n17945) );
  AOI21_X1 U21066 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n17945), .A(
        P3_REIP_REG_8__SCAN_IN), .ZN(n17940) );
  NAND2_X1 U21067 ( .A1(n13330), .A2(n17936), .ZN(n17949) );
  XNOR2_X1 U21068 ( .A(n17937), .B(n17949), .ZN(n17938) );
  OAI22_X1 U21069 ( .A1(n17940), .A2(n17939), .B1(n19631), .B2(n17938), .ZN(
        n17941) );
  AOI211_X1 U21070 ( .C1(n18032), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17942), .B(n17941), .ZN(n17943) );
  OAI211_X1 U21071 ( .C1(n17944), .C2(n18039), .A(n17943), .B(n19120), .ZN(
        P3_U2663) );
  INV_X1 U21072 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U21073 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17997), .B1(n17945), .B2(
        n19662), .ZN(n17957) );
  NAND2_X1 U21074 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17946), .ZN(
        n17973) );
  INV_X1 U21075 ( .A(n17973), .ZN(n17991) );
  NAND2_X1 U21076 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17991), .ZN(
        n17972) );
  NOR2_X1 U21077 ( .A1(n18864), .A2(n17972), .ZN(n17958) );
  OAI21_X1 U21078 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17958), .A(
        n17947), .ZN(n18855) );
  OAI21_X1 U21079 ( .B1(n17960), .B2(n18855), .A(n18025), .ZN(n17948) );
  AOI22_X1 U21080 ( .A1(n18855), .A2(n17949), .B1(n18029), .B2(n17948), .ZN(
        n17953) );
  OAI211_X1 U21081 ( .C1(n18371), .C2(n17962), .A(n17950), .B(n18011), .ZN(
        n17951) );
  INV_X1 U21082 ( .A(n17951), .ZN(n17952) );
  AOI211_X1 U21083 ( .C1(n18032), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n17953), .B(n17952), .ZN(n17956) );
  NOR3_X1 U21084 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18004), .A3(n17954), .ZN(
        n17964) );
  AOI21_X1 U21085 ( .B1(n17954), .B2(n18034), .A(n17983), .ZN(n17976) );
  INV_X1 U21086 ( .A(n17976), .ZN(n17967) );
  OAI21_X1 U21087 ( .B1(n17964), .B2(n17967), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n17955) );
  NAND4_X1 U21088 ( .A1(n17957), .A2(n17956), .A3(n19055), .A4(n17955), .ZN(
        P3_U2664) );
  AOI21_X1 U21089 ( .B1(n18864), .B2(n17972), .A(n17958), .ZN(n18866) );
  NOR3_X1 U21090 ( .A1(n18866), .A2(n17960), .A3(n17959), .ZN(n17961) );
  AOI21_X1 U21091 ( .B1(n17997), .B2(P3_EBX_REG_6__SCAN_IN), .A(n17961), .ZN(
        n17970) );
  AOI211_X1 U21092 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17978), .A(n17962), .B(
        n18038), .ZN(n17963) );
  AOI211_X1 U21093 ( .C1(n18032), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17964), .B(n17963), .ZN(n17969) );
  AOI21_X1 U21094 ( .B1(n13330), .B2(n17972), .A(n17965), .ZN(n17966) );
  AOI22_X1 U21095 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17967), .B1(n18866), 
        .B2(n17966), .ZN(n17968) );
  NAND4_X1 U21096 ( .A1(n17970), .A2(n17969), .A3(n17968), .A4(n19055), .ZN(
        P3_U2665) );
  INV_X1 U21097 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17982) );
  AOI21_X1 U21098 ( .B1(n18034), .B2(n17971), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n17975) );
  OAI21_X1 U21099 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17991), .A(
        n17972), .ZN(n18877) );
  OAI21_X1 U21100 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17973), .A(
        n13330), .ZN(n17992) );
  XNOR2_X1 U21101 ( .A(n18877), .B(n17992), .ZN(n17974) );
  OAI22_X1 U21102 ( .A1(n17976), .A2(n17975), .B1(n19631), .B2(n17974), .ZN(
        n17977) );
  AOI211_X1 U21103 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17997), .A(n19089), .B(
        n17977), .ZN(n17981) );
  OAI211_X1 U21104 ( .C1(n17984), .C2(n17979), .A(n18011), .B(n17978), .ZN(
        n17980) );
  OAI211_X1 U21105 ( .C1(n18015), .C2(n17982), .A(n17981), .B(n17980), .ZN(
        P3_U2666) );
  AOI21_X1 U21106 ( .B1(n18034), .B2(n17994), .A(n17983), .ZN(n18003) );
  AOI211_X1 U21107 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18010), .A(n17984), .B(
        n18038), .ZN(n17989) );
  NOR2_X1 U21108 ( .A1(n9560), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n17985) );
  OAI21_X1 U21109 ( .B1(n18046), .B2(n17985), .A(n19120), .ZN(n17986) );
  INV_X1 U21110 ( .A(n17986), .ZN(n17987) );
  OAI21_X1 U21111 ( .B1(n18015), .B2(n18882), .A(n17987), .ZN(n17988) );
  NOR2_X1 U21112 ( .A1(n17989), .A2(n17988), .ZN(n17999) );
  OR2_X1 U21113 ( .A1(n18020), .A2(n17990), .ZN(n18002) );
  AOI21_X1 U21114 ( .B1(n18882), .B2(n18002), .A(n17991), .ZN(n18885) );
  NOR2_X1 U21115 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17990), .ZN(
        n18878) );
  AOI22_X1 U21116 ( .A1(n18026), .A2(n18878), .B1(n18885), .B2(n18000), .ZN(
        n17993) );
  AOI221_X1 U21117 ( .B1(n18885), .B2(n17993), .C1(n17992), .C2(n17993), .A(
        n19631), .ZN(n17996) );
  NOR3_X1 U21118 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18004), .A3(n17994), .ZN(
        n17995) );
  AOI211_X1 U21119 ( .C1(n17997), .C2(P3_EBX_REG_4__SCAN_IN), .A(n17996), .B(
        n17995), .ZN(n17998) );
  OAI211_X1 U21120 ( .C1(n19656), .C2(n18003), .A(n17999), .B(n17998), .ZN(
        P3_U2667) );
  INV_X1 U21121 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21653) );
  INV_X1 U21122 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18907) );
  NOR2_X1 U21123 ( .A1(n18020), .A2(n18907), .ZN(n18019) );
  AOI21_X1 U21124 ( .B1(n18019), .B2(n18001), .A(n18000), .ZN(n18024) );
  OAI21_X1 U21125 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18019), .A(
        n18002), .ZN(n18896) );
  XNOR2_X1 U21126 ( .A(n18024), .B(n18896), .ZN(n18009) );
  NAND2_X1 U21127 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n18033) );
  AOI221_X1 U21128 ( .B1(n18004), .B2(n19655), .C1(n18033), .C2(n19655), .A(
        n18003), .ZN(n18008) );
  INV_X1 U21129 ( .A(n18005), .ZN(n18006) );
  OAI22_X1 U21130 ( .A1(n18046), .A2(n18006), .B1(n18012), .B2(n18039), .ZN(
        n18007) );
  AOI211_X1 U21131 ( .C1(n18025), .C2(n18009), .A(n18008), .B(n18007), .ZN(
        n18014) );
  OAI211_X1 U21132 ( .C1(n18017), .C2(n18012), .A(n18011), .B(n18010), .ZN(
        n18013) );
  OAI211_X1 U21133 ( .C1(n18015), .C2(n21653), .A(n18014), .B(n18013), .ZN(
        P3_U2668) );
  INV_X1 U21134 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n18037) );
  INV_X1 U21135 ( .A(n18016), .ZN(n18018) );
  AOI211_X1 U21136 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18018), .A(n18017), .B(
        n18038), .ZN(n18031) );
  AOI21_X1 U21137 ( .B1(n18020), .B2(n18907), .A(n18019), .ZN(n18021) );
  INV_X1 U21138 ( .A(n18021), .ZN(n18899) );
  OAI22_X1 U21139 ( .A1(n18046), .A2(n18022), .B1(n18042), .B2(n19653), .ZN(
        n18023) );
  INV_X1 U21140 ( .A(n18023), .ZN(n18028) );
  OAI211_X1 U21141 ( .C1(n18026), .C2(n18899), .A(n18025), .B(n18024), .ZN(
        n18027) );
  OAI211_X1 U21142 ( .C1(n18029), .C2(n18899), .A(n18028), .B(n18027), .ZN(
        n18030) );
  AOI211_X1 U21143 ( .C1(n18032), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n18031), .B(n18030), .ZN(n18036) );
  OAI211_X1 U21144 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n18034), .B(n18033), .ZN(n18035) );
  OAI211_X1 U21145 ( .C1(n18039), .C2(n18037), .A(n18036), .B(n18035), .ZN(
        P3_U2669) );
  NAND2_X1 U21146 ( .A1(n18039), .A2(n18038), .ZN(n18041) );
  AOI22_X1 U21147 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n18041), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n18040), .ZN(n18045) );
  NAND3_X1 U21148 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18043), .A3(
        n18042), .ZN(n18044) );
  OAI211_X1 U21149 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18046), .A(
        n18045), .B(n18044), .ZN(P3_U2671) );
  NOR4_X1 U21150 ( .A1(n18049), .A2(n18048), .A3(n18047), .A4(n21602), .ZN(
        n18050) );
  NAND4_X1 U21151 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18147), .A3(
        P3_EBX_REG_22__SCAN_IN), .A4(n18050), .ZN(n18084) );
  NOR2_X1 U21152 ( .A1(n18085), .A2(n18084), .ZN(n18053) );
  NAND2_X1 U21153 ( .A1(n9564), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18052) );
  NAND2_X1 U21154 ( .A1(n18053), .A2(n11836), .ZN(n18051) );
  OAI22_X1 U21155 ( .A1(n18053), .A2(n18052), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18051), .ZN(P3_U2672) );
  INV_X1 U21156 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18117) );
  AOI22_X1 U21157 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18056) );
  NAND2_X1 U21158 ( .A1(n18170), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n18055) );
  OAI211_X1 U21159 ( .C1(n11623), .C2(n18117), .A(n18056), .B(n18055), .ZN(
        n18057) );
  INV_X1 U21160 ( .A(n18057), .ZN(n18060) );
  AOI22_X1 U21161 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18059) );
  AOI22_X1 U21162 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9559), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18058) );
  NAND3_X1 U21163 ( .A1(n18060), .A2(n18059), .A3(n18058), .ZN(n18068) );
  AOI22_X1 U21164 ( .A1(n11684), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18061) );
  OAI21_X1 U21165 ( .B1(n18352), .B2(n18062), .A(n18061), .ZN(n18063) );
  AOI21_X1 U21166 ( .B1(n18345), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n18063), .ZN(n18066) );
  AOI22_X1 U21167 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18065) );
  AOI22_X1 U21168 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18064) );
  NAND3_X1 U21169 ( .A1(n18066), .A2(n18065), .A3(n18064), .ZN(n18067) );
  OR2_X1 U21170 ( .A1(n18068), .A2(n18067), .ZN(n18090) );
  NAND3_X1 U21171 ( .A1(n18089), .A2(n18088), .A3(n18090), .ZN(n18083) );
  INV_X1 U21172 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18069) );
  OAI22_X1 U21173 ( .A1(n18253), .A2(n18069), .B1(n18321), .B2(n21652), .ZN(
        n18072) );
  INV_X1 U21174 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18070) );
  OAI22_X1 U21175 ( .A1(n18255), .A2(n9567), .B1(n11799), .B2(n18070), .ZN(
        n18071) );
  AOI211_X1 U21176 ( .C1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n9560), .A(
        n18072), .B(n18071), .ZN(n18074) );
  AOI22_X1 U21177 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18330), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18073) );
  OAI211_X1 U21178 ( .C1(n18218), .C2(n18075), .A(n18074), .B(n18073), .ZN(
        n18081) );
  AOI22_X1 U21179 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17461), .B1(
        n18054), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U21180 ( .A1(n9582), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9561), .B1(n9556), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18077) );
  AOI22_X1 U21182 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11628), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18076) );
  NAND4_X1 U21183 ( .A1(n18079), .A2(n18078), .A3(n18077), .A4(n18076), .ZN(
        n18080) );
  NOR2_X1 U21184 ( .A1(n18081), .A2(n18080), .ZN(n18082) );
  XNOR2_X1 U21185 ( .A(n18083), .B(n18082), .ZN(n18403) );
  INV_X1 U21186 ( .A(n18084), .ZN(n18086) );
  OAI221_X1 U21187 ( .B1(P3_EBX_REG_30__SCAN_IN), .B2(n18086), .C1(n18085), 
        .C2(n18084), .A(n9564), .ZN(n18087) );
  OAI21_X1 U21188 ( .B1(n18403), .B2(n9564), .A(n18087), .ZN(P3_U2673) );
  NAND2_X1 U21189 ( .A1(n18089), .A2(n18088), .ZN(n18091) );
  XOR2_X1 U21190 ( .A(n18091), .B(n18090), .Z(n18407) );
  NAND3_X1 U21191 ( .A1(n18093), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n9564), .ZN(
        n18092) );
  OAI221_X1 U21192 ( .B1(n18093), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n9564), 
        .C2(n18407), .A(n18092), .ZN(P3_U2674) );
  AOI21_X1 U21193 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n9564), .A(n18101), .ZN(
        n18095) );
  XNOR2_X1 U21194 ( .A(n18094), .B(n18097), .ZN(n18416) );
  OAI22_X1 U21195 ( .A1(n18096), .A2(n18095), .B1(n9564), .B2(n18416), .ZN(
        P3_U2676) );
  AOI21_X1 U21196 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n9564), .A(n18105), .ZN(
        n18100) );
  OAI21_X1 U21197 ( .B1(n18099), .B2(n18098), .A(n18097), .ZN(n18420) );
  OAI22_X1 U21198 ( .A1(n18101), .A2(n18100), .B1(n9564), .B2(n18420), .ZN(
        P3_U2677) );
  AOI21_X1 U21199 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n9564), .A(n18102), .ZN(
        n18104) );
  XNOR2_X1 U21200 ( .A(n18103), .B(n18107), .ZN(n18425) );
  OAI22_X1 U21201 ( .A1(n18105), .A2(n18104), .B1(n9564), .B2(n18425), .ZN(
        P3_U2678) );
  NOR2_X1 U21202 ( .A1(n9658), .A2(n18106), .ZN(n18114) );
  AOI21_X1 U21203 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n9564), .A(n18114), .ZN(
        n18110) );
  OAI21_X1 U21204 ( .B1(n18109), .B2(n18108), .A(n18107), .ZN(n18430) );
  OAI22_X1 U21205 ( .A1(n18102), .A2(n18110), .B1(n9564), .B2(n18430), .ZN(
        P3_U2679) );
  INV_X1 U21206 ( .A(n9658), .ZN(n18131) );
  AOI21_X1 U21207 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n9564), .A(n18131), .ZN(
        n18113) );
  XNOR2_X1 U21208 ( .A(n18112), .B(n18111), .ZN(n18434) );
  OAI22_X1 U21209 ( .A1(n18114), .A2(n18113), .B1(n9564), .B2(n18434), .ZN(
        P3_U2680) );
  AOI21_X1 U21210 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n9564), .A(n18115), .ZN(
        n18130) );
  INV_X1 U21211 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18123) );
  INV_X1 U21212 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18116) );
  INV_X1 U21213 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18267) );
  OAI22_X1 U21214 ( .A1(n17408), .A2(n18116), .B1(n18321), .B2(n18267), .ZN(
        n18120) );
  INV_X1 U21215 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18118) );
  OAI22_X1 U21216 ( .A1(n18325), .A2(n18118), .B1(n11799), .B2(n18117), .ZN(
        n18119) );
  AOI211_X1 U21217 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n18120), .B(n18119), .ZN(n18122) );
  AOI22_X1 U21218 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9555), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18121) );
  OAI211_X1 U21219 ( .C1(n18218), .C2(n18123), .A(n18122), .B(n18121), .ZN(
        n18129) );
  AOI22_X1 U21220 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18127) );
  AOI22_X1 U21221 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18126) );
  AOI22_X1 U21222 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18125) );
  AOI22_X1 U21223 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9559), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18124) );
  NAND4_X1 U21224 ( .A1(n18127), .A2(n18126), .A3(n18125), .A4(n18124), .ZN(
        n18128) );
  NOR2_X1 U21225 ( .A1(n18129), .A2(n18128), .ZN(n18435) );
  OAI22_X1 U21226 ( .A1(n18131), .A2(n18130), .B1(n18435), .B2(n9564), .ZN(
        P3_U2681) );
  INV_X1 U21227 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18140) );
  INV_X1 U21228 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18132) );
  OAI22_X1 U21229 ( .A1(n11735), .A2(n18133), .B1(n11799), .B2(n18132), .ZN(
        n18137) );
  INV_X1 U21230 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18135) );
  OAI22_X1 U21231 ( .A1(n18327), .A2(n18135), .B1(n9567), .B2(n18134), .ZN(
        n18136) );
  AOI211_X1 U21232 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n18137), .B(n18136), .ZN(n18139) );
  AOI22_X1 U21233 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18138) );
  OAI211_X1 U21234 ( .C1(n18218), .C2(n18140), .A(n18139), .B(n18138), .ZN(
        n18146) );
  AOI22_X1 U21235 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18144) );
  AOI22_X1 U21236 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18143) );
  AOI22_X1 U21237 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18142) );
  AOI22_X1 U21238 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18141) );
  NAND4_X1 U21239 ( .A1(n18144), .A2(n18143), .A3(n18142), .A4(n18141), .ZN(
        n18145) );
  OR2_X1 U21240 ( .A1(n18146), .A2(n18145), .ZN(n18444) );
  NOR2_X1 U21241 ( .A1(n18385), .A2(n18147), .ZN(n18165) );
  AOI22_X1 U21242 ( .A1(n18385), .A2(n18444), .B1(P3_EBX_REG_21__SCAN_IN), 
        .B2(n18165), .ZN(n18148) );
  OAI21_X1 U21243 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18149), .A(n18148), .ZN(
        P3_U2682) );
  INV_X1 U21244 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18292) );
  AOI22_X1 U21245 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18150) );
  OAI21_X1 U21246 ( .B1(n11727), .B2(n18292), .A(n18150), .ZN(n18151) );
  AOI21_X1 U21247 ( .B1(n18345), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n18151), .ZN(n18154) );
  AOI22_X1 U21248 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18330), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18153) );
  AOI22_X1 U21249 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18152) );
  NAND3_X1 U21250 ( .A1(n18154), .A2(n18153), .A3(n18152), .ZN(n18163) );
  AOI22_X1 U21251 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18156) );
  NAND2_X1 U21252 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n18155) );
  OAI211_X1 U21253 ( .C1(n18157), .C2(n18323), .A(n18156), .B(n18155), .ZN(
        n18158) );
  INV_X1 U21254 ( .A(n18158), .ZN(n18161) );
  AOI22_X1 U21255 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18160) );
  AOI22_X1 U21256 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18159) );
  NAND3_X1 U21257 ( .A1(n18161), .A2(n18160), .A3(n18159), .ZN(n18162) );
  NOR2_X1 U21258 ( .A1(n18163), .A2(n18162), .ZN(n18448) );
  OAI21_X1 U21259 ( .B1(n18164), .B2(P3_EBX_REG_20__SCAN_IN), .A(n18165), .ZN(
        n18166) );
  OAI21_X1 U21260 ( .B1(n18448), .B2(n9564), .A(n18166), .ZN(P3_U2683) );
  AOI22_X1 U21261 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18167) );
  OAI21_X1 U21262 ( .B1(n11727), .B2(n18168), .A(n18167), .ZN(n18169) );
  AOI21_X1 U21263 ( .B1(n18345), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n18169), .ZN(n18173) );
  AOI22_X1 U21264 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18172) );
  AOI22_X1 U21265 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18171) );
  NAND3_X1 U21266 ( .A1(n18173), .A2(n18172), .A3(n18171), .ZN(n18182) );
  AOI22_X1 U21267 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18175) );
  NAND2_X1 U21268 ( .A1(n11628), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n18174) );
  OAI211_X1 U21269 ( .C1(n11623), .C2(n18302), .A(n18175), .B(n18174), .ZN(
        n18180) );
  INV_X1 U21270 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18176) );
  OAI22_X1 U21271 ( .A1(n18358), .A2(n18177), .B1(n18325), .B2(n18176), .ZN(
        n18179) );
  INV_X1 U21272 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18304) );
  INV_X1 U21273 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19156) );
  OAI22_X1 U21274 ( .A1(n18352), .A2(n18304), .B1(n18256), .B2(n19156), .ZN(
        n18178) );
  OR3_X1 U21275 ( .A1(n18180), .A2(n18179), .A3(n18178), .ZN(n18181) );
  NOR2_X1 U21276 ( .A1(n18182), .A2(n18181), .ZN(n18458) );
  INV_X1 U21277 ( .A(n18164), .ZN(n18183) );
  OAI21_X1 U21278 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18184), .A(n18183), .ZN(
        n18185) );
  AOI22_X1 U21279 ( .A1(n18385), .A2(n18458), .B1(n18185), .B2(n9564), .ZN(
        P3_U2684) );
  NAND2_X1 U21280 ( .A1(n9564), .A2(n18201), .ZN(n18225) );
  INV_X1 U21281 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18194) );
  INV_X1 U21282 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18187) );
  INV_X1 U21283 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18186) );
  OAI22_X1 U21284 ( .A1(n11735), .A2(n18187), .B1(n11799), .B2(n18186), .ZN(
        n18191) );
  INV_X1 U21285 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18189) );
  OAI22_X1 U21286 ( .A1(n18327), .A2(n18189), .B1(n9567), .B2(n18188), .ZN(
        n18190) );
  AOI211_X1 U21287 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n18191), .B(n18190), .ZN(n18193) );
  AOI22_X1 U21288 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18192) );
  OAI211_X1 U21289 ( .C1(n18218), .C2(n18194), .A(n18193), .B(n18192), .ZN(
        n18200) );
  AOI22_X1 U21290 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18198) );
  AOI22_X1 U21291 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18197) );
  AOI22_X1 U21292 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18196) );
  AOI22_X1 U21293 ( .A1(n9559), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18195) );
  NAND4_X1 U21294 ( .A1(n18198), .A2(n18197), .A3(n18196), .A4(n18195), .ZN(
        n18199) );
  OR2_X1 U21295 ( .A1(n18200), .A2(n18199), .ZN(n18459) );
  NOR3_X1 U21296 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18201), .A3(n19171), .ZN(
        n18202) );
  AOI21_X1 U21297 ( .B1(n18385), .B2(n18459), .A(n18202), .ZN(n18203) );
  OAI21_X1 U21298 ( .B1(n18204), .B2(n18225), .A(n18203), .ZN(P3_U2685) );
  NOR2_X1 U21299 ( .A1(n18205), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n18226) );
  NOR2_X1 U21300 ( .A1(n11623), .A2(n18206), .ZN(n18209) );
  INV_X1 U21301 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18357) );
  OAI22_X1 U21302 ( .A1(n18327), .A2(n18357), .B1(n9567), .B2(n18207), .ZN(
        n18208) );
  AOI211_X1 U21303 ( .C1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .C2(n18170), .A(
        n18209), .B(n18208), .ZN(n18212) );
  AOI22_X1 U21304 ( .A1(n9582), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18211) );
  AOI22_X1 U21305 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11628), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18210) );
  NAND3_X1 U21306 ( .A1(n18212), .A2(n18211), .A3(n18210), .ZN(n18224) );
  INV_X1 U21307 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19148) );
  NOR2_X1 U21308 ( .A1(n18256), .A2(n19148), .ZN(n18216) );
  OAI22_X1 U21309 ( .A1(n18358), .A2(n18343), .B1(n9557), .B2(n18213), .ZN(
        n18215) );
  AOI211_X1 U21310 ( .C1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .C2(n9561), .A(
        n18216), .B(n18215), .ZN(n18222) );
  AOI22_X1 U21311 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18221) );
  NAND2_X1 U21312 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n18220) );
  INV_X1 U21313 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18217) );
  OR2_X1 U21314 ( .A1(n18218), .A2(n18217), .ZN(n18219) );
  NAND4_X1 U21315 ( .A1(n18222), .A2(n18221), .A3(n18220), .A4(n18219), .ZN(
        n18223) );
  NOR2_X1 U21316 ( .A1(n18224), .A2(n18223), .ZN(n18468) );
  OAI22_X1 U21317 ( .A1(n18226), .A2(n18225), .B1(n18468), .B2(n9564), .ZN(
        P3_U2686) );
  INV_X1 U21318 ( .A(n18263), .ZN(n18227) );
  OAI21_X1 U21319 ( .B1(n18227), .B2(P3_EBX_REG_16__SCAN_IN), .A(n9564), .ZN(
        n18242) );
  OAI22_X1 U21320 ( .A1(n18325), .A2(n18229), .B1(n18253), .B2(n18228), .ZN(
        n18232) );
  INV_X1 U21321 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18230) );
  OAI22_X1 U21322 ( .A1(n18327), .A2(n21672), .B1(n11735), .B2(n18230), .ZN(
        n18231) );
  AOI211_X1 U21323 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n18232), .B(n18231), .ZN(n18234) );
  AOI22_X1 U21324 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18233) );
  OAI211_X1 U21325 ( .C1(n18218), .C2(n18235), .A(n18234), .B(n18233), .ZN(
        n18241) );
  AOI22_X1 U21326 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18239) );
  AOI22_X1 U21327 ( .A1(n9556), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18238) );
  AOI22_X1 U21328 ( .A1(n11684), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U21329 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11628), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18236) );
  NAND4_X1 U21330 ( .A1(n18239), .A2(n18238), .A3(n18237), .A4(n18236), .ZN(
        n18240) );
  NOR2_X1 U21331 ( .A1(n18241), .A2(n18240), .ZN(n18474) );
  OAI22_X1 U21332 ( .A1(n18205), .A2(n18242), .B1(n18474), .B2(n9564), .ZN(
        P3_U2687) );
  INV_X1 U21333 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18244) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18054), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18243) );
  OAI21_X1 U21335 ( .B1(n18244), .B2(n11727), .A(n18243), .ZN(n18245) );
  AOI21_X1 U21336 ( .B1(n9560), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(n18245), .ZN(n18248) );
  AOI22_X1 U21337 ( .A1(n17450), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18247) );
  AOI22_X1 U21338 ( .A1(n9556), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18246) );
  NAND3_X1 U21339 ( .A1(n18248), .A2(n18247), .A3(n18246), .ZN(n18262) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17461), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18250) );
  NAND2_X1 U21341 ( .A1(n18345), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n18249) );
  OAI211_X1 U21342 ( .C1(n18251), .C2(n18323), .A(n18250), .B(n18249), .ZN(
        n18260) );
  INV_X1 U21343 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18254) );
  OAI22_X1 U21344 ( .A1(n18358), .A2(n18254), .B1(n18253), .B2(n18252), .ZN(
        n18259) );
  INV_X1 U21345 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18257) );
  OAI22_X1 U21346 ( .A1(n18352), .A2(n18257), .B1(n18256), .B2(n18255), .ZN(
        n18258) );
  OR3_X1 U21347 ( .A1(n18260), .A2(n18259), .A3(n18258), .ZN(n18261) );
  NOR2_X1 U21348 ( .A1(n18262), .A2(n18261), .ZN(n18478) );
  OAI21_X1 U21349 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n18264), .A(n18263), .ZN(
        n18265) );
  AOI22_X1 U21350 ( .A1(n18385), .A2(n18478), .B1(n18265), .B2(n9564), .ZN(
        P3_U2688) );
  NAND2_X1 U21351 ( .A1(n9564), .A2(n18280), .ZN(n18283) );
  INV_X1 U21352 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19170) );
  INV_X1 U21353 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18266) );
  OAI22_X1 U21354 ( .A1(n11735), .A2(n18267), .B1(n11799), .B2(n18266), .ZN(
        n18271) );
  INV_X1 U21355 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18269) );
  INV_X1 U21356 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18268) );
  OAI22_X1 U21357 ( .A1(n18327), .A2(n18269), .B1(n9567), .B2(n18268), .ZN(
        n18270) );
  AOI211_X1 U21358 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n18271), .B(n18270), .ZN(n18273) );
  AOI22_X1 U21359 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18272) );
  OAI211_X1 U21360 ( .C1(n19170), .C2(n18218), .A(n18273), .B(n18272), .ZN(
        n18279) );
  AOI22_X1 U21361 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18277) );
  AOI22_X1 U21362 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18276) );
  AOI22_X1 U21363 ( .A1(n9582), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U21364 ( .A1(n11628), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18274) );
  NAND4_X1 U21365 ( .A1(n18277), .A2(n18276), .A3(n18275), .A4(n18274), .ZN(
        n18278) );
  OR2_X1 U21366 ( .A1(n18279), .A2(n18278), .ZN(n18481) );
  NOR3_X1 U21367 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18280), .A3(n19171), .ZN(
        n18281) );
  AOI21_X1 U21368 ( .B1(n18385), .B2(n18481), .A(n18281), .ZN(n18282) );
  OAI21_X1 U21369 ( .B1(n18284), .B2(n18283), .A(n18282), .ZN(P3_U2689) );
  OAI21_X1 U21370 ( .B1(n18317), .B2(P3_EBX_REG_12__SCAN_IN), .A(n9564), .ZN(
        n18300) );
  INV_X1 U21371 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18286) );
  AOI22_X1 U21372 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9582), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18285) );
  OAI21_X1 U21373 ( .B1(n18352), .B2(n18286), .A(n18285), .ZN(n18287) );
  AOI21_X1 U21374 ( .B1(n9560), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(n18287), .ZN(n18290) );
  AOI22_X1 U21375 ( .A1(n11606), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18289) );
  AOI22_X1 U21376 ( .A1(n18334), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11628), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18288) );
  NAND3_X1 U21377 ( .A1(n18290), .A2(n18289), .A3(n18288), .ZN(n18299) );
  AOI22_X1 U21378 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18291) );
  OAI21_X1 U21379 ( .B1(n17408), .B2(n18292), .A(n18291), .ZN(n18293) );
  AOI21_X1 U21380 ( .B1(n18345), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n18293), .ZN(n18297) );
  AOI22_X1 U21381 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U21382 ( .A1(n11784), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9555), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18295) );
  NAND3_X1 U21383 ( .A1(n18297), .A2(n18296), .A3(n18295), .ZN(n18298) );
  NOR2_X1 U21384 ( .A1(n18299), .A2(n18298), .ZN(n18491) );
  OAI22_X1 U21385 ( .A1(n18301), .A2(n18300), .B1(n18491), .B2(n9564), .ZN(
        P3_U2691) );
  OAI22_X1 U21386 ( .A1(n18325), .A2(n18303), .B1(n11799), .B2(n18302), .ZN(
        n18307) );
  INV_X1 U21387 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18305) );
  OAI22_X1 U21388 ( .A1(n11735), .A2(n18305), .B1(n9567), .B2(n18304), .ZN(
        n18306) );
  AOI211_X1 U21389 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n18307), .B(n18306), .ZN(n18309) );
  AOI22_X1 U21390 ( .A1(n11606), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9559), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18308) );
  OAI211_X1 U21391 ( .C1(n18218), .C2(n19156), .A(n18309), .B(n18308), .ZN(
        n18315) );
  AOI22_X1 U21392 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11784), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18313) );
  AOI22_X1 U21393 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9561), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U21394 ( .A1(n9555), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18311) );
  AOI22_X1 U21395 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18170), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18310) );
  NAND4_X1 U21396 ( .A1(n18313), .A2(n18312), .A3(n18311), .A4(n18310), .ZN(
        n18314) );
  NOR2_X1 U21397 ( .A1(n18315), .A2(n18314), .ZN(n18495) );
  INV_X1 U21398 ( .A(n18317), .ZN(n18318) );
  OAI21_X1 U21399 ( .B1(n18316), .B2(P3_EBX_REG_11__SCAN_IN), .A(n18318), .ZN(
        n18319) );
  AOI22_X1 U21400 ( .A1(n18385), .A2(n18495), .B1(n18319), .B2(n9564), .ZN(
        P3_U2692) );
  OAI21_X1 U21401 ( .B1(n18364), .B2(P3_EBX_REG_10__SCAN_IN), .A(n9564), .ZN(
        n18341) );
  INV_X1 U21402 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18333) );
  INV_X1 U21403 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18322) );
  INV_X1 U21404 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18320) );
  OAI22_X1 U21405 ( .A1(n18323), .A2(n18322), .B1(n18321), .B2(n18320), .ZN(
        n18329) );
  INV_X1 U21406 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18326) );
  OAI22_X1 U21407 ( .A1(n18327), .A2(n18326), .B1(n18325), .B2(n18324), .ZN(
        n18328) );
  AOI211_X1 U21408 ( .C1(n9560), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n18329), .B(n18328), .ZN(n18332) );
  AOI22_X1 U21409 ( .A1(n18330), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9556), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18331) );
  OAI211_X1 U21410 ( .C1(n18218), .C2(n18333), .A(n18332), .B(n18331), .ZN(
        n18340) );
  AOI22_X1 U21411 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18338) );
  AOI22_X1 U21412 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18337) );
  AOI22_X1 U21413 ( .A1(n9561), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18334), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18336) );
  AOI22_X1 U21414 ( .A1(n18349), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18335) );
  NAND4_X1 U21415 ( .A1(n18338), .A2(n18337), .A3(n18336), .A4(n18335), .ZN(
        n18339) );
  NOR2_X1 U21416 ( .A1(n18340), .A2(n18339), .ZN(n18499) );
  OAI22_X1 U21417 ( .A1(n18316), .A2(n18341), .B1(n18499), .B2(n9564), .ZN(
        P3_U2693) );
  AOI22_X1 U21418 ( .A1(n18054), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18342) );
  OAI21_X1 U21419 ( .B1(n18321), .B2(n18343), .A(n18342), .ZN(n18344) );
  AOI21_X1 U21420 ( .B1(n18345), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n18344), .ZN(n18348) );
  AOI22_X1 U21421 ( .A1(n9582), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11628), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18347) );
  AOI22_X1 U21422 ( .A1(n9556), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11606), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18346) );
  NAND3_X1 U21423 ( .A1(n18348), .A2(n18347), .A3(n18346), .ZN(n18363) );
  INV_X1 U21424 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18353) );
  AOI22_X1 U21425 ( .A1(n17461), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18349), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18351) );
  NAND2_X1 U21426 ( .A1(n9560), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n18350) );
  OAI211_X1 U21427 ( .C1(n18353), .C2(n18352), .A(n18351), .B(n18350), .ZN(
        n18361) );
  OAI22_X1 U21428 ( .A1(n17408), .A2(n18355), .B1(n18256), .B2(n18354), .ZN(
        n18360) );
  INV_X1 U21429 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18356) );
  OAI22_X1 U21430 ( .A1(n18358), .A2(n18357), .B1(n11727), .B2(n18356), .ZN(
        n18359) );
  OR3_X1 U21431 ( .A1(n18361), .A2(n18360), .A3(n18359), .ZN(n18362) );
  NOR2_X1 U21432 ( .A1(n18363), .A2(n18362), .ZN(n18504) );
  INV_X1 U21433 ( .A(n18364), .ZN(n18365) );
  OAI21_X1 U21434 ( .B1(n18366), .B2(P3_EBX_REG_9__SCAN_IN), .A(n18365), .ZN(
        n18367) );
  AOI22_X1 U21435 ( .A1(n18385), .A2(n18504), .B1(n18367), .B2(n9564), .ZN(
        P3_U2694) );
  NAND2_X1 U21436 ( .A1(n9564), .A2(n18368), .ZN(n18374) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18385), .B1(
        n18369), .B2(n18371), .ZN(n18370) );
  OAI21_X1 U21438 ( .B1(n18371), .B2(n18374), .A(n18370), .ZN(P3_U2696) );
  AND2_X1 U21439 ( .A1(n18373), .A2(n18372), .ZN(n18375) );
  OAI22_X1 U21440 ( .A1(n18375), .A2(n18374), .B1(n19170), .B2(n9564), .ZN(
        P3_U2697) );
  INV_X1 U21441 ( .A(n18376), .ZN(n18377) );
  OAI21_X1 U21442 ( .B1(n18377), .B2(P3_EBX_REG_5__SCAN_IN), .A(n9564), .ZN(
        n18378) );
  OAI22_X1 U21443 ( .A1(n14713), .A2(n18378), .B1(n19165), .B2(n9564), .ZN(
        P3_U2698) );
  INV_X1 U21444 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19160) );
  OAI21_X1 U21445 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18379), .A(n18376), .ZN(
        n18380) );
  AOI22_X1 U21446 ( .A1(n18385), .A2(n19160), .B1(n18380), .B2(n9564), .ZN(
        P3_U2699) );
  OAI21_X1 U21447 ( .B1(n10227), .B2(P3_EBX_REG_3__SCAN_IN), .A(n9564), .ZN(
        n18382) );
  OAI22_X1 U21448 ( .A1(n18379), .A2(n18382), .B1(n19156), .B2(n9564), .ZN(
        P3_U2700) );
  OAI21_X1 U21449 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n18383), .A(n18381), .ZN(
        n18384) );
  AOI22_X1 U21450 ( .A1(n18385), .A2(n18333), .B1(n18384), .B2(n9564), .ZN(
        P3_U2701) );
  OAI221_X1 U21451 ( .B1(n11836), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .C1(
        n19171), .C2(n18386), .A(n18389), .ZN(n18387) );
  OAI21_X1 U21452 ( .B1(n18389), .B2(n18388), .A(n18387), .ZN(P3_U2702) );
  INV_X1 U21453 ( .A(n18389), .ZN(n18390) );
  NOR2_X1 U21454 ( .A1(n19171), .A2(n18390), .ZN(n18392) );
  OAI21_X1 U21455 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18392), .A(n18391), .ZN(
        n18393) );
  OAI21_X1 U21456 ( .B1(n9564), .B2(n14698), .A(n18393), .ZN(P3_U2703) );
  INV_X1 U21457 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18600) );
  INV_X1 U21458 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18596) );
  INV_X1 U21459 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18591) );
  NAND2_X1 U21460 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n18514) );
  NAND4_X1 U21461 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n18394) );
  NOR4_X1 U21462 ( .A1(n18514), .A2(n18608), .A3(n18606), .A4(n18394), .ZN(
        n18513) );
  INV_X1 U21463 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18630) );
  INV_X1 U21464 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18628) );
  INV_X1 U21465 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18642) );
  AND4_X1 U21466 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n18437)
         );
  NAND2_X1 U21467 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18437), .ZN(n18443) );
  NAND2_X1 U21468 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18408), .ZN(n18404) );
  INV_X1 U21469 ( .A(n18404), .ZN(n18400) );
  NAND2_X1 U21470 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18400), .ZN(n18399) );
  NAND2_X1 U21471 ( .A1(n18399), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n18398) );
  NAND2_X1 U21472 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18469), .ZN(n18397) );
  OAI221_X1 U21473 ( .B1(n18399), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n18398), 
        .C2(n18533), .A(n18397), .ZN(P3_U2704) );
  AOI22_X1 U21474 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18469), .ZN(n18402) );
  OAI211_X1 U21475 ( .C1(n18400), .C2(P3_EAX_REG_30__SCAN_IN), .A(n18522), .B(
        n18399), .ZN(n18401) );
  OAI211_X1 U21476 ( .C1(n18403), .C2(n18525), .A(n18402), .B(n18401), .ZN(
        P3_U2705) );
  AOI22_X1 U21477 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18469), .ZN(n18406) );
  OAI211_X1 U21478 ( .C1(n18408), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18522), .B(
        n18404), .ZN(n18405) );
  OAI211_X1 U21479 ( .C1(n18525), .C2(n18407), .A(n18406), .B(n18405), .ZN(
        P3_U2706) );
  AOI22_X1 U21480 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18469), .ZN(n18411) );
  AOI211_X1 U21481 ( .C1(n18600), .C2(n18413), .A(n18408), .B(n18533), .ZN(
        n18409) );
  INV_X1 U21482 ( .A(n18409), .ZN(n18410) );
  OAI211_X1 U21483 ( .C1(n18525), .C2(n18412), .A(n18411), .B(n18410), .ZN(
        P3_U2707) );
  AOI22_X1 U21484 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18469), .ZN(n18415) );
  OAI211_X1 U21485 ( .C1(n9715), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18522), .B(
        n18413), .ZN(n18414) );
  OAI211_X1 U21486 ( .C1(n18525), .C2(n18416), .A(n18415), .B(n18414), .ZN(
        P3_U2708) );
  AOI22_X1 U21487 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18469), .ZN(n18419) );
  AOI211_X1 U21488 ( .C1(n18596), .C2(n18421), .A(n9715), .B(n18533), .ZN(
        n18417) );
  INV_X1 U21489 ( .A(n18417), .ZN(n18418) );
  OAI211_X1 U21490 ( .C1(n18525), .C2(n18420), .A(n18419), .B(n18418), .ZN(
        P3_U2709) );
  AOI22_X1 U21491 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18469), .ZN(n18424) );
  OAI211_X1 U21492 ( .C1(n18422), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18522), .B(
        n18421), .ZN(n18423) );
  OAI211_X1 U21493 ( .C1(n18525), .C2(n18425), .A(n18424), .B(n18423), .ZN(
        P3_U2710) );
  AOI22_X1 U21494 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18469), .ZN(n18429) );
  OAI211_X1 U21495 ( .C1(n18427), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18522), .B(
        n18426), .ZN(n18428) );
  OAI211_X1 U21496 ( .C1(n18525), .C2(n18430), .A(n18429), .B(n18428), .ZN(
        P3_U2711) );
  AOI22_X1 U21497 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18469), .ZN(n18433) );
  OAI211_X1 U21498 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n9729), .A(n18522), .B(
        n18431), .ZN(n18432) );
  OAI211_X1 U21499 ( .C1(n18525), .C2(n18434), .A(n18433), .B(n18432), .ZN(
        P3_U2712) );
  NAND2_X1 U21500 ( .A1(n18465), .A2(n18591), .ZN(n18442) );
  INV_X1 U21501 ( .A(n18435), .ZN(n18436) );
  AOI22_X1 U21502 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18469), .B1(n18530), .B2(
        n18436), .ZN(n18441) );
  NAND2_X1 U21503 ( .A1(n18437), .A2(n18465), .ZN(n18450) );
  NAND2_X1 U21504 ( .A1(n18522), .A2(n18450), .ZN(n18454) );
  OAI21_X1 U21505 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18438), .A(n18454), .ZN(
        n18439) );
  AOI22_X1 U21506 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18470), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n18439), .ZN(n18440) );
  OAI211_X1 U21507 ( .C1(n18443), .C2(n18442), .A(n18441), .B(n18440), .ZN(
        P3_U2713) );
  AOI22_X1 U21508 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18469), .B1(n18530), .B2(
        n18444), .ZN(n18447) );
  INV_X1 U21509 ( .A(n18454), .ZN(n18445) );
  AOI22_X1 U21510 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18470), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n18445), .ZN(n18446) );
  OAI211_X1 U21511 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n18450), .A(n18447), .B(
        n18446), .ZN(P3_U2714) );
  INV_X1 U21512 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18587) );
  INV_X1 U21513 ( .A(n18448), .ZN(n18449) );
  AOI22_X1 U21514 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18470), .B1(n18530), .B2(
        n18449), .ZN(n18453) );
  NAND2_X1 U21515 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18463), .ZN(n18455) );
  INV_X1 U21516 ( .A(n18455), .ZN(n18451) );
  AOI22_X1 U21517 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18469), .B1(n18451), .B2(
        n18450), .ZN(n18452) );
  OAI211_X1 U21518 ( .C1(n18587), .C2(n18454), .A(n18453), .B(n18452), .ZN(
        P3_U2715) );
  AOI22_X1 U21519 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18469), .ZN(n18457) );
  OAI211_X1 U21520 ( .C1(n18463), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18522), .B(
        n18455), .ZN(n18456) );
  OAI211_X1 U21521 ( .C1(n18458), .C2(n18525), .A(n18457), .B(n18456), .ZN(
        P3_U2716) );
  AOI22_X1 U21522 ( .A1(n18465), .A2(P3_EAX_REG_17__SCAN_IN), .B1(
        P3_EAX_REG_18__SCAN_IN), .B2(n18522), .ZN(n18462) );
  AOI22_X1 U21523 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n18469), .B1(n18530), .B2(
        n18459), .ZN(n18461) );
  NAND2_X1 U21524 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18470), .ZN(n18460) );
  OAI211_X1 U21525 ( .C1(n18463), .C2(n18462), .A(n18461), .B(n18460), .ZN(
        P3_U2717) );
  AOI22_X1 U21526 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18469), .ZN(n18467) );
  NAND2_X1 U21527 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n18465), .ZN(n18464) );
  OAI211_X1 U21528 ( .C1(n18465), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18522), .B(
        n18464), .ZN(n18466) );
  OAI211_X1 U21529 ( .C1(n18468), .C2(n18525), .A(n18467), .B(n18466), .ZN(
        P3_U2718) );
  AOI22_X1 U21530 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18470), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18469), .ZN(n18473) );
  OAI211_X1 U21531 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18475), .A(n18522), .B(
        n18471), .ZN(n18472) );
  OAI211_X1 U21532 ( .C1(n18474), .C2(n18525), .A(n18473), .B(n18472), .ZN(
        P3_U2719) );
  AOI211_X1 U21533 ( .C1(n18642), .C2(n18479), .A(n18533), .B(n18475), .ZN(
        n18476) );
  AOI21_X1 U21534 ( .B1(n18531), .B2(BUF2_REG_15__SCAN_IN), .A(n18476), .ZN(
        n18477) );
  OAI21_X1 U21535 ( .B1(n18478), .B2(n18525), .A(n18477), .ZN(P3_U2720) );
  INV_X1 U21536 ( .A(n18479), .ZN(n18484) );
  AOI22_X1 U21537 ( .A1(n11836), .A2(n18480), .B1(P3_EAX_REG_14__SCAN_IN), 
        .B2(n18522), .ZN(n18483) );
  AOI22_X1 U21538 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18531), .B1(n18530), .B2(
        n18481), .ZN(n18482) );
  OAI21_X1 U21539 ( .B1(n18484), .B2(n18483), .A(n18482), .ZN(P3_U2721) );
  INV_X1 U21540 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18626) );
  NAND3_X1 U21541 ( .A1(n18513), .A2(P3_EAX_REG_8__SCAN_IN), .A3(n18512), .ZN(
        n18503) );
  NOR2_X1 U21542 ( .A1(n18626), .A2(n18503), .ZN(n18506) );
  NAND2_X1 U21543 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18506), .ZN(n18498) );
  NOR2_X1 U21544 ( .A1(n18630), .A2(n18498), .ZN(n18490) );
  NAND2_X1 U21545 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18490), .ZN(n18489) );
  NAND2_X1 U21546 ( .A1(n18489), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n18488) );
  INV_X1 U21547 ( .A(n18485), .ZN(n18486) );
  AOI22_X1 U21548 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18531), .B1(n18530), .B2(
        n18486), .ZN(n18487) );
  OAI221_X1 U21549 ( .B1(n18489), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n18488), 
        .C2(n18533), .A(n18487), .ZN(P3_U2722) );
  INV_X1 U21550 ( .A(n18489), .ZN(n18493) );
  AOI21_X1 U21551 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18522), .A(n18490), .ZN(
        n18492) );
  OAI222_X1 U21552 ( .A1(n18528), .A2(n18494), .B1(n18493), .B2(n18492), .C1(
        n18525), .C2(n18491), .ZN(P3_U2723) );
  NAND2_X1 U21553 ( .A1(n18522), .A2(n18498), .ZN(n18501) );
  INV_X1 U21554 ( .A(n18495), .ZN(n18496) );
  AOI22_X1 U21555 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18531), .B1(n18530), .B2(
        n18496), .ZN(n18497) );
  OAI221_X1 U21556 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18498), .C1(n18630), 
        .C2(n18501), .A(n18497), .ZN(P3_U2724) );
  NOR2_X1 U21557 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18506), .ZN(n18500) );
  OAI222_X1 U21558 ( .A1(n18528), .A2(n18502), .B1(n18501), .B2(n18500), .C1(
        n18525), .C2(n18499), .ZN(P3_U2725) );
  INV_X1 U21559 ( .A(n18503), .ZN(n18507) );
  AOI21_X1 U21560 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18522), .A(n18507), .ZN(
        n18505) );
  OAI222_X1 U21561 ( .A1(n18528), .A2(n13851), .B1(n18506), .B2(n18505), .C1(
        n18525), .C2(n18504), .ZN(P3_U2726) );
  INV_X1 U21562 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18624) );
  AOI211_X1 U21563 ( .C1(n18508), .C2(n18624), .A(n18533), .B(n18507), .ZN(
        n18509) );
  AOI21_X1 U21564 ( .B1(n18531), .B2(BUF2_REG_8__SCAN_IN), .A(n18509), .ZN(
        n18510) );
  OAI21_X1 U21565 ( .B1(n18511), .B2(n18525), .A(n18510), .ZN(P3_U2727) );
  AND2_X1 U21566 ( .A1(n18513), .A2(n18512), .ZN(n18517) );
  NOR2_X1 U21567 ( .A1(n18514), .A2(n18535), .ZN(n18527) );
  AOI22_X1 U21568 ( .A1(n18527), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n18522), .ZN(n18516) );
  OAI222_X1 U21569 ( .A1(n18528), .A2(n13838), .B1(n18517), .B2(n18516), .C1(
        n18525), .C2(n18515), .ZN(P3_U2728) );
  INV_X1 U21570 ( .A(n18527), .ZN(n18521) );
  NAND2_X1 U21571 ( .A1(n18521), .A2(P3_EAX_REG_6__SCAN_IN), .ZN(n18520) );
  AOI22_X1 U21572 ( .A1(n18531), .A2(BUF2_REG_6__SCAN_IN), .B1(n18530), .B2(
        n18518), .ZN(n18519) );
  OAI221_X1 U21573 ( .B1(n18521), .B2(P3_EAX_REG_6__SCAN_IN), .C1(n18520), 
        .C2(n18533), .A(n18519), .ZN(P3_U2729) );
  AOI22_X1 U21574 ( .A1(n18523), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n18522), .ZN(n18526) );
  OAI222_X1 U21575 ( .A1(n13896), .A2(n18528), .B1(n18527), .B2(n18526), .C1(
        n18525), .C2(n18524), .ZN(P3_U2730) );
  NAND2_X1 U21576 ( .A1(n18535), .A2(P3_EAX_REG_4__SCAN_IN), .ZN(n18534) );
  AOI22_X1 U21577 ( .A1(n18531), .A2(BUF2_REG_4__SCAN_IN), .B1(n18530), .B2(
        n18529), .ZN(n18532) );
  OAI221_X1 U21578 ( .B1(n18535), .B2(P3_EAX_REG_4__SCAN_IN), .C1(n18534), 
        .C2(n18533), .A(n18532), .ZN(P3_U2731) );
  NOR2_X4 U21579 ( .A1(n18573), .A2(n18565), .ZN(n18567) );
  AND2_X1 U21580 ( .A1(n18567), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U21581 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18604) );
  NAND2_X1 U21582 ( .A1(n18565), .A2(n18538), .ZN(n18555) );
  AOI22_X1 U21583 ( .A1(n18573), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18539) );
  OAI21_X1 U21584 ( .B1(n18604), .B2(n18555), .A(n18539), .ZN(P3_U2737) );
  INV_X1 U21585 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18602) );
  AOI22_X1 U21586 ( .A1(n18573), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18540) );
  OAI21_X1 U21587 ( .B1(n18602), .B2(n18555), .A(n18540), .ZN(P3_U2738) );
  AOI22_X1 U21588 ( .A1(n18573), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18541) );
  OAI21_X1 U21589 ( .B1(n18600), .B2(n18555), .A(n18541), .ZN(P3_U2739) );
  INV_X1 U21590 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18598) );
  AOI22_X1 U21591 ( .A1(n18573), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18542) );
  OAI21_X1 U21592 ( .B1(n18598), .B2(n18555), .A(n18542), .ZN(P3_U2740) );
  INV_X2 U21593 ( .A(n19744), .ZN(n18573) );
  AOI22_X1 U21594 ( .A1(n18573), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18543) );
  OAI21_X1 U21595 ( .B1(n18596), .B2(n18555), .A(n18543), .ZN(P3_U2741) );
  AOI22_X1 U21596 ( .A1(n18573), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18544) );
  OAI21_X1 U21597 ( .B1(n10061), .B2(n18555), .A(n18544), .ZN(P3_U2742) );
  INV_X1 U21598 ( .A(P3_UWORD_REG_8__SCAN_IN), .ZN(n21643) );
  INV_X1 U21599 ( .A(n18555), .ZN(n18551) );
  AOI22_X1 U21600 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18551), .B1(n18567), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18545) );
  OAI21_X1 U21601 ( .B1(n19744), .B2(n21643), .A(n18545), .ZN(P3_U2743) );
  AOI22_X1 U21602 ( .A1(n18573), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18546) );
  OAI21_X1 U21603 ( .B1(n10059), .B2(n18555), .A(n18546), .ZN(P3_U2744) );
  AOI22_X1 U21604 ( .A1(n18573), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18547) );
  OAI21_X1 U21605 ( .B1(n18591), .B2(n18555), .A(n18547), .ZN(P3_U2745) );
  INV_X1 U21606 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18589) );
  AOI22_X1 U21607 ( .A1(n18573), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18548) );
  OAI21_X1 U21608 ( .B1(n18589), .B2(n18555), .A(n18548), .ZN(P3_U2746) );
  AOI22_X1 U21609 ( .A1(n18573), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18549) );
  OAI21_X1 U21610 ( .B1(n18587), .B2(n18555), .A(n18549), .ZN(P3_U2747) );
  INV_X1 U21611 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18585) );
  AOI22_X1 U21612 ( .A1(n18573), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18550) );
  OAI21_X1 U21613 ( .B1(n18585), .B2(n18555), .A(n18550), .ZN(P3_U2748) );
  INV_X1 U21614 ( .A(P3_UWORD_REG_2__SCAN_IN), .ZN(n21626) );
  AOI22_X1 U21615 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18551), .B1(n18567), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18552) );
  OAI21_X1 U21616 ( .B1(n19744), .B2(n21626), .A(n18552), .ZN(P3_U2749) );
  INV_X1 U21617 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18582) );
  AOI22_X1 U21618 ( .A1(n18573), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18553) );
  OAI21_X1 U21619 ( .B1(n18582), .B2(n18555), .A(n18553), .ZN(P3_U2750) );
  INV_X1 U21620 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18580) );
  AOI22_X1 U21621 ( .A1(n18573), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18554) );
  OAI21_X1 U21622 ( .B1(n18580), .B2(n18555), .A(n18554), .ZN(P3_U2751) );
  AOI22_X1 U21623 ( .A1(n18573), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18556) );
  OAI21_X1 U21624 ( .B1(n18642), .B2(n18575), .A(n18556), .ZN(P3_U2752) );
  INV_X1 U21625 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18637) );
  AOI22_X1 U21626 ( .A1(n18573), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18557) );
  OAI21_X1 U21627 ( .B1(n18637), .B2(n18575), .A(n18557), .ZN(P3_U2753) );
  INV_X1 U21628 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18635) );
  AOI22_X1 U21629 ( .A1(n18573), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18558) );
  OAI21_X1 U21630 ( .B1(n18635), .B2(n18575), .A(n18558), .ZN(P3_U2754) );
  INV_X1 U21631 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18632) );
  AOI22_X1 U21632 ( .A1(n18573), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18559) );
  OAI21_X1 U21633 ( .B1(n18632), .B2(n18575), .A(n18559), .ZN(P3_U2755) );
  AOI22_X1 U21634 ( .A1(n18573), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18560) );
  OAI21_X1 U21635 ( .B1(n18630), .B2(n18575), .A(n18560), .ZN(P3_U2756) );
  AOI22_X1 U21636 ( .A1(n18573), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18561) );
  OAI21_X1 U21637 ( .B1(n18628), .B2(n18575), .A(n18561), .ZN(P3_U2757) );
  AOI22_X1 U21638 ( .A1(n18573), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18562) );
  OAI21_X1 U21639 ( .B1(n18626), .B2(n18575), .A(n18562), .ZN(P3_U2758) );
  AOI22_X1 U21640 ( .A1(n18573), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18563) );
  OAI21_X1 U21641 ( .B1(n18624), .B2(n18575), .A(n18563), .ZN(P3_U2759) );
  INV_X1 U21642 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18621) );
  AOI22_X1 U21643 ( .A1(n18573), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18564) );
  OAI21_X1 U21644 ( .B1(n18621), .B2(n18575), .A(n18564), .ZN(P3_U2760) );
  INV_X1 U21645 ( .A(P3_LWORD_REG_6__SCAN_IN), .ZN(n21592) );
  AOI22_X1 U21646 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18565), .B1(n18567), .B2(
        P3_DATAO_REG_6__SCAN_IN), .ZN(n18566) );
  OAI21_X1 U21647 ( .B1(n19744), .B2(n21592), .A(n18566), .ZN(P3_U2761) );
  INV_X1 U21648 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18616) );
  AOI22_X1 U21649 ( .A1(n18573), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18568) );
  OAI21_X1 U21650 ( .B1(n18616), .B2(n18575), .A(n18568), .ZN(P3_U2762) );
  INV_X1 U21651 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18614) );
  AOI22_X1 U21652 ( .A1(n18573), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18569) );
  OAI21_X1 U21653 ( .B1(n18614), .B2(n18575), .A(n18569), .ZN(P3_U2763) );
  INV_X1 U21654 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18612) );
  AOI22_X1 U21655 ( .A1(n18573), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18570) );
  OAI21_X1 U21656 ( .B1(n18612), .B2(n18575), .A(n18570), .ZN(P3_U2764) );
  INV_X1 U21657 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18610) );
  AOI22_X1 U21658 ( .A1(n18573), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18571) );
  OAI21_X1 U21659 ( .B1(n18610), .B2(n18575), .A(n18571), .ZN(P3_U2765) );
  AOI22_X1 U21660 ( .A1(n18573), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18572) );
  OAI21_X1 U21661 ( .B1(n18608), .B2(n18575), .A(n18572), .ZN(P3_U2766) );
  AOI22_X1 U21662 ( .A1(n18573), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18567), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18574) );
  OAI21_X1 U21663 ( .B1(n18606), .B2(n18575), .A(n18574), .ZN(P3_U2767) );
  AOI22_X1 U21664 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18639), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18638), .ZN(n18579) );
  OAI21_X1 U21665 ( .B1(n18580), .B2(n18641), .A(n18579), .ZN(P3_U2768) );
  AOI22_X1 U21666 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18639), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18638), .ZN(n18581) );
  OAI21_X1 U21667 ( .B1(n18582), .B2(n18641), .A(n18581), .ZN(P3_U2769) );
  AOI22_X1 U21668 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18633), .B1(
        P3_EAX_REG_18__SCAN_IN), .B2(n18617), .ZN(n18583) );
  OAI21_X1 U21669 ( .B1(n18619), .B2(n21626), .A(n18583), .ZN(P3_U2770) );
  AOI22_X1 U21670 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18639), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18638), .ZN(n18584) );
  OAI21_X1 U21671 ( .B1(n18585), .B2(n18641), .A(n18584), .ZN(P3_U2771) );
  AOI22_X1 U21672 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18639), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18638), .ZN(n18586) );
  OAI21_X1 U21673 ( .B1(n18587), .B2(n18641), .A(n18586), .ZN(P3_U2772) );
  AOI22_X1 U21674 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18633), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18638), .ZN(n18588) );
  OAI21_X1 U21675 ( .B1(n18589), .B2(n18641), .A(n18588), .ZN(P3_U2773) );
  AOI22_X1 U21676 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18633), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18638), .ZN(n18590) );
  OAI21_X1 U21677 ( .B1(n18591), .B2(n18641), .A(n18590), .ZN(P3_U2774) );
  AOI22_X1 U21678 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18633), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18638), .ZN(n18592) );
  OAI21_X1 U21679 ( .B1(n10059), .B2(n18641), .A(n18592), .ZN(P3_U2775) );
  AOI22_X1 U21680 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18633), .B1(
        P3_EAX_REG_24__SCAN_IN), .B2(n18617), .ZN(n18593) );
  OAI21_X1 U21681 ( .B1(n18619), .B2(n21643), .A(n18593), .ZN(P3_U2776) );
  AOI22_X1 U21682 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18633), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18638), .ZN(n18594) );
  OAI21_X1 U21683 ( .B1(n10061), .B2(n18641), .A(n18594), .ZN(P3_U2777) );
  AOI22_X1 U21684 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18633), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18638), .ZN(n18595) );
  OAI21_X1 U21685 ( .B1(n18596), .B2(n18641), .A(n18595), .ZN(P3_U2778) );
  AOI22_X1 U21686 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18633), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18638), .ZN(n18597) );
  OAI21_X1 U21687 ( .B1(n18598), .B2(n18641), .A(n18597), .ZN(P3_U2779) );
  AOI22_X1 U21688 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18639), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18638), .ZN(n18599) );
  OAI21_X1 U21689 ( .B1(n18600), .B2(n18641), .A(n18599), .ZN(P3_U2780) );
  AOI22_X1 U21690 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18639), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18622), .ZN(n18601) );
  OAI21_X1 U21691 ( .B1(n18602), .B2(n18641), .A(n18601), .ZN(P3_U2781) );
  INV_X2 U21692 ( .A(n18617), .ZN(n18641) );
  AOI22_X1 U21693 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18639), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18622), .ZN(n18603) );
  OAI21_X1 U21694 ( .B1(n18604), .B2(n18641), .A(n18603), .ZN(P3_U2782) );
  AOI22_X1 U21695 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18622), .ZN(n18605) );
  OAI21_X1 U21696 ( .B1(n18606), .B2(n18641), .A(n18605), .ZN(P3_U2783) );
  AOI22_X1 U21697 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18622), .ZN(n18607) );
  OAI21_X1 U21698 ( .B1(n18608), .B2(n18641), .A(n18607), .ZN(P3_U2784) );
  AOI22_X1 U21699 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18622), .ZN(n18609) );
  OAI21_X1 U21700 ( .B1(n18610), .B2(n18641), .A(n18609), .ZN(P3_U2785) );
  AOI22_X1 U21701 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18622), .ZN(n18611) );
  OAI21_X1 U21702 ( .B1(n18612), .B2(n18641), .A(n18611), .ZN(P3_U2786) );
  AOI22_X1 U21703 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18622), .ZN(n18613) );
  OAI21_X1 U21704 ( .B1(n18614), .B2(n18641), .A(n18613), .ZN(P3_U2787) );
  AOI22_X1 U21705 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18622), .ZN(n18615) );
  OAI21_X1 U21706 ( .B1(n18616), .B2(n18641), .A(n18615), .ZN(P3_U2788) );
  AOI22_X1 U21707 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18639), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n18617), .ZN(n18618) );
  OAI21_X1 U21708 ( .B1(n18619), .B2(n21592), .A(n18618), .ZN(P3_U2789) );
  AOI22_X1 U21709 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18622), .ZN(n18620) );
  OAI21_X1 U21710 ( .B1(n18621), .B2(n18641), .A(n18620), .ZN(P3_U2790) );
  AOI22_X1 U21711 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18622), .ZN(n18623) );
  OAI21_X1 U21712 ( .B1(n18624), .B2(n18641), .A(n18623), .ZN(P3_U2791) );
  AOI22_X1 U21713 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18633), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18638), .ZN(n18625) );
  OAI21_X1 U21714 ( .B1(n18626), .B2(n18641), .A(n18625), .ZN(P3_U2792) );
  AOI22_X1 U21715 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18638), .ZN(n18627) );
  OAI21_X1 U21716 ( .B1(n18628), .B2(n18641), .A(n18627), .ZN(P3_U2793) );
  AOI22_X1 U21717 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18633), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18638), .ZN(n18629) );
  OAI21_X1 U21718 ( .B1(n18630), .B2(n18641), .A(n18629), .ZN(P3_U2794) );
  AOI22_X1 U21719 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18638), .ZN(n18631) );
  OAI21_X1 U21720 ( .B1(n18632), .B2(n18641), .A(n18631), .ZN(P3_U2795) );
  AOI22_X1 U21721 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18633), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18638), .ZN(n18634) );
  OAI21_X1 U21722 ( .B1(n18635), .B2(n18641), .A(n18634), .ZN(P3_U2796) );
  AOI22_X1 U21723 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18638), .ZN(n18636) );
  OAI21_X1 U21724 ( .B1(n18637), .B2(n18641), .A(n18636), .ZN(P3_U2797) );
  AOI22_X1 U21725 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18639), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18638), .ZN(n18640) );
  OAI21_X1 U21726 ( .B1(n18642), .B2(n18641), .A(n18640), .ZN(P3_U2798) );
  INV_X1 U21727 ( .A(n18713), .ZN(n18666) );
  NAND2_X1 U21728 ( .A1(n18666), .A2(n18911), .ZN(n18643) );
  XNOR2_X1 U21729 ( .A(n18643), .B(n11720), .ZN(n18915) );
  OAI21_X1 U21730 ( .B1(n18645), .B2(n18737), .A(n18906), .ZN(n18646) );
  AOI21_X1 U21731 ( .B1(n19515), .B2(n18644), .A(n18646), .ZN(n18683) );
  OAI21_X1 U21732 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18737), .A(
        n18683), .ZN(n18662) );
  NOR2_X1 U21733 ( .A1(n18739), .A2(n18644), .ZN(n18664) );
  OAI211_X1 U21734 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18664), .B(n18647), .ZN(n18648) );
  NAND2_X1 U21735 ( .A1(n19089), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18913) );
  OAI211_X1 U21736 ( .C1(n18749), .C2(n18649), .A(n18648), .B(n18913), .ZN(
        n18659) );
  NAND2_X1 U21737 ( .A1(n18911), .A2(n18665), .ZN(n18650) );
  XNOR2_X1 U21738 ( .A(n18650), .B(n11720), .ZN(n18920) );
  INV_X1 U21739 ( .A(n18651), .ZN(n18657) );
  NAND2_X1 U21740 ( .A1(n18652), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18655) );
  XNOR2_X1 U21741 ( .A(n18653), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18654) );
  MUX2_X1 U21742 ( .A(n18655), .B(n18654), .S(n18712), .Z(n18656) );
  OAI21_X1 U21743 ( .B1(n18657), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18656), .ZN(n18916) );
  OAI22_X1 U21744 ( .A1(n18811), .A2(n18920), .B1(n18829), .B2(n18916), .ZN(
        n18658) );
  AOI211_X1 U21745 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18662), .A(
        n18659), .B(n18658), .ZN(n18660) );
  OAI21_X1 U21746 ( .B1(n18810), .B2(n18915), .A(n18660), .ZN(P3_U2805) );
  AOI221_X1 U21747 ( .B1(n18664), .B2(n18663), .C1(n18662), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18661), .ZN(n18675) );
  OR2_X1 U21748 ( .A1(n18665), .A2(n18811), .ZN(n18668) );
  OR2_X1 U21749 ( .A1(n18810), .A2(n18666), .ZN(n18667) );
  NAND2_X1 U21750 ( .A1(n18668), .A2(n18667), .ZN(n18779) );
  AOI21_X1 U21751 ( .B1(n18780), .B2(n18669), .A(n18779), .ZN(n18680) );
  OAI22_X1 U21752 ( .A1(n18680), .A2(n17307), .B1(n18670), .B2(n18829), .ZN(
        n18671) );
  AOI21_X1 U21753 ( .B1(n18673), .B2(n18672), .A(n18671), .ZN(n18674) );
  OAI211_X1 U21754 ( .C1(n18749), .C2(n18676), .A(n18675), .B(n18674), .ZN(
        P3_U2806) );
  AND2_X1 U21755 ( .A1(n18711), .A2(n18716), .ZN(n18691) );
  NAND2_X1 U21756 ( .A1(n18712), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18678) );
  OAI211_X1 U21757 ( .C1(n9683), .C2(n18691), .A(n10321), .B(n18678), .ZN(
        n18679) );
  XNOR2_X1 U21758 ( .A(n18679), .B(n18921), .ZN(n18926) );
  AOI21_X1 U21759 ( .B1(n18921), .B2(n18681), .A(n18680), .ZN(n18685) );
  OAI22_X1 U21760 ( .A1(n18683), .A2(n18686), .B1(n18749), .B2(n18682), .ZN(
        n18684) );
  AOI211_X1 U21761 ( .C1(n19089), .C2(P3_REIP_REG_23__SCAN_IN), .A(n18685), 
        .B(n18684), .ZN(n18689) );
  NAND3_X1 U21762 ( .A1(n18687), .A2(n18818), .A3(n18686), .ZN(n18688) );
  OAI211_X1 U21763 ( .C1(n18829), .C2(n18926), .A(n18689), .B(n18688), .ZN(
        P3_U2807) );
  INV_X1 U21764 ( .A(n18937), .ZN(n18934) );
  NOR2_X1 U21765 ( .A1(n18713), .A2(n18934), .ZN(n18690) );
  OAI21_X1 U21766 ( .B1(n18691), .B2(n18690), .A(n10321), .ZN(n18693) );
  XNOR2_X1 U21767 ( .A(n18693), .B(n18692), .ZN(n18943) );
  INV_X1 U21768 ( .A(n18779), .ZN(n18694) );
  OAI21_X1 U21769 ( .B1(n18937), .B2(n18695), .A(n18694), .ZN(n18718) );
  OAI21_X1 U21770 ( .B1(n18697), .B2(n18737), .A(n18906), .ZN(n18698) );
  AOI21_X1 U21771 ( .B1(n18893), .B2(n18696), .A(n18698), .ZN(n18726) );
  OAI21_X1 U21772 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18725), .A(
        n18726), .ZN(n18708) );
  AOI22_X1 U21773 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18708), .B1(
        n18824), .B2(n18699), .ZN(n18702) );
  NOR2_X1 U21774 ( .A1(n18739), .A2(n18696), .ZN(n18709) );
  OAI211_X1 U21775 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18709), .B(n18700), .ZN(n18701) );
  OAI211_X1 U21776 ( .C1(n19691), .C2(n19055), .A(n18702), .B(n18701), .ZN(
        n18703) );
  AOI21_X1 U21777 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18718), .A(
        n18703), .ZN(n18705) );
  NAND3_X1 U21778 ( .A1(n18937), .A2(n18780), .A3(n18692), .ZN(n18704) );
  OAI211_X1 U21779 ( .C1(n18829), .C2(n18943), .A(n18705), .B(n18704), .ZN(
        P3_U2808) );
  NAND2_X1 U21780 ( .A1(n18952), .A2(n18716), .ZN(n18956) );
  NOR2_X1 U21781 ( .A1(n18973), .A2(n11713), .ZN(n18944) );
  NAND2_X1 U21782 ( .A1(n18780), .A2(n18944), .ZN(n18747) );
  OAI22_X1 U21783 ( .A1(n19120), .A2(n19690), .B1(n18749), .B2(n18706), .ZN(
        n18707) );
  AOI221_X1 U21784 ( .B1(n18709), .B2(n21596), .C1(n18708), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18707), .ZN(n18720) );
  INV_X1 U21785 ( .A(n18711), .ZN(n18715) );
  INV_X1 U21786 ( .A(n18952), .ZN(n18714) );
  OR4_X1 U21787 ( .A1(n18713), .A2(n11713), .A3(n18712), .A4(n18973), .ZN(
        n18735) );
  OAI22_X1 U21788 ( .A1(n18710), .A2(n18715), .B1(n18714), .B2(n18735), .ZN(
        n18717) );
  XNOR2_X1 U21789 ( .A(n18717), .B(n18716), .ZN(n18946) );
  AOI22_X1 U21790 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18718), .B1(
        n18846), .B2(n18946), .ZN(n18719) );
  OAI211_X1 U21791 ( .C1(n18956), .C2(n18747), .A(n18720), .B(n18719), .ZN(
        P3_U2809) );
  NAND2_X1 U21792 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18944), .ZN(
        n18957) );
  AOI21_X1 U21793 ( .B1(n18721), .B2(n18957), .A(n18779), .ZN(n18746) );
  INV_X1 U21794 ( .A(n18754), .ZN(n18723) );
  NAND2_X1 U21795 ( .A1(n18735), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18722) );
  OAI211_X1 U21796 ( .C1(n18723), .C2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10321), .B(n18722), .ZN(n18724) );
  XNOR2_X1 U21797 ( .A(n18724), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18960) );
  NAND2_X1 U21798 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18935), .ZN(
        n18964) );
  AOI221_X1 U21799 ( .B1(n18728), .B2(n18727), .C1(n19479), .C2(n18727), .A(
        n18726), .ZN(n18729) );
  AOI221_X1 U21800 ( .B1(n18824), .B2(n18731), .C1(n18730), .C2(n18731), .A(
        n18729), .ZN(n18732) );
  NAND2_X1 U21801 ( .A1(n19089), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18962) );
  OAI211_X1 U21802 ( .C1(n18964), .C2(n18747), .A(n18732), .B(n18962), .ZN(
        n18733) );
  AOI21_X1 U21803 ( .B1(n18846), .B2(n18960), .A(n18733), .ZN(n18734) );
  OAI21_X1 U21804 ( .B1(n18746), .B2(n18935), .A(n18734), .ZN(P3_U2810) );
  OR2_X1 U21805 ( .A1(n18710), .A2(n18754), .ZN(n18757) );
  NAND2_X1 U21806 ( .A1(n18757), .A2(n18735), .ZN(n18736) );
  XNOR2_X1 U21807 ( .A(n18736), .B(n18968), .ZN(n18965) );
  AOI21_X1 U21808 ( .B1(n18893), .B2(n9741), .A(n18880), .ZN(n18763) );
  OAI21_X1 U21809 ( .B1(n18738), .B2(n18737), .A(n18763), .ZN(n18751) );
  AOI22_X1 U21810 ( .A1(n19089), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18751), .ZN(n18742) );
  NOR2_X1 U21811 ( .A1(n18739), .A2(n9741), .ZN(n18753) );
  OAI211_X1 U21812 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18753), .B(n18740), .ZN(n18741) );
  OAI211_X1 U21813 ( .C1(n18749), .C2(n18743), .A(n18742), .B(n18741), .ZN(
        n18744) );
  AOI21_X1 U21814 ( .B1(n18846), .B2(n18965), .A(n18744), .ZN(n18745) );
  OAI221_X1 U21815 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18747), 
        .C1(n18968), .C2(n18746), .A(n18745), .ZN(P3_U2811) );
  AOI21_X1 U21816 ( .B1(n18780), .B2(n18973), .A(n18779), .ZN(n18769) );
  OAI22_X1 U21817 ( .A1(n19120), .A2(n19683), .B1(n18749), .B2(n18748), .ZN(
        n18750) );
  AOI221_X1 U21818 ( .B1(n18753), .B2(n18752), .C1(n18751), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18750), .ZN(n18760) );
  NAND2_X1 U21819 ( .A1(n10316), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18756) );
  NAND2_X1 U21820 ( .A1(n18756), .A2(n18754), .ZN(n18755) );
  MUX2_X1 U21821 ( .A(n18756), .B(n18755), .S(n18710), .Z(n18758) );
  NAND2_X1 U21822 ( .A1(n18758), .A2(n18757), .ZN(n18987) );
  NOR2_X1 U21823 ( .A1(n18973), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18986) );
  AOI22_X1 U21824 ( .A1(n18987), .A2(n18846), .B1(n18780), .B2(n18986), .ZN(
        n18759) );
  OAI211_X1 U21825 ( .C1(n18769), .C2(n11713), .A(n18760), .B(n18759), .ZN(
        P3_U2812) );
  AOI21_X1 U21826 ( .B1(n18761), .B2(n19515), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18762) );
  OAI22_X1 U21827 ( .A1(n18900), .A2(n18764), .B1(n18763), .B2(n18762), .ZN(
        n18765) );
  AOI21_X1 U21828 ( .B1(n19089), .B2(P3_REIP_REG_17__SCAN_IN), .A(n18765), 
        .ZN(n18768) );
  XNOR2_X1 U21829 ( .A(n18766), .B(n18979), .ZN(n18992) );
  INV_X1 U21830 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n19002) );
  NOR2_X1 U21831 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n19002), .ZN(
        n18991) );
  AOI22_X1 U21832 ( .A1(n18992), .A2(n18846), .B1(n18780), .B2(n18991), .ZN(
        n18767) );
  OAI211_X1 U21833 ( .C1(n18769), .C2(n18979), .A(n18768), .B(n18767), .ZN(
        P3_U2813) );
  OAI21_X1 U21834 ( .B1(n18985), .B2(n18833), .A(n18770), .ZN(n18771) );
  XNOR2_X1 U21835 ( .A(n18771), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n19007) );
  AOI22_X1 U21836 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18773), .B1(
        n18824), .B2(n18772), .ZN(n18777) );
  NAND2_X1 U21837 ( .A1(n19089), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n19005) );
  OAI211_X1 U21838 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18775), .B(n18774), .ZN(n18776) );
  NAND3_X1 U21839 ( .A1(n18777), .A2(n19005), .A3(n18776), .ZN(n18778) );
  AOI221_X1 U21840 ( .B1(n18780), .B2(n19002), .C1(n18779), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n18778), .ZN(n18781) );
  OAI21_X1 U21841 ( .B1(n19007), .B2(n18829), .A(n18781), .ZN(P3_U2814) );
  OAI21_X1 U21842 ( .B1(n9700), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18782), .ZN(n19043) );
  AOI21_X1 U21843 ( .B1(n18805), .B2(n18783), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18785) );
  OAI22_X1 U21844 ( .A1(n18900), .A2(n18786), .B1(n18785), .B2(n18784), .ZN(
        n18787) );
  AOI21_X1 U21845 ( .B1(n19089), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18787), 
        .ZN(n18793) );
  OAI21_X1 U21846 ( .B1(n18833), .B2(n19024), .A(n18788), .ZN(n18789) );
  XNOR2_X1 U21847 ( .A(n18789), .B(n19035), .ZN(n19040) );
  AOI21_X1 U21848 ( .B1(n14875), .B2(n19032), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18790) );
  OAI22_X1 U21849 ( .A1(n18790), .A2(n19010), .B1(n14875), .B2(n19035), .ZN(
        n19038) );
  AOI22_X1 U21850 ( .A1(n19040), .A2(n18846), .B1(n18791), .B2(n19038), .ZN(
        n18792) );
  OAI211_X1 U21851 ( .C1(n18811), .C2(n19043), .A(n18793), .B(n18792), .ZN(
        P3_U2816) );
  OR2_X1 U21852 ( .A1(n18794), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18816) );
  INV_X1 U21853 ( .A(n18816), .ZN(n18797) );
  OAI22_X1 U21854 ( .A1(n18795), .A2(n19045), .B1(n10316), .B2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18796) );
  OAI21_X1 U21855 ( .B1(n18797), .B2(n10316), .A(n18796), .ZN(n18798) );
  INV_X1 U21856 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n19022) );
  XNOR2_X1 U21857 ( .A(n18798), .B(n19022), .ZN(n19059) );
  NOR2_X1 U21858 ( .A1(n19120), .A2(n19673), .ZN(n18807) );
  OAI211_X1 U21859 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17232), .B(n18818), .ZN(n18804) );
  NOR2_X1 U21860 ( .A1(n17232), .A2(n18799), .ZN(n18800) );
  AOI211_X1 U21861 ( .C1(n18802), .C2(n18801), .A(n18880), .B(n18800), .ZN(
        n18819) );
  OAI22_X1 U21862 ( .A1(n18805), .A2(n18804), .B1(n18803), .B2(n18819), .ZN(
        n18806) );
  AOI211_X1 U21863 ( .C1(n18824), .C2(n18808), .A(n18807), .B(n18806), .ZN(
        n18815) );
  NOR2_X1 U21864 ( .A1(n18809), .A2(n19045), .ZN(n19047) );
  NOR2_X1 U21865 ( .A1(n18795), .A2(n19045), .ZN(n19049) );
  OAI22_X1 U21866 ( .A1(n19047), .A2(n18811), .B1(n18810), .B2(n19049), .ZN(
        n18826) );
  NOR2_X1 U21867 ( .A1(n18812), .A2(n19060), .ZN(n18825) );
  AOI22_X1 U21868 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18826), .B1(
        n18813), .B2(n18825), .ZN(n18814) );
  OAI211_X1 U21869 ( .C1(n18829), .C2(n19059), .A(n18815), .B(n18814), .ZN(
        P3_U2817) );
  OAI21_X1 U21870 ( .B1(n18833), .B2(n19060), .A(n18816), .ZN(n18817) );
  XNOR2_X1 U21871 ( .A(n18817), .B(n11705), .ZN(n19067) );
  INV_X1 U21872 ( .A(n19067), .ZN(n18830) );
  NAND2_X1 U21873 ( .A1(n17232), .A2(n18818), .ZN(n18821) );
  NAND2_X1 U21874 ( .A1(n19089), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n19068) );
  OAI221_X1 U21875 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18821), .C1(
        n18820), .C2(n18819), .A(n19068), .ZN(n18822) );
  AOI21_X1 U21876 ( .B1(n18824), .B2(n18823), .A(n18822), .ZN(n18828) );
  AOI22_X1 U21877 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18826), .B1(
        n18825), .B2(n11705), .ZN(n18827) );
  OAI211_X1 U21878 ( .C1(n18830), .C2(n18829), .A(n18828), .B(n18827), .ZN(
        P3_U2818) );
  AOI21_X1 U21879 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18860), .A(
        n18831), .ZN(n18848) );
  NOR2_X1 U21880 ( .A1(n18835), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18832) );
  OAI22_X1 U21881 ( .A1(n18832), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19080), .B2(n18833), .ZN(n18838) );
  INV_X1 U21882 ( .A(n18833), .ZN(n18834) );
  NAND3_X1 U21883 ( .A1(n18834), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n19080), .ZN(n18837) );
  NOR3_X1 U21884 ( .A1(n18835), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n19088), .ZN(n18836) );
  AOI21_X1 U21885 ( .B1(n18838), .B2(n18837), .A(n18836), .ZN(n19092) );
  INV_X1 U21886 ( .A(n18839), .ZN(n18844) );
  AOI21_X1 U21887 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18841), .A(
        n18840), .ZN(n18842) );
  OAI22_X1 U21888 ( .A1(n18900), .A2(n18844), .B1(n18843), .B2(n18842), .ZN(
        n18845) );
  AOI21_X1 U21889 ( .B1(n18846), .B2(n19092), .A(n18845), .ZN(n18847) );
  NAND2_X1 U21890 ( .A1(n19089), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n19094) );
  OAI211_X1 U21891 ( .C1(n18849), .C2(n18848), .A(n18847), .B(n19094), .ZN(
        P3_U2820) );
  AOI22_X1 U21892 ( .A1(n19089), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18850), .ZN(n18858) );
  NAND2_X1 U21893 ( .A1(n18852), .A2(n18851), .ZN(n18853) );
  XNOR2_X1 U21894 ( .A(n18853), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19110) );
  XNOR2_X1 U21895 ( .A(n18854), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19108) );
  OAI22_X1 U21896 ( .A1(n18900), .A2(n18855), .B1(n19108), .B2(n18897), .ZN(
        n18856) );
  AOI21_X1 U21897 ( .B1(n18904), .B2(n19110), .A(n18856), .ZN(n18857) );
  OAI211_X1 U21898 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18859), .A(
        n18858), .B(n18857), .ZN(P3_U2823) );
  INV_X1 U21899 ( .A(n18860), .ZN(n18861) );
  NOR2_X1 U21900 ( .A1(n18861), .A2(n18865), .ZN(n18874) );
  OAI22_X1 U21901 ( .A1(n18897), .A2(n18862), .B1(n19660), .B2(n19120), .ZN(
        n18863) );
  AOI221_X1 U21902 ( .B1(n18874), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C1(
        n18865), .C2(n18864), .A(n18863), .ZN(n18869) );
  AOI22_X1 U21903 ( .A1(n18904), .A2(n18867), .B1(n18866), .B2(n18884), .ZN(
        n18868) );
  NAND2_X1 U21904 ( .A1(n18869), .A2(n18868), .ZN(P3_U2824) );
  INV_X1 U21905 ( .A(n18870), .ZN(n18871) );
  INV_X1 U21906 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19658) );
  OAI22_X1 U21907 ( .A1(n18897), .A2(n18871), .B1(n19658), .B2(n19120), .ZN(
        n18872) );
  AOI21_X1 U21908 ( .B1(n18904), .B2(n18873), .A(n18872), .ZN(n18876) );
  OAI221_X1 U21909 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17946), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18906), .A(n18874), .ZN(n18875) );
  OAI211_X1 U21910 ( .C1(n18900), .C2(n18877), .A(n18876), .B(n18875), .ZN(
        P3_U2825) );
  AOI22_X1 U21911 ( .A1(n18904), .A2(n18879), .B1(n19515), .B2(n18878), .ZN(
        n18887) );
  AOI21_X1 U21912 ( .B1(n18893), .B2(n17990), .A(n18880), .ZN(n18889) );
  OAI22_X1 U21913 ( .A1(n18889), .A2(n18882), .B1(n18897), .B2(n18881), .ZN(
        n18883) );
  AOI21_X1 U21914 ( .B1(n18885), .B2(n18884), .A(n18883), .ZN(n18886) );
  OAI211_X1 U21915 ( .C1(n19055), .C2(n19656), .A(n18887), .B(n18886), .ZN(
        P3_U2826) );
  OAI22_X1 U21916 ( .A1(n18889), .A2(n21653), .B1(n18897), .B2(n18888), .ZN(
        n18890) );
  AOI211_X1 U21917 ( .C1(n18904), .C2(n18892), .A(n18891), .B(n18890), .ZN(
        n18895) );
  NAND4_X1 U21918 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18893), .A3(
        n18906), .A4(n21653), .ZN(n18894) );
  OAI211_X1 U21919 ( .C1(n18900), .C2(n18896), .A(n18895), .B(n18894), .ZN(
        P3_U2827) );
  OAI22_X1 U21920 ( .A1(n18900), .A2(n18899), .B1(n18898), .B2(n18897), .ZN(
        n18901) );
  AOI211_X1 U21921 ( .C1(n18904), .C2(n18903), .A(n18902), .B(n18901), .ZN(
        n18905) );
  OAI221_X1 U21922 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19479), .C1(
        n18907), .C2(n18906), .A(n18905), .ZN(P3_U2828) );
  OAI221_X1 U21923 ( .B1(n18971), .B2(n18972), .C1(n18971), .C2(n18911), .A(
        n18908), .ZN(n18912) );
  NOR2_X1 U21924 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18909), .ZN(
        n18910) );
  AOI22_X1 U21925 ( .A1(n18912), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18911), .B2(n18910), .ZN(n18914) );
  OAI21_X1 U21926 ( .B1(n19121), .B2(n18914), .A(n18913), .ZN(n18918) );
  OAI22_X1 U21927 ( .A1(n19058), .A2(n18916), .B1(n19037), .B2(n18915), .ZN(
        n18917) );
  AOI211_X1 U21928 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n19008), .A(
        n18918), .B(n18917), .ZN(n18919) );
  OAI21_X1 U21929 ( .B1(n19044), .B2(n18920), .A(n18919), .ZN(P3_U2837) );
  OAI21_X1 U21930 ( .B1(n19008), .B2(n18922), .A(n18921), .ZN(n18923) );
  OAI21_X1 U21931 ( .B1(n19058), .B2(n18926), .A(n18925), .ZN(P3_U2839) );
  AOI21_X1 U21932 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n19073), .A(
        n18927), .ZN(n18933) );
  INV_X1 U21933 ( .A(n18928), .ZN(n18930) );
  AOI21_X1 U21934 ( .B1(n18972), .B2(n18944), .A(n18971), .ZN(n18929) );
  AOI221_X1 U21935 ( .B1(n18930), .B2(n19122), .C1(n18957), .C2(n19122), .A(
        n18929), .ZN(n18950) );
  INV_X1 U21936 ( .A(n18950), .ZN(n18932) );
  OAI22_X1 U21937 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n19090), .B1(
        n18952), .B2(n18971), .ZN(n18931) );
  NOR4_X1 U21938 ( .A1(n18933), .A2(n18932), .A3(n18947), .A4(n18931), .ZN(
        n18939) );
  AOI22_X1 U21939 ( .A1(n19122), .A2(n18935), .B1(n18934), .B2(n18975), .ZN(
        n18951) );
  NAND2_X1 U21940 ( .A1(n18937), .A2(n18936), .ZN(n18938) );
  AOI22_X1 U21941 ( .A1(n18939), .A2(n18951), .B1(n18692), .B2(n18938), .ZN(
        n18940) );
  AOI22_X1 U21942 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19008), .B1(
        n19053), .B2(n18940), .ZN(n18942) );
  NAND2_X1 U21943 ( .A1(n19089), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18941) );
  OAI211_X1 U21944 ( .C1(n18943), .C2(n19058), .A(n18942), .B(n18941), .ZN(
        P3_U2840) );
  INV_X1 U21945 ( .A(n18944), .ZN(n18948) );
  AOI22_X1 U21946 ( .A1(n19089), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n19099), 
        .B2(n18946), .ZN(n18955) );
  OAI21_X1 U21947 ( .B1(n18999), .B2(n18948), .A(n18998), .ZN(n18949) );
  NAND3_X1 U21948 ( .A1(n19000), .A2(n18950), .A3(n18949), .ZN(n18958) );
  OAI21_X1 U21949 ( .B1(n19029), .B2(n18952), .A(n18951), .ZN(n18953) );
  OAI211_X1 U21950 ( .C1(n18958), .C2(n18953), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n19120), .ZN(n18954) );
  OAI211_X1 U21951 ( .C1(n18969), .C2(n18956), .A(n18955), .B(n18954), .ZN(
        P3_U2841) );
  NAND2_X1 U21952 ( .A1(n18968), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18959) );
  OAI221_X1 U21953 ( .B1(n18958), .B2(n18975), .C1(n18958), .C2(n18957), .A(
        n19120), .ZN(n18967) );
  OAI21_X1 U21954 ( .B1(n19029), .B2(n18959), .A(n18967), .ZN(n18961) );
  AOI22_X1 U21955 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18961), .B1(
        n19099), .B2(n18960), .ZN(n18963) );
  OAI211_X1 U21956 ( .C1(n18964), .C2(n18969), .A(n18963), .B(n18962), .ZN(
        P3_U2842) );
  AOI22_X1 U21957 ( .A1(n19089), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n19099), 
        .B2(n18965), .ZN(n18966) );
  OAI221_X1 U21958 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18969), 
        .C1(n18968), .C2(n18967), .A(n18966), .ZN(P3_U2843) );
  OAI21_X1 U21959 ( .B1(n19002), .B2(n18970), .A(n18978), .ZN(n18977) );
  NOR2_X1 U21960 ( .A1(n18972), .A2(n18971), .ZN(n18974) );
  OAI22_X1 U21961 ( .A1(n19586), .A2(n18975), .B1(n18974), .B2(n18973), .ZN(
        n18976) );
  NAND3_X1 U21962 ( .A1(n19000), .A2(n18977), .A3(n18976), .ZN(n18990) );
  OAI221_X1 U21963 ( .B1(n18990), .B2(n18979), .C1(n18990), .C2(n18978), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18989) );
  NOR2_X1 U21964 ( .A1(n18981), .A2(n18980), .ZN(n19104) );
  NAND2_X1 U21965 ( .A1(n18982), .A2(n19104), .ZN(n19009) );
  INV_X1 U21966 ( .A(n18983), .ZN(n18984) );
  OAI211_X1 U21967 ( .C1(n19048), .C2(n18795), .A(n19009), .B(n18984), .ZN(
        n19061) );
  NAND2_X1 U21968 ( .A1(n19053), .A2(n19061), .ZN(n19103) );
  NOR2_X1 U21969 ( .A1(n18985), .A2(n19103), .ZN(n19003) );
  AOI22_X1 U21970 ( .A1(n18987), .A2(n19099), .B1(n18986), .B2(n19003), .ZN(
        n18988) );
  OAI221_X1 U21971 ( .B1(n19089), .B2(n18989), .C1(n19055), .C2(n19683), .A(
        n18988), .ZN(P3_U2844) );
  NAND2_X1 U21972 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18990), .ZN(
        n18994) );
  AOI22_X1 U21973 ( .A1(n18992), .A2(n19099), .B1(n19003), .B2(n18991), .ZN(
        n18993) );
  OAI221_X1 U21974 ( .B1(n19089), .B2(n18994), .C1(n19055), .C2(n19681), .A(
        n18993), .ZN(P3_U2845) );
  INV_X1 U21975 ( .A(n18995), .ZN(n19001) );
  AOI22_X1 U21976 ( .A1(n19586), .A2(n19025), .B1(n19122), .B2(n19023), .ZN(
        n19071) );
  AOI21_X1 U21977 ( .B1(n19010), .B2(n19071), .A(n19090), .ZN(n18996) );
  AOI211_X1 U21978 ( .C1(n18999), .C2(n18998), .A(n18997), .B(n18996), .ZN(
        n19014) );
  AOI221_X1 U21979 ( .B1(n19001), .B2(n19000), .C1(n19014), .C2(n19000), .A(
        n19089), .ZN(n19004) );
  AOI22_X1 U21980 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19004), .B1(
        n19003), .B2(n19002), .ZN(n19006) );
  OAI211_X1 U21981 ( .C1(n19007), .C2(n19058), .A(n19006), .B(n19005), .ZN(
        P3_U2846) );
  AOI22_X1 U21982 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19008), .B1(
        n19089), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n19018) );
  INV_X1 U21983 ( .A(n19009), .ZN(n19031) );
  AOI21_X1 U21984 ( .B1(n19010), .B2(n19031), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19013) );
  AOI21_X1 U21985 ( .B1(n14875), .B2(n19010), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19012) );
  OAI22_X1 U21986 ( .A1(n19014), .A2(n19013), .B1(n19012), .B2(n19011), .ZN(
        n19016) );
  AOI22_X1 U21987 ( .A1(n19053), .A2(n19016), .B1(n19099), .B2(n19015), .ZN(
        n19017) );
  OAI211_X1 U21988 ( .C1(n19044), .C2(n19019), .A(n19018), .B(n19017), .ZN(
        P3_U2847) );
  NOR2_X1 U21989 ( .A1(n19020), .A2(n19023), .ZN(n19072) );
  AOI21_X1 U21990 ( .B1(n19021), .B2(n19072), .A(n19073), .ZN(n19052) );
  NOR2_X1 U21991 ( .A1(n19052), .A2(n19022), .ZN(n19028) );
  OAI21_X1 U21992 ( .B1(n19024), .B2(n19023), .A(n19122), .ZN(n19027) );
  OAI21_X1 U21993 ( .B1(n19045), .B2(n19025), .A(n19586), .ZN(n19026) );
  OAI211_X1 U21994 ( .C1(n19029), .C2(n19028), .A(n19027), .B(n19026), .ZN(
        n19030) );
  OAI21_X1 U21995 ( .B1(n19035), .B2(n19030), .A(n19053), .ZN(n19034) );
  NAND2_X1 U21996 ( .A1(n19032), .A2(n19031), .ZN(n19033) );
  AOI222_X1 U21997 ( .A1(n19035), .A2(n19034), .B1(n19035), .B2(n19033), .C1(
        n19034), .C2(n19114), .ZN(n19036) );
  AOI21_X1 U21998 ( .B1(n19089), .B2(P3_REIP_REG_14__SCAN_IN), .A(n19036), 
        .ZN(n19042) );
  INV_X1 U21999 ( .A(n19037), .ZN(n19039) );
  AOI22_X1 U22000 ( .A1(n19040), .A2(n19099), .B1(n19039), .B2(n19038), .ZN(
        n19041) );
  OAI211_X1 U22001 ( .C1(n19044), .C2(n19043), .A(n19042), .B(n19041), .ZN(
        P3_U2848) );
  NOR3_X1 U22002 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19045), .A3(
        n19103), .ZN(n19046) );
  AOI21_X1 U22003 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n19089), .A(n19046), 
        .ZN(n19057) );
  AOI21_X1 U22004 ( .B1(n19122), .B2(n19081), .A(n11705), .ZN(n19064) );
  AOI22_X1 U22005 ( .A1(n19586), .A2(n19060), .B1(n19122), .B2(n19080), .ZN(
        n19082) );
  OAI211_X1 U22006 ( .C1(n19047), .C2(n19077), .A(n19071), .B(n19082), .ZN(
        n19051) );
  NOR2_X1 U22007 ( .A1(n19049), .A2(n19048), .ZN(n19050) );
  NOR3_X1 U22008 ( .A1(n19052), .A2(n19051), .A3(n19050), .ZN(n19065) );
  OAI211_X1 U22009 ( .C1(n19090), .C2(n19064), .A(n19053), .B(n19065), .ZN(
        n19054) );
  NAND3_X1 U22010 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19055), .A3(
        n19054), .ZN(n19056) );
  OAI211_X1 U22011 ( .C1(n19059), .C2(n19058), .A(n19057), .B(n19056), .ZN(
        P3_U2849) );
  INV_X1 U22012 ( .A(n19060), .ZN(n19062) );
  AOI21_X1 U22013 ( .B1(n19062), .B2(n19061), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19063) );
  AOI211_X1 U22014 ( .C1(n19065), .C2(n19064), .A(n19063), .B(n19121), .ZN(
        n19066) );
  AOI21_X1 U22015 ( .B1(n19099), .B2(n19067), .A(n19066), .ZN(n19069) );
  OAI211_X1 U22016 ( .C1(n19114), .C2(n11705), .A(n19069), .B(n19068), .ZN(
        P3_U2850) );
  NAND2_X1 U22017 ( .A1(n19070), .A2(n19073), .ZN(n19079) );
  OAI211_X1 U22018 ( .C1(n19073), .C2(n19072), .A(n19071), .B(n19114), .ZN(
        n19074) );
  AOI21_X1 U22019 ( .B1(n19075), .B2(n18795), .A(n19074), .ZN(n19076) );
  OAI21_X1 U22020 ( .B1(n19078), .B2(n19077), .A(n19076), .ZN(n19097) );
  AOI21_X1 U22021 ( .B1(n19080), .B2(n19079), .A(n19097), .ZN(n19091) );
  AOI211_X1 U22022 ( .C1(n19082), .C2(n19091), .A(n19089), .B(n19081), .ZN(
        n19083) );
  AOI211_X1 U22023 ( .C1(n19099), .C2(n19085), .A(n19084), .B(n19083), .ZN(
        n19086) );
  OAI21_X1 U22024 ( .B1(n19103), .B2(n19087), .A(n19086), .ZN(P3_U2851) );
  NAND2_X1 U22025 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n19088), .ZN(
        n19096) );
  AOI221_X1 U22026 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19091), .C1(
        n19090), .C2(n19091), .A(n19089), .ZN(n19093) );
  AOI22_X1 U22027 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n19093), .B1(
        n19099), .B2(n19092), .ZN(n19095) );
  OAI211_X1 U22028 ( .C1(n19096), .C2(n19103), .A(n19095), .B(n19094), .ZN(
        P3_U2852) );
  NAND2_X1 U22029 ( .A1(n19097), .A2(n19055), .ZN(n19101) );
  AOI22_X1 U22030 ( .A1(n19089), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n19099), 
        .B2(n19098), .ZN(n19100) );
  OAI221_X1 U22031 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19103), .C1(
        n19102), .C2(n19101), .A(n19100), .ZN(P3_U2853) );
  AOI21_X1 U22032 ( .B1(n19104), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19105) );
  OR3_X1 U22033 ( .A1(n19106), .A2(n19105), .A3(n19121), .ZN(n19107) );
  OAI21_X1 U22034 ( .B1(n19108), .B2(n19115), .A(n19107), .ZN(n19109) );
  AOI21_X1 U22035 ( .B1(n19119), .B2(n19110), .A(n19109), .ZN(n19112) );
  NAND2_X1 U22036 ( .A1(n19089), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n19111) );
  OAI211_X1 U22037 ( .C1(n19114), .C2(n19113), .A(n19112), .B(n19111), .ZN(
        P3_U2855) );
  NOR2_X1 U22038 ( .A1(n19115), .A2(n19118), .ZN(n19116) );
  AOI211_X1 U22039 ( .C1(n19119), .C2(n19118), .A(n19117), .B(n19116), .ZN(
        n19125) );
  OAI211_X1 U22040 ( .C1(n19122), .C2(n19121), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n19120), .ZN(n19123) );
  NAND3_X1 U22041 ( .A1(n19125), .A2(n19124), .A3(n19123), .ZN(P3_U2862) );
  INV_X1 U22042 ( .A(n19126), .ZN(n19129) );
  AOI21_X1 U22043 ( .B1(n19129), .B2(n19128), .A(n19127), .ZN(n19618) );
  OAI21_X1 U22044 ( .B1(n19618), .B2(n19130), .A(n19135), .ZN(n19131) );
  OAI221_X1 U22045 ( .B1(n11865), .B2(n19742), .C1(n11865), .C2(n19135), .A(
        n19131), .ZN(P3_U2863) );
  NOR2_X1 U22046 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11856), .ZN(
        n19316) );
  NOR2_X1 U22047 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19609), .ZN(
        n19360) );
  NOR2_X1 U22048 ( .A1(n19316), .A2(n19360), .ZN(n19133) );
  OAI22_X1 U22049 ( .A1(n19134), .A2(n19609), .B1(n19133), .B2(n19132), .ZN(
        P3_U2866) );
  NOR2_X1 U22050 ( .A1(n11859), .A2(n19135), .ZN(P3_U2867) );
  NOR2_X1 U22051 ( .A1(n19609), .A2(n19288), .ZN(n19513) );
  INV_X1 U22052 ( .A(n19513), .ZN(n19508) );
  NOR2_X2 U22053 ( .A1(n11865), .A2(n19508), .ZN(n19546) );
  NAND2_X1 U22054 ( .A1(n11853), .A2(n11865), .ZN(n19575) );
  NOR2_X1 U22055 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19225) );
  INV_X1 U22056 ( .A(n19225), .ZN(n19179) );
  OR2_X1 U22057 ( .A1(n19575), .A2(n19179), .ZN(n19216) );
  NOR2_X1 U22058 ( .A1(n19546), .A2(n19241), .ZN(n19201) );
  OAI21_X1 U22059 ( .B1(n11865), .B2(n19723), .A(n19384), .ZN(n19202) );
  NOR2_X2 U22060 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19508), .ZN(
        n19496) );
  NOR2_X1 U22061 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n11865), .ZN(
        n19359) );
  INV_X1 U22062 ( .A(n19359), .ZN(n19136) );
  NAND2_X1 U22063 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19452) );
  NOR2_X2 U22064 ( .A1(n19136), .A2(n19452), .ZN(n19560) );
  OAI21_X1 U22065 ( .B1(n19496), .B2(n19560), .A(n19384), .ZN(n19478) );
  OAI22_X1 U22066 ( .A1(n19201), .A2(n19202), .B1(n19381), .B2(n19478), .ZN(
        n19175) );
  NAND2_X1 U22067 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19515), .ZN(n19485) );
  INV_X1 U22068 ( .A(n19485), .ZN(n19511) );
  NOR2_X2 U22069 ( .A1(n19428), .A2(n19137), .ZN(n19510) );
  NOR2_X1 U22070 ( .A1(n19509), .A2(n19201), .ZN(n19174) );
  AOI22_X1 U22071 ( .A1(n19511), .A2(n19560), .B1(n19510), .B2(n19174), .ZN(
        n19142) );
  NOR2_X1 U22072 ( .A1(n19139), .A2(n19138), .ZN(n19172) );
  INV_X1 U22073 ( .A(n19172), .ZN(n19161) );
  NOR2_X1 U22074 ( .A1(n19140), .A2(n19161), .ZN(n19482) );
  AND2_X1 U22075 ( .A1(n19515), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19516) );
  AOI22_X1 U22076 ( .A1(n19482), .A2(n19241), .B1(n19516), .B2(n19496), .ZN(
        n19141) );
  OAI211_X1 U22077 ( .C1(n14698), .C2(n19175), .A(n19142), .B(n19141), .ZN(
        P3_U2868) );
  NOR2_X2 U22078 ( .A1(n19428), .A2(n19143), .ZN(n19520) );
  NOR2_X2 U22079 ( .A1(n19857), .A2(n19479), .ZN(n19522) );
  AOI22_X1 U22080 ( .A1(n19520), .A2(n19174), .B1(n19522), .B2(n19560), .ZN(
        n19147) );
  NOR2_X2 U22081 ( .A1(n19479), .A2(n19144), .ZN(n19521) );
  NAND2_X1 U22082 ( .A1(n19172), .A2(n19736), .ZN(n19525) );
  INV_X1 U22083 ( .A(n19525), .ZN(n19145) );
  AOI22_X1 U22084 ( .A1(n19521), .A2(n19496), .B1(n19145), .B2(n19241), .ZN(
        n19146) );
  OAI211_X1 U22085 ( .C1(n19148), .C2(n19175), .A(n19147), .B(n19146), .ZN(
        P3_U2869) );
  AND2_X1 U22086 ( .A1(n19515), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19527) );
  NOR2_X2 U22087 ( .A1(n19428), .A2(n19149), .ZN(n19526) );
  AOI22_X1 U22088 ( .A1(n19527), .A2(n19496), .B1(n19526), .B2(n19174), .ZN(
        n19151) );
  NAND2_X1 U22089 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19515), .ZN(n19531) );
  INV_X1 U22090 ( .A(n19531), .ZN(n19461) );
  NOR2_X1 U22091 ( .A1(n9695), .A2(n19161), .ZN(n19528) );
  AOI22_X1 U22092 ( .A1(n19461), .A2(n19560), .B1(n19528), .B2(n19241), .ZN(
        n19150) );
  OAI211_X1 U22093 ( .C1(n18333), .C2(n19175), .A(n19151), .B(n19150), .ZN(
        P3_U2870) );
  NOR2_X2 U22094 ( .A1(n19428), .A2(n19152), .ZN(n19533) );
  AND2_X1 U22095 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19515), .ZN(n19532) );
  AOI22_X1 U22096 ( .A1(n19533), .A2(n19174), .B1(n19532), .B2(n19560), .ZN(
        n19155) );
  NOR2_X2 U22097 ( .A1(n19479), .A2(n19867), .ZN(n19534) );
  NOR2_X1 U22098 ( .A1(n19161), .A2(n19153), .ZN(n19187) );
  AOI22_X1 U22099 ( .A1(n19534), .A2(n19496), .B1(n19187), .B2(n19241), .ZN(
        n19154) );
  OAI211_X1 U22100 ( .C1(n19156), .C2(n19175), .A(n19155), .B(n19154), .ZN(
        P3_U2871) );
  AND2_X1 U22101 ( .A1(n19515), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19540) );
  AND2_X1 U22102 ( .A1(n19384), .A2(BUF2_REG_4__SCAN_IN), .ZN(n19539) );
  AOI22_X1 U22103 ( .A1(n19540), .A2(n19496), .B1(n19539), .B2(n19174), .ZN(
        n19159) );
  NOR2_X1 U22104 ( .A1(n19161), .A2(n19157), .ZN(n19190) );
  NOR2_X2 U22105 ( .A1(n19874), .A2(n19479), .ZN(n19538) );
  AOI22_X1 U22106 ( .A1(n19190), .A2(n19241), .B1(n19538), .B2(n19560), .ZN(
        n19158) );
  OAI211_X1 U22107 ( .C1(n19160), .C2(n19175), .A(n19159), .B(n19158), .ZN(
        P3_U2872) );
  NOR2_X2 U22108 ( .A1(n19428), .A2(n13896), .ZN(n19545) );
  NAND2_X1 U22109 ( .A1(n19515), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19499) );
  INV_X1 U22110 ( .A(n19499), .ZN(n19544) );
  AOI22_X1 U22111 ( .A1(n19545), .A2(n19174), .B1(n19544), .B2(n19496), .ZN(
        n19164) );
  NAND2_X1 U22112 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19515), .ZN(n19551) );
  NOR2_X2 U22113 ( .A1(n19162), .A2(n19161), .ZN(n19547) );
  AOI22_X1 U22114 ( .A1(n19495), .A2(n19560), .B1(n19547), .B2(n19241), .ZN(
        n19163) );
  OAI211_X1 U22115 ( .C1(n19165), .C2(n19175), .A(n19164), .B(n19163), .ZN(
        P3_U2873) );
  NOR2_X2 U22116 ( .A1(n19428), .A2(n13881), .ZN(n19552) );
  NOR2_X2 U22117 ( .A1(n19884), .A2(n19479), .ZN(n19554) );
  AOI22_X1 U22118 ( .A1(n19552), .A2(n19174), .B1(n19554), .B2(n19560), .ZN(
        n19169) );
  AND2_X1 U22119 ( .A1(n19515), .A2(BUF2_REG_22__SCAN_IN), .ZN(n19553) );
  NAND2_X1 U22120 ( .A1(n19172), .A2(n19166), .ZN(n19557) );
  INV_X1 U22121 ( .A(n19557), .ZN(n19167) );
  AOI22_X1 U22122 ( .A1(n19553), .A2(n19496), .B1(n19167), .B2(n19241), .ZN(
        n19168) );
  OAI211_X1 U22123 ( .C1(n19170), .C2(n19175), .A(n19169), .B(n19168), .ZN(
        P3_U2874) );
  NAND2_X1 U22124 ( .A1(n19172), .A2(n19171), .ZN(n19568) );
  NOR2_X2 U22125 ( .A1(n19479), .A2(n19173), .ZN(n19563) );
  NOR2_X2 U22126 ( .A1(n13838), .A2(n19428), .ZN(n19559) );
  AOI22_X1 U22127 ( .A1(n19563), .A2(n19560), .B1(n19559), .B2(n19174), .ZN(
        n19178) );
  INV_X1 U22128 ( .A(n19175), .ZN(n19176) );
  NOR2_X2 U22129 ( .A1(n16490), .A2(n19479), .ZN(n19561) );
  AOI22_X1 U22130 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19176), .B1(
        n19561), .B2(n19496), .ZN(n19177) );
  OAI211_X1 U22131 ( .C1(n19568), .C2(n19216), .A(n19178), .B(n19177), .ZN(
        P3_U2875) );
  NAND2_X1 U22132 ( .A1(n19225), .A2(n19359), .ZN(n19259) );
  INV_X1 U22133 ( .A(n19509), .ZN(n19626) );
  NAND2_X1 U22134 ( .A1(n11853), .A2(n19626), .ZN(n19451) );
  NOR2_X1 U22135 ( .A1(n19179), .A2(n19451), .ZN(n19197) );
  AOI22_X1 U22136 ( .A1(n19511), .A2(n19496), .B1(n19510), .B2(n19197), .ZN(
        n19182) );
  NAND2_X1 U22137 ( .A1(n19384), .A2(n19180), .ZN(n19405) );
  NOR2_X1 U22138 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19405), .ZN(
        n19453) );
  AOI22_X1 U22139 ( .A1(n19515), .A2(n19513), .B1(n19225), .B2(n19453), .ZN(
        n19198) );
  AOI22_X1 U22140 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19198), .B1(
        n19516), .B2(n19546), .ZN(n19181) );
  OAI211_X1 U22141 ( .C1(n19259), .C2(n19519), .A(n19182), .B(n19181), .ZN(
        P3_U2876) );
  AOI22_X1 U22142 ( .A1(n19521), .A2(n19546), .B1(n19520), .B2(n19197), .ZN(
        n19184) );
  AOI22_X1 U22143 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19198), .B1(
        n19522), .B2(n19496), .ZN(n19183) );
  OAI211_X1 U22144 ( .C1(n19259), .C2(n19525), .A(n19184), .B(n19183), .ZN(
        P3_U2877) );
  AOI22_X1 U22145 ( .A1(n19461), .A2(n19496), .B1(n19526), .B2(n19197), .ZN(
        n19186) );
  AOI22_X1 U22146 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19198), .B1(
        n19527), .B2(n19546), .ZN(n19185) );
  OAI211_X1 U22147 ( .C1(n19259), .C2(n19464), .A(n19186), .B(n19185), .ZN(
        P3_U2878) );
  AOI22_X1 U22148 ( .A1(n19534), .A2(n19546), .B1(n19533), .B2(n19197), .ZN(
        n19189) );
  AOI22_X1 U22149 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19198), .B1(
        n19532), .B2(n19496), .ZN(n19188) );
  OAI211_X1 U22150 ( .C1(n19259), .C2(n19537), .A(n19189), .B(n19188), .ZN(
        P3_U2879) );
  INV_X1 U22151 ( .A(n19190), .ZN(n19543) );
  AOI22_X1 U22152 ( .A1(n19539), .A2(n19197), .B1(n19538), .B2(n19496), .ZN(
        n19192) );
  AOI22_X1 U22153 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19198), .B1(
        n19540), .B2(n19546), .ZN(n19191) );
  OAI211_X1 U22154 ( .C1(n19259), .C2(n19543), .A(n19192), .B(n19191), .ZN(
        P3_U2880) );
  INV_X1 U22155 ( .A(n19496), .ZN(n19507) );
  AOI22_X1 U22156 ( .A1(n19545), .A2(n19197), .B1(n19544), .B2(n19546), .ZN(
        n19194) );
  AOI22_X1 U22157 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19198), .B1(
        n19263), .B2(n19547), .ZN(n19193) );
  OAI211_X1 U22158 ( .C1(n19551), .C2(n19507), .A(n19194), .B(n19193), .ZN(
        P3_U2881) );
  AOI22_X1 U22159 ( .A1(n19553), .A2(n19546), .B1(n19552), .B2(n19197), .ZN(
        n19196) );
  AOI22_X1 U22160 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19198), .B1(
        n19554), .B2(n19496), .ZN(n19195) );
  OAI211_X1 U22161 ( .C1(n19259), .C2(n19557), .A(n19196), .B(n19195), .ZN(
        P3_U2882) );
  AOI22_X1 U22162 ( .A1(n19561), .A2(n19546), .B1(n19559), .B2(n19197), .ZN(
        n19200) );
  AOI22_X1 U22163 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19198), .B1(
        n19563), .B2(n19496), .ZN(n19199) );
  OAI211_X1 U22164 ( .C1(n19259), .C2(n19568), .A(n19200), .B(n19199), .ZN(
        P3_U2883) );
  NAND2_X1 U22165 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19225), .ZN(
        n19224) );
  NOR2_X2 U22166 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19224), .ZN(
        n19284) );
  INV_X1 U22167 ( .A(n19284), .ZN(n19223) );
  NOR2_X1 U22168 ( .A1(n19284), .A2(n19263), .ZN(n19245) );
  NOR2_X1 U22169 ( .A1(n19509), .A2(n19245), .ZN(n19219) );
  AOI22_X1 U22170 ( .A1(n19511), .A2(n19546), .B1(n19510), .B2(n19219), .ZN(
        n19205) );
  OAI21_X1 U22171 ( .B1(n19381), .B2(n19201), .A(n19245), .ZN(n19203) );
  INV_X1 U22172 ( .A(n19202), .ZN(n19289) );
  NAND2_X1 U22173 ( .A1(n19203), .A2(n19289), .ZN(n19220) );
  AOI22_X1 U22174 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19220), .B1(
        n19516), .B2(n19241), .ZN(n19204) );
  OAI211_X1 U22175 ( .C1(n19223), .C2(n19519), .A(n19205), .B(n19204), .ZN(
        P3_U2884) );
  AOI22_X1 U22176 ( .A1(n19521), .A2(n19241), .B1(n19520), .B2(n19219), .ZN(
        n19207) );
  AOI22_X1 U22177 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19220), .B1(
        n19522), .B2(n19546), .ZN(n19206) );
  OAI211_X1 U22178 ( .C1(n19223), .C2(n19525), .A(n19207), .B(n19206), .ZN(
        P3_U2885) );
  AOI22_X1 U22179 ( .A1(n19461), .A2(n19546), .B1(n19526), .B2(n19219), .ZN(
        n19209) );
  AOI22_X1 U22180 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19220), .B1(
        n19527), .B2(n19241), .ZN(n19208) );
  OAI211_X1 U22181 ( .C1(n19223), .C2(n19464), .A(n19209), .B(n19208), .ZN(
        P3_U2886) );
  AOI22_X1 U22182 ( .A1(n19533), .A2(n19219), .B1(n19532), .B2(n19546), .ZN(
        n19211) );
  AOI22_X1 U22183 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19220), .B1(
        n19534), .B2(n19241), .ZN(n19210) );
  OAI211_X1 U22184 ( .C1(n19223), .C2(n19537), .A(n19211), .B(n19210), .ZN(
        P3_U2887) );
  AOI22_X1 U22185 ( .A1(n19539), .A2(n19219), .B1(n19538), .B2(n19546), .ZN(
        n19213) );
  AOI22_X1 U22186 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19220), .B1(
        n19540), .B2(n19241), .ZN(n19212) );
  OAI211_X1 U22187 ( .C1(n19223), .C2(n19543), .A(n19213), .B(n19212), .ZN(
        P3_U2888) );
  AOI22_X1 U22188 ( .A1(n19495), .A2(n19546), .B1(n19545), .B2(n19219), .ZN(
        n19215) );
  AOI22_X1 U22189 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19220), .B1(
        n19284), .B2(n19547), .ZN(n19214) );
  OAI211_X1 U22190 ( .C1(n19499), .C2(n19216), .A(n19215), .B(n19214), .ZN(
        P3_U2889) );
  AOI22_X1 U22191 ( .A1(n19553), .A2(n19241), .B1(n19552), .B2(n19219), .ZN(
        n19218) );
  AOI22_X1 U22192 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19220), .B1(
        n19554), .B2(n19546), .ZN(n19217) );
  OAI211_X1 U22193 ( .C1(n19223), .C2(n19557), .A(n19218), .B(n19217), .ZN(
        P3_U2890) );
  AOI22_X1 U22194 ( .A1(n19561), .A2(n19241), .B1(n19559), .B2(n19219), .ZN(
        n19222) );
  AOI22_X1 U22195 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19220), .B1(
        n19563), .B2(n19546), .ZN(n19221) );
  OAI211_X1 U22196 ( .C1(n19223), .C2(n19568), .A(n19222), .B(n19221), .ZN(
        P3_U2891) );
  INV_X1 U22197 ( .A(n19224), .ZN(n19268) );
  NAND2_X1 U22198 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19268), .ZN(
        n19295) );
  NOR2_X1 U22199 ( .A1(n19509), .A2(n19224), .ZN(n19240) );
  AOI22_X1 U22200 ( .A1(n19263), .A2(n19516), .B1(n19510), .B2(n19240), .ZN(
        n19227) );
  AOI21_X1 U22201 ( .B1(n11853), .B2(n19381), .A(n19405), .ZN(n19315) );
  NAND2_X1 U22202 ( .A1(n19225), .A2(n19315), .ZN(n19242) );
  AOI22_X1 U22203 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19242), .B1(
        n19511), .B2(n19241), .ZN(n19226) );
  OAI211_X1 U22204 ( .C1(n19295), .C2(n19519), .A(n19227), .B(n19226), .ZN(
        P3_U2892) );
  AOI22_X1 U22205 ( .A1(n19263), .A2(n19521), .B1(n19520), .B2(n19240), .ZN(
        n19229) );
  AOI22_X1 U22206 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19242), .B1(
        n19522), .B2(n19241), .ZN(n19228) );
  OAI211_X1 U22207 ( .C1(n19295), .C2(n19525), .A(n19229), .B(n19228), .ZN(
        P3_U2893) );
  AOI22_X1 U22208 ( .A1(n19461), .A2(n19241), .B1(n19526), .B2(n19240), .ZN(
        n19231) );
  AOI22_X1 U22209 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19242), .B1(
        n19263), .B2(n19527), .ZN(n19230) );
  OAI211_X1 U22210 ( .C1(n19295), .C2(n19464), .A(n19231), .B(n19230), .ZN(
        P3_U2894) );
  AOI22_X1 U22211 ( .A1(n19533), .A2(n19240), .B1(n19532), .B2(n19241), .ZN(
        n19233) );
  AOI22_X1 U22212 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19242), .B1(
        n19263), .B2(n19534), .ZN(n19232) );
  OAI211_X1 U22213 ( .C1(n19295), .C2(n19537), .A(n19233), .B(n19232), .ZN(
        P3_U2895) );
  AOI22_X1 U22214 ( .A1(n19263), .A2(n19540), .B1(n19539), .B2(n19240), .ZN(
        n19235) );
  AOI22_X1 U22215 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19242), .B1(
        n19538), .B2(n19241), .ZN(n19234) );
  OAI211_X1 U22216 ( .C1(n19295), .C2(n19543), .A(n19235), .B(n19234), .ZN(
        P3_U2896) );
  AOI22_X1 U22217 ( .A1(n19495), .A2(n19241), .B1(n19545), .B2(n19240), .ZN(
        n19237) );
  INV_X1 U22218 ( .A(n19295), .ZN(n19310) );
  AOI22_X1 U22219 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19242), .B1(
        n19310), .B2(n19547), .ZN(n19236) );
  OAI211_X1 U22220 ( .C1(n19259), .C2(n19499), .A(n19237), .B(n19236), .ZN(
        P3_U2897) );
  AOI22_X1 U22221 ( .A1(n19263), .A2(n19553), .B1(n19552), .B2(n19240), .ZN(
        n19239) );
  AOI22_X1 U22222 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19242), .B1(
        n19554), .B2(n19241), .ZN(n19238) );
  OAI211_X1 U22223 ( .C1(n19295), .C2(n19557), .A(n19239), .B(n19238), .ZN(
        P3_U2898) );
  AOI22_X1 U22224 ( .A1(n19263), .A2(n19561), .B1(n19559), .B2(n19240), .ZN(
        n19244) );
  AOI22_X1 U22225 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19242), .B1(
        n19563), .B2(n19241), .ZN(n19243) );
  OAI211_X1 U22226 ( .C1(n19295), .C2(n19568), .A(n19244), .B(n19243), .ZN(
        P3_U2899) );
  INV_X1 U22227 ( .A(n19575), .ZN(n19427) );
  NAND2_X1 U22228 ( .A1(n19427), .A2(n19316), .ZN(n19306) );
  AOI21_X1 U22229 ( .B1(n19306), .B2(n19295), .A(n19509), .ZN(n19262) );
  AOI22_X1 U22230 ( .A1(n19284), .A2(n19516), .B1(n19510), .B2(n19262), .ZN(
        n19248) );
  AOI221_X1 U22231 ( .B1(n19245), .B2(n19295), .C1(n19381), .C2(n19295), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19246) );
  OAI21_X1 U22232 ( .B1(n19332), .B2(n19246), .A(n19384), .ZN(n19264) );
  AOI22_X1 U22233 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19264), .B1(
        n19332), .B2(n19482), .ZN(n19247) );
  OAI211_X1 U22234 ( .C1(n19259), .C2(n19485), .A(n19248), .B(n19247), .ZN(
        P3_U2900) );
  AOI22_X1 U22235 ( .A1(n19263), .A2(n19522), .B1(n19262), .B2(n19520), .ZN(
        n19250) );
  AOI22_X1 U22236 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19264), .B1(
        n19284), .B2(n19521), .ZN(n19249) );
  OAI211_X1 U22237 ( .C1(n19306), .C2(n19525), .A(n19250), .B(n19249), .ZN(
        P3_U2901) );
  AOI22_X1 U22238 ( .A1(n19284), .A2(n19527), .B1(n19262), .B2(n19526), .ZN(
        n19252) );
  AOI22_X1 U22239 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19264), .B1(
        n19332), .B2(n19528), .ZN(n19251) );
  OAI211_X1 U22240 ( .C1(n19259), .C2(n19531), .A(n19252), .B(n19251), .ZN(
        P3_U2902) );
  AOI22_X1 U22241 ( .A1(n19263), .A2(n19532), .B1(n19262), .B2(n19533), .ZN(
        n19254) );
  AOI22_X1 U22242 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19264), .B1(
        n19284), .B2(n19534), .ZN(n19253) );
  OAI211_X1 U22243 ( .C1(n19306), .C2(n19537), .A(n19254), .B(n19253), .ZN(
        P3_U2903) );
  AOI22_X1 U22244 ( .A1(n19263), .A2(n19538), .B1(n19262), .B2(n19539), .ZN(
        n19256) );
  AOI22_X1 U22245 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19264), .B1(
        n19284), .B2(n19540), .ZN(n19255) );
  OAI211_X1 U22246 ( .C1(n19306), .C2(n19543), .A(n19256), .B(n19255), .ZN(
        P3_U2904) );
  AOI22_X1 U22247 ( .A1(n19284), .A2(n19544), .B1(n19262), .B2(n19545), .ZN(
        n19258) );
  AOI22_X1 U22248 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19264), .B1(
        n19332), .B2(n19547), .ZN(n19257) );
  OAI211_X1 U22249 ( .C1(n19259), .C2(n19551), .A(n19258), .B(n19257), .ZN(
        P3_U2905) );
  AOI22_X1 U22250 ( .A1(n19263), .A2(n19554), .B1(n19262), .B2(n19552), .ZN(
        n19261) );
  AOI22_X1 U22251 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19264), .B1(
        n19284), .B2(n19553), .ZN(n19260) );
  OAI211_X1 U22252 ( .C1(n19306), .C2(n19557), .A(n19261), .B(n19260), .ZN(
        P3_U2906) );
  AOI22_X1 U22253 ( .A1(n19263), .A2(n19563), .B1(n19262), .B2(n19559), .ZN(
        n19266) );
  AOI22_X1 U22254 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19264), .B1(
        n19284), .B2(n19561), .ZN(n19265) );
  OAI211_X1 U22255 ( .C1(n19306), .C2(n19568), .A(n19266), .B(n19265), .ZN(
        P3_U2907) );
  NAND2_X1 U22256 ( .A1(n19316), .A2(n19359), .ZN(n19344) );
  INV_X1 U22257 ( .A(n19316), .ZN(n19267) );
  NOR2_X1 U22258 ( .A1(n19267), .A2(n19451), .ZN(n19283) );
  AOI22_X1 U22259 ( .A1(n19310), .A2(n19516), .B1(n19510), .B2(n19283), .ZN(
        n19270) );
  AOI22_X1 U22260 ( .A1(n19515), .A2(n19268), .B1(n19316), .B2(n19453), .ZN(
        n19285) );
  AOI22_X1 U22261 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19511), .ZN(n19269) );
  OAI211_X1 U22262 ( .C1(n19519), .C2(n19344), .A(n19270), .B(n19269), .ZN(
        P3_U2908) );
  AOI22_X1 U22263 ( .A1(n19310), .A2(n19521), .B1(n19520), .B2(n19283), .ZN(
        n19272) );
  AOI22_X1 U22264 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19522), .ZN(n19271) );
  OAI211_X1 U22265 ( .C1(n19525), .C2(n19344), .A(n19272), .B(n19271), .ZN(
        P3_U2909) );
  AOI22_X1 U22266 ( .A1(n19310), .A2(n19527), .B1(n19526), .B2(n19283), .ZN(
        n19274) );
  AOI22_X1 U22267 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19461), .ZN(n19273) );
  OAI211_X1 U22268 ( .C1(n19464), .C2(n19344), .A(n19274), .B(n19273), .ZN(
        P3_U2910) );
  AOI22_X1 U22269 ( .A1(n19284), .A2(n19532), .B1(n19533), .B2(n19283), .ZN(
        n19276) );
  AOI22_X1 U22270 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19285), .B1(
        n19310), .B2(n19534), .ZN(n19275) );
  OAI211_X1 U22271 ( .C1(n19537), .C2(n19344), .A(n19276), .B(n19275), .ZN(
        P3_U2911) );
  AOI22_X1 U22272 ( .A1(n19284), .A2(n19538), .B1(n19539), .B2(n19283), .ZN(
        n19278) );
  AOI22_X1 U22273 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19285), .B1(
        n19310), .B2(n19540), .ZN(n19277) );
  OAI211_X1 U22274 ( .C1(n19543), .C2(n19344), .A(n19278), .B(n19277), .ZN(
        P3_U2912) );
  AOI22_X1 U22275 ( .A1(n19284), .A2(n19495), .B1(n19545), .B2(n19283), .ZN(
        n19280) );
  AOI22_X1 U22276 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19285), .B1(
        n19547), .B2(n19355), .ZN(n19279) );
  OAI211_X1 U22277 ( .C1(n19295), .C2(n19499), .A(n19280), .B(n19279), .ZN(
        P3_U2913) );
  AOI22_X1 U22278 ( .A1(n19284), .A2(n19554), .B1(n19552), .B2(n19283), .ZN(
        n19282) );
  AOI22_X1 U22279 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19285), .B1(
        n19310), .B2(n19553), .ZN(n19281) );
  OAI211_X1 U22280 ( .C1(n19557), .C2(n19344), .A(n19282), .B(n19281), .ZN(
        P3_U2914) );
  AOI22_X1 U22281 ( .A1(n19310), .A2(n19561), .B1(n19559), .B2(n19283), .ZN(
        n19287) );
  AOI22_X1 U22282 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19563), .ZN(n19286) );
  OAI211_X1 U22283 ( .C1(n19568), .C2(n19344), .A(n19287), .B(n19286), .ZN(
        P3_U2915) );
  NOR2_X1 U22284 ( .A1(n19288), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19361) );
  INV_X1 U22285 ( .A(n19361), .ZN(n19314) );
  NOR2_X2 U22286 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19314), .ZN(
        n19376) );
  NOR2_X1 U22287 ( .A1(n19355), .A2(n19376), .ZN(n19336) );
  NOR2_X1 U22288 ( .A1(n19509), .A2(n19336), .ZN(n19309) );
  AOI22_X1 U22289 ( .A1(n19332), .A2(n19516), .B1(n19510), .B2(n19309), .ZN(
        n19294) );
  INV_X1 U22290 ( .A(n19336), .ZN(n19292) );
  NAND2_X1 U22291 ( .A1(n19306), .A2(n19295), .ZN(n19290) );
  OAI221_X1 U22292 ( .B1(n19292), .B2(n19291), .C1(n19292), .C2(n19290), .A(
        n19289), .ZN(n19311) );
  AOI22_X1 U22293 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19311), .B1(
        n19482), .B2(n19376), .ZN(n19293) );
  OAI211_X1 U22294 ( .C1(n19295), .C2(n19485), .A(n19294), .B(n19293), .ZN(
        P3_U2916) );
  INV_X1 U22295 ( .A(n19376), .ZN(n19351) );
  AOI22_X1 U22296 ( .A1(n19332), .A2(n19521), .B1(n19520), .B2(n19309), .ZN(
        n19297) );
  AOI22_X1 U22297 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19311), .B1(
        n19310), .B2(n19522), .ZN(n19296) );
  OAI211_X1 U22298 ( .C1(n19525), .C2(n19351), .A(n19297), .B(n19296), .ZN(
        P3_U2917) );
  AOI22_X1 U22299 ( .A1(n19310), .A2(n19461), .B1(n19526), .B2(n19309), .ZN(
        n19299) );
  AOI22_X1 U22300 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19311), .B1(
        n19332), .B2(n19527), .ZN(n19298) );
  OAI211_X1 U22301 ( .C1(n19464), .C2(n19351), .A(n19299), .B(n19298), .ZN(
        P3_U2918) );
  AOI22_X1 U22302 ( .A1(n19310), .A2(n19532), .B1(n19533), .B2(n19309), .ZN(
        n19301) );
  AOI22_X1 U22303 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19311), .B1(
        n19332), .B2(n19534), .ZN(n19300) );
  OAI211_X1 U22304 ( .C1(n19537), .C2(n19351), .A(n19301), .B(n19300), .ZN(
        P3_U2919) );
  AOI22_X1 U22305 ( .A1(n19332), .A2(n19540), .B1(n19539), .B2(n19309), .ZN(
        n19303) );
  AOI22_X1 U22306 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19311), .B1(
        n19310), .B2(n19538), .ZN(n19302) );
  OAI211_X1 U22307 ( .C1(n19543), .C2(n19351), .A(n19303), .B(n19302), .ZN(
        P3_U2920) );
  AOI22_X1 U22308 ( .A1(n19310), .A2(n19495), .B1(n19545), .B2(n19309), .ZN(
        n19305) );
  AOI22_X1 U22309 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19311), .B1(
        n19547), .B2(n19376), .ZN(n19304) );
  OAI211_X1 U22310 ( .C1(n19306), .C2(n19499), .A(n19305), .B(n19304), .ZN(
        P3_U2921) );
  AOI22_X1 U22311 ( .A1(n19332), .A2(n19553), .B1(n19552), .B2(n19309), .ZN(
        n19308) );
  AOI22_X1 U22312 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19311), .B1(
        n19310), .B2(n19554), .ZN(n19307) );
  OAI211_X1 U22313 ( .C1(n19557), .C2(n19351), .A(n19308), .B(n19307), .ZN(
        P3_U2922) );
  AOI22_X1 U22314 ( .A1(n19310), .A2(n19563), .B1(n19559), .B2(n19309), .ZN(
        n19313) );
  AOI22_X1 U22315 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19311), .B1(
        n19332), .B2(n19561), .ZN(n19312) );
  OAI211_X1 U22316 ( .C1(n19568), .C2(n19351), .A(n19313), .B(n19312), .ZN(
        P3_U2923) );
  NAND2_X1 U22317 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19361), .ZN(
        n19397) );
  NOR2_X1 U22318 ( .A1(n19509), .A2(n19314), .ZN(n19331) );
  AOI22_X1 U22319 ( .A1(n19332), .A2(n19511), .B1(n19510), .B2(n19331), .ZN(
        n19318) );
  NAND2_X1 U22320 ( .A1(n19316), .A2(n19315), .ZN(n19333) );
  AOI22_X1 U22321 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19333), .B1(
        n19516), .B2(n19355), .ZN(n19317) );
  OAI211_X1 U22322 ( .C1(n19519), .C2(n19397), .A(n19318), .B(n19317), .ZN(
        P3_U2924) );
  AOI22_X1 U22323 ( .A1(n19332), .A2(n19522), .B1(n19520), .B2(n19331), .ZN(
        n19320) );
  AOI22_X1 U22324 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19333), .B1(
        n19521), .B2(n19355), .ZN(n19319) );
  OAI211_X1 U22325 ( .C1(n19525), .C2(n19397), .A(n19320), .B(n19319), .ZN(
        P3_U2925) );
  AOI22_X1 U22326 ( .A1(n19527), .A2(n19355), .B1(n19526), .B2(n19331), .ZN(
        n19322) );
  AOI22_X1 U22327 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19333), .B1(
        n19332), .B2(n19461), .ZN(n19321) );
  OAI211_X1 U22328 ( .C1(n19464), .C2(n19397), .A(n19322), .B(n19321), .ZN(
        P3_U2926) );
  AOI22_X1 U22329 ( .A1(n19332), .A2(n19532), .B1(n19533), .B2(n19331), .ZN(
        n19324) );
  AOI22_X1 U22330 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19333), .B1(
        n19534), .B2(n19355), .ZN(n19323) );
  OAI211_X1 U22331 ( .C1(n19537), .C2(n19397), .A(n19324), .B(n19323), .ZN(
        P3_U2927) );
  AOI22_X1 U22332 ( .A1(n19540), .A2(n19355), .B1(n19539), .B2(n19331), .ZN(
        n19326) );
  AOI22_X1 U22333 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19333), .B1(
        n19332), .B2(n19538), .ZN(n19325) );
  OAI211_X1 U22334 ( .C1(n19543), .C2(n19397), .A(n19326), .B(n19325), .ZN(
        P3_U2928) );
  AOI22_X1 U22335 ( .A1(n19332), .A2(n19495), .B1(n19545), .B2(n19331), .ZN(
        n19328) );
  AOI22_X1 U22336 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19333), .B1(
        n19547), .B2(n19401), .ZN(n19327) );
  OAI211_X1 U22337 ( .C1(n19499), .C2(n19344), .A(n19328), .B(n19327), .ZN(
        P3_U2929) );
  AOI22_X1 U22338 ( .A1(n19332), .A2(n19554), .B1(n19552), .B2(n19331), .ZN(
        n19330) );
  AOI22_X1 U22339 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19333), .B1(
        n19553), .B2(n19355), .ZN(n19329) );
  OAI211_X1 U22340 ( .C1(n19557), .C2(n19397), .A(n19330), .B(n19329), .ZN(
        P3_U2930) );
  AOI22_X1 U22341 ( .A1(n19332), .A2(n19563), .B1(n19559), .B2(n19331), .ZN(
        n19335) );
  AOI22_X1 U22342 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19333), .B1(
        n19561), .B2(n19355), .ZN(n19334) );
  OAI211_X1 U22343 ( .C1(n19568), .C2(n19397), .A(n19335), .B(n19334), .ZN(
        P3_U2931) );
  NAND2_X1 U22344 ( .A1(n19427), .A2(n19360), .ZN(n19413) );
  NOR2_X1 U22345 ( .A1(n19401), .A2(n19423), .ZN(n19382) );
  NOR2_X1 U22346 ( .A1(n19509), .A2(n19382), .ZN(n19354) );
  AOI22_X1 U22347 ( .A1(n19516), .A2(n19376), .B1(n19510), .B2(n19354), .ZN(
        n19339) );
  OAI21_X1 U22348 ( .B1(n19336), .B2(n19381), .A(n19382), .ZN(n19337) );
  OAI211_X1 U22349 ( .C1(n19423), .C2(n19723), .A(n19384), .B(n19337), .ZN(
        n19356) );
  AOI22_X1 U22350 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19356), .B1(
        n19511), .B2(n19355), .ZN(n19338) );
  OAI211_X1 U22351 ( .C1(n19519), .C2(n19413), .A(n19339), .B(n19338), .ZN(
        P3_U2932) );
  AOI22_X1 U22352 ( .A1(n19521), .A2(n19376), .B1(n19520), .B2(n19354), .ZN(
        n19341) );
  AOI22_X1 U22353 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19356), .B1(
        n19522), .B2(n19355), .ZN(n19340) );
  OAI211_X1 U22354 ( .C1(n19525), .C2(n19413), .A(n19341), .B(n19340), .ZN(
        P3_U2933) );
  AOI22_X1 U22355 ( .A1(n19527), .A2(n19376), .B1(n19526), .B2(n19354), .ZN(
        n19343) );
  AOI22_X1 U22356 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19356), .B1(
        n19528), .B2(n19423), .ZN(n19342) );
  OAI211_X1 U22357 ( .C1(n19531), .C2(n19344), .A(n19343), .B(n19342), .ZN(
        P3_U2934) );
  AOI22_X1 U22358 ( .A1(n19534), .A2(n19376), .B1(n19533), .B2(n19354), .ZN(
        n19346) );
  AOI22_X1 U22359 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19356), .B1(
        n19532), .B2(n19355), .ZN(n19345) );
  OAI211_X1 U22360 ( .C1(n19537), .C2(n19413), .A(n19346), .B(n19345), .ZN(
        P3_U2935) );
  AOI22_X1 U22361 ( .A1(n19539), .A2(n19354), .B1(n19538), .B2(n19355), .ZN(
        n19348) );
  AOI22_X1 U22362 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19356), .B1(
        n19540), .B2(n19376), .ZN(n19347) );
  OAI211_X1 U22363 ( .C1(n19543), .C2(n19413), .A(n19348), .B(n19347), .ZN(
        P3_U2936) );
  AOI22_X1 U22364 ( .A1(n19495), .A2(n19355), .B1(n19545), .B2(n19354), .ZN(
        n19350) );
  AOI22_X1 U22365 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19356), .B1(
        n19547), .B2(n19423), .ZN(n19349) );
  OAI211_X1 U22366 ( .C1(n19499), .C2(n19351), .A(n19350), .B(n19349), .ZN(
        P3_U2937) );
  AOI22_X1 U22367 ( .A1(n19553), .A2(n19376), .B1(n19552), .B2(n19354), .ZN(
        n19353) );
  AOI22_X1 U22368 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19356), .B1(
        n19554), .B2(n19355), .ZN(n19352) );
  OAI211_X1 U22369 ( .C1(n19557), .C2(n19413), .A(n19353), .B(n19352), .ZN(
        P3_U2938) );
  AOI22_X1 U22370 ( .A1(n19561), .A2(n19376), .B1(n19559), .B2(n19354), .ZN(
        n19358) );
  AOI22_X1 U22371 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19356), .B1(
        n19563), .B2(n19355), .ZN(n19357) );
  OAI211_X1 U22372 ( .C1(n19568), .C2(n19413), .A(n19358), .B(n19357), .ZN(
        P3_U2939) );
  NAND2_X1 U22373 ( .A1(n19359), .A2(n19360), .ZN(n19443) );
  INV_X1 U22374 ( .A(n19360), .ZN(n19380) );
  NOR2_X1 U22375 ( .A1(n19380), .A2(n19451), .ZN(n19406) );
  AOI22_X1 U22376 ( .A1(n19516), .A2(n19401), .B1(n19510), .B2(n19406), .ZN(
        n19363) );
  AOI22_X1 U22377 ( .A1(n19515), .A2(n19361), .B1(n19360), .B2(n19453), .ZN(
        n19377) );
  AOI22_X1 U22378 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19377), .B1(
        n19511), .B2(n19376), .ZN(n19362) );
  OAI211_X1 U22379 ( .C1(n19519), .C2(n19443), .A(n19363), .B(n19362), .ZN(
        P3_U2940) );
  AOI22_X1 U22380 ( .A1(n19520), .A2(n19406), .B1(n19522), .B2(n19376), .ZN(
        n19365) );
  AOI22_X1 U22381 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19377), .B1(
        n19521), .B2(n19401), .ZN(n19364) );
  OAI211_X1 U22382 ( .C1(n19525), .C2(n19443), .A(n19365), .B(n19364), .ZN(
        P3_U2941) );
  AOI22_X1 U22383 ( .A1(n19527), .A2(n19401), .B1(n19526), .B2(n19406), .ZN(
        n19367) );
  AOI22_X1 U22384 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19377), .B1(
        n19461), .B2(n19376), .ZN(n19366) );
  OAI211_X1 U22385 ( .C1(n19464), .C2(n19443), .A(n19367), .B(n19366), .ZN(
        P3_U2942) );
  AOI22_X1 U22386 ( .A1(n19534), .A2(n19401), .B1(n19533), .B2(n19406), .ZN(
        n19369) );
  AOI22_X1 U22387 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19377), .B1(
        n19532), .B2(n19376), .ZN(n19368) );
  OAI211_X1 U22388 ( .C1(n19537), .C2(n19443), .A(n19369), .B(n19368), .ZN(
        P3_U2943) );
  AOI22_X1 U22389 ( .A1(n19540), .A2(n19401), .B1(n19539), .B2(n19406), .ZN(
        n19371) );
  AOI22_X1 U22390 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19377), .B1(
        n19538), .B2(n19376), .ZN(n19370) );
  OAI211_X1 U22391 ( .C1(n19543), .C2(n19443), .A(n19371), .B(n19370), .ZN(
        P3_U2944) );
  AOI22_X1 U22392 ( .A1(n19495), .A2(n19376), .B1(n19545), .B2(n19406), .ZN(
        n19373) );
  AOI22_X1 U22393 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19377), .B1(
        n19547), .B2(n19447), .ZN(n19372) );
  OAI211_X1 U22394 ( .C1(n19499), .C2(n19397), .A(n19373), .B(n19372), .ZN(
        P3_U2945) );
  AOI22_X1 U22395 ( .A1(n19552), .A2(n19406), .B1(n19554), .B2(n19376), .ZN(
        n19375) );
  AOI22_X1 U22396 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19377), .B1(
        n19553), .B2(n19401), .ZN(n19374) );
  OAI211_X1 U22397 ( .C1(n19557), .C2(n19443), .A(n19375), .B(n19374), .ZN(
        P3_U2946) );
  AOI22_X1 U22398 ( .A1(n19563), .A2(n19376), .B1(n19559), .B2(n19406), .ZN(
        n19379) );
  AOI22_X1 U22399 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19377), .B1(
        n19561), .B2(n19401), .ZN(n19378) );
  OAI211_X1 U22400 ( .C1(n19568), .C2(n19443), .A(n19379), .B(n19378), .ZN(
        P3_U2947) );
  NOR2_X1 U22401 ( .A1(n11853), .A2(n19380), .ZN(n19455) );
  NAND2_X1 U22402 ( .A1(n11865), .A2(n19455), .ZN(n19458) );
  INV_X1 U22403 ( .A(n19458), .ZN(n19473) );
  NOR2_X1 U22404 ( .A1(n19447), .A2(n19473), .ZN(n19429) );
  NOR2_X1 U22405 ( .A1(n19509), .A2(n19429), .ZN(n19400) );
  AOI22_X1 U22406 ( .A1(n19516), .A2(n19423), .B1(n19510), .B2(n19400), .ZN(
        n19386) );
  OAI21_X1 U22407 ( .B1(n19382), .B2(n19381), .A(n19429), .ZN(n19383) );
  OAI211_X1 U22408 ( .C1(n19473), .C2(n19723), .A(n19384), .B(n19383), .ZN(
        n19402) );
  AOI22_X1 U22409 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19402), .B1(
        n19482), .B2(n19473), .ZN(n19385) );
  OAI211_X1 U22410 ( .C1(n19485), .C2(n19397), .A(n19386), .B(n19385), .ZN(
        P3_U2948) );
  AOI22_X1 U22411 ( .A1(n19520), .A2(n19400), .B1(n19522), .B2(n19401), .ZN(
        n19388) );
  AOI22_X1 U22412 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19402), .B1(
        n19521), .B2(n19423), .ZN(n19387) );
  OAI211_X1 U22413 ( .C1(n19525), .C2(n19458), .A(n19388), .B(n19387), .ZN(
        P3_U2949) );
  AOI22_X1 U22414 ( .A1(n19527), .A2(n19423), .B1(n19526), .B2(n19400), .ZN(
        n19390) );
  AOI22_X1 U22415 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19402), .B1(
        n19528), .B2(n19473), .ZN(n19389) );
  OAI211_X1 U22416 ( .C1(n19531), .C2(n19397), .A(n19390), .B(n19389), .ZN(
        P3_U2950) );
  AOI22_X1 U22417 ( .A1(n19534), .A2(n19423), .B1(n19533), .B2(n19400), .ZN(
        n19392) );
  AOI22_X1 U22418 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19402), .B1(
        n19532), .B2(n19401), .ZN(n19391) );
  OAI211_X1 U22419 ( .C1(n19537), .C2(n19458), .A(n19392), .B(n19391), .ZN(
        P3_U2951) );
  AOI22_X1 U22420 ( .A1(n19540), .A2(n19423), .B1(n19539), .B2(n19400), .ZN(
        n19394) );
  AOI22_X1 U22421 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19402), .B1(
        n19538), .B2(n19401), .ZN(n19393) );
  OAI211_X1 U22422 ( .C1(n19543), .C2(n19458), .A(n19394), .B(n19393), .ZN(
        P3_U2952) );
  AOI22_X1 U22423 ( .A1(n19545), .A2(n19400), .B1(n19544), .B2(n19423), .ZN(
        n19396) );
  AOI22_X1 U22424 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19402), .B1(
        n19547), .B2(n19473), .ZN(n19395) );
  OAI211_X1 U22425 ( .C1(n19551), .C2(n19397), .A(n19396), .B(n19395), .ZN(
        P3_U2953) );
  AOI22_X1 U22426 ( .A1(n19552), .A2(n19400), .B1(n19554), .B2(n19401), .ZN(
        n19399) );
  AOI22_X1 U22427 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19402), .B1(
        n19553), .B2(n19423), .ZN(n19398) );
  OAI211_X1 U22428 ( .C1(n19557), .C2(n19458), .A(n19399), .B(n19398), .ZN(
        P3_U2954) );
  AOI22_X1 U22429 ( .A1(n19563), .A2(n19401), .B1(n19559), .B2(n19400), .ZN(
        n19404) );
  AOI22_X1 U22430 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19402), .B1(
        n19561), .B2(n19423), .ZN(n19403) );
  OAI211_X1 U22431 ( .C1(n19568), .C2(n19458), .A(n19404), .B(n19403), .ZN(
        P3_U2955) );
  AND2_X1 U22432 ( .A1(n19626), .A2(n19455), .ZN(n19422) );
  AOI22_X1 U22433 ( .A1(n19516), .A2(n19447), .B1(n19510), .B2(n19422), .ZN(
        n19408) );
  INV_X1 U22434 ( .A(n19405), .ZN(n19512) );
  AOI22_X1 U22435 ( .A1(n19515), .A2(n19406), .B1(n19512), .B2(n19455), .ZN(
        n19424) );
  NAND2_X1 U22436 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19455), .ZN(
        n19490) );
  INV_X1 U22437 ( .A(n19490), .ZN(n19503) );
  AOI22_X1 U22438 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19424), .B1(
        n19482), .B2(n19503), .ZN(n19407) );
  OAI211_X1 U22439 ( .C1(n19485), .C2(n19413), .A(n19408), .B(n19407), .ZN(
        P3_U2956) );
  AOI22_X1 U22440 ( .A1(n19521), .A2(n19447), .B1(n19520), .B2(n19422), .ZN(
        n19410) );
  AOI22_X1 U22441 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19424), .B1(
        n19522), .B2(n19423), .ZN(n19409) );
  OAI211_X1 U22442 ( .C1(n19525), .C2(n19490), .A(n19410), .B(n19409), .ZN(
        P3_U2957) );
  AOI22_X1 U22443 ( .A1(n19527), .A2(n19447), .B1(n19526), .B2(n19422), .ZN(
        n19412) );
  AOI22_X1 U22444 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19424), .B1(
        n19528), .B2(n19503), .ZN(n19411) );
  OAI211_X1 U22445 ( .C1(n19531), .C2(n19413), .A(n19412), .B(n19411), .ZN(
        P3_U2958) );
  AOI22_X1 U22446 ( .A1(n19534), .A2(n19447), .B1(n19533), .B2(n19422), .ZN(
        n19415) );
  AOI22_X1 U22447 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19424), .B1(
        n19532), .B2(n19423), .ZN(n19414) );
  OAI211_X1 U22448 ( .C1(n19537), .C2(n19490), .A(n19415), .B(n19414), .ZN(
        P3_U2959) );
  AOI22_X1 U22449 ( .A1(n19539), .A2(n19422), .B1(n19538), .B2(n19423), .ZN(
        n19417) );
  AOI22_X1 U22450 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19424), .B1(
        n19540), .B2(n19447), .ZN(n19416) );
  OAI211_X1 U22451 ( .C1(n19543), .C2(n19490), .A(n19417), .B(n19416), .ZN(
        P3_U2960) );
  AOI22_X1 U22452 ( .A1(n19495), .A2(n19423), .B1(n19545), .B2(n19422), .ZN(
        n19419) );
  AOI22_X1 U22453 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19424), .B1(
        n19547), .B2(n19503), .ZN(n19418) );
  OAI211_X1 U22454 ( .C1(n19499), .C2(n19443), .A(n19419), .B(n19418), .ZN(
        P3_U2961) );
  AOI22_X1 U22455 ( .A1(n19553), .A2(n19447), .B1(n19552), .B2(n19422), .ZN(
        n19421) );
  AOI22_X1 U22456 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19424), .B1(
        n19554), .B2(n19423), .ZN(n19420) );
  OAI211_X1 U22457 ( .C1(n19557), .C2(n19490), .A(n19421), .B(n19420), .ZN(
        P3_U2962) );
  AOI22_X1 U22458 ( .A1(n19561), .A2(n19447), .B1(n19559), .B2(n19422), .ZN(
        n19426) );
  AOI22_X1 U22459 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19424), .B1(
        n19563), .B2(n19423), .ZN(n19425) );
  OAI211_X1 U22460 ( .C1(n19568), .C2(n19490), .A(n19426), .B(n19425), .ZN(
        P3_U2963) );
  INV_X1 U22461 ( .A(n19452), .ZN(n19454) );
  NAND2_X1 U22462 ( .A1(n19427), .A2(n19454), .ZN(n19550) );
  INV_X1 U22463 ( .A(n19550), .ZN(n19562) );
  NOR2_X1 U22464 ( .A1(n19503), .A2(n19562), .ZN(n19480) );
  NOR2_X1 U22465 ( .A1(n19509), .A2(n19480), .ZN(n19446) );
  AOI22_X1 U22466 ( .A1(n19511), .A2(n19447), .B1(n19510), .B2(n19446), .ZN(
        n19432) );
  OAI22_X1 U22467 ( .A1(n19429), .A2(n19479), .B1(n19480), .B2(n19428), .ZN(
        n19430) );
  OAI21_X1 U22468 ( .B1(n19562), .B2(n19723), .A(n19430), .ZN(n19448) );
  AOI22_X1 U22469 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19448), .B1(
        n19516), .B2(n19473), .ZN(n19431) );
  OAI211_X1 U22470 ( .C1(n19519), .C2(n19550), .A(n19432), .B(n19431), .ZN(
        P3_U2964) );
  AOI22_X1 U22471 ( .A1(n19520), .A2(n19446), .B1(n19522), .B2(n19447), .ZN(
        n19434) );
  AOI22_X1 U22472 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19448), .B1(
        n19521), .B2(n19473), .ZN(n19433) );
  OAI211_X1 U22473 ( .C1(n19525), .C2(n19550), .A(n19434), .B(n19433), .ZN(
        P3_U2965) );
  AOI22_X1 U22474 ( .A1(n19461), .A2(n19447), .B1(n19526), .B2(n19446), .ZN(
        n19436) );
  AOI22_X1 U22475 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19448), .B1(
        n19527), .B2(n19473), .ZN(n19435) );
  OAI211_X1 U22476 ( .C1(n19464), .C2(n19550), .A(n19436), .B(n19435), .ZN(
        P3_U2966) );
  AOI22_X1 U22477 ( .A1(n19534), .A2(n19473), .B1(n19533), .B2(n19446), .ZN(
        n19438) );
  AOI22_X1 U22478 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19448), .B1(
        n19532), .B2(n19447), .ZN(n19437) );
  OAI211_X1 U22479 ( .C1(n19537), .C2(n19550), .A(n19438), .B(n19437), .ZN(
        P3_U2967) );
  AOI22_X1 U22480 ( .A1(n19540), .A2(n19473), .B1(n19539), .B2(n19446), .ZN(
        n19440) );
  AOI22_X1 U22481 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19448), .B1(
        n19538), .B2(n19447), .ZN(n19439) );
  OAI211_X1 U22482 ( .C1(n19543), .C2(n19550), .A(n19440), .B(n19439), .ZN(
        P3_U2968) );
  AOI22_X1 U22483 ( .A1(n19545), .A2(n19446), .B1(n19544), .B2(n19473), .ZN(
        n19442) );
  AOI22_X1 U22484 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19448), .B1(
        n19547), .B2(n19562), .ZN(n19441) );
  OAI211_X1 U22485 ( .C1(n19551), .C2(n19443), .A(n19442), .B(n19441), .ZN(
        P3_U2969) );
  AOI22_X1 U22486 ( .A1(n19553), .A2(n19473), .B1(n19552), .B2(n19446), .ZN(
        n19445) );
  AOI22_X1 U22487 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19448), .B1(
        n19554), .B2(n19447), .ZN(n19444) );
  OAI211_X1 U22488 ( .C1(n19557), .C2(n19550), .A(n19445), .B(n19444), .ZN(
        P3_U2970) );
  AOI22_X1 U22489 ( .A1(n19563), .A2(n19447), .B1(n19559), .B2(n19446), .ZN(
        n19450) );
  AOI22_X1 U22490 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19448), .B1(
        n19561), .B2(n19473), .ZN(n19449) );
  OAI211_X1 U22491 ( .C1(n19568), .C2(n19550), .A(n19450), .B(n19449), .ZN(
        P3_U2971) );
  NOR2_X1 U22492 ( .A1(n19452), .A2(n19451), .ZN(n19514) );
  AOI22_X1 U22493 ( .A1(n19516), .A2(n19503), .B1(n19510), .B2(n19514), .ZN(
        n19457) );
  AOI22_X1 U22494 ( .A1(n19515), .A2(n19455), .B1(n19454), .B2(n19453), .ZN(
        n19474) );
  AOI22_X1 U22495 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19474), .B1(
        n19482), .B2(n19560), .ZN(n19456) );
  OAI211_X1 U22496 ( .C1(n19485), .C2(n19458), .A(n19457), .B(n19456), .ZN(
        P3_U2972) );
  INV_X1 U22497 ( .A(n19560), .ZN(n19477) );
  AOI22_X1 U22498 ( .A1(n19520), .A2(n19514), .B1(n19522), .B2(n19473), .ZN(
        n19460) );
  AOI22_X1 U22499 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19474), .B1(
        n19521), .B2(n19503), .ZN(n19459) );
  OAI211_X1 U22500 ( .C1(n19525), .C2(n19477), .A(n19460), .B(n19459), .ZN(
        P3_U2973) );
  AOI22_X1 U22501 ( .A1(n19461), .A2(n19473), .B1(n19526), .B2(n19514), .ZN(
        n19463) );
  AOI22_X1 U22502 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19474), .B1(
        n19527), .B2(n19503), .ZN(n19462) );
  OAI211_X1 U22503 ( .C1(n19464), .C2(n19477), .A(n19463), .B(n19462), .ZN(
        P3_U2974) );
  AOI22_X1 U22504 ( .A1(n19533), .A2(n19514), .B1(n19532), .B2(n19473), .ZN(
        n19466) );
  AOI22_X1 U22505 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19474), .B1(
        n19534), .B2(n19503), .ZN(n19465) );
  OAI211_X1 U22506 ( .C1(n19537), .C2(n19477), .A(n19466), .B(n19465), .ZN(
        P3_U2975) );
  AOI22_X1 U22507 ( .A1(n19539), .A2(n19514), .B1(n19538), .B2(n19473), .ZN(
        n19468) );
  AOI22_X1 U22508 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19474), .B1(
        n19540), .B2(n19503), .ZN(n19467) );
  OAI211_X1 U22509 ( .C1(n19543), .C2(n19477), .A(n19468), .B(n19467), .ZN(
        P3_U2976) );
  AOI22_X1 U22510 ( .A1(n19495), .A2(n19473), .B1(n19545), .B2(n19514), .ZN(
        n19470) );
  AOI22_X1 U22511 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19474), .B1(
        n19547), .B2(n19560), .ZN(n19469) );
  OAI211_X1 U22512 ( .C1(n19499), .C2(n19490), .A(n19470), .B(n19469), .ZN(
        P3_U2977) );
  AOI22_X1 U22513 ( .A1(n19553), .A2(n19503), .B1(n19552), .B2(n19514), .ZN(
        n19472) );
  AOI22_X1 U22514 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19474), .B1(
        n19554), .B2(n19473), .ZN(n19471) );
  OAI211_X1 U22515 ( .C1(n19557), .C2(n19477), .A(n19472), .B(n19471), .ZN(
        P3_U2978) );
  AOI22_X1 U22516 ( .A1(n19561), .A2(n19503), .B1(n19559), .B2(n19514), .ZN(
        n19476) );
  AOI22_X1 U22517 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19474), .B1(
        n19563), .B2(n19473), .ZN(n19475) );
  OAI211_X1 U22518 ( .C1(n19568), .C2(n19477), .A(n19476), .B(n19475), .ZN(
        P3_U2979) );
  AOI21_X1 U22519 ( .B1(n19507), .B2(n19477), .A(n19509), .ZN(n19502) );
  AOI22_X1 U22520 ( .A1(n19516), .A2(n19562), .B1(n19510), .B2(n19502), .ZN(
        n19484) );
  OAI21_X1 U22521 ( .B1(n19480), .B2(n19479), .A(n19478), .ZN(n19481) );
  OAI21_X1 U22522 ( .B1(n19496), .B2(n19723), .A(n19481), .ZN(n19504) );
  AOI22_X1 U22523 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19504), .B1(
        n19482), .B2(n19496), .ZN(n19483) );
  OAI211_X1 U22524 ( .C1(n19485), .C2(n19490), .A(n19484), .B(n19483), .ZN(
        P3_U2980) );
  AOI22_X1 U22525 ( .A1(n19521), .A2(n19562), .B1(n19520), .B2(n19502), .ZN(
        n19487) );
  AOI22_X1 U22526 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19504), .B1(
        n19522), .B2(n19503), .ZN(n19486) );
  OAI211_X1 U22527 ( .C1(n19525), .C2(n19507), .A(n19487), .B(n19486), .ZN(
        P3_U2981) );
  AOI22_X1 U22528 ( .A1(n19527), .A2(n19562), .B1(n19526), .B2(n19502), .ZN(
        n19489) );
  AOI22_X1 U22529 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19504), .B1(
        n19528), .B2(n19496), .ZN(n19488) );
  OAI211_X1 U22530 ( .C1(n19531), .C2(n19490), .A(n19489), .B(n19488), .ZN(
        P3_U2982) );
  AOI22_X1 U22531 ( .A1(n19534), .A2(n19562), .B1(n19533), .B2(n19502), .ZN(
        n19492) );
  AOI22_X1 U22532 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19504), .B1(
        n19532), .B2(n19503), .ZN(n19491) );
  OAI211_X1 U22533 ( .C1(n19537), .C2(n19507), .A(n19492), .B(n19491), .ZN(
        P3_U2983) );
  AOI22_X1 U22534 ( .A1(n19540), .A2(n19562), .B1(n19539), .B2(n19502), .ZN(
        n19494) );
  AOI22_X1 U22535 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19504), .B1(
        n19538), .B2(n19503), .ZN(n19493) );
  OAI211_X1 U22536 ( .C1(n19543), .C2(n19507), .A(n19494), .B(n19493), .ZN(
        P3_U2984) );
  AOI22_X1 U22537 ( .A1(n19495), .A2(n19503), .B1(n19545), .B2(n19502), .ZN(
        n19498) );
  AOI22_X1 U22538 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19504), .B1(
        n19547), .B2(n19496), .ZN(n19497) );
  OAI211_X1 U22539 ( .C1(n19499), .C2(n19550), .A(n19498), .B(n19497), .ZN(
        P3_U2985) );
  AOI22_X1 U22540 ( .A1(n19553), .A2(n19562), .B1(n19552), .B2(n19502), .ZN(
        n19501) );
  AOI22_X1 U22541 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19504), .B1(
        n19554), .B2(n19503), .ZN(n19500) );
  OAI211_X1 U22542 ( .C1(n19557), .C2(n19507), .A(n19501), .B(n19500), .ZN(
        P3_U2986) );
  AOI22_X1 U22543 ( .A1(n19561), .A2(n19562), .B1(n19559), .B2(n19502), .ZN(
        n19506) );
  AOI22_X1 U22544 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19504), .B1(
        n19563), .B2(n19503), .ZN(n19505) );
  OAI211_X1 U22545 ( .C1(n19568), .C2(n19507), .A(n19506), .B(n19505), .ZN(
        P3_U2987) );
  INV_X1 U22546 ( .A(n19546), .ZN(n19567) );
  NOR2_X1 U22547 ( .A1(n19509), .A2(n19508), .ZN(n19558) );
  AOI22_X1 U22548 ( .A1(n19511), .A2(n19562), .B1(n19510), .B2(n19558), .ZN(
        n19518) );
  AOI22_X1 U22549 ( .A1(n19515), .A2(n19514), .B1(n19513), .B2(n19512), .ZN(
        n19564) );
  AOI22_X1 U22550 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19564), .B1(
        n19516), .B2(n19560), .ZN(n19517) );
  OAI211_X1 U22551 ( .C1(n19519), .C2(n19567), .A(n19518), .B(n19517), .ZN(
        P3_U2988) );
  AOI22_X1 U22552 ( .A1(n19521), .A2(n19560), .B1(n19520), .B2(n19558), .ZN(
        n19524) );
  AOI22_X1 U22553 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19564), .B1(
        n19522), .B2(n19562), .ZN(n19523) );
  OAI211_X1 U22554 ( .C1(n19525), .C2(n19567), .A(n19524), .B(n19523), .ZN(
        P3_U2989) );
  AOI22_X1 U22555 ( .A1(n19527), .A2(n19560), .B1(n19526), .B2(n19558), .ZN(
        n19530) );
  AOI22_X1 U22556 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19564), .B1(
        n19528), .B2(n19546), .ZN(n19529) );
  OAI211_X1 U22557 ( .C1(n19531), .C2(n19550), .A(n19530), .B(n19529), .ZN(
        P3_U2990) );
  AOI22_X1 U22558 ( .A1(n19533), .A2(n19558), .B1(n19532), .B2(n19562), .ZN(
        n19536) );
  AOI22_X1 U22559 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19564), .B1(
        n19534), .B2(n19560), .ZN(n19535) );
  OAI211_X1 U22560 ( .C1(n19537), .C2(n19567), .A(n19536), .B(n19535), .ZN(
        P3_U2991) );
  AOI22_X1 U22561 ( .A1(n19539), .A2(n19558), .B1(n19538), .B2(n19562), .ZN(
        n19542) );
  AOI22_X1 U22562 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19564), .B1(
        n19540), .B2(n19560), .ZN(n19541) );
  OAI211_X1 U22563 ( .C1(n19543), .C2(n19567), .A(n19542), .B(n19541), .ZN(
        P3_U2992) );
  AOI22_X1 U22564 ( .A1(n19545), .A2(n19558), .B1(n19544), .B2(n19560), .ZN(
        n19549) );
  AOI22_X1 U22565 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19564), .B1(
        n19547), .B2(n19546), .ZN(n19548) );
  OAI211_X1 U22566 ( .C1(n19551), .C2(n19550), .A(n19549), .B(n19548), .ZN(
        P3_U2993) );
  AOI22_X1 U22567 ( .A1(n19553), .A2(n19560), .B1(n19552), .B2(n19558), .ZN(
        n19556) );
  AOI22_X1 U22568 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19564), .B1(
        n19554), .B2(n19562), .ZN(n19555) );
  OAI211_X1 U22569 ( .C1(n19557), .C2(n19567), .A(n19556), .B(n19555), .ZN(
        P3_U2994) );
  AOI22_X1 U22570 ( .A1(n19561), .A2(n19560), .B1(n19559), .B2(n19558), .ZN(
        n19566) );
  AOI22_X1 U22571 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19564), .B1(
        n19563), .B2(n19562), .ZN(n19565) );
  OAI211_X1 U22572 ( .C1(n19568), .C2(n19567), .A(n19566), .B(n19565), .ZN(
        P3_U2995) );
  INV_X1 U22573 ( .A(n19602), .ZN(n19598) );
  NOR2_X1 U22574 ( .A1(n19598), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n19569) );
  AOI21_X1 U22575 ( .B1(n19570), .B2(n19598), .A(n19569), .ZN(n19597) );
  INV_X1 U22576 ( .A(n19597), .ZN(n19579) );
  NAND3_X1 U22577 ( .A1(n19571), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19573) );
  AOI22_X1 U22578 ( .A1(n19574), .A2(n19573), .B1(n11853), .B2(n19572), .ZN(
        n19576) );
  OAI21_X1 U22579 ( .B1(n19576), .B2(n19602), .A(n19575), .ZN(n19577) );
  AOI21_X1 U22580 ( .B1(n19597), .B2(n11856), .A(n19577), .ZN(n19578) );
  AOI211_X1 U22581 ( .C1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n19579), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n19578), .ZN(n19610) );
  INV_X1 U22582 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19609) );
  OAI21_X1 U22583 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19580), .ZN(n19581) );
  OAI211_X1 U22584 ( .C1(n19583), .C2(n19598), .A(n19582), .B(n19581), .ZN(
        n19596) );
  INV_X1 U22585 ( .A(n19584), .ZN(n19594) );
  NOR2_X1 U22586 ( .A1(n19585), .A2(n19586), .ZN(n19591) );
  AND2_X1 U22587 ( .A1(n19588), .A2(n19587), .ZN(n19590) );
  OAI222_X1 U22588 ( .A1(n19594), .A2(n19593), .B1(n19592), .B2(n19591), .C1(
        n19590), .C2(n19589), .ZN(n19734) );
  INV_X1 U22589 ( .A(n19610), .ZN(n19606) );
  AOI21_X1 U22590 ( .B1(n19609), .B2(n11859), .A(n19597), .ZN(n19605) );
  AND2_X1 U22591 ( .A1(n19599), .A2(n19598), .ZN(n19603) );
  NAND2_X1 U22592 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19600), .ZN(
        n19601) );
  OAI22_X1 U22593 ( .A1(n19603), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19602), .B2(n19601), .ZN(n19604) );
  AOI21_X1 U22594 ( .B1(n19606), .B2(n19605), .A(n19604), .ZN(n19607) );
  INV_X1 U22595 ( .A(n19739), .ZN(n19611) );
  INV_X1 U22596 ( .A(n19617), .ZN(n19745) );
  AOI22_X1 U22597 ( .A1(n19612), .A2(n19611), .B1(n19745), .B2(n18573), .ZN(
        n19613) );
  INV_X1 U22598 ( .A(n19613), .ZN(n19620) );
  INV_X1 U22599 ( .A(n19614), .ZN(n19616) );
  OAI211_X1 U22600 ( .C1(n19616), .C2(n19615), .A(n19743), .B(n19624), .ZN(
        n19722) );
  OAI21_X1 U22601 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19617), .A(n19722), 
        .ZN(n19625) );
  NOR2_X1 U22602 ( .A1(n19618), .A2(n19625), .ZN(n19619) );
  MUX2_X1 U22603 ( .A(n19620), .B(n19619), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19622) );
  OAI211_X1 U22604 ( .C1(n19624), .C2(n19623), .A(n19622), .B(n19621), .ZN(
        P3_U2996) );
  NAND2_X1 U22605 ( .A1(n19745), .A2(n18573), .ZN(n19630) );
  NAND4_X1 U22606 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19745), .A4(n19737), .ZN(n19632) );
  INV_X1 U22607 ( .A(n19625), .ZN(n19627) );
  NAND3_X1 U22608 ( .A1(n19628), .A2(n19627), .A3(n19626), .ZN(n19629) );
  NAND4_X1 U22609 ( .A1(n19631), .A2(n19630), .A3(n19632), .A4(n19629), .ZN(
        P3_U2997) );
  AND4_X1 U22610 ( .A1(n19739), .A2(n19633), .A3(n19632), .A4(n19721), .ZN(
        P3_U2998) );
  AND2_X1 U22611 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19717), .ZN(
        P3_U2999) );
  AND2_X1 U22612 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19717), .ZN(
        P3_U3000) );
  AND2_X1 U22613 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19717), .ZN(
        P3_U3001) );
  AND2_X1 U22614 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19717), .ZN(
        P3_U3002) );
  AND2_X1 U22615 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19717), .ZN(
        P3_U3003) );
  AND2_X1 U22616 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19717), .ZN(
        P3_U3004) );
  AND2_X1 U22617 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19717), .ZN(
        P3_U3005) );
  AND2_X1 U22618 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19717), .ZN(
        P3_U3006) );
  AND2_X1 U22619 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19717), .ZN(
        P3_U3007) );
  AND2_X1 U22620 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19717), .ZN(
        P3_U3008) );
  AND2_X1 U22621 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19717), .ZN(
        P3_U3009) );
  AND2_X1 U22622 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19717), .ZN(
        P3_U3010) );
  AND2_X1 U22623 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19717), .ZN(
        P3_U3011) );
  AND2_X1 U22624 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19717), .ZN(
        P3_U3012) );
  AND2_X1 U22625 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19717), .ZN(
        P3_U3013) );
  AND2_X1 U22626 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19717), .ZN(
        P3_U3014) );
  AND2_X1 U22627 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19717), .ZN(
        P3_U3015) );
  AND2_X1 U22628 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19717), .ZN(
        P3_U3016) );
  AND2_X1 U22629 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19717), .ZN(
        P3_U3017) );
  INV_X1 U22630 ( .A(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21630) );
  NOR2_X1 U22631 ( .A1(n21630), .A2(n19720), .ZN(P3_U3018) );
  AND2_X1 U22632 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19717), .ZN(
        P3_U3019) );
  AND2_X1 U22633 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19717), .ZN(
        P3_U3020) );
  AND2_X1 U22634 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19717), .ZN(P3_U3021) );
  AND2_X1 U22635 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19717), .ZN(P3_U3022) );
  AND2_X1 U22636 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19717), .ZN(P3_U3023) );
  AND2_X1 U22637 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19717), .ZN(P3_U3024) );
  AND2_X1 U22638 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19717), .ZN(P3_U3025) );
  AND2_X1 U22639 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19717), .ZN(P3_U3026) );
  AND2_X1 U22640 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19717), .ZN(P3_U3027) );
  AND2_X1 U22641 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19717), .ZN(P3_U3028) );
  NOR2_X1 U22642 ( .A1(n19650), .A2(n21441), .ZN(n19645) );
  INV_X1 U22643 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19637) );
  AOI211_X1 U22644 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n19645), .B(
        n19637), .ZN(n19636) );
  NAND2_X1 U22645 ( .A1(n19745), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19643) );
  AND2_X1 U22646 ( .A1(n19643), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19649) );
  INV_X1 U22647 ( .A(NA), .ZN(n21446) );
  OAI21_X1 U22648 ( .B1(n21446), .B2(n19634), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19648) );
  INV_X1 U22649 ( .A(n19648), .ZN(n19635) );
  OAI22_X1 U22650 ( .A1(n19749), .A2(n19636), .B1(n19649), .B2(n19635), .ZN(
        P3_U3029) );
  NOR2_X1 U22651 ( .A1(n19645), .A2(n19637), .ZN(n19640) );
  NOR2_X1 U22652 ( .A1(n19638), .A2(n21441), .ZN(n19639) );
  AOI22_X1 U22653 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19640), .B1(n19639), 
        .B2(n19650), .ZN(n19642) );
  NAND3_X1 U22654 ( .A1(n19642), .A2(n19641), .A3(n19643), .ZN(P3_U3030) );
  OAI22_X1 U22655 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19643), .ZN(n19644) );
  OAI22_X1 U22656 ( .A1(n19645), .A2(n19644), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19646) );
  OAI22_X1 U22657 ( .A1(n19649), .A2(n19648), .B1(n19647), .B2(n19646), .ZN(
        P3_U3031) );
  OAI222_X1 U22658 ( .A1(n19652), .A2(n19708), .B1(n19651), .B2(n19749), .C1(
        n19653), .C2(n19706), .ZN(P3_U3032) );
  OAI222_X1 U22659 ( .A1(n19706), .A2(n19655), .B1(n19654), .B2(n19749), .C1(
        n19653), .C2(n19708), .ZN(P3_U3033) );
  OAI222_X1 U22660 ( .A1(n19706), .A2(n19656), .B1(n21637), .B2(n19749), .C1(
        n19655), .C2(n19708), .ZN(P3_U3034) );
  OAI222_X1 U22661 ( .A1(n19706), .A2(n19658), .B1(n19657), .B2(n19749), .C1(
        n19656), .C2(n19708), .ZN(P3_U3035) );
  OAI222_X1 U22662 ( .A1(n19706), .A2(n19660), .B1(n19659), .B2(n19749), .C1(
        n19658), .C2(n19708), .ZN(P3_U3036) );
  OAI222_X1 U22663 ( .A1(n19706), .A2(n19662), .B1(n19661), .B2(n19749), .C1(
        n19660), .C2(n19708), .ZN(P3_U3037) );
  INV_X1 U22664 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19664) );
  OAI222_X1 U22665 ( .A1(n19706), .A2(n19664), .B1(n19663), .B2(n19749), .C1(
        n19662), .C2(n19708), .ZN(P3_U3038) );
  OAI222_X1 U22666 ( .A1(n19706), .A2(n19666), .B1(n19665), .B2(n19749), .C1(
        n19664), .C2(n19708), .ZN(P3_U3039) );
  INV_X1 U22667 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19668) );
  OAI222_X1 U22668 ( .A1(n19706), .A2(n19668), .B1(n19667), .B2(n19749), .C1(
        n19666), .C2(n19708), .ZN(P3_U3040) );
  OAI222_X1 U22669 ( .A1(n19706), .A2(n19670), .B1(n19669), .B2(n19749), .C1(
        n19668), .C2(n19708), .ZN(P3_U3041) );
  INV_X1 U22670 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19672) );
  OAI222_X1 U22671 ( .A1(n19706), .A2(n19672), .B1(n19671), .B2(n19749), .C1(
        n19670), .C2(n19708), .ZN(P3_U3042) );
  OAI222_X1 U22672 ( .A1(n19706), .A2(n19673), .B1(n21658), .B2(n19749), .C1(
        n19672), .C2(n19708), .ZN(P3_U3043) );
  OAI222_X1 U22673 ( .A1(n19706), .A2(n19675), .B1(n19674), .B2(n19749), .C1(
        n19673), .C2(n19708), .ZN(P3_U3044) );
  OAI222_X1 U22674 ( .A1(n19706), .A2(n19677), .B1(n19676), .B2(n19749), .C1(
        n19675), .C2(n19708), .ZN(P3_U3045) );
  INV_X1 U22675 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19679) );
  OAI222_X1 U22676 ( .A1(n19706), .A2(n19679), .B1(n19678), .B2(n19749), .C1(
        n19677), .C2(n19708), .ZN(P3_U3046) );
  OAI222_X1 U22677 ( .A1(n19706), .A2(n19681), .B1(n19680), .B2(n19749), .C1(
        n19679), .C2(n19708), .ZN(P3_U3047) );
  OAI222_X1 U22678 ( .A1(n19706), .A2(n19683), .B1(n19682), .B2(n19749), .C1(
        n19681), .C2(n19708), .ZN(P3_U3048) );
  OAI222_X1 U22679 ( .A1(n19706), .A2(n19686), .B1(n19684), .B2(n19749), .C1(
        n19683), .C2(n19708), .ZN(P3_U3049) );
  INV_X1 U22680 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19687) );
  OAI222_X1 U22681 ( .A1(n19686), .A2(n19708), .B1(n19685), .B2(n19749), .C1(
        n19687), .C2(n19706), .ZN(P3_U3050) );
  OAI222_X1 U22682 ( .A1(n19706), .A2(n19690), .B1(n19688), .B2(n19749), .C1(
        n19687), .C2(n19708), .ZN(P3_U3051) );
  OAI222_X1 U22683 ( .A1(n19690), .A2(n19708), .B1(n19689), .B2(n19749), .C1(
        n19691), .C2(n19706), .ZN(P3_U3052) );
  OAI222_X1 U22684 ( .A1(n19706), .A2(n19694), .B1(n19692), .B2(n19749), .C1(
        n19691), .C2(n19708), .ZN(P3_U3053) );
  OAI222_X1 U22685 ( .A1(n19694), .A2(n19708), .B1(n19693), .B2(n19749), .C1(
        n19695), .C2(n19706), .ZN(P3_U3054) );
  OAI222_X1 U22686 ( .A1(n19706), .A2(n19697), .B1(n19696), .B2(n19749), .C1(
        n19695), .C2(n19708), .ZN(P3_U3055) );
  OAI222_X1 U22687 ( .A1(n19706), .A2(n19699), .B1(n19698), .B2(n19749), .C1(
        n19697), .C2(n19708), .ZN(P3_U3056) );
  OAI222_X1 U22688 ( .A1(n19706), .A2(n17190), .B1(n19700), .B2(n19749), .C1(
        n19699), .C2(n19708), .ZN(P3_U3057) );
  OAI222_X1 U22689 ( .A1(n19706), .A2(n19703), .B1(n19701), .B2(n19749), .C1(
        n17190), .C2(n19708), .ZN(P3_U3058) );
  OAI222_X1 U22690 ( .A1(n19703), .A2(n19708), .B1(n19702), .B2(n19749), .C1(
        n19704), .C2(n19706), .ZN(P3_U3059) );
  OAI222_X1 U22691 ( .A1(n19706), .A2(n11958), .B1(n19705), .B2(n19749), .C1(
        n19704), .C2(n19708), .ZN(P3_U3060) );
  OAI222_X1 U22692 ( .A1(n19708), .A2(n11958), .B1(n21675), .B2(n19749), .C1(
        n19707), .C2(n19706), .ZN(P3_U3061) );
  INV_X1 U22693 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19709) );
  AOI22_X1 U22694 ( .A1(n19749), .A2(n19710), .B1(n19709), .B2(n19731), .ZN(
        P3_U3274) );
  INV_X1 U22695 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19725) );
  INV_X1 U22696 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19711) );
  AOI22_X1 U22697 ( .A1(n19749), .A2(n19725), .B1(n19711), .B2(n19731), .ZN(
        P3_U3275) );
  INV_X1 U22698 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19712) );
  AOI22_X1 U22699 ( .A1(n19749), .A2(n19713), .B1(n19712), .B2(n19731), .ZN(
        P3_U3276) );
  INV_X1 U22700 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19728) );
  INV_X1 U22701 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19714) );
  AOI22_X1 U22702 ( .A1(n19749), .A2(n19728), .B1(n19714), .B2(n19731), .ZN(
        P3_U3277) );
  INV_X1 U22703 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19716) );
  INV_X1 U22704 ( .A(n19718), .ZN(n19715) );
  AOI21_X1 U22705 ( .B1(n19717), .B2(n19716), .A(n19715), .ZN(P3_U3280) );
  OAI21_X1 U22706 ( .B1(n19720), .B2(n19719), .A(n19718), .ZN(P3_U3281) );
  OAI221_X1 U22707 ( .B1(n19723), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19723), 
        .C2(n19722), .A(n19721), .ZN(P3_U3282) );
  AOI211_X1 U22708 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19724) );
  AOI21_X1 U22709 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19724), .ZN(n19726) );
  AOI22_X1 U22710 ( .A1(n19730), .A2(n19726), .B1(n19725), .B2(n19727), .ZN(
        P3_U3292) );
  NOR2_X1 U22711 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n19729) );
  AOI22_X1 U22712 ( .A1(n19730), .A2(n19729), .B1(n19728), .B2(n19727), .ZN(
        P3_U3293) );
  INV_X1 U22713 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19732) );
  AOI22_X1 U22714 ( .A1(n19749), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19732), 
        .B2(n19731), .ZN(P3_U3294) );
  MUX2_X1 U22715 ( .A(P3_MORE_REG_SCAN_IN), .B(n19734), .S(n19733), .Z(
        P3_U3295) );
  OAI21_X1 U22716 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19736), .A(n19735), 
        .ZN(n19738) );
  AOI211_X1 U22717 ( .C1(n19752), .C2(n19738), .A(n19745), .B(n19737), .ZN(
        n19741) );
  OAI21_X1 U22718 ( .B1(n19741), .B2(n19740), .A(n19739), .ZN(n19748) );
  OAI22_X1 U22719 ( .A1(n19745), .A2(n19744), .B1(n19743), .B2(n19742), .ZN(
        n19746) );
  NOR2_X1 U22720 ( .A1(n19756), .A2(n19746), .ZN(n19747) );
  MUX2_X1 U22721 ( .A(n19748), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n19747), 
        .Z(P3_U3296) );
  MUX2_X1 U22722 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n19749), .Z(P3_U3297) );
  OAI21_X1 U22723 ( .B1(P3_READREQUEST_REG_SCAN_IN), .B2(n19753), .A(n19751), 
        .ZN(n19750) );
  OAI21_X1 U22724 ( .B1(n19752), .B2(n19751), .A(n19750), .ZN(P3_U3298) );
  NOR2_X1 U22725 ( .A1(n19753), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19755)
         );
  OAI21_X1 U22726 ( .B1(n19756), .B2(n19755), .A(n19754), .ZN(P3_U3299) );
  INV_X1 U22727 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20476) );
  INV_X1 U22728 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19757) );
  NAND2_X1 U22729 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20493), .ZN(n20483) );
  NAND2_X1 U22730 ( .A1(n20476), .A2(n20475), .ZN(n20480) );
  OAI21_X1 U22731 ( .B1(n20476), .B2(n20483), .A(n20480), .ZN(n20560) );
  OAI21_X1 U22732 ( .B1(n20476), .B2(n19757), .A(n20474), .ZN(P2_U2815) );
  NAND2_X1 U22733 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20476), .ZN(n20593) );
  INV_X2 U22734 ( .A(n20593), .ZN(n20542) );
  AOI21_X1 U22735 ( .B1(n20476), .B2(n20493), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19758) );
  AOI22_X1 U22736 ( .A1(n20542), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19758), 
        .B2(n20593), .ZN(P2_U2817) );
  OAI21_X1 U22737 ( .B1(n20487), .B2(BS16), .A(n20560), .ZN(n20558) );
  OAI21_X1 U22738 ( .B1(n20560), .B2(n20615), .A(n20558), .ZN(P2_U2818) );
  NOR4_X1 U22739 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19762) );
  NOR4_X1 U22740 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19761) );
  NOR4_X1 U22741 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19760) );
  NOR4_X1 U22742 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19759) );
  NAND4_X1 U22743 ( .A1(n19762), .A2(n19761), .A3(n19760), .A4(n19759), .ZN(
        n19768) );
  NOR4_X1 U22744 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19766) );
  AOI211_X1 U22745 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19765) );
  NOR4_X1 U22746 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19764) );
  NOR4_X1 U22747 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19763) );
  NAND4_X1 U22748 ( .A1(n19766), .A2(n19765), .A3(n19764), .A4(n19763), .ZN(
        n19767) );
  NOR2_X1 U22749 ( .A1(n19768), .A2(n19767), .ZN(n19776) );
  INV_X1 U22750 ( .A(n19776), .ZN(n19775) );
  NOR2_X1 U22751 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19775), .ZN(n19769) );
  INV_X1 U22752 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20556) );
  AOI22_X1 U22753 ( .A1(n19769), .A2(n19770), .B1(n19775), .B2(n20556), .ZN(
        P2_U2820) );
  OR3_X1 U22754 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19774) );
  INV_X1 U22755 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20554) );
  AOI22_X1 U22756 ( .A1(n19769), .A2(n19774), .B1(n19775), .B2(n20554), .ZN(
        P2_U2821) );
  INV_X1 U22757 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20559) );
  NAND2_X1 U22758 ( .A1(n19769), .A2(n20559), .ZN(n19773) );
  OAI21_X1 U22759 ( .B1(n20494), .B2(n19770), .A(n19776), .ZN(n19771) );
  OAI21_X1 U22760 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19776), .A(n19771), 
        .ZN(n19772) );
  OAI221_X1 U22761 ( .B1(n19773), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19773), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19772), .ZN(P2_U2822) );
  INV_X1 U22762 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20551) );
  OAI221_X1 U22763 ( .B1(n19776), .B2(n20551), .C1(n19775), .C2(n19774), .A(
        n19773), .ZN(P2_U2823) );
  AOI22_X1 U22764 ( .A1(n19777), .A2(n19797), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19796), .ZN(n19782) );
  XOR2_X1 U22765 ( .A(n19779), .B(n19778), .Z(n19780) );
  NAND2_X1 U22766 ( .A1(n19780), .A2(n19798), .ZN(n19781) );
  OAI211_X1 U22767 ( .C1(n19877), .C2(n19803), .A(n19782), .B(n19781), .ZN(
        P2_U2915) );
  INV_X1 U22768 ( .A(n20565), .ZN(n19783) );
  AOI22_X1 U22769 ( .A1(n19783), .A2(n19797), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19796), .ZN(n19788) );
  XNOR2_X1 U22770 ( .A(n19785), .B(n19784), .ZN(n19786) );
  NAND2_X1 U22771 ( .A1(n19786), .A2(n19798), .ZN(n19787) );
  OAI211_X1 U22772 ( .C1(n19871), .C2(n19803), .A(n19788), .B(n19787), .ZN(
        P2_U2916) );
  INV_X1 U22773 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n21642) );
  OAI21_X1 U22774 ( .B1(n19791), .B2(n19790), .A(n19789), .ZN(n19792) );
  AOI222_X1 U22775 ( .A1(n19793), .A2(n19864), .B1(n20576), .B2(n19797), .C1(
        n19792), .C2(n19798), .ZN(n19794) );
  OAI21_X1 U22776 ( .B1(n19795), .B2(n21642), .A(n19794), .ZN(P2_U2917) );
  AOI22_X1 U22777 ( .A1(n19797), .A2(n19800), .B1(n19796), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19802) );
  OAI211_X1 U22778 ( .C1(n19840), .C2(n19800), .A(n19799), .B(n19798), .ZN(
        n19801) );
  OAI211_X1 U22779 ( .C1(n19849), .C2(n19803), .A(n19802), .B(n19801), .ZN(
        P2_U2919) );
  NOR2_X1 U22780 ( .A1(n21639), .A2(n19828), .ZN(P2_U2920) );
  AOI22_X1 U22781 ( .A1(n19833), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19804) );
  OAI21_X1 U22782 ( .B1(n19836), .B2(n13835), .A(n19804), .ZN(P2_U2936) );
  AOI22_X1 U22783 ( .A1(n19833), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19805) );
  OAI21_X1 U22784 ( .B1(n19836), .B2(n19806), .A(n19805), .ZN(P2_U2937) );
  AOI22_X1 U22785 ( .A1(n19833), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19807) );
  OAI21_X1 U22786 ( .B1(n19836), .B2(n19808), .A(n19807), .ZN(P2_U2938) );
  AOI22_X1 U22787 ( .A1(n19833), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19809) );
  OAI21_X1 U22788 ( .B1(n19836), .B2(n19810), .A(n19809), .ZN(P2_U2939) );
  AOI22_X1 U22789 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n19832), .B1(n19833), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n19811) );
  OAI21_X1 U22790 ( .B1(n19836), .B2(n19812), .A(n19811), .ZN(P2_U2940) );
  AOI22_X1 U22791 ( .A1(n19833), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19813) );
  OAI21_X1 U22792 ( .B1(n19836), .B2(n19814), .A(n19813), .ZN(P2_U2941) );
  AOI22_X1 U22793 ( .A1(n19833), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19815) );
  OAI21_X1 U22794 ( .B1(n19836), .B2(n19816), .A(n19815), .ZN(P2_U2942) );
  AOI22_X1 U22795 ( .A1(n19833), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19817) );
  OAI21_X1 U22796 ( .B1(n19836), .B2(n19818), .A(n19817), .ZN(P2_U2943) );
  AOI22_X1 U22797 ( .A1(n19833), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19819) );
  OAI21_X1 U22798 ( .B1(n19836), .B2(n19820), .A(n19819), .ZN(P2_U2944) );
  AOI22_X1 U22799 ( .A1(n19833), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19821) );
  OAI21_X1 U22800 ( .B1(n19836), .B2(n19822), .A(n19821), .ZN(P2_U2945) );
  INV_X1 U22801 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n21674) );
  AOI22_X1 U22802 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19826), .B1(n19832), .B2(
        P2_DATAO_REG_5__SCAN_IN), .ZN(n19823) );
  OAI21_X1 U22803 ( .B1(n21674), .B2(n20611), .A(n19823), .ZN(P2_U2946) );
  INV_X1 U22804 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U22805 ( .A1(n19833), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19824) );
  OAI21_X1 U22806 ( .B1(n19836), .B2(n19825), .A(n19824), .ZN(P2_U2947) );
  AOI22_X1 U22807 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n19826), .B1(n19833), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n19827) );
  OAI21_X1 U22808 ( .B1(n21655), .B2(n19828), .A(n19827), .ZN(P2_U2948) );
  AOI22_X1 U22809 ( .A1(n19833), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19829) );
  OAI21_X1 U22810 ( .B1(n19836), .B2(n21642), .A(n19829), .ZN(P2_U2949) );
  INV_X1 U22811 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19831) );
  AOI22_X1 U22812 ( .A1(n19833), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19830) );
  OAI21_X1 U22813 ( .B1(n19836), .B2(n19831), .A(n19830), .ZN(P2_U2950) );
  INV_X1 U22814 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19835) );
  AOI22_X1 U22815 ( .A1(n19833), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19832), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19834) );
  OAI21_X1 U22816 ( .B1(n19836), .B2(n19835), .A(n19834), .ZN(P2_U2951) );
  AOI22_X1 U22817 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19892), .ZN(n20374) );
  AOI22_X1 U22818 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19892), .ZN(n20424) );
  AND2_X1 U22819 ( .A1(n10578), .A2(n19894), .ZN(n20411) );
  INV_X1 U22820 ( .A(n20411), .ZN(n20242) );
  NOR2_X1 U22821 ( .A1(n20137), .A2(n19970), .ZN(n19850) );
  INV_X1 U22822 ( .A(n19850), .ZN(n19896) );
  OAI22_X1 U22823 ( .A1(n20472), .A2(n20424), .B1(n20242), .B2(n19896), .ZN(
        n19841) );
  INV_X1 U22824 ( .A(n19841), .ZN(n19856) );
  INV_X1 U22825 ( .A(n19940), .ZN(n19842) );
  OAI21_X1 U22826 ( .B1(n20452), .B2(n19842), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19843) );
  NAND2_X1 U22827 ( .A1(n19843), .A2(n20606), .ZN(n19854) );
  INV_X1 U22828 ( .A(n19844), .ZN(n19845) );
  AND2_X1 U22829 ( .A1(n19845), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20463) );
  NOR2_X1 U22830 ( .A1(n20463), .A2(n19850), .ZN(n19853) );
  INV_X1 U22831 ( .A(n19853), .ZN(n19848) );
  INV_X1 U22832 ( .A(n19851), .ZN(n19846) );
  INV_X1 U22833 ( .A(n20606), .ZN(n20570) );
  OAI211_X1 U22834 ( .C1(n19846), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19896), 
        .B(n20570), .ZN(n19847) );
  OAI211_X2 U22835 ( .C1(n19854), .C2(n19848), .A(n20419), .B(n19847), .ZN(
        n19900) );
  OR2_X1 U22836 ( .A1(n19849), .A2(n20328), .ZN(n20243) );
  OAI21_X1 U22837 ( .B1(n19851), .B2(n19850), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19852) );
  OAI21_X2 U22838 ( .B1(n19854), .B2(n19853), .A(n19852), .ZN(n19899) );
  AOI22_X1 U22839 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19900), .B1(
        n20412), .B2(n19899), .ZN(n19855) );
  OAI211_X1 U22840 ( .C1(n20374), .C2(n19940), .A(n19856), .B(n19855), .ZN(
        P2_U3048) );
  INV_X1 U22841 ( .A(n19892), .ZN(n19891) );
  OAI22_X1 U22842 ( .A1(n19857), .A2(n19891), .B1(n16476), .B2(n19889), .ZN(
        n20427) );
  INV_X1 U22843 ( .A(n20425), .ZN(n20254) );
  OAI22_X1 U22844 ( .A1(n20472), .A2(n20341), .B1(n20254), .B2(n19896), .ZN(
        n19858) );
  INV_X1 U22845 ( .A(n19858), .ZN(n19861) );
  AOI22_X1 U22846 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19900), .B1(
        n20426), .B2(n19899), .ZN(n19860) );
  OAI211_X1 U22847 ( .C1(n20430), .C2(n19940), .A(n19861), .B(n19860), .ZN(
        P2_U3049) );
  OAI22_X1 U22848 ( .A1(n16467), .A2(n19891), .B1(n21580), .B2(n19889), .ZN(
        n20433) );
  NAND2_X1 U22849 ( .A1(n19862), .A2(n19894), .ZN(n20377) );
  OAI22_X1 U22850 ( .A1(n20472), .A2(n20381), .B1(n20377), .B2(n19896), .ZN(
        n19863) );
  INV_X1 U22851 ( .A(n19863), .ZN(n19866) );
  AOI22_X1 U22852 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19900), .B1(
        n20432), .B2(n19899), .ZN(n19865) );
  OAI211_X1 U22853 ( .C1(n20436), .C2(n19940), .A(n19866), .B(n19865), .ZN(
        P2_U3050) );
  OAI22_X1 U22854 ( .A1(n19868), .A2(n19889), .B1(n19867), .B2(n19891), .ZN(
        n20439) );
  INV_X1 U22855 ( .A(n20439), .ZN(n20385) );
  AOI22_X1 U22856 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19892), .ZN(n20442) );
  AND2_X1 U22857 ( .A1(n19869), .A2(n19894), .ZN(n20437) );
  INV_X1 U22858 ( .A(n20437), .ZN(n20263) );
  OAI22_X1 U22859 ( .A1(n20472), .A2(n20442), .B1(n20263), .B2(n19896), .ZN(
        n19870) );
  INV_X1 U22860 ( .A(n19870), .ZN(n19873) );
  OR2_X1 U22861 ( .A1(n19871), .A2(n20328), .ZN(n20264) );
  AOI22_X1 U22862 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19900), .B1(
        n20438), .B2(n19899), .ZN(n19872) );
  OAI211_X1 U22863 ( .C1(n20385), .C2(n19940), .A(n19873), .B(n19872), .ZN(
        P2_U3051) );
  AOI22_X1 U22864 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19892), .ZN(n20387) );
  OAI22_X1 U22865 ( .A1(n19874), .A2(n19891), .B1(n16452), .B2(n19889), .ZN(
        n20309) );
  NAND2_X1 U22866 ( .A1(n19875), .A2(n19894), .ZN(n20386) );
  OAI22_X1 U22867 ( .A1(n20472), .A2(n20448), .B1(n20386), .B2(n19896), .ZN(
        n19876) );
  INV_X1 U22868 ( .A(n19876), .ZN(n19879) );
  OR2_X1 U22869 ( .A1(n19877), .A2(n20328), .ZN(n20268) );
  AOI22_X1 U22870 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19900), .B1(
        n20444), .B2(n19899), .ZN(n19878) );
  OAI211_X1 U22871 ( .C1(n20387), .C2(n19940), .A(n19879), .B(n19878), .ZN(
        P2_U3052) );
  AOI22_X1 U22872 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19892), .ZN(n20456) );
  NAND2_X1 U22873 ( .A1(n9594), .A2(n19894), .ZN(n20391) );
  OAI22_X1 U22874 ( .A1(n20472), .A2(n20456), .B1(n20391), .B2(n19896), .ZN(
        n19880) );
  INV_X1 U22875 ( .A(n19880), .ZN(n19883) );
  AOI22_X1 U22876 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19900), .B1(
        n20450), .B2(n19899), .ZN(n19882) );
  OAI211_X1 U22877 ( .C1(n20392), .C2(n19940), .A(n19883), .B(n19882), .ZN(
        P2_U3053) );
  AOI22_X2 U22878 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19892), .ZN(n20462) );
  OAI22_X1 U22879 ( .A1(n19884), .A2(n19891), .B1(n13724), .B2(n19889), .ZN(
        n20459) );
  AND2_X1 U22880 ( .A1(n13347), .A2(n19894), .ZN(n20457) );
  INV_X1 U22881 ( .A(n20457), .ZN(n20277) );
  OAI22_X1 U22882 ( .A1(n20472), .A2(n20354), .B1(n20277), .B2(n19896), .ZN(
        n19885) );
  INV_X1 U22883 ( .A(n19885), .ZN(n19888) );
  AOI22_X1 U22884 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19900), .B1(
        n20458), .B2(n19899), .ZN(n19887) );
  OAI211_X1 U22885 ( .C1(n20462), .C2(n19940), .A(n19888), .B(n19887), .ZN(
        P2_U3054) );
  OAI22_X1 U22886 ( .A1(n16490), .A2(n19891), .B1(n19890), .B2(n19889), .ZN(
        n20356) );
  INV_X1 U22887 ( .A(n20356), .ZN(n20473) );
  AOI22_X1 U22888 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19893), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19892), .ZN(n20408) );
  NAND2_X1 U22889 ( .A1(n19895), .A2(n19894), .ZN(n20401) );
  OAI22_X1 U22890 ( .A1(n20472), .A2(n20408), .B1(n20401), .B2(n19896), .ZN(
        n19897) );
  INV_X1 U22891 ( .A(n19897), .ZN(n19902) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19900), .B1(
        n20465), .B2(n19899), .ZN(n19901) );
  OAI211_X1 U22893 ( .C1(n20473), .C2(n19940), .A(n19902), .B(n19901), .ZN(
        P2_U3055) );
  NAND2_X1 U22894 ( .A1(n19941), .A2(n20591), .ZN(n19909) );
  NOR2_X1 U22895 ( .A1(n20291), .A2(n19909), .ZN(n19912) );
  AND2_X1 U22896 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19934), .ZN(n19903) );
  INV_X1 U22897 ( .A(n19909), .ZN(n19905) );
  AOI21_X1 U22898 ( .B1(n20607), .B2(n19905), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19906) );
  OAI22_X1 U22899 ( .A1(n19935), .A2(n20243), .B1(n20242), .B2(n19934), .ZN(
        n19907) );
  INV_X1 U22900 ( .A(n19907), .ZN(n19915) );
  OR2_X1 U22901 ( .A1(n20567), .A2(n20615), .ZN(n20110) );
  INV_X1 U22902 ( .A(n20110), .ZN(n19973) );
  NAND2_X1 U22903 ( .A1(n19973), .A2(n20136), .ZN(n19910) );
  AOI21_X1 U22904 ( .B1(n19910), .B2(n19909), .A(n19908), .ZN(n19911) );
  INV_X1 U22905 ( .A(n20115), .ZN(n19913) );
  NAND2_X1 U22906 ( .A1(n20136), .A2(n19913), .ZN(n19945) );
  INV_X1 U22907 ( .A(n20374), .ZN(n20421) );
  AOI22_X1 U22908 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19937), .B1(
        n19966), .B2(n20421), .ZN(n19914) );
  OAI211_X1 U22909 ( .C1(n20424), .C2(n19940), .A(n19915), .B(n19914), .ZN(
        P2_U3056) );
  INV_X1 U22910 ( .A(n20426), .ZN(n20255) );
  OAI22_X1 U22911 ( .A1(n19935), .A2(n20255), .B1(n20254), .B2(n19934), .ZN(
        n19916) );
  INV_X1 U22912 ( .A(n19916), .ZN(n19918) );
  INV_X1 U22913 ( .A(n20430), .ZN(n20338) );
  AOI22_X1 U22914 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19937), .B1(
        n19966), .B2(n20338), .ZN(n19917) );
  OAI211_X1 U22915 ( .C1(n20341), .C2(n19940), .A(n19918), .B(n19917), .ZN(
        P2_U3057) );
  INV_X1 U22916 ( .A(n20432), .ZN(n20259) );
  OAI22_X1 U22917 ( .A1(n19935), .A2(n20259), .B1(n20377), .B2(n19934), .ZN(
        n19919) );
  INV_X1 U22918 ( .A(n19919), .ZN(n19921) );
  INV_X1 U22919 ( .A(n20436), .ZN(n20342) );
  AOI22_X1 U22920 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19937), .B1(
        n19966), .B2(n20342), .ZN(n19920) );
  OAI211_X1 U22921 ( .C1(n20381), .C2(n19940), .A(n19921), .B(n19920), .ZN(
        P2_U3058) );
  OAI22_X1 U22922 ( .A1(n19935), .A2(n20264), .B1(n20263), .B2(n19934), .ZN(
        n19922) );
  INV_X1 U22923 ( .A(n19922), .ZN(n19924) );
  AOI22_X1 U22924 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19937), .B1(
        n19966), .B2(n20439), .ZN(n19923) );
  OAI211_X1 U22925 ( .C1(n20442), .C2(n19940), .A(n19924), .B(n19923), .ZN(
        P2_U3059) );
  OAI22_X1 U22926 ( .A1(n19935), .A2(n20268), .B1(n20386), .B2(n19934), .ZN(
        n19925) );
  INV_X1 U22927 ( .A(n19925), .ZN(n19927) );
  INV_X1 U22928 ( .A(n20387), .ZN(n20445) );
  AOI22_X1 U22929 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19937), .B1(
        n19966), .B2(n20445), .ZN(n19926) );
  OAI211_X1 U22930 ( .C1(n20448), .C2(n19940), .A(n19927), .B(n19926), .ZN(
        P2_U3060) );
  INV_X1 U22931 ( .A(n20450), .ZN(n20273) );
  OAI22_X1 U22932 ( .A1(n19935), .A2(n20273), .B1(n20391), .B2(n19934), .ZN(
        n19928) );
  INV_X1 U22933 ( .A(n19928), .ZN(n19930) );
  INV_X1 U22934 ( .A(n20392), .ZN(n20451) );
  AOI22_X1 U22935 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19937), .B1(
        n19966), .B2(n20451), .ZN(n19929) );
  OAI211_X1 U22936 ( .C1(n20456), .C2(n19940), .A(n19930), .B(n19929), .ZN(
        P2_U3061) );
  INV_X1 U22937 ( .A(n20458), .ZN(n20278) );
  OAI22_X1 U22938 ( .A1(n19935), .A2(n20278), .B1(n20277), .B2(n19934), .ZN(
        n19931) );
  INV_X1 U22939 ( .A(n19931), .ZN(n19933) );
  INV_X1 U22940 ( .A(n20462), .ZN(n20351) );
  AOI22_X1 U22941 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19937), .B1(
        n19966), .B2(n20351), .ZN(n19932) );
  OAI211_X1 U22942 ( .C1(n20354), .C2(n19940), .A(n19933), .B(n19932), .ZN(
        P2_U3062) );
  INV_X1 U22943 ( .A(n20465), .ZN(n20283) );
  OAI22_X1 U22944 ( .A1(n19935), .A2(n20283), .B1(n20401), .B2(n19934), .ZN(
        n19936) );
  INV_X1 U22945 ( .A(n19936), .ZN(n19939) );
  AOI22_X1 U22946 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19937), .B1(
        n19966), .B2(n20356), .ZN(n19938) );
  OAI211_X1 U22947 ( .C1(n20408), .C2(n19940), .A(n19939), .B(n19938), .ZN(
        P2_U3063) );
  NAND2_X1 U22948 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19941), .ZN(
        n19980) );
  NOR2_X1 U22949 ( .A1(n19980), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19964) );
  INV_X1 U22950 ( .A(n19964), .ZN(n19946) );
  INV_X1 U22951 ( .A(n20211), .ZN(n19942) );
  NAND2_X1 U22952 ( .A1(n19942), .A2(n19941), .ZN(n19944) );
  AOI22_X1 U22953 ( .A1(n19965), .A2(n20412), .B1(n20411), .B2(n19964), .ZN(
        n19951) );
  OAI221_X1 U22954 ( .B1(n20615), .B2(n20003), .C1(n20615), .C2(n19945), .A(
        n19944), .ZN(n19949) );
  OAI211_X1 U22955 ( .C1(n19947), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19946), 
        .B(n20570), .ZN(n19948) );
  INV_X1 U22956 ( .A(n20424), .ZN(n20363) );
  AOI22_X1 U22957 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n20363), .ZN(n19950) );
  OAI211_X1 U22958 ( .C1(n20374), .C2(n20003), .A(n19951), .B(n19950), .ZN(
        P2_U3064) );
  AOI22_X1 U22959 ( .A1(n19965), .A2(n20426), .B1(n20425), .B2(n19964), .ZN(
        n19953) );
  AOI22_X1 U22960 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n20427), .ZN(n19952) );
  OAI211_X1 U22961 ( .C1(n20430), .C2(n20003), .A(n19953), .B(n19952), .ZN(
        P2_U3065) );
  INV_X1 U22962 ( .A(n20377), .ZN(n20431) );
  AOI22_X1 U22963 ( .A1(n19965), .A2(n20432), .B1(n20431), .B2(n19964), .ZN(
        n19955) );
  AOI22_X1 U22964 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n20433), .ZN(n19954) );
  OAI211_X1 U22965 ( .C1(n20436), .C2(n20003), .A(n19955), .B(n19954), .ZN(
        P2_U3066) );
  AOI22_X1 U22966 ( .A1(n19965), .A2(n20438), .B1(n20437), .B2(n19964), .ZN(
        n19957) );
  INV_X1 U22967 ( .A(n20442), .ZN(n20382) );
  AOI22_X1 U22968 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n20382), .ZN(n19956) );
  OAI211_X1 U22969 ( .C1(n20385), .C2(n20003), .A(n19957), .B(n19956), .ZN(
        P2_U3067) );
  INV_X1 U22970 ( .A(n20386), .ZN(n20443) );
  AOI22_X1 U22971 ( .A1(n19965), .A2(n20444), .B1(n20443), .B2(n19964), .ZN(
        n19959) );
  AOI22_X1 U22972 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n20309), .ZN(n19958) );
  OAI211_X1 U22973 ( .C1(n20387), .C2(n20003), .A(n19959), .B(n19958), .ZN(
        P2_U3068) );
  INV_X1 U22974 ( .A(n20391), .ZN(n20449) );
  AOI22_X1 U22975 ( .A1(n19965), .A2(n20450), .B1(n20449), .B2(n19964), .ZN(
        n19961) );
  INV_X1 U22976 ( .A(n20456), .ZN(n20312) );
  AOI22_X1 U22977 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n20312), .ZN(n19960) );
  OAI211_X1 U22978 ( .C1(n20392), .C2(n20003), .A(n19961), .B(n19960), .ZN(
        P2_U3069) );
  AOI22_X1 U22979 ( .A1(n19965), .A2(n20458), .B1(n20457), .B2(n19964), .ZN(
        n19963) );
  AOI22_X1 U22980 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n20459), .ZN(n19962) );
  OAI211_X1 U22981 ( .C1(n20462), .C2(n20003), .A(n19963), .B(n19962), .ZN(
        P2_U3070) );
  INV_X1 U22982 ( .A(n20401), .ZN(n20464) );
  AOI22_X1 U22983 ( .A1(n19965), .A2(n20465), .B1(n20464), .B2(n19964), .ZN(
        n19969) );
  INV_X1 U22984 ( .A(n20408), .ZN(n20467) );
  AOI22_X1 U22985 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19967), .B1(
        n19966), .B2(n20467), .ZN(n19968) );
  OAI211_X1 U22986 ( .C1(n20473), .C2(n20003), .A(n19969), .B(n19968), .ZN(
        P2_U3071) );
  NOR2_X1 U22987 ( .A1(n20235), .A2(n19970), .ZN(n19977) );
  INV_X1 U22988 ( .A(n19977), .ZN(n20002) );
  OAI22_X1 U22989 ( .A1(n20014), .A2(n20374), .B1(n20002), .B2(n20242), .ZN(
        n19971) );
  INV_X1 U22990 ( .A(n19971), .ZN(n19983) );
  INV_X1 U22991 ( .A(n19978), .ZN(n19972) );
  AOI21_X1 U22992 ( .B1(n19972), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19975) );
  AOI21_X1 U22993 ( .B1(n19973), .B2(n20250), .A(n20570), .ZN(n19976) );
  NAND2_X1 U22994 ( .A1(n19976), .A2(n19980), .ZN(n19974) );
  INV_X1 U22995 ( .A(n19976), .ZN(n19981) );
  OAI21_X1 U22996 ( .B1(n19978), .B2(n19977), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19979) );
  AOI22_X1 U22997 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20006), .B1(
        n20412), .B2(n20005), .ZN(n19982) );
  OAI211_X1 U22998 ( .C1(n20424), .C2(n20003), .A(n19983), .B(n19982), .ZN(
        P2_U3072) );
  OAI22_X1 U22999 ( .A1(n20003), .A2(n20341), .B1(n20002), .B2(n20254), .ZN(
        n19984) );
  INV_X1 U23000 ( .A(n19984), .ZN(n19986) );
  AOI22_X1 U23001 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20006), .B1(
        n20426), .B2(n20005), .ZN(n19985) );
  OAI211_X1 U23002 ( .C1(n20430), .C2(n20014), .A(n19986), .B(n19985), .ZN(
        P2_U3073) );
  OAI22_X1 U23003 ( .A1(n20014), .A2(n20436), .B1(n20002), .B2(n20377), .ZN(
        n19987) );
  INV_X1 U23004 ( .A(n19987), .ZN(n19989) );
  AOI22_X1 U23005 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20006), .B1(
        n20432), .B2(n20005), .ZN(n19988) );
  OAI211_X1 U23006 ( .C1(n20381), .C2(n20003), .A(n19989), .B(n19988), .ZN(
        P2_U3074) );
  OAI22_X1 U23007 ( .A1(n20003), .A2(n20442), .B1(n20002), .B2(n20263), .ZN(
        n19990) );
  INV_X1 U23008 ( .A(n19990), .ZN(n19992) );
  AOI22_X1 U23009 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20006), .B1(
        n20438), .B2(n20005), .ZN(n19991) );
  OAI211_X1 U23010 ( .C1(n20385), .C2(n20014), .A(n19992), .B(n19991), .ZN(
        P2_U3075) );
  OAI22_X1 U23011 ( .A1(n20014), .A2(n20387), .B1(n20002), .B2(n20386), .ZN(
        n19993) );
  INV_X1 U23012 ( .A(n19993), .ZN(n19995) );
  AOI22_X1 U23013 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20006), .B1(
        n20444), .B2(n20005), .ZN(n19994) );
  OAI211_X1 U23014 ( .C1(n20448), .C2(n20003), .A(n19995), .B(n19994), .ZN(
        P2_U3076) );
  OAI22_X1 U23015 ( .A1(n20014), .A2(n20392), .B1(n20002), .B2(n20391), .ZN(
        n19996) );
  INV_X1 U23016 ( .A(n19996), .ZN(n19998) );
  AOI22_X1 U23017 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20006), .B1(
        n20450), .B2(n20005), .ZN(n19997) );
  OAI211_X1 U23018 ( .C1(n20456), .C2(n20003), .A(n19998), .B(n19997), .ZN(
        P2_U3077) );
  OAI22_X1 U23019 ( .A1(n20014), .A2(n20462), .B1(n20002), .B2(n20277), .ZN(
        n19999) );
  INV_X1 U23020 ( .A(n19999), .ZN(n20001) );
  AOI22_X1 U23021 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20006), .B1(
        n20458), .B2(n20005), .ZN(n20000) );
  OAI211_X1 U23022 ( .C1(n20354), .C2(n20003), .A(n20001), .B(n20000), .ZN(
        P2_U3078) );
  OAI22_X1 U23023 ( .A1(n20003), .A2(n20408), .B1(n20002), .B2(n20401), .ZN(
        n20004) );
  INV_X1 U23024 ( .A(n20004), .ZN(n20008) );
  AOI22_X1 U23025 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20006), .B1(
        n20465), .B2(n20005), .ZN(n20007) );
  OAI211_X1 U23026 ( .C1(n20473), .C2(n20014), .A(n20008), .B(n20007), .ZN(
        P2_U3079) );
  AND2_X1 U23027 ( .A1(n20012), .A2(n20011), .ZN(n20299) );
  NAND2_X1 U23028 ( .A1(n20299), .A2(n20574), .ZN(n20019) );
  NOR2_X1 U23029 ( .A1(n20079), .A2(n20137), .ZN(n20035) );
  OAI21_X1 U23030 ( .B1(n20016), .B2(n20035), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20013) );
  AOI22_X1 U23031 ( .A1(n20036), .A2(n20412), .B1(n20411), .B2(n20035), .ZN(
        n20022) );
  INV_X1 U23032 ( .A(n20076), .ZN(n20015) );
  OAI21_X1 U23033 ( .B1(n20037), .B2(n20015), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20018) );
  AOI211_X1 U23034 ( .C1(n20019), .C2(n20018), .A(n20328), .B(n20017), .ZN(
        n20020) );
  AOI22_X1 U23035 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20038), .B1(
        n20037), .B2(n20363), .ZN(n20021) );
  OAI211_X1 U23036 ( .C1(n20374), .C2(n20076), .A(n20022), .B(n20021), .ZN(
        P2_U3080) );
  AOI22_X1 U23037 ( .A1(n20036), .A2(n20426), .B1(n20425), .B2(n20035), .ZN(
        n20024) );
  AOI22_X1 U23038 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20038), .B1(
        n20037), .B2(n20427), .ZN(n20023) );
  OAI211_X1 U23039 ( .C1(n20430), .C2(n20076), .A(n20024), .B(n20023), .ZN(
        P2_U3081) );
  AOI22_X1 U23040 ( .A1(n20036), .A2(n20432), .B1(n20431), .B2(n20035), .ZN(
        n20026) );
  AOI22_X1 U23041 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20038), .B1(
        n20037), .B2(n20433), .ZN(n20025) );
  OAI211_X1 U23042 ( .C1(n20436), .C2(n20076), .A(n20026), .B(n20025), .ZN(
        P2_U3082) );
  AOI22_X1 U23043 ( .A1(n20036), .A2(n20438), .B1(n20437), .B2(n20035), .ZN(
        n20028) );
  AOI22_X1 U23044 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20038), .B1(
        n20037), .B2(n20382), .ZN(n20027) );
  OAI211_X1 U23045 ( .C1(n20385), .C2(n20076), .A(n20028), .B(n20027), .ZN(
        P2_U3083) );
  AOI22_X1 U23046 ( .A1(n20036), .A2(n20444), .B1(n20443), .B2(n20035), .ZN(
        n20030) );
  AOI22_X1 U23047 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20038), .B1(
        n20037), .B2(n20309), .ZN(n20029) );
  OAI211_X1 U23048 ( .C1(n20387), .C2(n20076), .A(n20030), .B(n20029), .ZN(
        P2_U3084) );
  AOI22_X1 U23049 ( .A1(n20036), .A2(n20450), .B1(n20449), .B2(n20035), .ZN(
        n20032) );
  AOI22_X1 U23050 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20038), .B1(
        n20037), .B2(n20312), .ZN(n20031) );
  OAI211_X1 U23051 ( .C1(n20392), .C2(n20076), .A(n20032), .B(n20031), .ZN(
        P2_U3085) );
  AOI22_X1 U23052 ( .A1(n20036), .A2(n20458), .B1(n20457), .B2(n20035), .ZN(
        n20034) );
  AOI22_X1 U23053 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20038), .B1(
        n20037), .B2(n20459), .ZN(n20033) );
  OAI211_X1 U23054 ( .C1(n20462), .C2(n20076), .A(n20034), .B(n20033), .ZN(
        P2_U3086) );
  AOI22_X1 U23055 ( .A1(n20036), .A2(n20465), .B1(n20464), .B2(n20035), .ZN(
        n20040) );
  AOI22_X1 U23056 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20038), .B1(
        n20037), .B2(n20467), .ZN(n20039) );
  OAI211_X1 U23057 ( .C1(n20473), .C2(n20076), .A(n20040), .B(n20039), .ZN(
        P2_U3087) );
  NOR2_X1 U23058 ( .A1(n20079), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20044) );
  INV_X1 U23059 ( .A(n20044), .ZN(n20048) );
  NOR2_X1 U23060 ( .A1(n20291), .A2(n20048), .ZN(n20045) );
  INV_X1 U23061 ( .A(n20045), .ZN(n20070) );
  OAI22_X1 U23062 ( .A1(n20087), .A2(n20374), .B1(n20070), .B2(n20242), .ZN(
        n20041) );
  INV_X1 U23063 ( .A(n20041), .ZN(n20051) );
  OAI21_X1 U23064 ( .B1(n20334), .B2(n20110), .A(n20606), .ZN(n20049) );
  OAI21_X1 U23065 ( .B1(n20046), .B2(n20326), .A(n20607), .ZN(n20042) );
  NAND2_X1 U23066 ( .A1(n20042), .A2(n20070), .ZN(n20043) );
  OAI21_X1 U23067 ( .B1(n20046), .B2(n20045), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20047) );
  AOI22_X1 U23068 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20073), .B1(
        n20412), .B2(n20072), .ZN(n20050) );
  OAI211_X1 U23069 ( .C1(n20424), .C2(n20076), .A(n20051), .B(n20050), .ZN(
        P2_U3088) );
  OAI22_X1 U23070 ( .A1(n20076), .A2(n20341), .B1(n20254), .B2(n20070), .ZN(
        n20052) );
  INV_X1 U23071 ( .A(n20052), .ZN(n20054) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20073), .B1(
        n20426), .B2(n20072), .ZN(n20053) );
  OAI211_X1 U23073 ( .C1(n20430), .C2(n20087), .A(n20054), .B(n20053), .ZN(
        P2_U3089) );
  OAI22_X1 U23074 ( .A1(n20076), .A2(n20381), .B1(n20070), .B2(n20377), .ZN(
        n20055) );
  INV_X1 U23075 ( .A(n20055), .ZN(n20057) );
  AOI22_X1 U23076 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20073), .B1(
        n20432), .B2(n20072), .ZN(n20056) );
  OAI211_X1 U23077 ( .C1(n20436), .C2(n20087), .A(n20057), .B(n20056), .ZN(
        P2_U3090) );
  OAI22_X1 U23078 ( .A1(n20076), .A2(n20442), .B1(n20263), .B2(n20070), .ZN(
        n20058) );
  INV_X1 U23079 ( .A(n20058), .ZN(n20060) );
  AOI22_X1 U23080 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20073), .B1(
        n20438), .B2(n20072), .ZN(n20059) );
  OAI211_X1 U23081 ( .C1(n20385), .C2(n20087), .A(n20060), .B(n20059), .ZN(
        P2_U3091) );
  OAI22_X1 U23082 ( .A1(n20076), .A2(n20448), .B1(n20070), .B2(n20386), .ZN(
        n20061) );
  INV_X1 U23083 ( .A(n20061), .ZN(n20063) );
  AOI22_X1 U23084 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20073), .B1(
        n20444), .B2(n20072), .ZN(n20062) );
  OAI211_X1 U23085 ( .C1(n20387), .C2(n20087), .A(n20063), .B(n20062), .ZN(
        P2_U3092) );
  OAI22_X1 U23086 ( .A1(n20076), .A2(n20456), .B1(n20070), .B2(n20391), .ZN(
        n20064) );
  INV_X1 U23087 ( .A(n20064), .ZN(n20066) );
  AOI22_X1 U23088 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20073), .B1(
        n20450), .B2(n20072), .ZN(n20065) );
  OAI211_X1 U23089 ( .C1(n20392), .C2(n20087), .A(n20066), .B(n20065), .ZN(
        P2_U3093) );
  OAI22_X1 U23090 ( .A1(n20087), .A2(n20462), .B1(n20070), .B2(n20277), .ZN(
        n20067) );
  INV_X1 U23091 ( .A(n20067), .ZN(n20069) );
  AOI22_X1 U23092 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20073), .B1(
        n20458), .B2(n20072), .ZN(n20068) );
  OAI211_X1 U23093 ( .C1(n20354), .C2(n20076), .A(n20069), .B(n20068), .ZN(
        P2_U3094) );
  OAI22_X1 U23094 ( .A1(n20087), .A2(n20473), .B1(n20401), .B2(n20070), .ZN(
        n20071) );
  INV_X1 U23095 ( .A(n20071), .ZN(n20075) );
  AOI22_X1 U23096 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20073), .B1(
        n20465), .B2(n20072), .ZN(n20074) );
  OAI211_X1 U23097 ( .C1(n20408), .C2(n20076), .A(n20075), .B(n20074), .ZN(
        P2_U3095) );
  NOR3_X2 U23098 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20413), .ZN(n20102) );
  OAI21_X1 U23099 ( .B1(n10798), .B2(n20102), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20078) );
  AOI22_X1 U23100 ( .A1(n20103), .A2(n20412), .B1(n20411), .B2(n20102), .ZN(
        n20089) );
  INV_X1 U23101 ( .A(n10798), .ZN(n20080) );
  AOI21_X1 U23102 ( .B1(n20080), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20086) );
  AOI21_X1 U23103 ( .B1(n20087), .B2(n20135), .A(n20615), .ZN(n20081) );
  AOI21_X1 U23104 ( .B1(n20083), .B2(n20082), .A(n20081), .ZN(n20084) );
  INV_X1 U23105 ( .A(n20084), .ZN(n20085) );
  AOI22_X1 U23106 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20105), .B1(
        n20104), .B2(n20363), .ZN(n20088) );
  OAI211_X1 U23107 ( .C1(n20374), .C2(n20135), .A(n20089), .B(n20088), .ZN(
        P2_U3096) );
  AOI22_X1 U23108 ( .A1(n20103), .A2(n20426), .B1(n20425), .B2(n20102), .ZN(
        n20091) );
  AOI22_X1 U23109 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20105), .B1(
        n20104), .B2(n20427), .ZN(n20090) );
  OAI211_X1 U23110 ( .C1(n20430), .C2(n20135), .A(n20091), .B(n20090), .ZN(
        P2_U3097) );
  AOI22_X1 U23111 ( .A1(n20103), .A2(n20432), .B1(n20431), .B2(n20102), .ZN(
        n20093) );
  AOI22_X1 U23112 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20105), .B1(
        n20104), .B2(n20433), .ZN(n20092) );
  OAI211_X1 U23113 ( .C1(n20436), .C2(n20135), .A(n20093), .B(n20092), .ZN(
        P2_U3098) );
  AOI22_X1 U23114 ( .A1(n20103), .A2(n20438), .B1(n20437), .B2(n20102), .ZN(
        n20095) );
  AOI22_X1 U23115 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20105), .B1(
        n20104), .B2(n20382), .ZN(n20094) );
  OAI211_X1 U23116 ( .C1(n20385), .C2(n20135), .A(n20095), .B(n20094), .ZN(
        P2_U3099) );
  AOI22_X1 U23117 ( .A1(n20103), .A2(n20444), .B1(n20443), .B2(n20102), .ZN(
        n20097) );
  AOI22_X1 U23118 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20105), .B1(
        n20104), .B2(n20309), .ZN(n20096) );
  OAI211_X1 U23119 ( .C1(n20387), .C2(n20135), .A(n20097), .B(n20096), .ZN(
        P2_U3100) );
  AOI22_X1 U23120 ( .A1(n20103), .A2(n20450), .B1(n20449), .B2(n20102), .ZN(
        n20099) );
  AOI22_X1 U23121 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20105), .B1(
        n20104), .B2(n20312), .ZN(n20098) );
  OAI211_X1 U23122 ( .C1(n20392), .C2(n20135), .A(n20099), .B(n20098), .ZN(
        P2_U3101) );
  AOI22_X1 U23123 ( .A1(n20103), .A2(n20458), .B1(n20457), .B2(n20102), .ZN(
        n20101) );
  AOI22_X1 U23124 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20105), .B1(
        n20104), .B2(n20459), .ZN(n20100) );
  OAI211_X1 U23125 ( .C1(n20462), .C2(n20135), .A(n20101), .B(n20100), .ZN(
        P2_U3102) );
  AOI22_X1 U23126 ( .A1(n20103), .A2(n20465), .B1(n20464), .B2(n20102), .ZN(
        n20107) );
  AOI22_X1 U23127 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20105), .B1(
        n20104), .B2(n20467), .ZN(n20106) );
  OAI211_X1 U23128 ( .C1(n20473), .C2(n20135), .A(n20107), .B(n20106), .ZN(
        P2_U3103) );
  NOR2_X1 U23129 ( .A1(n20413), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20113) );
  INV_X1 U23130 ( .A(n20113), .ZN(n20109) );
  INV_X1 U23131 ( .A(n20142), .ZN(n20145) );
  AOI22_X1 U23132 ( .A1(n20130), .A2(n20412), .B1(n20145), .B2(n20411), .ZN(
        n20117) );
  INV_X1 U23133 ( .A(n20361), .ZN(n20414) );
  OR2_X1 U23134 ( .A1(n20110), .A2(n20414), .ZN(n20571) );
  INV_X1 U23135 ( .A(n20571), .ZN(n20114) );
  OAI211_X1 U23136 ( .C1(n20111), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20142), 
        .B(n20570), .ZN(n20112) );
  AOI22_X1 U23137 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20132), .B1(
        n20131), .B2(n20421), .ZN(n20116) );
  OAI211_X1 U23138 ( .C1(n20424), .C2(n20135), .A(n20117), .B(n20116), .ZN(
        P2_U3104) );
  AOI22_X1 U23139 ( .A1(n20130), .A2(n20426), .B1(n20145), .B2(n20425), .ZN(
        n20119) );
  AOI22_X1 U23140 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20132), .B1(
        n20131), .B2(n20338), .ZN(n20118) );
  OAI211_X1 U23141 ( .C1(n20341), .C2(n20135), .A(n20119), .B(n20118), .ZN(
        P2_U3105) );
  AOI22_X1 U23142 ( .A1(n20130), .A2(n20432), .B1(n20145), .B2(n20431), .ZN(
        n20121) );
  AOI22_X1 U23143 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20132), .B1(
        n20131), .B2(n20342), .ZN(n20120) );
  OAI211_X1 U23144 ( .C1(n20381), .C2(n20135), .A(n20121), .B(n20120), .ZN(
        P2_U3106) );
  AOI22_X1 U23145 ( .A1(n20130), .A2(n20438), .B1(n20145), .B2(n20437), .ZN(
        n20123) );
  AOI22_X1 U23146 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20132), .B1(
        n20131), .B2(n20439), .ZN(n20122) );
  OAI211_X1 U23147 ( .C1(n20442), .C2(n20135), .A(n20123), .B(n20122), .ZN(
        P2_U3107) );
  AOI22_X1 U23148 ( .A1(n20130), .A2(n20444), .B1(n20145), .B2(n20443), .ZN(
        n20125) );
  AOI22_X1 U23149 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20132), .B1(
        n20131), .B2(n20445), .ZN(n20124) );
  OAI211_X1 U23150 ( .C1(n20448), .C2(n20135), .A(n20125), .B(n20124), .ZN(
        P2_U3108) );
  AOI22_X1 U23151 ( .A1(n20130), .A2(n20450), .B1(n20145), .B2(n20449), .ZN(
        n20127) );
  AOI22_X1 U23152 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20132), .B1(
        n20131), .B2(n20451), .ZN(n20126) );
  OAI211_X1 U23153 ( .C1(n20456), .C2(n20135), .A(n20127), .B(n20126), .ZN(
        P2_U3109) );
  AOI22_X1 U23154 ( .A1(n20130), .A2(n20458), .B1(n20145), .B2(n20457), .ZN(
        n20129) );
  AOI22_X1 U23155 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20132), .B1(
        n20131), .B2(n20351), .ZN(n20128) );
  OAI211_X1 U23156 ( .C1(n20354), .C2(n20135), .A(n20129), .B(n20128), .ZN(
        P2_U3110) );
  AOI22_X1 U23157 ( .A1(n20130), .A2(n20465), .B1(n20145), .B2(n20464), .ZN(
        n20134) );
  AOI22_X1 U23158 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20132), .B1(
        n20131), .B2(n20356), .ZN(n20133) );
  OAI211_X1 U23159 ( .C1(n20408), .C2(n20135), .A(n20134), .B(n20133), .ZN(
        P2_U3111) );
  NAND2_X1 U23160 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20582), .ZN(
        n20238) );
  NOR2_X1 U23161 ( .A1(n20137), .A2(n20238), .ZN(n20157) );
  INV_X1 U23162 ( .A(n20157), .ZN(n20170) );
  OAI22_X1 U23163 ( .A1(n20176), .A2(n20424), .B1(n20242), .B2(n20170), .ZN(
        n20138) );
  INV_X1 U23164 ( .A(n20138), .ZN(n20150) );
  AOI21_X1 U23165 ( .B1(n20176), .B2(n20208), .A(n20615), .ZN(n20139) );
  NOR2_X1 U23166 ( .A1(n20139), .A2(n20570), .ZN(n20144) );
  INV_X1 U23167 ( .A(n20140), .ZN(n20146) );
  OAI21_X1 U23168 ( .B1(n20146), .B2(n20326), .A(n20607), .ZN(n20141) );
  AOI21_X1 U23169 ( .B1(n20144), .B2(n20142), .A(n20141), .ZN(n20143) );
  OAI21_X2 U23170 ( .B1(n20157), .B2(n20143), .A(n20419), .ZN(n20173) );
  OAI21_X1 U23171 ( .B1(n20145), .B2(n20157), .A(n20144), .ZN(n20148) );
  OAI21_X1 U23172 ( .B1(n20146), .B2(n20157), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20147) );
  AOI22_X1 U23173 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20173), .B1(
        n20412), .B2(n20172), .ZN(n20149) );
  OAI211_X1 U23174 ( .C1(n20374), .C2(n20208), .A(n20150), .B(n20149), .ZN(
        P2_U3112) );
  OAI22_X1 U23175 ( .A1(n20176), .A2(n20341), .B1(n20254), .B2(n20170), .ZN(
        n20151) );
  INV_X1 U23176 ( .A(n20151), .ZN(n20153) );
  AOI22_X1 U23177 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20173), .B1(
        n20426), .B2(n20172), .ZN(n20152) );
  OAI211_X1 U23178 ( .C1(n20430), .C2(n20208), .A(n20153), .B(n20152), .ZN(
        P2_U3113) );
  OAI22_X1 U23179 ( .A1(n20176), .A2(n20381), .B1(n20377), .B2(n20170), .ZN(
        n20154) );
  INV_X1 U23180 ( .A(n20154), .ZN(n20156) );
  AOI22_X1 U23181 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20173), .B1(
        n20432), .B2(n20172), .ZN(n20155) );
  OAI211_X1 U23182 ( .C1(n20436), .C2(n20208), .A(n20156), .B(n20155), .ZN(
        P2_U3114) );
  INV_X1 U23183 ( .A(n20208), .ZN(n20158) );
  AOI22_X1 U23184 ( .A1(n20158), .A2(n20439), .B1(n20437), .B2(n20157), .ZN(
        n20160) );
  AOI22_X1 U23185 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20173), .B1(
        n20438), .B2(n20172), .ZN(n20159) );
  OAI211_X1 U23186 ( .C1(n20442), .C2(n20176), .A(n20160), .B(n20159), .ZN(
        P2_U3115) );
  OAI22_X1 U23187 ( .A1(n20176), .A2(n20448), .B1(n20386), .B2(n20170), .ZN(
        n20161) );
  INV_X1 U23188 ( .A(n20161), .ZN(n20163) );
  AOI22_X1 U23189 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20173), .B1(
        n20444), .B2(n20172), .ZN(n20162) );
  OAI211_X1 U23190 ( .C1(n20387), .C2(n20208), .A(n20163), .B(n20162), .ZN(
        P2_U3116) );
  OAI22_X1 U23191 ( .A1(n20208), .A2(n20392), .B1(n20391), .B2(n20170), .ZN(
        n20164) );
  INV_X1 U23192 ( .A(n20164), .ZN(n20166) );
  AOI22_X1 U23193 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20173), .B1(
        n20450), .B2(n20172), .ZN(n20165) );
  OAI211_X1 U23194 ( .C1(n20456), .C2(n20176), .A(n20166), .B(n20165), .ZN(
        P2_U3117) );
  OAI22_X1 U23195 ( .A1(n20176), .A2(n20354), .B1(n20170), .B2(n20277), .ZN(
        n20167) );
  INV_X1 U23196 ( .A(n20167), .ZN(n20169) );
  AOI22_X1 U23197 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20173), .B1(
        n20458), .B2(n20172), .ZN(n20168) );
  OAI211_X1 U23198 ( .C1(n20462), .C2(n20208), .A(n20169), .B(n20168), .ZN(
        P2_U3118) );
  OAI22_X1 U23199 ( .A1(n20208), .A2(n20473), .B1(n20401), .B2(n20170), .ZN(
        n20171) );
  INV_X1 U23200 ( .A(n20171), .ZN(n20175) );
  AOI22_X1 U23201 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20173), .B1(
        n20465), .B2(n20172), .ZN(n20174) );
  OAI211_X1 U23202 ( .C1(n20408), .C2(n20176), .A(n20175), .B(n20174), .ZN(
        P2_U3119) );
  NOR3_X2 U23203 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20291), .A3(
        n20238), .ZN(n20212) );
  AOI22_X1 U23204 ( .A1(n20231), .A2(n20421), .B1(n20411), .B2(n20212), .ZN(
        n20187) );
  INV_X1 U23205 ( .A(n20331), .ZN(n20415) );
  OAI21_X1 U23206 ( .B1(n20415), .B2(n20178), .A(n20606), .ZN(n20185) );
  NOR2_X1 U23207 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20238), .ZN(
        n20181) );
  OAI21_X1 U23208 ( .B1(n20182), .B2(n20326), .A(n20607), .ZN(n20179) );
  INV_X1 U23209 ( .A(n20212), .ZN(n20199) );
  NAND2_X1 U23210 ( .A1(n20179), .A2(n20199), .ZN(n20180) );
  INV_X1 U23211 ( .A(n20181), .ZN(n20184) );
  OAI21_X1 U23212 ( .B1(n20182), .B2(n20212), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20183) );
  AOI22_X1 U23213 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20205), .B1(
        n20412), .B2(n20204), .ZN(n20186) );
  OAI211_X1 U23214 ( .C1(n20424), .C2(n20208), .A(n20187), .B(n20186), .ZN(
        P2_U3120) );
  AOI22_X1 U23215 ( .A1(n20231), .A2(n20338), .B1(n20425), .B2(n20212), .ZN(
        n20189) );
  AOI22_X1 U23216 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20205), .B1(
        n20426), .B2(n20204), .ZN(n20188) );
  OAI211_X1 U23217 ( .C1(n20341), .C2(n20208), .A(n20189), .B(n20188), .ZN(
        P2_U3121) );
  AOI22_X1 U23218 ( .A1(n20231), .A2(n20342), .B1(n20431), .B2(n20212), .ZN(
        n20191) );
  AOI22_X1 U23219 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20205), .B1(
        n20432), .B2(n20204), .ZN(n20190) );
  OAI211_X1 U23220 ( .C1(n20381), .C2(n20208), .A(n20191), .B(n20190), .ZN(
        P2_U3122) );
  AOI22_X1 U23221 ( .A1(n20231), .A2(n20439), .B1(n20437), .B2(n20212), .ZN(
        n20193) );
  AOI22_X1 U23222 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20205), .B1(
        n20438), .B2(n20204), .ZN(n20192) );
  OAI211_X1 U23223 ( .C1(n20442), .C2(n20208), .A(n20193), .B(n20192), .ZN(
        P2_U3123) );
  AOI22_X1 U23224 ( .A1(n20231), .A2(n20445), .B1(n20443), .B2(n20212), .ZN(
        n20195) );
  AOI22_X1 U23225 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20205), .B1(
        n20444), .B2(n20204), .ZN(n20194) );
  OAI211_X1 U23226 ( .C1(n20448), .C2(n20208), .A(n20195), .B(n20194), .ZN(
        P2_U3124) );
  INV_X1 U23227 ( .A(n20231), .ZN(n20203) );
  OAI22_X1 U23228 ( .A1(n20208), .A2(n20456), .B1(n20391), .B2(n20199), .ZN(
        n20196) );
  INV_X1 U23229 ( .A(n20196), .ZN(n20198) );
  AOI22_X1 U23230 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20205), .B1(
        n20450), .B2(n20204), .ZN(n20197) );
  OAI211_X1 U23231 ( .C1(n20392), .C2(n20203), .A(n20198), .B(n20197), .ZN(
        P2_U3125) );
  OAI22_X1 U23232 ( .A1(n20208), .A2(n20354), .B1(n20277), .B2(n20199), .ZN(
        n20200) );
  INV_X1 U23233 ( .A(n20200), .ZN(n20202) );
  AOI22_X1 U23234 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20205), .B1(
        n20458), .B2(n20204), .ZN(n20201) );
  OAI211_X1 U23235 ( .C1(n20462), .C2(n20203), .A(n20202), .B(n20201), .ZN(
        P2_U3126) );
  AOI22_X1 U23236 ( .A1(n20231), .A2(n20356), .B1(n20464), .B2(n20212), .ZN(
        n20207) );
  AOI22_X1 U23237 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20205), .B1(
        n20465), .B2(n20204), .ZN(n20206) );
  OAI211_X1 U23238 ( .C1(n20408), .C2(n20208), .A(n20207), .B(n20206), .ZN(
        P2_U3127) );
  NOR3_X2 U23239 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20591), .A3(
        n20238), .ZN(n20229) );
  OAI21_X1 U23240 ( .B1(n20209), .B2(n20229), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20210) );
  AOI22_X1 U23241 ( .A1(n20230), .A2(n20412), .B1(n20411), .B2(n20229), .ZN(
        n20216) );
  AOI221_X1 U23242 ( .B1(n20286), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20231), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n20212), .ZN(n20213) );
  OAI21_X2 U23243 ( .B1(n20214), .B2(n20229), .A(n20419), .ZN(n20232) );
  AOI22_X1 U23244 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20232), .B1(
        n20231), .B2(n20363), .ZN(n20215) );
  OAI211_X1 U23245 ( .C1(n20374), .C2(n20272), .A(n20216), .B(n20215), .ZN(
        P2_U3128) );
  AOI22_X1 U23246 ( .A1(n20230), .A2(n20426), .B1(n20425), .B2(n20229), .ZN(
        n20218) );
  AOI22_X1 U23247 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20232), .B1(
        n20231), .B2(n20427), .ZN(n20217) );
  OAI211_X1 U23248 ( .C1(n20430), .C2(n20272), .A(n20218), .B(n20217), .ZN(
        P2_U3129) );
  AOI22_X1 U23249 ( .A1(n20230), .A2(n20432), .B1(n20431), .B2(n20229), .ZN(
        n20220) );
  AOI22_X1 U23250 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20232), .B1(
        n20231), .B2(n20433), .ZN(n20219) );
  OAI211_X1 U23251 ( .C1(n20436), .C2(n20272), .A(n20220), .B(n20219), .ZN(
        P2_U3130) );
  AOI22_X1 U23252 ( .A1(n20230), .A2(n20438), .B1(n20437), .B2(n20229), .ZN(
        n20222) );
  AOI22_X1 U23253 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20232), .B1(
        n20231), .B2(n20382), .ZN(n20221) );
  OAI211_X1 U23254 ( .C1(n20385), .C2(n20272), .A(n20222), .B(n20221), .ZN(
        P2_U3131) );
  AOI22_X1 U23255 ( .A1(n20230), .A2(n20444), .B1(n20443), .B2(n20229), .ZN(
        n20224) );
  AOI22_X1 U23256 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20232), .B1(
        n20231), .B2(n20309), .ZN(n20223) );
  OAI211_X1 U23257 ( .C1(n20387), .C2(n20272), .A(n20224), .B(n20223), .ZN(
        P2_U3132) );
  AOI22_X1 U23258 ( .A1(n20230), .A2(n20450), .B1(n20449), .B2(n20229), .ZN(
        n20226) );
  AOI22_X1 U23259 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20232), .B1(
        n20231), .B2(n20312), .ZN(n20225) );
  OAI211_X1 U23260 ( .C1(n20392), .C2(n20272), .A(n20226), .B(n20225), .ZN(
        P2_U3133) );
  AOI22_X1 U23261 ( .A1(n20230), .A2(n20458), .B1(n20457), .B2(n20229), .ZN(
        n20228) );
  AOI22_X1 U23262 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20232), .B1(
        n20231), .B2(n20459), .ZN(n20227) );
  OAI211_X1 U23263 ( .C1(n20462), .C2(n20272), .A(n20228), .B(n20227), .ZN(
        P2_U3134) );
  AOI22_X1 U23264 ( .A1(n20230), .A2(n20465), .B1(n20464), .B2(n20229), .ZN(
        n20234) );
  AOI22_X1 U23265 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20232), .B1(
        n20231), .B2(n20467), .ZN(n20233) );
  OAI211_X1 U23266 ( .C1(n20473), .C2(n20272), .A(n20234), .B(n20233), .ZN(
        P2_U3135) );
  NOR2_X1 U23267 ( .A1(n20235), .A2(n20238), .ZN(n20249) );
  OR2_X1 U23268 ( .A1(n20249), .A2(n20326), .ZN(n20236) );
  INV_X1 U23269 ( .A(n20238), .ZN(n20239) );
  NAND2_X1 U23270 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20239), .ZN(
        n20246) );
  OAI21_X1 U23271 ( .B1(n20246), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20326), 
        .ZN(n20240) );
  INV_X1 U23272 ( .A(n20240), .ZN(n20241) );
  INV_X1 U23273 ( .A(n20249), .ZN(n20282) );
  OAI22_X1 U23274 ( .A1(n20284), .A2(n20243), .B1(n20242), .B2(n20282), .ZN(
        n20244) );
  INV_X1 U23275 ( .A(n20244), .ZN(n20253) );
  NAND2_X1 U23276 ( .A1(n20331), .A2(n20250), .ZN(n20247) );
  AOI21_X1 U23277 ( .B1(n20247), .B2(n20246), .A(n20245), .ZN(n20248) );
  AOI22_X1 U23278 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20287), .B1(
        n20319), .B2(n20421), .ZN(n20252) );
  OAI211_X1 U23279 ( .C1(n20424), .C2(n20272), .A(n20253), .B(n20252), .ZN(
        P2_U3136) );
  OAI22_X1 U23280 ( .A1(n20284), .A2(n20255), .B1(n20254), .B2(n20282), .ZN(
        n20256) );
  INV_X1 U23281 ( .A(n20256), .ZN(n20258) );
  AOI22_X1 U23282 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20287), .B1(
        n20286), .B2(n20427), .ZN(n20257) );
  OAI211_X1 U23283 ( .C1(n20430), .C2(n20295), .A(n20258), .B(n20257), .ZN(
        P2_U3137) );
  OAI22_X1 U23284 ( .A1(n20284), .A2(n20259), .B1(n20377), .B2(n20282), .ZN(
        n20260) );
  INV_X1 U23285 ( .A(n20260), .ZN(n20262) );
  AOI22_X1 U23286 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20287), .B1(
        n20286), .B2(n20433), .ZN(n20261) );
  OAI211_X1 U23287 ( .C1(n20436), .C2(n20295), .A(n20262), .B(n20261), .ZN(
        P2_U3138) );
  OAI22_X1 U23288 ( .A1(n20284), .A2(n20264), .B1(n20263), .B2(n20282), .ZN(
        n20265) );
  INV_X1 U23289 ( .A(n20265), .ZN(n20267) );
  AOI22_X1 U23290 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20287), .B1(
        n20319), .B2(n20439), .ZN(n20266) );
  OAI211_X1 U23291 ( .C1(n20442), .C2(n20272), .A(n20267), .B(n20266), .ZN(
        P2_U3139) );
  OAI22_X1 U23292 ( .A1(n20284), .A2(n20268), .B1(n20386), .B2(n20282), .ZN(
        n20269) );
  INV_X1 U23293 ( .A(n20269), .ZN(n20271) );
  AOI22_X1 U23294 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20287), .B1(
        n20319), .B2(n20445), .ZN(n20270) );
  OAI211_X1 U23295 ( .C1(n20448), .C2(n20272), .A(n20271), .B(n20270), .ZN(
        P2_U3140) );
  OAI22_X1 U23296 ( .A1(n20284), .A2(n20273), .B1(n20391), .B2(n20282), .ZN(
        n20274) );
  INV_X1 U23297 ( .A(n20274), .ZN(n20276) );
  AOI22_X1 U23298 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20287), .B1(
        n20286), .B2(n20312), .ZN(n20275) );
  OAI211_X1 U23299 ( .C1(n20392), .C2(n20295), .A(n20276), .B(n20275), .ZN(
        P2_U3141) );
  OAI22_X1 U23300 ( .A1(n20284), .A2(n20278), .B1(n20277), .B2(n20282), .ZN(
        n20279) );
  INV_X1 U23301 ( .A(n20279), .ZN(n20281) );
  AOI22_X1 U23302 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20287), .B1(
        n20286), .B2(n20459), .ZN(n20280) );
  OAI211_X1 U23303 ( .C1(n20462), .C2(n20295), .A(n20281), .B(n20280), .ZN(
        P2_U3142) );
  OAI22_X1 U23304 ( .A1(n20284), .A2(n20283), .B1(n20401), .B2(n20282), .ZN(
        n20285) );
  INV_X1 U23305 ( .A(n20285), .ZN(n20289) );
  AOI22_X1 U23306 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20287), .B1(
        n20286), .B2(n20467), .ZN(n20288) );
  OAI211_X1 U23307 ( .C1(n20473), .C2(n20295), .A(n20289), .B(n20288), .ZN(
        P2_U3143) );
  NOR3_X1 U23308 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20582), .A3(
        n20574), .ZN(n20333) );
  NAND2_X1 U23309 ( .A1(n20333), .A2(n20291), .ZN(n20296) );
  AND2_X1 U23310 ( .A1(n20290), .A2(n20296), .ZN(n20294) );
  NAND3_X1 U23311 ( .A1(n20292), .A2(n20606), .A3(n20299), .ZN(n20293) );
  INV_X1 U23312 ( .A(n20296), .ZN(n20317) );
  AOI22_X1 U23313 ( .A1(n20318), .A2(n20412), .B1(n20411), .B2(n20317), .ZN(
        n20302) );
  AOI21_X1 U23314 ( .B1(n20295), .B2(n20360), .A(n20615), .ZN(n20300) );
  OAI211_X1 U23315 ( .C1(n20290), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20296), 
        .B(n20570), .ZN(n20297) );
  AND2_X1 U23316 ( .A1(n20297), .A2(n20419), .ZN(n20298) );
  OAI211_X1 U23317 ( .C1(n20300), .C2(n20299), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n20298), .ZN(n20320) );
  AOI22_X1 U23318 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20363), .ZN(n20301) );
  OAI211_X1 U23319 ( .C1(n20374), .C2(n20360), .A(n20302), .B(n20301), .ZN(
        P2_U3144) );
  AOI22_X1 U23320 ( .A1(n20318), .A2(n20426), .B1(n20425), .B2(n20317), .ZN(
        n20304) );
  AOI22_X1 U23321 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20427), .ZN(n20303) );
  OAI211_X1 U23322 ( .C1(n20430), .C2(n20360), .A(n20304), .B(n20303), .ZN(
        P2_U3145) );
  AOI22_X1 U23323 ( .A1(n20318), .A2(n20432), .B1(n20431), .B2(n20317), .ZN(
        n20306) );
  AOI22_X1 U23324 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20433), .ZN(n20305) );
  OAI211_X1 U23325 ( .C1(n20436), .C2(n20360), .A(n20306), .B(n20305), .ZN(
        P2_U3146) );
  AOI22_X1 U23326 ( .A1(n20318), .A2(n20438), .B1(n20437), .B2(n20317), .ZN(
        n20308) );
  AOI22_X1 U23327 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20382), .ZN(n20307) );
  OAI211_X1 U23328 ( .C1(n20385), .C2(n20360), .A(n20308), .B(n20307), .ZN(
        P2_U3147) );
  AOI22_X1 U23329 ( .A1(n20318), .A2(n20444), .B1(n20443), .B2(n20317), .ZN(
        n20311) );
  AOI22_X1 U23330 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20309), .ZN(n20310) );
  OAI211_X1 U23331 ( .C1(n20387), .C2(n20360), .A(n20311), .B(n20310), .ZN(
        P2_U3148) );
  AOI22_X1 U23332 ( .A1(n20318), .A2(n20450), .B1(n20449), .B2(n20317), .ZN(
        n20314) );
  AOI22_X1 U23333 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20312), .ZN(n20313) );
  OAI211_X1 U23334 ( .C1(n20392), .C2(n20360), .A(n20314), .B(n20313), .ZN(
        P2_U3149) );
  AOI22_X1 U23335 ( .A1(n20318), .A2(n20458), .B1(n20457), .B2(n20317), .ZN(
        n20316) );
  AOI22_X1 U23336 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20459), .ZN(n20315) );
  OAI211_X1 U23337 ( .C1(n20462), .C2(n20360), .A(n20316), .B(n20315), .ZN(
        P2_U3150) );
  AOI22_X1 U23338 ( .A1(n20318), .A2(n20465), .B1(n20464), .B2(n20317), .ZN(
        n20322) );
  AOI22_X1 U23339 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20320), .B1(
        n20319), .B2(n20467), .ZN(n20321) );
  OAI211_X1 U23340 ( .C1(n20473), .C2(n20360), .A(n20322), .B(n20321), .ZN(
        P2_U3151) );
  INV_X1 U23341 ( .A(n20333), .ZN(n20323) );
  OR2_X1 U23342 ( .A1(n20323), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20325) );
  NAND2_X1 U23343 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20333), .ZN(
        n20329) );
  AOI22_X1 U23344 ( .A1(n20355), .A2(n20412), .B1(n20411), .B2(n20365), .ZN(
        n20337) );
  AOI211_X1 U23345 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20329), .A(n20328), 
        .B(n20327), .ZN(n20330) );
  OAI221_X1 U23346 ( .B1(n20333), .B2(n20332), .C1(n20333), .C2(n20331), .A(
        n20330), .ZN(n20357) );
  AOI22_X1 U23347 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20357), .B1(
        n20397), .B2(n20421), .ZN(n20336) );
  OAI211_X1 U23348 ( .C1(n20424), .C2(n20360), .A(n20337), .B(n20336), .ZN(
        P2_U3152) );
  AOI22_X1 U23349 ( .A1(n20355), .A2(n20426), .B1(n20425), .B2(n20365), .ZN(
        n20340) );
  AOI22_X1 U23350 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20357), .B1(
        n20397), .B2(n20338), .ZN(n20339) );
  OAI211_X1 U23351 ( .C1(n20341), .C2(n20360), .A(n20340), .B(n20339), .ZN(
        P2_U3153) );
  AOI22_X1 U23352 ( .A1(n20355), .A2(n20432), .B1(n20431), .B2(n20365), .ZN(
        n20344) );
  AOI22_X1 U23353 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20357), .B1(
        n20397), .B2(n20342), .ZN(n20343) );
  OAI211_X1 U23354 ( .C1(n20381), .C2(n20360), .A(n20344), .B(n20343), .ZN(
        P2_U3154) );
  AOI22_X1 U23355 ( .A1(n20355), .A2(n20438), .B1(n20437), .B2(n20365), .ZN(
        n20346) );
  AOI22_X1 U23356 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20357), .B1(
        n20397), .B2(n20439), .ZN(n20345) );
  OAI211_X1 U23357 ( .C1(n20442), .C2(n20360), .A(n20346), .B(n20345), .ZN(
        P2_U3155) );
  AOI22_X1 U23358 ( .A1(n20355), .A2(n20444), .B1(n20443), .B2(n20365), .ZN(
        n20348) );
  AOI22_X1 U23359 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20357), .B1(
        n20397), .B2(n20445), .ZN(n20347) );
  OAI211_X1 U23360 ( .C1(n20448), .C2(n20360), .A(n20348), .B(n20347), .ZN(
        P2_U3156) );
  AOI22_X1 U23361 ( .A1(n20355), .A2(n20450), .B1(n20449), .B2(n20365), .ZN(
        n20350) );
  AOI22_X1 U23362 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20357), .B1(
        n20397), .B2(n20451), .ZN(n20349) );
  OAI211_X1 U23363 ( .C1(n20456), .C2(n20360), .A(n20350), .B(n20349), .ZN(
        P2_U3157) );
  AOI22_X1 U23364 ( .A1(n20355), .A2(n20458), .B1(n20457), .B2(n20365), .ZN(
        n20353) );
  AOI22_X1 U23365 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20357), .B1(
        n20397), .B2(n20351), .ZN(n20352) );
  OAI211_X1 U23366 ( .C1(n20354), .C2(n20360), .A(n20353), .B(n20352), .ZN(
        P2_U3158) );
  AOI22_X1 U23367 ( .A1(n20355), .A2(n20465), .B1(n20464), .B2(n20365), .ZN(
        n20359) );
  AOI22_X1 U23368 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20357), .B1(
        n20397), .B2(n20356), .ZN(n20358) );
  OAI211_X1 U23369 ( .C1(n20408), .C2(n20360), .A(n20359), .B(n20358), .ZN(
        P2_U3159) );
  NOR3_X1 U23370 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20574), .A3(
        n20413), .ZN(n20396) );
  AOI22_X1 U23371 ( .A1(n20397), .A2(n20363), .B1(n20411), .B2(n20396), .ZN(
        n20373) );
  OAI21_X1 U23372 ( .B1(n20397), .B2(n20468), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20364) );
  NAND2_X1 U23373 ( .A1(n20364), .A2(n20606), .ZN(n20371) );
  NOR2_X1 U23374 ( .A1(n20396), .A2(n20365), .ZN(n20370) );
  INV_X1 U23375 ( .A(n20370), .ZN(n20368) );
  INV_X1 U23376 ( .A(n20396), .ZN(n20400) );
  OAI211_X1 U23377 ( .C1(n20366), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20400), 
        .B(n20570), .ZN(n20367) );
  OAI21_X1 U23378 ( .B1(n10716), .B2(n20396), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20369) );
  AOI22_X1 U23379 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20404), .B1(
        n20412), .B2(n20403), .ZN(n20372) );
  OAI211_X1 U23380 ( .C1(n20374), .C2(n20455), .A(n20373), .B(n20372), .ZN(
        P2_U3160) );
  AOI22_X1 U23381 ( .A1(n20397), .A2(n20427), .B1(n20425), .B2(n20396), .ZN(
        n20376) );
  AOI22_X1 U23382 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20404), .B1(
        n20426), .B2(n20403), .ZN(n20375) );
  OAI211_X1 U23383 ( .C1(n20430), .C2(n20455), .A(n20376), .B(n20375), .ZN(
        P2_U3161) );
  INV_X1 U23384 ( .A(n20397), .ZN(n20407) );
  OAI22_X1 U23385 ( .A1(n20455), .A2(n20436), .B1(n20377), .B2(n20400), .ZN(
        n20378) );
  INV_X1 U23386 ( .A(n20378), .ZN(n20380) );
  AOI22_X1 U23387 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20404), .B1(
        n20432), .B2(n20403), .ZN(n20379) );
  OAI211_X1 U23388 ( .C1(n20381), .C2(n20407), .A(n20380), .B(n20379), .ZN(
        P2_U3162) );
  AOI22_X1 U23389 ( .A1(n20397), .A2(n20382), .B1(n20437), .B2(n20396), .ZN(
        n20384) );
  AOI22_X1 U23390 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20404), .B1(
        n20438), .B2(n20403), .ZN(n20383) );
  OAI211_X1 U23391 ( .C1(n20385), .C2(n20455), .A(n20384), .B(n20383), .ZN(
        P2_U3163) );
  OAI22_X1 U23392 ( .A1(n20455), .A2(n20387), .B1(n20386), .B2(n20400), .ZN(
        n20388) );
  INV_X1 U23393 ( .A(n20388), .ZN(n20390) );
  AOI22_X1 U23394 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20404), .B1(
        n20444), .B2(n20403), .ZN(n20389) );
  OAI211_X1 U23395 ( .C1(n20448), .C2(n20407), .A(n20390), .B(n20389), .ZN(
        P2_U3164) );
  OAI22_X1 U23396 ( .A1(n20455), .A2(n20392), .B1(n20391), .B2(n20400), .ZN(
        n20393) );
  INV_X1 U23397 ( .A(n20393), .ZN(n20395) );
  AOI22_X1 U23398 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20404), .B1(
        n20450), .B2(n20403), .ZN(n20394) );
  OAI211_X1 U23399 ( .C1(n20456), .C2(n20407), .A(n20395), .B(n20394), .ZN(
        P2_U3165) );
  AOI22_X1 U23400 ( .A1(n20397), .A2(n20459), .B1(n20457), .B2(n20396), .ZN(
        n20399) );
  AOI22_X1 U23401 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20404), .B1(
        n20458), .B2(n20403), .ZN(n20398) );
  OAI211_X1 U23402 ( .C1(n20462), .C2(n20455), .A(n20399), .B(n20398), .ZN(
        P2_U3166) );
  OAI22_X1 U23403 ( .A1(n20455), .A2(n20473), .B1(n20401), .B2(n20400), .ZN(
        n20402) );
  INV_X1 U23404 ( .A(n20402), .ZN(n20406) );
  AOI22_X1 U23405 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20404), .B1(
        n20465), .B2(n20403), .ZN(n20405) );
  OAI211_X1 U23406 ( .C1(n20408), .C2(n20407), .A(n20406), .B(n20405), .ZN(
        P2_U3167) );
  OR2_X1 U23407 ( .A1(n20574), .A2(n20413), .ZN(n20410) );
  OAI21_X1 U23408 ( .B1(n10779), .B2(n20463), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20409) );
  AOI22_X1 U23409 ( .A1(n20466), .A2(n20412), .B1(n20411), .B2(n20463), .ZN(
        n20423) );
  OAI22_X1 U23410 ( .A1(n20415), .A2(n20414), .B1(n20413), .B2(n20574), .ZN(
        n20420) );
  INV_X1 U23411 ( .A(n20463), .ZN(n20416) );
  OAI211_X1 U23412 ( .C1(n20417), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20416), 
        .B(n20570), .ZN(n20418) );
  NAND3_X1 U23413 ( .A1(n20420), .A2(n20419), .A3(n20418), .ZN(n20469) );
  AOI22_X1 U23414 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20469), .B1(
        n20452), .B2(n20421), .ZN(n20422) );
  OAI211_X1 U23415 ( .C1(n20424), .C2(n20455), .A(n20423), .B(n20422), .ZN(
        P2_U3168) );
  AOI22_X1 U23416 ( .A1(n20466), .A2(n20426), .B1(n20425), .B2(n20463), .ZN(
        n20429) );
  AOI22_X1 U23417 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20469), .B1(
        n20468), .B2(n20427), .ZN(n20428) );
  OAI211_X1 U23418 ( .C1(n20430), .C2(n20472), .A(n20429), .B(n20428), .ZN(
        P2_U3169) );
  AOI22_X1 U23419 ( .A1(n20466), .A2(n20432), .B1(n20431), .B2(n20463), .ZN(
        n20435) );
  AOI22_X1 U23420 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20469), .B1(
        n20468), .B2(n20433), .ZN(n20434) );
  OAI211_X1 U23421 ( .C1(n20436), .C2(n20472), .A(n20435), .B(n20434), .ZN(
        P2_U3170) );
  AOI22_X1 U23422 ( .A1(n20466), .A2(n20438), .B1(n20437), .B2(n20463), .ZN(
        n20441) );
  AOI22_X1 U23423 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20469), .B1(
        n20452), .B2(n20439), .ZN(n20440) );
  OAI211_X1 U23424 ( .C1(n20442), .C2(n20455), .A(n20441), .B(n20440), .ZN(
        P2_U3171) );
  AOI22_X1 U23425 ( .A1(n20466), .A2(n20444), .B1(n20443), .B2(n20463), .ZN(
        n20447) );
  AOI22_X1 U23426 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20469), .B1(
        n20452), .B2(n20445), .ZN(n20446) );
  OAI211_X1 U23427 ( .C1(n20448), .C2(n20455), .A(n20447), .B(n20446), .ZN(
        P2_U3172) );
  AOI22_X1 U23428 ( .A1(n20466), .A2(n20450), .B1(n20449), .B2(n20463), .ZN(
        n20454) );
  AOI22_X1 U23429 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20469), .B1(
        n20452), .B2(n20451), .ZN(n20453) );
  OAI211_X1 U23430 ( .C1(n20456), .C2(n20455), .A(n20454), .B(n20453), .ZN(
        P2_U3173) );
  AOI22_X1 U23431 ( .A1(n20466), .A2(n20458), .B1(n20457), .B2(n20463), .ZN(
        n20461) );
  AOI22_X1 U23432 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20469), .B1(
        n20468), .B2(n20459), .ZN(n20460) );
  OAI211_X1 U23433 ( .C1(n20462), .C2(n20472), .A(n20461), .B(n20460), .ZN(
        P2_U3174) );
  AOI22_X1 U23434 ( .A1(n20466), .A2(n20465), .B1(n20464), .B2(n20463), .ZN(
        n20471) );
  AOI22_X1 U23435 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20469), .B1(
        n20468), .B2(n20467), .ZN(n20470) );
  OAI211_X1 U23436 ( .C1(n20473), .C2(n20472), .A(n20471), .B(n20470), .ZN(
        P2_U3175) );
  AND2_X1 U23437 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20474), .ZN(
        P2_U3179) );
  AND2_X1 U23438 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20474), .ZN(
        P2_U3180) );
  AND2_X1 U23439 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20474), .ZN(
        P2_U3181) );
  AND2_X1 U23440 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20474), .ZN(
        P2_U3182) );
  AND2_X1 U23441 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20474), .ZN(
        P2_U3183) );
  AND2_X1 U23442 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20474), .ZN(
        P2_U3184) );
  AND2_X1 U23443 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20474), .ZN(
        P2_U3185) );
  AND2_X1 U23444 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20474), .ZN(
        P2_U3186) );
  AND2_X1 U23445 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20474), .ZN(
        P2_U3187) );
  AND2_X1 U23446 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20474), .ZN(
        P2_U3188) );
  AND2_X1 U23447 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20474), .ZN(
        P2_U3189) );
  AND2_X1 U23448 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20474), .ZN(
        P2_U3190) );
  AND2_X1 U23449 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20474), .ZN(
        P2_U3191) );
  AND2_X1 U23450 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20474), .ZN(
        P2_U3192) );
  AND2_X1 U23451 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20474), .ZN(
        P2_U3193) );
  AND2_X1 U23452 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20474), .ZN(
        P2_U3194) );
  AND2_X1 U23453 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20474), .ZN(
        P2_U3195) );
  AND2_X1 U23454 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20474), .ZN(
        P2_U3196) );
  AND2_X1 U23455 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20474), .ZN(
        P2_U3197) );
  AND2_X1 U23456 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20474), .ZN(
        P2_U3198) );
  AND2_X1 U23457 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20474), .ZN(
        P2_U3199) );
  AND2_X1 U23458 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20474), .ZN(
        P2_U3200) );
  AND2_X1 U23459 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20474), .ZN(P2_U3201) );
  AND2_X1 U23460 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20474), .ZN(P2_U3202) );
  AND2_X1 U23461 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20474), .ZN(P2_U3203) );
  AND2_X1 U23462 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20474), .ZN(P2_U3204) );
  AND2_X1 U23463 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20474), .ZN(P2_U3205) );
  AND2_X1 U23464 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20474), .ZN(P2_U3206) );
  AND2_X1 U23465 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20474), .ZN(P2_U3207) );
  AND2_X1 U23466 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20474), .ZN(P2_U3208) );
  NOR2_X1 U23467 ( .A1(n20475), .A2(n20613), .ZN(n20486) );
  INV_X1 U23468 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20626) );
  OR3_X1 U23469 ( .A1(n20486), .A2(n20626), .A3(n20476), .ZN(n20478) );
  AOI211_X1 U23470 ( .C1(n21441), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n20487), .B(n20542), .ZN(n20477) );
  NOR2_X1 U23471 ( .A1(n21446), .A2(n20480), .ZN(n20492) );
  AOI211_X1 U23472 ( .C1(n20493), .C2(n20478), .A(n20477), .B(n20492), .ZN(
        n20479) );
  INV_X1 U23473 ( .A(n20479), .ZN(P2_U3209) );
  AOI21_X1 U23474 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21441), .A(n20493), 
        .ZN(n20484) );
  NOR2_X1 U23475 ( .A1(n20626), .A2(n20484), .ZN(n20481) );
  AOI21_X1 U23476 ( .B1(n20481), .B2(n20480), .A(n20486), .ZN(n20482) );
  OAI211_X1 U23477 ( .C1(n21441), .C2(n20483), .A(n20482), .B(n20618), .ZN(
        P2_U3210) );
  AOI21_X1 U23478 ( .B1(n20612), .B2(n20485), .A(n20484), .ZN(n20491) );
  AOI22_X1 U23479 ( .A1(n20626), .A2(n20487), .B1(n21446), .B2(n20486), .ZN(
        n20488) );
  INV_X1 U23480 ( .A(n20488), .ZN(n20489) );
  OAI211_X1 U23481 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20489), .ZN(n20490) );
  OAI21_X1 U23482 ( .B1(n20492), .B2(n20491), .A(n20490), .ZN(P2_U3211) );
  NAND2_X1 U23483 ( .A1(n20542), .A2(n20493), .ZN(n20549) );
  CLKBUF_X1 U23484 ( .A(n20549), .Z(n20544) );
  NAND2_X2 U23485 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20542), .ZN(n20545) );
  OAI222_X1 U23486 ( .A1(n20544), .A2(n20496), .B1(n20495), .B2(n20542), .C1(
        n20494), .C2(n20545), .ZN(P2_U3212) );
  OAI222_X1 U23487 ( .A1(n20549), .A2(n20498), .B1(n20497), .B2(n20542), .C1(
        n20496), .C2(n20545), .ZN(P2_U3213) );
  OAI222_X1 U23488 ( .A1(n20549), .A2(n20500), .B1(n20499), .B2(n20542), .C1(
        n20498), .C2(n20545), .ZN(P2_U3214) );
  OAI222_X1 U23489 ( .A1(n20549), .A2(n16279), .B1(n20501), .B2(n20542), .C1(
        n20500), .C2(n20545), .ZN(P2_U3215) );
  OAI222_X1 U23490 ( .A1(n20549), .A2(n20503), .B1(n20502), .B2(n20542), .C1(
        n16279), .C2(n20545), .ZN(P2_U3216) );
  OAI222_X1 U23491 ( .A1(n20549), .A2(n20505), .B1(n20504), .B2(n20542), .C1(
        n20503), .C2(n20545), .ZN(P2_U3217) );
  INV_X1 U23492 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n21646) );
  OAI222_X1 U23493 ( .A1(n20544), .A2(n21646), .B1(n20506), .B2(n20542), .C1(
        n20505), .C2(n20545), .ZN(P2_U3218) );
  OAI222_X1 U23494 ( .A1(n20544), .A2(n20508), .B1(n20507), .B2(n20542), .C1(
        n21646), .C2(n20545), .ZN(P2_U3219) );
  OAI222_X1 U23495 ( .A1(n20544), .A2(n20510), .B1(n20509), .B2(n20542), .C1(
        n20508), .C2(n20545), .ZN(P2_U3220) );
  OAI222_X1 U23496 ( .A1(n20544), .A2(n16746), .B1(n20511), .B2(n20542), .C1(
        n20510), .C2(n20545), .ZN(P2_U3221) );
  OAI222_X1 U23497 ( .A1(n20544), .A2(n16731), .B1(n20512), .B2(n20542), .C1(
        n16746), .C2(n20545), .ZN(P2_U3222) );
  OAI222_X1 U23498 ( .A1(n20544), .A2(n16718), .B1(n20513), .B2(n20542), .C1(
        n16731), .C2(n20545), .ZN(P2_U3223) );
  OAI222_X1 U23499 ( .A1(n20549), .A2(n16706), .B1(n20514), .B2(n20542), .C1(
        n16718), .C2(n20545), .ZN(P2_U3224) );
  OAI222_X1 U23500 ( .A1(n20549), .A2(n16692), .B1(n20515), .B2(n20542), .C1(
        n16706), .C2(n20545), .ZN(P2_U3225) );
  INV_X1 U23501 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20517) );
  OAI222_X1 U23502 ( .A1(n20549), .A2(n20517), .B1(n20516), .B2(n20542), .C1(
        n16692), .C2(n20545), .ZN(P2_U3226) );
  OAI222_X1 U23503 ( .A1(n20549), .A2(n20519), .B1(n20518), .B2(n20542), .C1(
        n20517), .C2(n20545), .ZN(P2_U3227) );
  OAI222_X1 U23504 ( .A1(n20549), .A2(n20521), .B1(n20520), .B2(n20542), .C1(
        n20519), .C2(n20545), .ZN(P2_U3228) );
  OAI222_X1 U23505 ( .A1(n20549), .A2(n20523), .B1(n20522), .B2(n20542), .C1(
        n20521), .C2(n20545), .ZN(P2_U3229) );
  INV_X1 U23506 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20525) );
  OAI222_X1 U23507 ( .A1(n20544), .A2(n20525), .B1(n20524), .B2(n20542), .C1(
        n20523), .C2(n20545), .ZN(P2_U3230) );
  OAI222_X1 U23508 ( .A1(n20544), .A2(n20527), .B1(n20526), .B2(n20542), .C1(
        n20525), .C2(n20545), .ZN(P2_U3231) );
  OAI222_X1 U23509 ( .A1(n20544), .A2(n20529), .B1(n20528), .B2(n20542), .C1(
        n20527), .C2(n20545), .ZN(P2_U3232) );
  OAI222_X1 U23510 ( .A1(n20544), .A2(n20531), .B1(n20530), .B2(n20542), .C1(
        n20529), .C2(n20545), .ZN(P2_U3233) );
  OAI222_X1 U23511 ( .A1(n20544), .A2(n16619), .B1(n20532), .B2(n20542), .C1(
        n20531), .C2(n20545), .ZN(P2_U3234) );
  OAI222_X1 U23512 ( .A1(n20544), .A2(n20534), .B1(n20533), .B2(n20542), .C1(
        n16619), .C2(n20545), .ZN(P2_U3235) );
  OAI222_X1 U23513 ( .A1(n20544), .A2(n20536), .B1(n20535), .B2(n20542), .C1(
        n20534), .C2(n20545), .ZN(P2_U3236) );
  OAI222_X1 U23514 ( .A1(n20544), .A2(n20538), .B1(n20537), .B2(n20542), .C1(
        n20536), .C2(n20545), .ZN(P2_U3237) );
  OAI222_X1 U23515 ( .A1(n20545), .A2(n20538), .B1(n21636), .B2(n20542), .C1(
        n20539), .C2(n20544), .ZN(P2_U3238) );
  OAI222_X1 U23516 ( .A1(n20544), .A2(n20541), .B1(n20540), .B2(n20542), .C1(
        n20539), .C2(n20545), .ZN(P2_U3239) );
  OAI222_X1 U23517 ( .A1(n20544), .A2(n20546), .B1(n20543), .B2(n20542), .C1(
        n20541), .C2(n20545), .ZN(P2_U3240) );
  OAI222_X1 U23518 ( .A1(n20549), .A2(n20548), .B1(n20547), .B2(n20542), .C1(
        n20546), .C2(n20545), .ZN(P2_U3241) );
  INV_X1 U23519 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20550) );
  AOI22_X1 U23520 ( .A1(n20542), .A2(n20551), .B1(n20550), .B2(n20593), .ZN(
        P2_U3585) );
  INV_X1 U23521 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20552) );
  AOI22_X1 U23522 ( .A1(n20542), .A2(n20552), .B1(n21590), .B2(n20593), .ZN(
        P2_U3586) );
  INV_X1 U23523 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20553) );
  AOI22_X1 U23524 ( .A1(n20542), .A2(n20554), .B1(n20553), .B2(n20593), .ZN(
        P2_U3587) );
  INV_X1 U23525 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20555) );
  AOI22_X1 U23526 ( .A1(n20542), .A2(n20556), .B1(n20555), .B2(n20593), .ZN(
        P2_U3588) );
  OAI21_X1 U23527 ( .B1(n20560), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20558), 
        .ZN(n20557) );
  INV_X1 U23528 ( .A(n20557), .ZN(P2_U3591) );
  OAI21_X1 U23529 ( .B1(n20560), .B2(n20559), .A(n20558), .ZN(P2_U3592) );
  INV_X1 U23530 ( .A(n20587), .ZN(n20561) );
  OR2_X1 U23531 ( .A1(n20562), .A2(n20561), .ZN(n20580) );
  NAND3_X1 U23532 ( .A1(n20585), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20563), 
        .ZN(n20564) );
  NAND2_X1 U23533 ( .A1(n20564), .A2(n20583), .ZN(n20575) );
  NAND2_X1 U23534 ( .A1(n20580), .A2(n20575), .ZN(n20568) );
  NOR2_X1 U23535 ( .A1(n20565), .A2(n20607), .ZN(n20566) );
  AOI21_X1 U23536 ( .B1(n20568), .B2(n20567), .A(n20566), .ZN(n20569) );
  OAI21_X1 U23537 ( .B1(n20571), .B2(n20570), .A(n20569), .ZN(n20572) );
  INV_X1 U23538 ( .A(n20572), .ZN(n20573) );
  AOI22_X1 U23539 ( .A1(n20592), .A2(n20574), .B1(n20573), .B2(n21695), .ZN(
        P2_U3602) );
  INV_X1 U23540 ( .A(n20575), .ZN(n20577) );
  AOI22_X1 U23541 ( .A1(n20578), .A2(n20577), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20576), .ZN(n20579) );
  AND2_X1 U23542 ( .A1(n20580), .A2(n20579), .ZN(n20581) );
  AOI22_X1 U23543 ( .A1(n20592), .A2(n20582), .B1(n20581), .B2(n21695), .ZN(
        P2_U3603) );
  INV_X1 U23544 ( .A(n20583), .ZN(n21691) );
  AND2_X1 U23545 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20584) );
  NOR2_X1 U23546 ( .A1(n21691), .A2(n20584), .ZN(n20586) );
  MUX2_X1 U23547 ( .A(n20587), .B(n20586), .S(n20585), .Z(n20588) );
  AOI21_X1 U23548 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20589), .A(n20588), 
        .ZN(n20590) );
  AOI22_X1 U23549 ( .A1(n20592), .A2(n20591), .B1(n20590), .B2(n21695), .ZN(
        P2_U3604) );
  AOI22_X1 U23550 ( .A1(n20542), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20594), 
        .B2(n20593), .ZN(P2_U3608) );
  INV_X1 U23551 ( .A(n20595), .ZN(n20596) );
  AOI21_X1 U23552 ( .B1(n20598), .B2(n20597), .A(n20596), .ZN(n20600) );
  AOI211_X1 U23553 ( .C1(n20602), .C2(n20601), .A(n20600), .B(n20599), .ZN(
        n20603) );
  INV_X1 U23554 ( .A(n20603), .ZN(n20605) );
  MUX2_X1 U23555 ( .A(P2_MORE_REG_SCAN_IN), .B(n20605), .S(n20604), .Z(
        P2_U3609) );
  AOI21_X1 U23556 ( .B1(n20608), .B2(n20607), .A(n20606), .ZN(n20609) );
  OAI211_X1 U23557 ( .C1(n20612), .C2(n20611), .A(n20610), .B(n20609), .ZN(
        n20627) );
  AOI22_X1 U23558 ( .A1(n20614), .A2(n13189), .B1(n20613), .B2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n20624) );
  NOR2_X1 U23559 ( .A1(n20615), .A2(n20618), .ZN(n20616) );
  NOR2_X1 U23560 ( .A1(n20617), .A2(n20616), .ZN(n20622) );
  AND3_X1 U23561 ( .A1(n20619), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20618), 
        .ZN(n20621) );
  MUX2_X1 U23562 ( .A(n20622), .B(n20621), .S(n17491), .Z(n20623) );
  OAI21_X1 U23563 ( .B1(n20624), .B2(n20623), .A(n20627), .ZN(n20625) );
  OAI21_X1 U23564 ( .B1(n20627), .B2(n20626), .A(n20625), .ZN(P2_U3610) );
  MUX2_X1 U23565 ( .A(P2_M_IO_N_REG_SCAN_IN), .B(P2_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20542), .Z(P2_U3611) );
  NAND2_X1 U23566 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21452), .ZN(n21444) );
  AND2_X1 U23567 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21444), .ZN(n20630) );
  INV_X1 U23568 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20629) );
  INV_X2 U23569 ( .A(n21532), .ZN(n21531) );
  AOI21_X1 U23570 ( .B1(n20630), .B2(n20629), .A(n21531), .ZN(P1_U2802) );
  NOR2_X1 U23571 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20632) );
  OAI21_X1 U23572 ( .B1(n20632), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21532), .ZN(
        n20631) );
  OAI21_X1 U23573 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21532), .A(n20631), 
        .ZN(P1_U2804) );
  AOI21_X1 U23574 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21444), .A(n21531), 
        .ZN(n21510) );
  OAI21_X1 U23575 ( .B1(BS16), .B2(n20632), .A(n21510), .ZN(n21508) );
  OAI21_X1 U23576 ( .B1(n21510), .B2(n21050), .A(n21508), .ZN(P1_U2805) );
  OAI21_X1 U23577 ( .B1(n20635), .B2(n20634), .A(n20633), .ZN(P1_U2806) );
  NOR4_X1 U23578 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20645) );
  NOR4_X1 U23579 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20644) );
  AOI211_X1 U23580 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_3__SCAN_IN), .B(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20636) );
  INV_X1 U23581 ( .A(P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n21586) );
  INV_X1 U23582 ( .A(P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n21613) );
  NAND3_X1 U23583 ( .A1(n20636), .A2(n21586), .A3(n21613), .ZN(n20642) );
  NOR4_X1 U23584 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20640) );
  NOR4_X1 U23585 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20639) );
  NOR4_X1 U23586 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20638) );
  NOR4_X1 U23587 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20637) );
  NAND4_X1 U23588 ( .A1(n20640), .A2(n20639), .A3(n20638), .A4(n20637), .ZN(
        n20641) );
  NOR4_X1 U23589 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(n20642), .A4(n20641), .ZN(n20643) );
  NAND3_X1 U23590 ( .A1(n20645), .A2(n20644), .A3(n20643), .ZN(n21513) );
  NOR2_X1 U23591 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n21513), .ZN(n20647) );
  INV_X1 U23592 ( .A(n21513), .ZN(n21518) );
  NOR2_X1 U23593 ( .A1(n21518), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20646)
         );
  NOR2_X1 U23594 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(n21513), .ZN(n21511) );
  INV_X1 U23595 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21515) );
  INV_X1 U23596 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21509) );
  NAND3_X1 U23597 ( .A1(n21511), .A2(n21515), .A3(n21509), .ZN(n20648) );
  OAI21_X1 U23598 ( .B1(n20647), .B2(n20646), .A(n20648), .ZN(P1_U2807) );
  INV_X1 U23599 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21505) );
  NAND2_X1 U23600 ( .A1(n20647), .A2(n21509), .ZN(n21516) );
  OAI211_X1 U23601 ( .C1(n21518), .C2(n21505), .A(n20648), .B(n21516), .ZN(
        P1_U2808) );
  NAND2_X1 U23602 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20649) );
  NOR3_X1 U23603 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20649), .A3(n20688), .ZN(
        n20657) );
  INV_X1 U23604 ( .A(n20649), .ZN(n20650) );
  NAND2_X1 U23605 ( .A1(n20684), .A2(n20650), .ZN(n20662) );
  NAND3_X1 U23606 ( .A1(n20662), .A2(P1_REIP_REG_7__SCAN_IN), .A3(n20673), 
        .ZN(n20654) );
  NAND2_X1 U23607 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n20651) );
  NAND2_X1 U23608 ( .A1(n20651), .A2(n20771), .ZN(n20652) );
  AOI21_X1 U23609 ( .B1(n20681), .B2(P1_EBX_REG_7__SCAN_IN), .A(n20652), .ZN(
        n20653) );
  OAI211_X1 U23610 ( .C1(n20655), .C2(n20678), .A(n20654), .B(n20653), .ZN(
        n20656) );
  NOR2_X1 U23611 ( .A1(n20657), .A2(n20656), .ZN(n20660) );
  NAND2_X1 U23612 ( .A1(n20658), .A2(n20668), .ZN(n20659) );
  OAI211_X1 U23613 ( .C1(n9558), .C2(n20661), .A(n20660), .B(n20659), .ZN(
        P1_U2833) );
  NAND3_X1 U23614 ( .A1(n20662), .A2(P1_REIP_REG_6__SCAN_IN), .A3(n20673), 
        .ZN(n20664) );
  AOI22_X1 U23615 ( .A1(n20693), .A2(n10459), .B1(n20691), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n20663) );
  NAND2_X1 U23616 ( .A1(n20664), .A2(n20663), .ZN(n20665) );
  AOI211_X1 U23617 ( .C1(n20674), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20666), .B(n20665), .ZN(n20670) );
  NOR2_X1 U23618 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20688), .ZN(n20667) );
  AOI22_X1 U23619 ( .A1(n20709), .A2(n20668), .B1(n20667), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20669) );
  OAI211_X1 U23620 ( .C1(n20671), .C2(n9558), .A(n20670), .B(n20669), .ZN(
        P1_U2834) );
  INV_X1 U23621 ( .A(n20672), .ZN(n20702) );
  NAND2_X1 U23622 ( .A1(n20673), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n20683) );
  NAND2_X1 U23623 ( .A1(n20674), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n20675) );
  OAI211_X1 U23624 ( .C1(n9558), .C2(n20676), .A(n20771), .B(n20675), .ZN(
        n20680) );
  NOR2_X1 U23625 ( .A1(n20678), .A2(n20677), .ZN(n20679) );
  AOI211_X1 U23626 ( .C1(n20681), .C2(P1_EBX_REG_5__SCAN_IN), .A(n20680), .B(
        n20679), .ZN(n20682) );
  OAI21_X1 U23627 ( .B1(n20684), .B2(n20683), .A(n20682), .ZN(n20685) );
  AOI21_X1 U23628 ( .B1(n20686), .B2(n20702), .A(n20685), .ZN(n20687) );
  OAI21_X1 U23629 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20688), .A(n20687), .ZN(
        P1_U2835) );
  AOI21_X1 U23630 ( .B1(n20690), .B2(n15246), .A(n20689), .ZN(n20706) );
  INV_X1 U23631 ( .A(n20807), .ZN(n20692) );
  AOI22_X1 U23632 ( .A1(n20693), .A2(n20692), .B1(n20691), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n20705) );
  OAI22_X1 U23633 ( .A1(n9558), .A2(n20696), .B1(n20695), .B2(n20694), .ZN(
        n20697) );
  AOI21_X1 U23634 ( .B1(n20844), .B2(n20698), .A(n20697), .ZN(n20699) );
  OAI21_X1 U23635 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n20700), .A(n20699), .ZN(
        n20701) );
  AOI21_X1 U23636 ( .B1(n20703), .B2(n20702), .A(n20701), .ZN(n20704) );
  OAI211_X1 U23637 ( .C1(n20706), .C2(n14260), .A(n20705), .B(n20704), .ZN(
        P1_U2838) );
  AOI22_X1 U23638 ( .A1(n20709), .A2(n20708), .B1(n20707), .B2(n10459), .ZN(
        n20710) );
  OAI21_X1 U23639 ( .B1(n20712), .B2(n20711), .A(n20710), .ZN(P1_U2866) );
  INV_X1 U23640 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n21671) );
  INV_X1 U23641 ( .A(n20713), .ZN(n20716) );
  AOI22_X1 U23642 ( .A1(n20716), .A2(P1_EAX_REG_24__SCAN_IN), .B1(n21524), 
        .B2(P1_UWORD_REG_8__SCAN_IN), .ZN(n20714) );
  OAI21_X1 U23643 ( .B1(n21671), .B2(n20732), .A(n20714), .ZN(P1_U2912) );
  INV_X1 U23644 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n21561) );
  AOI22_X1 U23645 ( .A1(n20716), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n21524), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n20715) );
  OAI21_X1 U23646 ( .B1(n21561), .B2(n20732), .A(n20715), .ZN(P1_U2914) );
  AOI22_X1 U23647 ( .A1(n20716), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n21524), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n20717) );
  OAI21_X1 U23648 ( .B1(n21560), .B2(n20732), .A(n20717), .ZN(P1_U2919) );
  AOI22_X1 U23649 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20721), .B1(n20736), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20718) );
  OAI21_X1 U23650 ( .B1(n20719), .B2(n20735), .A(n20718), .ZN(P1_U2921) );
  AOI22_X1 U23651 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20720) );
  OAI21_X1 U23652 ( .B1(n15398), .B2(n20741), .A(n20720), .ZN(P1_U2922) );
  INV_X1 U23653 ( .A(P1_LWORD_REG_13__SCAN_IN), .ZN(n21606) );
  AOI22_X1 U23654 ( .A1(P1_EAX_REG_13__SCAN_IN), .A2(n20721), .B1(n20736), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20722) );
  OAI21_X1 U23655 ( .B1(n21606), .B2(n20735), .A(n20722), .ZN(P1_U2923) );
  AOI22_X1 U23656 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20723) );
  OAI21_X1 U23657 ( .B1(n15404), .B2(n20741), .A(n20723), .ZN(P1_U2924) );
  AOI22_X1 U23658 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20724) );
  OAI21_X1 U23659 ( .B1(n21575), .B2(n20741), .A(n20724), .ZN(P1_U2925) );
  INV_X1 U23660 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20726) );
  AOI22_X1 U23661 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20725) );
  OAI21_X1 U23662 ( .B1(n20726), .B2(n20741), .A(n20725), .ZN(P1_U2926) );
  AOI22_X1 U23663 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20727) );
  OAI21_X1 U23664 ( .B1(n15409), .B2(n20741), .A(n20727), .ZN(P1_U2927) );
  AOI22_X1 U23665 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20728) );
  OAI21_X1 U23666 ( .B1(n15410), .B2(n20741), .A(n20728), .ZN(P1_U2928) );
  AOI22_X1 U23667 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20729) );
  OAI21_X1 U23668 ( .B1(n12333), .B2(n20741), .A(n20729), .ZN(P1_U2929) );
  AOI22_X1 U23669 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20730) );
  OAI21_X1 U23670 ( .B1(n21595), .B2(n20741), .A(n20730), .ZN(P1_U2930) );
  INV_X1 U23671 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n21603) );
  OAI222_X1 U23672 ( .A1(n20735), .A2(n21603), .B1(n20741), .B2(n12303), .C1(
        n20732), .C2(n20731), .ZN(P1_U2931) );
  INV_X1 U23673 ( .A(P1_LWORD_REG_4__SCAN_IN), .ZN(n20734) );
  OAI222_X1 U23674 ( .A1(n20735), .A2(n20734), .B1(n20741), .B2(n20733), .C1(
        n21587), .C2(n20732), .ZN(P1_U2932) );
  AOI22_X1 U23675 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20737) );
  OAI21_X1 U23676 ( .B1(n12259), .B2(n20741), .A(n20737), .ZN(P1_U2933) );
  AOI22_X1 U23677 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20738) );
  OAI21_X1 U23678 ( .B1(n12207), .B2(n20741), .A(n20738), .ZN(P1_U2934) );
  AOI22_X1 U23679 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20739) );
  OAI21_X1 U23680 ( .B1(n12211), .B2(n20741), .A(n20739), .ZN(P1_U2935) );
  AOI22_X1 U23681 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21524), .B1(n20736), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20740) );
  OAI21_X1 U23682 ( .B1(n20742), .B2(n20741), .A(n20740), .ZN(P1_U2936) );
  AOI22_X1 U23683 ( .A1(n14493), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20768), .ZN(n20745) );
  INV_X1 U23684 ( .A(n20743), .ZN(n20744) );
  NAND2_X1 U23685 ( .A1(n20756), .A2(n20744), .ZN(n20758) );
  NAND2_X1 U23686 ( .A1(n20745), .A2(n20758), .ZN(P1_U2945) );
  AOI22_X1 U23687 ( .A1(n14493), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20748) );
  INV_X1 U23688 ( .A(n20746), .ZN(n20747) );
  NAND2_X1 U23689 ( .A1(n20756), .A2(n20747), .ZN(n20762) );
  NAND2_X1 U23690 ( .A1(n20748), .A2(n20762), .ZN(P1_U2947) );
  AOI22_X1 U23691 ( .A1(n14493), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20751) );
  INV_X1 U23692 ( .A(n20749), .ZN(n20750) );
  NAND2_X1 U23693 ( .A1(n20756), .A2(n20750), .ZN(n20764) );
  NAND2_X1 U23694 ( .A1(n20751), .A2(n20764), .ZN(P1_U2949) );
  AOI22_X1 U23695 ( .A1(n14493), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20753) );
  NAND2_X1 U23696 ( .A1(n20756), .A2(n20752), .ZN(n20766) );
  NAND2_X1 U23697 ( .A1(n20753), .A2(n20766), .ZN(P1_U2950) );
  AOI22_X1 U23698 ( .A1(n14493), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20768), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20757) );
  INV_X1 U23699 ( .A(n20754), .ZN(n20755) );
  NAND2_X1 U23700 ( .A1(n20756), .A2(n20755), .ZN(n20769) );
  NAND2_X1 U23701 ( .A1(n20757), .A2(n20769), .ZN(P1_U2951) );
  AOI22_X1 U23702 ( .A1(n14493), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20759) );
  NAND2_X1 U23703 ( .A1(n20759), .A2(n20758), .ZN(P1_U2960) );
  AOI22_X1 U23704 ( .A1(n14493), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20768), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20761) );
  NAND2_X1 U23705 ( .A1(n20761), .A2(n20760), .ZN(P1_U2961) );
  AOI22_X1 U23706 ( .A1(n14493), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20768), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20763) );
  NAND2_X1 U23707 ( .A1(n20763), .A2(n20762), .ZN(P1_U2962) );
  AOI22_X1 U23708 ( .A1(n14493), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20768), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20765) );
  NAND2_X1 U23709 ( .A1(n20765), .A2(n20764), .ZN(P1_U2964) );
  AOI22_X1 U23710 ( .A1(n14493), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20768), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20767) );
  NAND2_X1 U23711 ( .A1(n20767), .A2(n20766), .ZN(P1_U2965) );
  AOI22_X1 U23712 ( .A1(n14493), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20768), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20770) );
  NAND2_X1 U23713 ( .A1(n20770), .A2(n20769), .ZN(P1_U2966) );
  NOR2_X1 U23714 ( .A1(n20771), .A2(n21457), .ZN(n20788) );
  AOI21_X1 U23715 ( .B1(n20772), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20788), .ZN(n20781) );
  AOI21_X1 U23716 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14520), .A(
        n20773), .ZN(n20776) );
  XNOR2_X1 U23717 ( .A(n20774), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20775) );
  XNOR2_X1 U23718 ( .A(n20776), .B(n20775), .ZN(n20793) );
  AOI22_X1 U23719 ( .A1(n20793), .A2(n20779), .B1(n20778), .B2(n20777), .ZN(
        n20780) );
  OAI211_X1 U23720 ( .C1(n20783), .C2(n20782), .A(n20781), .B(n20780), .ZN(
        P1_U2995) );
  AOI21_X1 U23721 ( .B1(n21660), .B2(n20785), .A(n20784), .ZN(n20786) );
  INV_X1 U23722 ( .A(n20786), .ZN(n20796) );
  INV_X1 U23723 ( .A(n20787), .ZN(n20789) );
  AOI21_X1 U23724 ( .B1(n20823), .B2(n20789), .A(n20788), .ZN(n20795) );
  INV_X1 U23725 ( .A(n20790), .ZN(n20791) );
  NAND2_X1 U23726 ( .A1(n20811), .A2(n20791), .ZN(n20806) );
  NAND2_X1 U23727 ( .A1(n20792), .A2(n20806), .ZN(n20799) );
  AOI22_X1 U23728 ( .A1(n20793), .A2(n20828), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20799), .ZN(n20794) );
  OAI211_X1 U23729 ( .C1(n20803), .C2(n20796), .A(n20795), .B(n20794), .ZN(
        P1_U3027) );
  AOI21_X1 U23730 ( .B1(n20823), .B2(n20798), .A(n20797), .ZN(n20802) );
  AOI22_X1 U23731 ( .A1(n20800), .A2(n20828), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20799), .ZN(n20801) );
  OAI211_X1 U23732 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20803), .A(
        n20802), .B(n20801), .ZN(P1_U3028) );
  NAND2_X1 U23733 ( .A1(n20804), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20805) );
  OAI211_X1 U23734 ( .C1(n20808), .C2(n20807), .A(n20806), .B(n20805), .ZN(
        n20809) );
  INV_X1 U23735 ( .A(n20809), .ZN(n20818) );
  INV_X1 U23736 ( .A(n20810), .ZN(n20816) );
  NAND3_X1 U23737 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n20811), .ZN(n20812) );
  OAI211_X1 U23738 ( .C1(n20814), .C2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20813), .B(n20812), .ZN(n20815) );
  AOI22_X1 U23739 ( .A1(n20816), .A2(n20828), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20815), .ZN(n20817) );
  OAI211_X1 U23740 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n20819), .A(
        n20818), .B(n20817), .ZN(P1_U3029) );
  INV_X1 U23741 ( .A(n20820), .ZN(n20821) );
  AOI21_X1 U23742 ( .B1(n20823), .B2(n20822), .A(n20821), .ZN(n20831) );
  INV_X1 U23743 ( .A(n20824), .ZN(n20829) );
  AND2_X1 U23744 ( .A1(n20825), .A2(n20832), .ZN(n20827) );
  AOI22_X1 U23745 ( .A1(n20829), .A2(n20828), .B1(n20827), .B2(n20826), .ZN(
        n20830) );
  OAI211_X1 U23746 ( .C1(n20833), .C2(n20832), .A(n20831), .B(n20830), .ZN(
        P1_U3030) );
  NOR2_X1 U23747 ( .A1(n20835), .A2(n20834), .ZN(P1_U3032) );
  AOI22_X1 U23748 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20883), .B1(DATAI_24_), 
        .B2(n20839), .ZN(n21388) );
  NOR2_X1 U23749 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20956) );
  INV_X1 U23750 ( .A(n21240), .ZN(n20841) );
  NAND2_X1 U23751 ( .A1(n20956), .A2(n20841), .ZN(n20886) );
  OAI22_X1 U23752 ( .A1(n21413), .A2(n21388), .B1(n21241), .B2(n20886), .ZN(
        n20842) );
  INV_X1 U23753 ( .A(n20842), .ZN(n20853) );
  OAI21_X1 U23754 ( .B1(n20916), .B2(n21432), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20843) );
  NAND2_X1 U23755 ( .A1(n20843), .A2(n21210), .ZN(n20851) );
  OR2_X1 U23756 ( .A1(n21119), .A2(n20844), .ZN(n20961) );
  NOR2_X1 U23757 ( .A1(n20961), .A2(n21329), .ZN(n20848) );
  AND2_X1 U23758 ( .A1(n20849), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21239) );
  INV_X1 U23759 ( .A(n20845), .ZN(n21122) );
  NAND2_X1 U23760 ( .A1(n21122), .A2(n21179), .ZN(n20997) );
  AOI22_X1 U23761 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20997), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20886), .ZN(n20846) );
  OR2_X1 U23762 ( .A1(n20847), .A2(n21000), .ZN(n21253) );
  INV_X1 U23763 ( .A(n20848), .ZN(n20850) );
  NOR2_X1 U23764 ( .A1(n20849), .A2(n21373), .ZN(n21174) );
  INV_X1 U23765 ( .A(n21174), .ZN(n21123) );
  AOI22_X1 U23766 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20890), .B1(
        n21376), .B2(n20889), .ZN(n20852) );
  OAI211_X1 U23767 ( .C1(n21341), .C2(n20913), .A(n20853), .B(n20852), .ZN(
        P1_U3033) );
  AOI22_X1 U23768 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20883), .B1(DATAI_17_), 
        .B2(n20839), .ZN(n21394) );
  AOI22_X1 U23769 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20883), .B1(DATAI_25_), 
        .B2(n20839), .ZN(n21307) );
  OAI22_X1 U23770 ( .A1(n21413), .A2(n21307), .B1(n21254), .B2(n20886), .ZN(
        n20855) );
  INV_X1 U23771 ( .A(n20855), .ZN(n20858) );
  INV_X1 U23772 ( .A(n21000), .ZN(n20865) );
  AOI22_X1 U23773 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20890), .B1(
        n21390), .B2(n20889), .ZN(n20857) );
  OAI211_X1 U23774 ( .C1(n21394), .C2(n20913), .A(n20858), .B(n20857), .ZN(
        P1_U3034) );
  AOI22_X1 U23775 ( .A1(DATAI_18_), .A2(n20839), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20883), .ZN(n21347) );
  AOI22_X1 U23776 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20883), .B1(DATAI_26_), 
        .B2(n20839), .ZN(n21400) );
  OAI22_X1 U23777 ( .A1(n21413), .A2(n21400), .B1(n21259), .B2(n20886), .ZN(
        n20860) );
  INV_X1 U23778 ( .A(n20860), .ZN(n20863) );
  OR2_X1 U23779 ( .A1(n20861), .A2(n21000), .ZN(n21263) );
  AOI22_X1 U23780 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20890), .B1(
        n21396), .B2(n20889), .ZN(n20862) );
  OAI211_X1 U23781 ( .C1(n21347), .C2(n20913), .A(n20863), .B(n20862), .ZN(
        P1_U3035) );
  AOI22_X1 U23782 ( .A1(DATAI_19_), .A2(n20839), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20883), .ZN(n21406) );
  AOI22_X1 U23783 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20883), .B1(DATAI_27_), 
        .B2(n20839), .ZN(n21313) );
  OAI22_X1 U23784 ( .A1(n21413), .A2(n21313), .B1(n21264), .B2(n20886), .ZN(
        n20864) );
  INV_X1 U23785 ( .A(n20864), .ZN(n20868) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20890), .B1(
        n21402), .B2(n20889), .ZN(n20867) );
  OAI211_X1 U23787 ( .C1(n21406), .C2(n20913), .A(n20868), .B(n20867), .ZN(
        P1_U3036) );
  AOI22_X1 U23788 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20883), .B1(DATAI_28_), 
        .B2(n20839), .ZN(n21317) );
  OAI22_X1 U23789 ( .A1(n21413), .A2(n21317), .B1(n21269), .B2(n20886), .ZN(
        n20870) );
  INV_X1 U23790 ( .A(n20870), .ZN(n20873) );
  OR2_X1 U23791 ( .A1(n20871), .A2(n21000), .ZN(n21273) );
  AOI22_X1 U23792 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20890), .B1(
        n21408), .B2(n20889), .ZN(n20872) );
  OAI211_X1 U23793 ( .C1(n21414), .C2(n20913), .A(n20873), .B(n20872), .ZN(
        P1_U3037) );
  AOI22_X1 U23794 ( .A1(DATAI_21_), .A2(n20839), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20883), .ZN(n21355) );
  AOI22_X1 U23795 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20883), .B1(DATAI_29_), 
        .B2(n20839), .ZN(n21420) );
  OAI22_X1 U23796 ( .A1(n21413), .A2(n21420), .B1(n21274), .B2(n20886), .ZN(
        n20874) );
  INV_X1 U23797 ( .A(n20874), .ZN(n20877) );
  OR2_X1 U23798 ( .A1(n20875), .A2(n21000), .ZN(n21278) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20890), .B1(
        n21416), .B2(n20889), .ZN(n20876) );
  OAI211_X1 U23800 ( .C1(n21355), .C2(n20913), .A(n20877), .B(n20876), .ZN(
        P1_U3038) );
  AOI22_X1 U23801 ( .A1(DATAI_22_), .A2(n20839), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20883), .ZN(n21359) );
  AOI22_X1 U23802 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20883), .B1(DATAI_30_), 
        .B2(n20839), .ZN(n21426) );
  OAI22_X1 U23803 ( .A1(n21413), .A2(n21426), .B1(n21279), .B2(n20886), .ZN(
        n20879) );
  INV_X1 U23804 ( .A(n20879), .ZN(n20882) );
  OR2_X1 U23805 ( .A1(n20880), .A2(n21000), .ZN(n21283) );
  AOI22_X1 U23806 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20890), .B1(
        n21422), .B2(n20889), .ZN(n20881) );
  OAI211_X1 U23807 ( .C1(n21359), .C2(n20913), .A(n20882), .B(n20881), .ZN(
        P1_U3039) );
  AOI22_X1 U23808 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20883), .B1(DATAI_23_), 
        .B2(n20839), .ZN(n21367) );
  AOI22_X1 U23809 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20883), .B1(DATAI_31_), 
        .B2(n20839), .ZN(n21437) );
  OAI22_X1 U23810 ( .A1(n21413), .A2(n21437), .B1(n21285), .B2(n20886), .ZN(
        n20887) );
  INV_X1 U23811 ( .A(n20887), .ZN(n20892) );
  OR2_X1 U23812 ( .A1(n20888), .A2(n21000), .ZN(n21291) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20890), .B1(
        n21429), .B2(n20889), .ZN(n20891) );
  OAI211_X1 U23814 ( .C1(n21367), .C2(n20913), .A(n20892), .B(n20891), .ZN(
        P1_U3040) );
  INV_X1 U23815 ( .A(n20961), .ZN(n20894) );
  INV_X1 U23816 ( .A(n20893), .ZN(n21295) );
  NAND2_X1 U23817 ( .A1(n20956), .A2(n21372), .ZN(n20895) );
  NOR2_X1 U23818 ( .A1(n21294), .A2(n20895), .ZN(n20914) );
  AOI21_X1 U23819 ( .B1(n20894), .B2(n21295), .A(n20914), .ZN(n20896) );
  OAI22_X1 U23820 ( .A1(n20896), .A2(n21382), .B1(n20895), .B2(n21373), .ZN(
        n20915) );
  AOI22_X1 U23821 ( .A1(n20915), .A2(n21376), .B1(n21375), .B2(n20914), .ZN(
        n20900) );
  INV_X1 U23822 ( .A(n20895), .ZN(n20898) );
  OAI211_X1 U23823 ( .C1(n20958), .C2(n21149), .A(n21210), .B(n20896), .ZN(
        n20897) );
  OAI211_X1 U23824 ( .C1(n21384), .C2(n20898), .A(n21380), .B(n20897), .ZN(
        n20917) );
  INV_X1 U23825 ( .A(n21388), .ZN(n21338) );
  AOI22_X1 U23826 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20917), .B1(
        n20916), .B2(n21338), .ZN(n20899) );
  OAI211_X1 U23827 ( .C1(n21341), .C2(n20954), .A(n20900), .B(n20899), .ZN(
        P1_U3041) );
  AOI22_X1 U23828 ( .A1(n20915), .A2(n21390), .B1(n21389), .B2(n20914), .ZN(
        n20902) );
  INV_X1 U23829 ( .A(n21394), .ZN(n21304) );
  AOI22_X1 U23830 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20917), .B1(
        n20921), .B2(n21304), .ZN(n20901) );
  OAI211_X1 U23831 ( .C1(n21307), .C2(n20913), .A(n20902), .B(n20901), .ZN(
        P1_U3042) );
  AOI22_X1 U23832 ( .A1(n20915), .A2(n21396), .B1(n21395), .B2(n20914), .ZN(
        n20904) );
  INV_X1 U23833 ( .A(n21400), .ZN(n21344) );
  AOI22_X1 U23834 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20917), .B1(
        n20916), .B2(n21344), .ZN(n20903) );
  OAI211_X1 U23835 ( .C1(n21347), .C2(n20954), .A(n20904), .B(n20903), .ZN(
        P1_U3043) );
  AOI22_X1 U23836 ( .A1(n20915), .A2(n21402), .B1(n21401), .B2(n20914), .ZN(
        n20906) );
  INV_X1 U23837 ( .A(n21406), .ZN(n21310) );
  AOI22_X1 U23838 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20917), .B1(
        n20921), .B2(n21310), .ZN(n20905) );
  OAI211_X1 U23839 ( .C1(n21313), .C2(n20913), .A(n20906), .B(n20905), .ZN(
        P1_U3044) );
  AOI22_X1 U23840 ( .A1(n20915), .A2(n21408), .B1(n21407), .B2(n20914), .ZN(
        n20908) );
  INV_X1 U23841 ( .A(n21414), .ZN(n21314) );
  AOI22_X1 U23842 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20917), .B1(
        n20921), .B2(n21314), .ZN(n20907) );
  OAI211_X1 U23843 ( .C1(n21317), .C2(n20913), .A(n20908), .B(n20907), .ZN(
        P1_U3045) );
  AOI22_X1 U23844 ( .A1(n20915), .A2(n21416), .B1(n21415), .B2(n20914), .ZN(
        n20910) );
  INV_X1 U23845 ( .A(n21420), .ZN(n21352) );
  AOI22_X1 U23846 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20917), .B1(
        n20916), .B2(n21352), .ZN(n20909) );
  OAI211_X1 U23847 ( .C1(n21355), .C2(n20954), .A(n20910), .B(n20909), .ZN(
        P1_U3046) );
  AOI22_X1 U23848 ( .A1(n20915), .A2(n21422), .B1(n21421), .B2(n20914), .ZN(
        n20912) );
  INV_X1 U23849 ( .A(n21359), .ZN(n21423) );
  AOI22_X1 U23850 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20917), .B1(
        n20921), .B2(n21423), .ZN(n20911) );
  OAI211_X1 U23851 ( .C1(n21426), .C2(n20913), .A(n20912), .B(n20911), .ZN(
        P1_U3047) );
  AOI22_X1 U23852 ( .A1(n20915), .A2(n21429), .B1(n21427), .B2(n20914), .ZN(
        n20919) );
  INV_X1 U23853 ( .A(n21437), .ZN(n21362) );
  AOI22_X1 U23854 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20917), .B1(
        n20916), .B2(n21362), .ZN(n20918) );
  OAI211_X1 U23855 ( .C1(n21367), .C2(n20954), .A(n20919), .B(n20918), .ZN(
        P1_U3048) );
  NAND2_X1 U23856 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20956), .ZN(
        n20965) );
  OR2_X1 U23857 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20965), .ZN(
        n20948) );
  OAI22_X1 U23858 ( .A1(n20954), .A2(n21388), .B1(n20948), .B2(n21241), .ZN(
        n20920) );
  INV_X1 U23859 ( .A(n20920), .ZN(n20929) );
  INV_X1 U23860 ( .A(n20994), .ZN(n20922) );
  OAI21_X1 U23861 ( .B1(n20922), .B2(n20921), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20923) );
  NAND2_X1 U23862 ( .A1(n20923), .A2(n21210), .ZN(n20927) );
  NOR2_X1 U23863 ( .A1(n20961), .A2(n15284), .ZN(n20925) );
  OR2_X1 U23864 ( .A1(n21179), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21056) );
  AND2_X1 U23865 ( .A1(n21056), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21052) );
  AOI21_X1 U23866 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20948), .A(n21052), 
        .ZN(n20924) );
  INV_X1 U23867 ( .A(n20925), .ZN(n20926) );
  AOI22_X1 U23868 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20951), .B1(
        n21376), .B2(n20950), .ZN(n20928) );
  OAI211_X1 U23869 ( .C1(n21341), .C2(n20994), .A(n20929), .B(n20928), .ZN(
        P1_U3049) );
  OAI22_X1 U23870 ( .A1(n20994), .A2(n21394), .B1(n21254), .B2(n20948), .ZN(
        n20930) );
  INV_X1 U23871 ( .A(n20930), .ZN(n20932) );
  AOI22_X1 U23872 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20951), .B1(
        n21390), .B2(n20950), .ZN(n20931) );
  OAI211_X1 U23873 ( .C1(n21307), .C2(n20954), .A(n20932), .B(n20931), .ZN(
        P1_U3050) );
  OAI22_X1 U23874 ( .A1(n20994), .A2(n21347), .B1(n20948), .B2(n21259), .ZN(
        n20933) );
  INV_X1 U23875 ( .A(n20933), .ZN(n20935) );
  AOI22_X1 U23876 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20951), .B1(
        n21396), .B2(n20950), .ZN(n20934) );
  OAI211_X1 U23877 ( .C1(n21400), .C2(n20954), .A(n20935), .B(n20934), .ZN(
        P1_U3051) );
  OAI22_X1 U23878 ( .A1(n20994), .A2(n21406), .B1(n20948), .B2(n21264), .ZN(
        n20936) );
  INV_X1 U23879 ( .A(n20936), .ZN(n20938) );
  AOI22_X1 U23880 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20951), .B1(
        n21402), .B2(n20950), .ZN(n20937) );
  OAI211_X1 U23881 ( .C1(n21313), .C2(n20954), .A(n20938), .B(n20937), .ZN(
        P1_U3052) );
  OAI22_X1 U23882 ( .A1(n20994), .A2(n21414), .B1(n20948), .B2(n21269), .ZN(
        n20939) );
  INV_X1 U23883 ( .A(n20939), .ZN(n20941) );
  AOI22_X1 U23884 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20951), .B1(
        n21408), .B2(n20950), .ZN(n20940) );
  OAI211_X1 U23885 ( .C1(n21317), .C2(n20954), .A(n20941), .B(n20940), .ZN(
        P1_U3053) );
  OAI22_X1 U23886 ( .A1(n20994), .A2(n21355), .B1(n20948), .B2(n21274), .ZN(
        n20942) );
  INV_X1 U23887 ( .A(n20942), .ZN(n20944) );
  AOI22_X1 U23888 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20951), .B1(
        n21416), .B2(n20950), .ZN(n20943) );
  OAI211_X1 U23889 ( .C1(n21420), .C2(n20954), .A(n20944), .B(n20943), .ZN(
        P1_U3054) );
  OAI22_X1 U23890 ( .A1(n20994), .A2(n21359), .B1(n20948), .B2(n21279), .ZN(
        n20945) );
  INV_X1 U23891 ( .A(n20945), .ZN(n20947) );
  AOI22_X1 U23892 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20951), .B1(
        n21422), .B2(n20950), .ZN(n20946) );
  OAI211_X1 U23893 ( .C1(n21426), .C2(n20954), .A(n20947), .B(n20946), .ZN(
        P1_U3055) );
  OAI22_X1 U23894 ( .A1(n20994), .A2(n21367), .B1(n20948), .B2(n21285), .ZN(
        n20949) );
  INV_X1 U23895 ( .A(n20949), .ZN(n20953) );
  AOI22_X1 U23896 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20951), .B1(
        n21429), .B2(n20950), .ZN(n20952) );
  OAI211_X1 U23897 ( .C1(n21437), .C2(n20954), .A(n20953), .B(n20952), .ZN(
        P1_U3056) );
  NAND2_X1 U23898 ( .A1(n20956), .A2(n20955), .ZN(n20988) );
  OAI22_X1 U23899 ( .A1(n20994), .A2(n21388), .B1(n21241), .B2(n20988), .ZN(
        n20957) );
  INV_X1 U23900 ( .A(n20957), .ZN(n20969) );
  OAI21_X1 U23901 ( .B1(n20958), .B2(n21378), .A(n21210), .ZN(n20967) );
  AND2_X1 U23902 ( .A1(n20959), .A2(n12223), .ZN(n21369) );
  INV_X1 U23903 ( .A(n21369), .ZN(n20960) );
  OR2_X1 U23904 ( .A1(n20961), .A2(n20960), .ZN(n20962) );
  INV_X1 U23905 ( .A(n20966), .ZN(n20964) );
  NAND2_X1 U23906 ( .A1(n21382), .A2(n20965), .ZN(n20963) );
  OAI211_X1 U23907 ( .C1(n20967), .C2(n20964), .A(n21380), .B(n20963), .ZN(
        n20991) );
  OAI22_X1 U23908 ( .A1(n20967), .A2(n20966), .B1(n21373), .B2(n20965), .ZN(
        n20990) );
  AOI22_X1 U23909 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20991), .B1(
        n21376), .B2(n20990), .ZN(n20968) );
  OAI211_X1 U23910 ( .C1(n21341), .C2(n21021), .A(n20969), .B(n20968), .ZN(
        P1_U3057) );
  OAI22_X1 U23911 ( .A1(n21021), .A2(n21394), .B1(n21254), .B2(n20988), .ZN(
        n20970) );
  INV_X1 U23912 ( .A(n20970), .ZN(n20972) );
  AOI22_X1 U23913 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20991), .B1(
        n21390), .B2(n20990), .ZN(n20971) );
  OAI211_X1 U23914 ( .C1(n21307), .C2(n20994), .A(n20972), .B(n20971), .ZN(
        P1_U3058) );
  OAI22_X1 U23915 ( .A1(n20994), .A2(n21400), .B1(n21259), .B2(n20988), .ZN(
        n20973) );
  INV_X1 U23916 ( .A(n20973), .ZN(n20975) );
  AOI22_X1 U23917 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20991), .B1(
        n21396), .B2(n20990), .ZN(n20974) );
  OAI211_X1 U23918 ( .C1(n21347), .C2(n21021), .A(n20975), .B(n20974), .ZN(
        P1_U3059) );
  OAI22_X1 U23919 ( .A1(n20994), .A2(n21313), .B1(n21264), .B2(n20988), .ZN(
        n20976) );
  INV_X1 U23920 ( .A(n20976), .ZN(n20978) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20991), .B1(
        n21402), .B2(n20990), .ZN(n20977) );
  OAI211_X1 U23922 ( .C1(n21406), .C2(n21021), .A(n20978), .B(n20977), .ZN(
        P1_U3060) );
  OAI22_X1 U23923 ( .A1(n20994), .A2(n21317), .B1(n21269), .B2(n20988), .ZN(
        n20979) );
  INV_X1 U23924 ( .A(n20979), .ZN(n20981) );
  AOI22_X1 U23925 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20991), .B1(
        n21408), .B2(n20990), .ZN(n20980) );
  OAI211_X1 U23926 ( .C1(n21414), .C2(n21021), .A(n20981), .B(n20980), .ZN(
        P1_U3061) );
  OAI22_X1 U23927 ( .A1(n21021), .A2(n21355), .B1(n21274), .B2(n20988), .ZN(
        n20982) );
  INV_X1 U23928 ( .A(n20982), .ZN(n20984) );
  AOI22_X1 U23929 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20991), .B1(
        n21416), .B2(n20990), .ZN(n20983) );
  OAI211_X1 U23930 ( .C1(n21420), .C2(n20994), .A(n20984), .B(n20983), .ZN(
        P1_U3062) );
  OAI22_X1 U23931 ( .A1(n20994), .A2(n21426), .B1(n21279), .B2(n20988), .ZN(
        n20985) );
  INV_X1 U23932 ( .A(n20985), .ZN(n20987) );
  AOI22_X1 U23933 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20991), .B1(
        n21422), .B2(n20990), .ZN(n20986) );
  OAI211_X1 U23934 ( .C1(n21359), .C2(n21021), .A(n20987), .B(n20986), .ZN(
        P1_U3063) );
  OAI22_X1 U23935 ( .A1(n21021), .A2(n21367), .B1(n21285), .B2(n20988), .ZN(
        n20989) );
  INV_X1 U23936 ( .A(n20989), .ZN(n20993) );
  AOI22_X1 U23937 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20991), .B1(
        n21429), .B2(n20990), .ZN(n20992) );
  OAI211_X1 U23938 ( .C1(n21437), .C2(n20994), .A(n20993), .B(n20992), .ZN(
        P1_U3064) );
  INV_X1 U23939 ( .A(n21239), .ZN(n21331) );
  NOR2_X1 U23940 ( .A1(n14332), .A2(n20995), .ZN(n21089) );
  NAND3_X1 U23941 ( .A1(n21089), .A2(n21210), .A3(n15284), .ZN(n20996) );
  OAI21_X1 U23942 ( .B1(n20997), .B2(n21331), .A(n20996), .ZN(n21017) );
  AOI22_X1 U23943 ( .A1(n21017), .A2(n21376), .B1(n21375), .B2(n10477), .ZN(
        n21004) );
  AOI21_X1 U23944 ( .B1(n21021), .B2(n21047), .A(n21050), .ZN(n20998) );
  AOI21_X1 U23945 ( .B1(n21089), .B2(n15284), .A(n20998), .ZN(n20999) );
  NOR2_X1 U23946 ( .A1(n20999), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21001) );
  INV_X1 U23947 ( .A(n21021), .ZN(n21002) );
  AOI22_X1 U23948 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n21018), .B1(
        n21002), .B2(n21338), .ZN(n21003) );
  OAI211_X1 U23949 ( .C1(n21341), .C2(n21047), .A(n21004), .B(n21003), .ZN(
        P1_U3065) );
  AOI22_X1 U23950 ( .A1(n21017), .A2(n21390), .B1(n21389), .B2(n10477), .ZN(
        n21006) );
  AOI22_X1 U23951 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n21018), .B1(
        n21038), .B2(n21304), .ZN(n21005) );
  OAI211_X1 U23952 ( .C1(n21307), .C2(n21021), .A(n21006), .B(n21005), .ZN(
        P1_U3066) );
  AOI22_X1 U23953 ( .A1(n21017), .A2(n21396), .B1(n21395), .B2(n10477), .ZN(
        n21008) );
  INV_X1 U23954 ( .A(n21347), .ZN(n21397) );
  AOI22_X1 U23955 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n21018), .B1(
        n21038), .B2(n21397), .ZN(n21007) );
  OAI211_X1 U23956 ( .C1(n21400), .C2(n21021), .A(n21008), .B(n21007), .ZN(
        P1_U3067) );
  AOI22_X1 U23957 ( .A1(n21017), .A2(n21402), .B1(n21401), .B2(n10477), .ZN(
        n21010) );
  AOI22_X1 U23958 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n21018), .B1(
        n21038), .B2(n21310), .ZN(n21009) );
  OAI211_X1 U23959 ( .C1(n21313), .C2(n21021), .A(n21010), .B(n21009), .ZN(
        P1_U3068) );
  AOI22_X1 U23960 ( .A1(n21017), .A2(n21408), .B1(n21407), .B2(n10477), .ZN(
        n21012) );
  AOI22_X1 U23961 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n21018), .B1(
        n21038), .B2(n21314), .ZN(n21011) );
  OAI211_X1 U23962 ( .C1(n21317), .C2(n21021), .A(n21012), .B(n21011), .ZN(
        P1_U3069) );
  AOI22_X1 U23963 ( .A1(n21017), .A2(n21416), .B1(n21415), .B2(n10477), .ZN(
        n21014) );
  INV_X1 U23964 ( .A(n21355), .ZN(n21417) );
  AOI22_X1 U23965 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n21018), .B1(
        n21038), .B2(n21417), .ZN(n21013) );
  OAI211_X1 U23966 ( .C1(n21420), .C2(n21021), .A(n21014), .B(n21013), .ZN(
        P1_U3070) );
  AOI22_X1 U23967 ( .A1(n21017), .A2(n21422), .B1(n21421), .B2(n10477), .ZN(
        n21016) );
  AOI22_X1 U23968 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n21018), .B1(
        n21038), .B2(n21423), .ZN(n21015) );
  OAI211_X1 U23969 ( .C1(n21426), .C2(n21021), .A(n21016), .B(n21015), .ZN(
        P1_U3071) );
  AOI22_X1 U23970 ( .A1(n21017), .A2(n21429), .B1(n21427), .B2(n10477), .ZN(
        n21020) );
  INV_X1 U23971 ( .A(n21367), .ZN(n21431) );
  AOI22_X1 U23972 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n21018), .B1(
        n21038), .B2(n21431), .ZN(n21019) );
  OAI211_X1 U23973 ( .C1(n21437), .C2(n21021), .A(n21020), .B(n21019), .ZN(
        P1_U3072) );
  NOR2_X1 U23974 ( .A1(n21048), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21025) );
  INV_X1 U23975 ( .A(n21025), .ZN(n21022) );
  NOR2_X1 U23976 ( .A1(n21294), .A2(n21022), .ZN(n21041) );
  AOI21_X1 U23977 ( .B1(n21089), .B2(n21295), .A(n21041), .ZN(n21023) );
  OAI22_X1 U23978 ( .A1(n21023), .A2(n21382), .B1(n21022), .B2(n21373), .ZN(
        n21042) );
  AOI22_X1 U23979 ( .A1(n21042), .A2(n21376), .B1(n21375), .B2(n21041), .ZN(
        n21027) );
  OAI211_X1 U23980 ( .C1(n21087), .C2(n21149), .A(n21210), .B(n21023), .ZN(
        n21024) );
  OAI211_X1 U23981 ( .C1(n21384), .C2(n21025), .A(n21380), .B(n21024), .ZN(
        n21044) );
  INV_X1 U23982 ( .A(n21085), .ZN(n21043) );
  INV_X1 U23983 ( .A(n21341), .ZN(n21385) );
  AOI22_X1 U23984 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21044), .B1(
        n21043), .B2(n21385), .ZN(n21026) );
  OAI211_X1 U23985 ( .C1(n21388), .C2(n21047), .A(n21027), .B(n21026), .ZN(
        P1_U3073) );
  AOI22_X1 U23986 ( .A1(n21042), .A2(n21390), .B1(n21389), .B2(n21041), .ZN(
        n21029) );
  INV_X1 U23987 ( .A(n21307), .ZN(n21391) );
  AOI22_X1 U23988 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21044), .B1(
        n21038), .B2(n21391), .ZN(n21028) );
  OAI211_X1 U23989 ( .C1(n21394), .C2(n21085), .A(n21029), .B(n21028), .ZN(
        P1_U3074) );
  AOI22_X1 U23990 ( .A1(n21042), .A2(n21396), .B1(n21395), .B2(n21041), .ZN(
        n21031) );
  AOI22_X1 U23991 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21044), .B1(
        n21038), .B2(n21344), .ZN(n21030) );
  OAI211_X1 U23992 ( .C1(n21347), .C2(n21085), .A(n21031), .B(n21030), .ZN(
        P1_U3075) );
  AOI22_X1 U23993 ( .A1(n21042), .A2(n21402), .B1(n21401), .B2(n21041), .ZN(
        n21033) );
  AOI22_X1 U23994 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21044), .B1(
        n21043), .B2(n21310), .ZN(n21032) );
  OAI211_X1 U23995 ( .C1(n21313), .C2(n21047), .A(n21033), .B(n21032), .ZN(
        P1_U3076) );
  AOI22_X1 U23996 ( .A1(n21042), .A2(n21408), .B1(n21407), .B2(n21041), .ZN(
        n21035) );
  INV_X1 U23997 ( .A(n21317), .ZN(n21409) );
  AOI22_X1 U23998 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21044), .B1(
        n21038), .B2(n21409), .ZN(n21034) );
  OAI211_X1 U23999 ( .C1(n21414), .C2(n21085), .A(n21035), .B(n21034), .ZN(
        P1_U3077) );
  AOI22_X1 U24000 ( .A1(n21042), .A2(n21416), .B1(n21415), .B2(n21041), .ZN(
        n21037) );
  AOI22_X1 U24001 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21044), .B1(
        n21038), .B2(n21352), .ZN(n21036) );
  OAI211_X1 U24002 ( .C1(n21355), .C2(n21085), .A(n21037), .B(n21036), .ZN(
        P1_U3078) );
  AOI22_X1 U24003 ( .A1(n21042), .A2(n21422), .B1(n21421), .B2(n21041), .ZN(
        n21040) );
  INV_X1 U24004 ( .A(n21426), .ZN(n21356) );
  AOI22_X1 U24005 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21044), .B1(
        n21038), .B2(n21356), .ZN(n21039) );
  OAI211_X1 U24006 ( .C1(n21359), .C2(n21085), .A(n21040), .B(n21039), .ZN(
        P1_U3079) );
  AOI22_X1 U24007 ( .A1(n21042), .A2(n21429), .B1(n21427), .B2(n21041), .ZN(
        n21046) );
  AOI22_X1 U24008 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21044), .B1(
        n21043), .B2(n21431), .ZN(n21045) );
  OAI211_X1 U24009 ( .C1(n21437), .C2(n21047), .A(n21046), .B(n21045), .ZN(
        P1_U3080) );
  NOR2_X1 U24010 ( .A1(n21372), .A2(n21048), .ZN(n21095) );
  INV_X1 U24011 ( .A(n21095), .ZN(n21090) );
  NOR2_X1 U24012 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21090), .ZN(
        n21054) );
  INV_X1 U24013 ( .A(n21054), .ZN(n21079) );
  OAI22_X1 U24014 ( .A1(n21085), .A2(n21388), .B1(n21241), .B2(n21079), .ZN(
        n21049) );
  INV_X1 U24015 ( .A(n21049), .ZN(n21060) );
  NAND3_X1 U24016 ( .A1(n21117), .A2(n21085), .A3(n21384), .ZN(n21051) );
  NAND2_X1 U24017 ( .A1(n21210), .A2(n21050), .ZN(n21235) );
  NAND2_X1 U24018 ( .A1(n21051), .A2(n21235), .ZN(n21055) );
  NAND2_X1 U24019 ( .A1(n21089), .A2(n21329), .ZN(n21057) );
  AOI21_X1 U24020 ( .B1(n21055), .B2(n21057), .A(n21052), .ZN(n21053) );
  INV_X1 U24021 ( .A(n21055), .ZN(n21058) );
  AOI22_X1 U24022 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n21082), .B1(
        n21376), .B2(n21081), .ZN(n21059) );
  OAI211_X1 U24023 ( .C1(n21341), .C2(n21117), .A(n21060), .B(n21059), .ZN(
        P1_U3081) );
  OAI22_X1 U24024 ( .A1(n21085), .A2(n21307), .B1(n21254), .B2(n21079), .ZN(
        n21061) );
  INV_X1 U24025 ( .A(n21061), .ZN(n21063) );
  AOI22_X1 U24026 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n21082), .B1(
        n21390), .B2(n21081), .ZN(n21062) );
  OAI211_X1 U24027 ( .C1(n21394), .C2(n21117), .A(n21063), .B(n21062), .ZN(
        P1_U3082) );
  OAI22_X1 U24028 ( .A1(n21085), .A2(n21400), .B1(n21259), .B2(n21079), .ZN(
        n21064) );
  INV_X1 U24029 ( .A(n21064), .ZN(n21066) );
  AOI22_X1 U24030 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n21082), .B1(
        n21396), .B2(n21081), .ZN(n21065) );
  OAI211_X1 U24031 ( .C1(n21347), .C2(n21117), .A(n21066), .B(n21065), .ZN(
        P1_U3083) );
  OAI22_X1 U24032 ( .A1(n21085), .A2(n21313), .B1(n21264), .B2(n21079), .ZN(
        n21067) );
  INV_X1 U24033 ( .A(n21067), .ZN(n21069) );
  AOI22_X1 U24034 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n21082), .B1(
        n21402), .B2(n21081), .ZN(n21068) );
  OAI211_X1 U24035 ( .C1(n21406), .C2(n21117), .A(n21069), .B(n21068), .ZN(
        P1_U3084) );
  OAI22_X1 U24036 ( .A1(n21117), .A2(n21414), .B1(n21269), .B2(n21079), .ZN(
        n21070) );
  INV_X1 U24037 ( .A(n21070), .ZN(n21072) );
  AOI22_X1 U24038 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n21082), .B1(
        n21408), .B2(n21081), .ZN(n21071) );
  OAI211_X1 U24039 ( .C1(n21317), .C2(n21085), .A(n21072), .B(n21071), .ZN(
        P1_U3085) );
  OAI22_X1 U24040 ( .A1(n21085), .A2(n21420), .B1(n21274), .B2(n21079), .ZN(
        n21073) );
  INV_X1 U24041 ( .A(n21073), .ZN(n21075) );
  AOI22_X1 U24042 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n21082), .B1(
        n21416), .B2(n21081), .ZN(n21074) );
  OAI211_X1 U24043 ( .C1(n21355), .C2(n21117), .A(n21075), .B(n21074), .ZN(
        P1_U3086) );
  OAI22_X1 U24044 ( .A1(n21085), .A2(n21426), .B1(n21279), .B2(n21079), .ZN(
        n21076) );
  INV_X1 U24045 ( .A(n21076), .ZN(n21078) );
  AOI22_X1 U24046 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n21082), .B1(
        n21422), .B2(n21081), .ZN(n21077) );
  OAI211_X1 U24047 ( .C1(n21359), .C2(n21117), .A(n21078), .B(n21077), .ZN(
        P1_U3087) );
  OAI22_X1 U24048 ( .A1(n21117), .A2(n21367), .B1(n21285), .B2(n21079), .ZN(
        n21080) );
  INV_X1 U24049 ( .A(n21080), .ZN(n21084) );
  AOI22_X1 U24050 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n21082), .B1(
        n21429), .B2(n21081), .ZN(n21083) );
  OAI211_X1 U24051 ( .C1(n21437), .C2(n21085), .A(n21084), .B(n21083), .ZN(
        P1_U3088) );
  INV_X1 U24052 ( .A(n21088), .ZN(n21112) );
  AOI21_X1 U24053 ( .B1(n21089), .B2(n21369), .A(n21112), .ZN(n21092) );
  OAI22_X1 U24054 ( .A1(n21092), .A2(n21382), .B1(n21090), .B2(n21373), .ZN(
        n21113) );
  AOI22_X1 U24055 ( .A1(n21113), .A2(n21376), .B1(n21112), .B2(n21375), .ZN(
        n21097) );
  INV_X1 U24056 ( .A(n21091), .ZN(n21093) );
  NAND3_X1 U24057 ( .A1(n21093), .A2(n21384), .A3(n21092), .ZN(n21094) );
  OAI211_X1 U24058 ( .C1(n21384), .C2(n21095), .A(n21380), .B(n21094), .ZN(
        n21114) );
  INV_X1 U24059 ( .A(n21117), .ZN(n21104) );
  AOI22_X1 U24060 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n21114), .B1(
        n21104), .B2(n21338), .ZN(n21096) );
  OAI211_X1 U24061 ( .C1(n21341), .C2(n21107), .A(n21097), .B(n21096), .ZN(
        P1_U3089) );
  AOI22_X1 U24062 ( .A1(n21113), .A2(n21390), .B1(n21112), .B2(n21389), .ZN(
        n21099) );
  AOI22_X1 U24063 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n21114), .B1(
        n21143), .B2(n21304), .ZN(n21098) );
  OAI211_X1 U24064 ( .C1(n21307), .C2(n21117), .A(n21099), .B(n21098), .ZN(
        P1_U3090) );
  AOI22_X1 U24065 ( .A1(n21113), .A2(n21396), .B1(n21112), .B2(n21395), .ZN(
        n21101) );
  AOI22_X1 U24066 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n21114), .B1(
        n21143), .B2(n21397), .ZN(n21100) );
  OAI211_X1 U24067 ( .C1(n21400), .C2(n21117), .A(n21101), .B(n21100), .ZN(
        P1_U3091) );
  AOI22_X1 U24068 ( .A1(n21113), .A2(n21402), .B1(n21112), .B2(n21401), .ZN(
        n21103) );
  INV_X1 U24069 ( .A(n21313), .ZN(n21403) );
  AOI22_X1 U24070 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n21114), .B1(
        n21104), .B2(n21403), .ZN(n21102) );
  OAI211_X1 U24071 ( .C1(n21406), .C2(n21107), .A(n21103), .B(n21102), .ZN(
        P1_U3092) );
  AOI22_X1 U24072 ( .A1(n21113), .A2(n21408), .B1(n21112), .B2(n21407), .ZN(
        n21106) );
  AOI22_X1 U24073 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n21114), .B1(
        n21104), .B2(n21409), .ZN(n21105) );
  OAI211_X1 U24074 ( .C1(n21414), .C2(n21107), .A(n21106), .B(n21105), .ZN(
        P1_U3093) );
  AOI22_X1 U24075 ( .A1(n21113), .A2(n21416), .B1(n21112), .B2(n21415), .ZN(
        n21109) );
  AOI22_X1 U24076 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n21114), .B1(
        n21143), .B2(n21417), .ZN(n21108) );
  OAI211_X1 U24077 ( .C1(n21420), .C2(n21117), .A(n21109), .B(n21108), .ZN(
        P1_U3094) );
  AOI22_X1 U24078 ( .A1(n21113), .A2(n21422), .B1(n21112), .B2(n21421), .ZN(
        n21111) );
  AOI22_X1 U24079 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n21114), .B1(
        n21143), .B2(n21423), .ZN(n21110) );
  OAI211_X1 U24080 ( .C1(n21426), .C2(n21117), .A(n21111), .B(n21110), .ZN(
        P1_U3095) );
  AOI22_X1 U24081 ( .A1(n21113), .A2(n21429), .B1(n21112), .B2(n21427), .ZN(
        n21116) );
  AOI22_X1 U24082 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n21114), .B1(
        n21143), .B2(n21431), .ZN(n21115) );
  OAI211_X1 U24083 ( .C1(n21437), .C2(n21117), .A(n21116), .B(n21115), .ZN(
        P1_U3096) );
  AND2_X1 U24084 ( .A1(n21119), .A2(n14332), .ZN(n21207) );
  NAND2_X1 U24085 ( .A1(n21120), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21205) );
  AOI21_X1 U24086 ( .B1(n21207), .B2(n15284), .A(n10472), .ZN(n21125) );
  NOR2_X1 U24087 ( .A1(n21122), .A2(n21121), .ZN(n21238) );
  INV_X1 U24088 ( .A(n21238), .ZN(n21244) );
  OAI22_X1 U24089 ( .A1(n21125), .A2(n21382), .B1(n21123), .B2(n21244), .ZN(
        n21142) );
  AOI22_X1 U24090 ( .A1(n21142), .A2(n21376), .B1(n10472), .B2(n21375), .ZN(
        n21129) );
  INV_X1 U24091 ( .A(n21171), .ZN(n21124) );
  OAI21_X1 U24092 ( .B1(n21124), .B2(n21143), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21126) );
  NAND2_X1 U24093 ( .A1(n21126), .A2(n21125), .ZN(n21127) );
  AOI22_X1 U24094 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n21144), .B1(
        n21143), .B2(n21338), .ZN(n21128) );
  OAI211_X1 U24095 ( .C1(n21341), .C2(n21171), .A(n21129), .B(n21128), .ZN(
        P1_U3097) );
  AOI22_X1 U24096 ( .A1(n21142), .A2(n21390), .B1(n10472), .B2(n21389), .ZN(
        n21131) );
  AOI22_X1 U24097 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21144), .B1(
        n21143), .B2(n21391), .ZN(n21130) );
  OAI211_X1 U24098 ( .C1(n21394), .C2(n21171), .A(n21131), .B(n21130), .ZN(
        P1_U3098) );
  AOI22_X1 U24099 ( .A1(n21142), .A2(n21396), .B1(n10472), .B2(n21395), .ZN(
        n21133) );
  AOI22_X1 U24100 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n21144), .B1(
        n21143), .B2(n21344), .ZN(n21132) );
  OAI211_X1 U24101 ( .C1(n21347), .C2(n21171), .A(n21133), .B(n21132), .ZN(
        P1_U3099) );
  AOI22_X1 U24102 ( .A1(n21142), .A2(n21402), .B1(n10472), .B2(n21401), .ZN(
        n21135) );
  AOI22_X1 U24103 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n21144), .B1(
        n21143), .B2(n21403), .ZN(n21134) );
  OAI211_X1 U24104 ( .C1(n21406), .C2(n21171), .A(n21135), .B(n21134), .ZN(
        P1_U3100) );
  AOI22_X1 U24105 ( .A1(n21142), .A2(n21408), .B1(n10472), .B2(n21407), .ZN(
        n21137) );
  AOI22_X1 U24106 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n21144), .B1(
        n21143), .B2(n21409), .ZN(n21136) );
  OAI211_X1 U24107 ( .C1(n21414), .C2(n21171), .A(n21137), .B(n21136), .ZN(
        P1_U3101) );
  AOI22_X1 U24108 ( .A1(n21142), .A2(n21416), .B1(n10472), .B2(n21415), .ZN(
        n21139) );
  AOI22_X1 U24109 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n21144), .B1(
        n21143), .B2(n21352), .ZN(n21138) );
  OAI211_X1 U24110 ( .C1(n21355), .C2(n21171), .A(n21139), .B(n21138), .ZN(
        P1_U3102) );
  AOI22_X1 U24111 ( .A1(n21142), .A2(n21422), .B1(n10472), .B2(n21421), .ZN(
        n21141) );
  AOI22_X1 U24112 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n21144), .B1(
        n21143), .B2(n21356), .ZN(n21140) );
  OAI211_X1 U24113 ( .C1(n21359), .C2(n21171), .A(n21141), .B(n21140), .ZN(
        P1_U3103) );
  AOI22_X1 U24114 ( .A1(n21142), .A2(n21429), .B1(n10472), .B2(n21427), .ZN(
        n21146) );
  AOI22_X1 U24115 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n21144), .B1(
        n21143), .B2(n21362), .ZN(n21145) );
  OAI211_X1 U24116 ( .C1(n21367), .C2(n21171), .A(n21146), .B(n21145), .ZN(
        P1_U3104) );
  NOR2_X1 U24117 ( .A1(n21205), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21151) );
  INV_X1 U24118 ( .A(n21151), .ZN(n21147) );
  NOR2_X1 U24119 ( .A1(n21294), .A2(n21147), .ZN(n21166) );
  AOI21_X1 U24120 ( .B1(n21207), .B2(n21295), .A(n21166), .ZN(n21148) );
  OAI22_X1 U24121 ( .A1(n21148), .A2(n21382), .B1(n21147), .B2(n21373), .ZN(
        n21167) );
  AOI22_X1 U24122 ( .A1(n21167), .A2(n21376), .B1(n21375), .B2(n21166), .ZN(
        n21153) );
  OAI211_X1 U24123 ( .C1(n21211), .C2(n21149), .A(n21210), .B(n21148), .ZN(
        n21150) );
  OAI211_X1 U24124 ( .C1(n21384), .C2(n21151), .A(n21380), .B(n21150), .ZN(
        n21168) );
  AOI22_X1 U24125 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21168), .B1(
        n21198), .B2(n21385), .ZN(n21152) );
  OAI211_X1 U24126 ( .C1(n21388), .C2(n21171), .A(n21153), .B(n21152), .ZN(
        P1_U3105) );
  AOI22_X1 U24127 ( .A1(n21167), .A2(n21390), .B1(n21389), .B2(n21166), .ZN(
        n21155) );
  AOI22_X1 U24128 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21168), .B1(
        n21198), .B2(n21304), .ZN(n21154) );
  OAI211_X1 U24129 ( .C1(n21307), .C2(n21171), .A(n21155), .B(n21154), .ZN(
        P1_U3106) );
  AOI22_X1 U24130 ( .A1(n21167), .A2(n21396), .B1(n21395), .B2(n21166), .ZN(
        n21157) );
  AOI22_X1 U24131 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21168), .B1(
        n21198), .B2(n21397), .ZN(n21156) );
  OAI211_X1 U24132 ( .C1(n21400), .C2(n21171), .A(n21157), .B(n21156), .ZN(
        P1_U3107) );
  AOI22_X1 U24133 ( .A1(n21167), .A2(n21402), .B1(n21401), .B2(n21166), .ZN(
        n21159) );
  AOI22_X1 U24134 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21168), .B1(
        n21198), .B2(n21310), .ZN(n21158) );
  OAI211_X1 U24135 ( .C1(n21313), .C2(n21171), .A(n21159), .B(n21158), .ZN(
        P1_U3108) );
  AOI22_X1 U24136 ( .A1(n21167), .A2(n21408), .B1(n21407), .B2(n21166), .ZN(
        n21161) );
  AOI22_X1 U24137 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21168), .B1(
        n21198), .B2(n21314), .ZN(n21160) );
  OAI211_X1 U24138 ( .C1(n21317), .C2(n21171), .A(n21161), .B(n21160), .ZN(
        P1_U3109) );
  AOI22_X1 U24139 ( .A1(n21167), .A2(n21416), .B1(n21415), .B2(n21166), .ZN(
        n21163) );
  AOI22_X1 U24140 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21168), .B1(
        n21198), .B2(n21417), .ZN(n21162) );
  OAI211_X1 U24141 ( .C1(n21420), .C2(n21171), .A(n21163), .B(n21162), .ZN(
        P1_U3110) );
  AOI22_X1 U24142 ( .A1(n21167), .A2(n21422), .B1(n21421), .B2(n21166), .ZN(
        n21165) );
  AOI22_X1 U24143 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21168), .B1(
        n21198), .B2(n21423), .ZN(n21164) );
  OAI211_X1 U24144 ( .C1(n21426), .C2(n21171), .A(n21165), .B(n21164), .ZN(
        P1_U3111) );
  AOI22_X1 U24145 ( .A1(n21167), .A2(n21429), .B1(n21427), .B2(n21166), .ZN(
        n21170) );
  AOI22_X1 U24146 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21168), .B1(
        n21198), .B2(n21431), .ZN(n21169) );
  OAI211_X1 U24147 ( .C1(n21437), .C2(n21171), .A(n21170), .B(n21169), .ZN(
        P1_U3112) );
  INV_X1 U24148 ( .A(n21198), .ZN(n21172) );
  NAND2_X1 U24149 ( .A1(n21172), .A2(n21210), .ZN(n21173) );
  NOR2_X1 U24150 ( .A1(n21179), .A2(n21180), .ZN(n21330) );
  NOR2_X1 U24151 ( .A1(n21372), .A2(n21205), .ZN(n21213) );
  INV_X1 U24152 ( .A(n21213), .ZN(n21208) );
  NOR2_X1 U24153 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21208), .ZN(
        n21197) );
  AOI22_X1 U24154 ( .A1(n21230), .A2(n21385), .B1(n21375), .B2(n21197), .ZN(
        n21184) );
  INV_X1 U24155 ( .A(n21175), .ZN(n21177) );
  INV_X1 U24156 ( .A(n21197), .ZN(n21176) );
  AOI22_X1 U24157 ( .A1(n21178), .A2(n21177), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21176), .ZN(n21181) );
  OAI21_X1 U24158 ( .B1(n21180), .B2(n21179), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n21335) );
  NAND3_X1 U24159 ( .A1(n21182), .A2(n21181), .A3(n21335), .ZN(n21199) );
  AOI22_X1 U24160 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21199), .B1(
        n21198), .B2(n21338), .ZN(n21183) );
  OAI211_X1 U24161 ( .C1(n21202), .C2(n21253), .A(n21184), .B(n21183), .ZN(
        P1_U3113) );
  INV_X1 U24162 ( .A(n21390), .ZN(n21258) );
  AOI22_X1 U24163 ( .A1(n21230), .A2(n21304), .B1(n21389), .B2(n21197), .ZN(
        n21186) );
  AOI22_X1 U24164 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21199), .B1(
        n21198), .B2(n21391), .ZN(n21185) );
  OAI211_X1 U24165 ( .C1(n21202), .C2(n21258), .A(n21186), .B(n21185), .ZN(
        P1_U3114) );
  AOI22_X1 U24166 ( .A1(n21198), .A2(n21344), .B1(n21395), .B2(n21197), .ZN(
        n21188) );
  AOI22_X1 U24167 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21199), .B1(
        n21230), .B2(n21397), .ZN(n21187) );
  OAI211_X1 U24168 ( .C1(n21202), .C2(n21263), .A(n21188), .B(n21187), .ZN(
        P1_U3115) );
  INV_X1 U24169 ( .A(n21402), .ZN(n21268) );
  AOI22_X1 U24170 ( .A1(n21198), .A2(n21403), .B1(n21401), .B2(n21197), .ZN(
        n21190) );
  AOI22_X1 U24171 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21199), .B1(
        n21230), .B2(n21310), .ZN(n21189) );
  OAI211_X1 U24172 ( .C1(n21202), .C2(n21268), .A(n21190), .B(n21189), .ZN(
        P1_U3116) );
  AOI22_X1 U24173 ( .A1(n21230), .A2(n21314), .B1(n21407), .B2(n21197), .ZN(
        n21192) );
  AOI22_X1 U24174 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21199), .B1(
        n21198), .B2(n21409), .ZN(n21191) );
  OAI211_X1 U24175 ( .C1(n21202), .C2(n21273), .A(n21192), .B(n21191), .ZN(
        P1_U3117) );
  AOI22_X1 U24176 ( .A1(n21230), .A2(n21417), .B1(n21415), .B2(n21197), .ZN(
        n21194) );
  AOI22_X1 U24177 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21199), .B1(
        n21198), .B2(n21352), .ZN(n21193) );
  OAI211_X1 U24178 ( .C1(n21202), .C2(n21278), .A(n21194), .B(n21193), .ZN(
        P1_U3118) );
  AOI22_X1 U24179 ( .A1(n21230), .A2(n21423), .B1(n21421), .B2(n21197), .ZN(
        n21196) );
  AOI22_X1 U24180 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21199), .B1(
        n21198), .B2(n21356), .ZN(n21195) );
  OAI211_X1 U24181 ( .C1(n21202), .C2(n21283), .A(n21196), .B(n21195), .ZN(
        P1_U3119) );
  AOI22_X1 U24182 ( .A1(n21198), .A2(n21362), .B1(n21427), .B2(n21197), .ZN(
        n21201) );
  AOI22_X1 U24183 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21199), .B1(
        n21230), .B2(n21431), .ZN(n21200) );
  OAI211_X1 U24184 ( .C1(n21202), .C2(n21291), .A(n21201), .B(n21200), .ZN(
        P1_U3120) );
  NOR2_X1 U24185 ( .A1(n21206), .A2(n21205), .ZN(n21228) );
  AOI21_X1 U24186 ( .B1(n21207), .B2(n21369), .A(n21228), .ZN(n21209) );
  OAI22_X1 U24187 ( .A1(n21209), .A2(n21382), .B1(n21208), .B2(n21373), .ZN(
        n21229) );
  AOI22_X1 U24188 ( .A1(n21229), .A2(n21376), .B1(n21375), .B2(n21228), .ZN(
        n21215) );
  OAI211_X1 U24189 ( .C1(n21211), .C2(n21378), .A(n21210), .B(n21209), .ZN(
        n21212) );
  OAI211_X1 U24190 ( .C1(n21384), .C2(n21213), .A(n21380), .B(n21212), .ZN(
        n21231) );
  AOI22_X1 U24191 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21231), .B1(
        n21230), .B2(n21338), .ZN(n21214) );
  OAI211_X1 U24192 ( .C1(n21341), .C2(n21250), .A(n21215), .B(n21214), .ZN(
        P1_U3121) );
  AOI22_X1 U24193 ( .A1(n21229), .A2(n21390), .B1(n21389), .B2(n21228), .ZN(
        n21217) );
  AOI22_X1 U24194 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21231), .B1(
        n21230), .B2(n21391), .ZN(n21216) );
  OAI211_X1 U24195 ( .C1(n21394), .C2(n21250), .A(n21217), .B(n21216), .ZN(
        P1_U3122) );
  AOI22_X1 U24196 ( .A1(n21229), .A2(n21396), .B1(n21395), .B2(n21228), .ZN(
        n21219) );
  AOI22_X1 U24197 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21231), .B1(
        n21230), .B2(n21344), .ZN(n21218) );
  OAI211_X1 U24198 ( .C1(n21347), .C2(n21250), .A(n21219), .B(n21218), .ZN(
        P1_U3123) );
  AOI22_X1 U24199 ( .A1(n21229), .A2(n21402), .B1(n21401), .B2(n21228), .ZN(
        n21221) );
  AOI22_X1 U24200 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21231), .B1(
        n21230), .B2(n21403), .ZN(n21220) );
  OAI211_X1 U24201 ( .C1(n21406), .C2(n21250), .A(n21221), .B(n21220), .ZN(
        P1_U3124) );
  AOI22_X1 U24202 ( .A1(n21229), .A2(n21408), .B1(n21407), .B2(n21228), .ZN(
        n21223) );
  AOI22_X1 U24203 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21231), .B1(
        n21230), .B2(n21409), .ZN(n21222) );
  OAI211_X1 U24204 ( .C1(n21414), .C2(n21250), .A(n21223), .B(n21222), .ZN(
        P1_U3125) );
  AOI22_X1 U24205 ( .A1(n21229), .A2(n21416), .B1(n21415), .B2(n21228), .ZN(
        n21225) );
  AOI22_X1 U24206 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21231), .B1(
        n21230), .B2(n21352), .ZN(n21224) );
  OAI211_X1 U24207 ( .C1(n21355), .C2(n21250), .A(n21225), .B(n21224), .ZN(
        P1_U3126) );
  AOI22_X1 U24208 ( .A1(n21229), .A2(n21422), .B1(n21421), .B2(n21228), .ZN(
        n21227) );
  AOI22_X1 U24209 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21231), .B1(
        n21230), .B2(n21356), .ZN(n21226) );
  OAI211_X1 U24210 ( .C1(n21359), .C2(n21250), .A(n21227), .B(n21226), .ZN(
        P1_U3127) );
  AOI22_X1 U24211 ( .A1(n21229), .A2(n21429), .B1(n21427), .B2(n21228), .ZN(
        n21233) );
  AOI22_X1 U24212 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21231), .B1(
        n21230), .B2(n21362), .ZN(n21232) );
  OAI211_X1 U24213 ( .C1(n21367), .C2(n21250), .A(n21233), .B(n21232), .ZN(
        P1_U3128) );
  NAND3_X1 U24214 ( .A1(n21250), .A2(n21384), .A3(n21327), .ZN(n21236) );
  NAND2_X1 U24215 ( .A1(n21236), .A2(n21235), .ZN(n21246) );
  OR2_X1 U24216 ( .A1(n14332), .A2(n21237), .ZN(n21293) );
  NOR2_X1 U24217 ( .A1(n21293), .A2(n21329), .ZN(n21243) );
  OR2_X1 U24218 ( .A1(n21240), .A2(n21371), .ZN(n21284) );
  OAI22_X1 U24219 ( .A1(n21327), .A2(n21341), .B1(n21241), .B2(n21284), .ZN(
        n21242) );
  INV_X1 U24220 ( .A(n21242), .ZN(n21252) );
  INV_X1 U24221 ( .A(n21284), .ZN(n21249) );
  INV_X1 U24222 ( .A(n21243), .ZN(n21245) );
  AOI22_X1 U24223 ( .A1(n21246), .A2(n21245), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21244), .ZN(n21247) );
  AOI22_X1 U24224 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21288), .B1(
        n21287), .B2(n21338), .ZN(n21251) );
  OAI211_X1 U24225 ( .C1(n21292), .C2(n21253), .A(n21252), .B(n21251), .ZN(
        P1_U3129) );
  OAI22_X1 U24226 ( .A1(n21327), .A2(n21394), .B1(n21254), .B2(n21284), .ZN(
        n21255) );
  INV_X1 U24227 ( .A(n21255), .ZN(n21257) );
  AOI22_X1 U24228 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21288), .B1(
        n21287), .B2(n21391), .ZN(n21256) );
  OAI211_X1 U24229 ( .C1(n21292), .C2(n21258), .A(n21257), .B(n21256), .ZN(
        P1_U3130) );
  OAI22_X1 U24230 ( .A1(n21327), .A2(n21347), .B1(n21259), .B2(n21284), .ZN(
        n21260) );
  INV_X1 U24231 ( .A(n21260), .ZN(n21262) );
  AOI22_X1 U24232 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21288), .B1(
        n21287), .B2(n21344), .ZN(n21261) );
  OAI211_X1 U24233 ( .C1(n21292), .C2(n21263), .A(n21262), .B(n21261), .ZN(
        P1_U3131) );
  OAI22_X1 U24234 ( .A1(n21327), .A2(n21406), .B1(n21264), .B2(n21284), .ZN(
        n21265) );
  INV_X1 U24235 ( .A(n21265), .ZN(n21267) );
  AOI22_X1 U24236 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21288), .B1(
        n21287), .B2(n21403), .ZN(n21266) );
  OAI211_X1 U24237 ( .C1(n21292), .C2(n21268), .A(n21267), .B(n21266), .ZN(
        P1_U3132) );
  OAI22_X1 U24238 ( .A1(n21327), .A2(n21414), .B1(n21269), .B2(n21284), .ZN(
        n21270) );
  INV_X1 U24239 ( .A(n21270), .ZN(n21272) );
  AOI22_X1 U24240 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21288), .B1(
        n21287), .B2(n21409), .ZN(n21271) );
  OAI211_X1 U24241 ( .C1(n21292), .C2(n21273), .A(n21272), .B(n21271), .ZN(
        P1_U3133) );
  OAI22_X1 U24242 ( .A1(n21327), .A2(n21355), .B1(n21274), .B2(n21284), .ZN(
        n21275) );
  INV_X1 U24243 ( .A(n21275), .ZN(n21277) );
  AOI22_X1 U24244 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21288), .B1(
        n21287), .B2(n21352), .ZN(n21276) );
  OAI211_X1 U24245 ( .C1(n21292), .C2(n21278), .A(n21277), .B(n21276), .ZN(
        P1_U3134) );
  OAI22_X1 U24246 ( .A1(n21327), .A2(n21359), .B1(n21279), .B2(n21284), .ZN(
        n21280) );
  INV_X1 U24247 ( .A(n21280), .ZN(n21282) );
  AOI22_X1 U24248 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21288), .B1(
        n21287), .B2(n21356), .ZN(n21281) );
  OAI211_X1 U24249 ( .C1(n21292), .C2(n21283), .A(n21282), .B(n21281), .ZN(
        P1_U3135) );
  OAI22_X1 U24250 ( .A1(n21327), .A2(n21367), .B1(n21285), .B2(n21284), .ZN(
        n21286) );
  INV_X1 U24251 ( .A(n21286), .ZN(n21290) );
  AOI22_X1 U24252 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21288), .B1(
        n21287), .B2(n21362), .ZN(n21289) );
  OAI211_X1 U24253 ( .C1(n21292), .C2(n21291), .A(n21290), .B(n21289), .ZN(
        P1_U3136) );
  NOR3_X2 U24254 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21294), .A3(
        n21371), .ZN(n21322) );
  AOI21_X1 U24255 ( .B1(n21370), .B2(n21295), .A(n21322), .ZN(n21297) );
  NOR2_X1 U24256 ( .A1(n21371), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21299) );
  INV_X1 U24257 ( .A(n21299), .ZN(n21296) );
  OAI22_X1 U24258 ( .A1(n21297), .A2(n21382), .B1(n21296), .B2(n21373), .ZN(
        n21323) );
  AOI22_X1 U24259 ( .A1(n21323), .A2(n21376), .B1(n21375), .B2(n21322), .ZN(
        n21303) );
  INV_X1 U24260 ( .A(n21298), .ZN(n21300) );
  AOI22_X1 U24261 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21324), .B1(
        n21363), .B2(n21385), .ZN(n21302) );
  OAI211_X1 U24262 ( .C1(n21388), .C2(n21327), .A(n21303), .B(n21302), .ZN(
        P1_U3137) );
  AOI22_X1 U24263 ( .A1(n21323), .A2(n21390), .B1(n21389), .B2(n21322), .ZN(
        n21306) );
  AOI22_X1 U24264 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21324), .B1(
        n21363), .B2(n21304), .ZN(n21305) );
  OAI211_X1 U24265 ( .C1(n21307), .C2(n21327), .A(n21306), .B(n21305), .ZN(
        P1_U3138) );
  AOI22_X1 U24266 ( .A1(n21323), .A2(n21396), .B1(n21395), .B2(n21322), .ZN(
        n21309) );
  AOI22_X1 U24267 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21324), .B1(
        n21363), .B2(n21397), .ZN(n21308) );
  OAI211_X1 U24268 ( .C1(n21400), .C2(n21327), .A(n21309), .B(n21308), .ZN(
        P1_U3139) );
  AOI22_X1 U24269 ( .A1(n21323), .A2(n21402), .B1(n21401), .B2(n21322), .ZN(
        n21312) );
  AOI22_X1 U24270 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21324), .B1(
        n21363), .B2(n21310), .ZN(n21311) );
  OAI211_X1 U24271 ( .C1(n21313), .C2(n21327), .A(n21312), .B(n21311), .ZN(
        P1_U3140) );
  AOI22_X1 U24272 ( .A1(n21323), .A2(n21408), .B1(n21407), .B2(n21322), .ZN(
        n21316) );
  AOI22_X1 U24273 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21324), .B1(
        n21363), .B2(n21314), .ZN(n21315) );
  OAI211_X1 U24274 ( .C1(n21317), .C2(n21327), .A(n21316), .B(n21315), .ZN(
        P1_U3141) );
  AOI22_X1 U24275 ( .A1(n21323), .A2(n21416), .B1(n21415), .B2(n21322), .ZN(
        n21319) );
  AOI22_X1 U24276 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21324), .B1(
        n21363), .B2(n21417), .ZN(n21318) );
  OAI211_X1 U24277 ( .C1(n21420), .C2(n21327), .A(n21319), .B(n21318), .ZN(
        P1_U3142) );
  AOI22_X1 U24278 ( .A1(n21323), .A2(n21422), .B1(n21421), .B2(n21322), .ZN(
        n21321) );
  AOI22_X1 U24279 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21324), .B1(
        n21363), .B2(n21423), .ZN(n21320) );
  OAI211_X1 U24280 ( .C1(n21426), .C2(n21327), .A(n21321), .B(n21320), .ZN(
        P1_U3143) );
  AOI22_X1 U24281 ( .A1(n21323), .A2(n21429), .B1(n21427), .B2(n21322), .ZN(
        n21326) );
  AOI22_X1 U24282 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21324), .B1(
        n21363), .B2(n21431), .ZN(n21325) );
  OAI211_X1 U24283 ( .C1(n21437), .C2(n21327), .A(n21326), .B(n21325), .ZN(
        P1_U3144) );
  NAND2_X1 U24284 ( .A1(n21370), .A2(n21329), .ZN(n21333) );
  INV_X1 U24285 ( .A(n21330), .ZN(n21332) );
  OAI22_X1 U24286 ( .A1(n21333), .A2(n21382), .B1(n21332), .B2(n21331), .ZN(
        n21361) );
  NOR3_X2 U24287 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21372), .A3(
        n21371), .ZN(n21360) );
  AOI22_X1 U24288 ( .A1(n21361), .A2(n21376), .B1(n21375), .B2(n21360), .ZN(
        n21340) );
  OAI21_X1 U24289 ( .B1(n21363), .B2(n21410), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21334) );
  AOI21_X1 U24290 ( .B1(n21334), .B2(n21333), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21337) );
  AOI22_X1 U24291 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21338), .ZN(n21339) );
  OAI211_X1 U24292 ( .C1(n21341), .C2(n21436), .A(n21340), .B(n21339), .ZN(
        P1_U3145) );
  AOI22_X1 U24293 ( .A1(n21361), .A2(n21390), .B1(n21389), .B2(n21360), .ZN(
        n21343) );
  AOI22_X1 U24294 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21391), .ZN(n21342) );
  OAI211_X1 U24295 ( .C1(n21394), .C2(n21436), .A(n21343), .B(n21342), .ZN(
        P1_U3146) );
  AOI22_X1 U24296 ( .A1(n21361), .A2(n21396), .B1(n21395), .B2(n21360), .ZN(
        n21346) );
  AOI22_X1 U24297 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21344), .ZN(n21345) );
  OAI211_X1 U24298 ( .C1(n21347), .C2(n21436), .A(n21346), .B(n21345), .ZN(
        P1_U3147) );
  AOI22_X1 U24299 ( .A1(n21361), .A2(n21402), .B1(n21401), .B2(n21360), .ZN(
        n21349) );
  AOI22_X1 U24300 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21403), .ZN(n21348) );
  OAI211_X1 U24301 ( .C1(n21406), .C2(n21436), .A(n21349), .B(n21348), .ZN(
        P1_U3148) );
  AOI22_X1 U24302 ( .A1(n21361), .A2(n21408), .B1(n21407), .B2(n21360), .ZN(
        n21351) );
  AOI22_X1 U24303 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21409), .ZN(n21350) );
  OAI211_X1 U24304 ( .C1(n21414), .C2(n21436), .A(n21351), .B(n21350), .ZN(
        P1_U3149) );
  AOI22_X1 U24305 ( .A1(n21361), .A2(n21416), .B1(n21415), .B2(n21360), .ZN(
        n21354) );
  AOI22_X1 U24306 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21352), .ZN(n21353) );
  OAI211_X1 U24307 ( .C1(n21355), .C2(n21436), .A(n21354), .B(n21353), .ZN(
        P1_U3150) );
  AOI22_X1 U24308 ( .A1(n21361), .A2(n21422), .B1(n21421), .B2(n21360), .ZN(
        n21358) );
  AOI22_X1 U24309 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21356), .ZN(n21357) );
  OAI211_X1 U24310 ( .C1(n21359), .C2(n21436), .A(n21358), .B(n21357), .ZN(
        P1_U3151) );
  AOI22_X1 U24311 ( .A1(n21361), .A2(n21429), .B1(n21427), .B2(n21360), .ZN(
        n21366) );
  AOI22_X1 U24312 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21362), .ZN(n21365) );
  OAI211_X1 U24313 ( .C1(n21367), .C2(n21436), .A(n21366), .B(n21365), .ZN(
        P1_U3152) );
  INV_X1 U24314 ( .A(n21368), .ZN(n21428) );
  AOI21_X1 U24315 ( .B1(n21370), .B2(n21369), .A(n21428), .ZN(n21377) );
  NOR2_X1 U24316 ( .A1(n21372), .A2(n21371), .ZN(n21383) );
  INV_X1 U24317 ( .A(n21383), .ZN(n21374) );
  OAI22_X1 U24318 ( .A1(n21377), .A2(n21382), .B1(n21374), .B2(n21373), .ZN(
        n21430) );
  AOI22_X1 U24319 ( .A1(n21430), .A2(n21376), .B1(n21428), .B2(n21375), .ZN(
        n21387) );
  OAI21_X1 U24320 ( .B1(n21379), .B2(n21378), .A(n21377), .ZN(n21381) );
  OAI221_X1 U24321 ( .B1(n21384), .B2(n21383), .C1(n21382), .C2(n21381), .A(
        n21380), .ZN(n21433) );
  AOI22_X1 U24322 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21433), .B1(
        n21432), .B2(n21385), .ZN(n21386) );
  OAI211_X1 U24323 ( .C1(n21388), .C2(n21436), .A(n21387), .B(n21386), .ZN(
        P1_U3153) );
  AOI22_X1 U24324 ( .A1(n21430), .A2(n21390), .B1(n21428), .B2(n21389), .ZN(
        n21393) );
  AOI22_X1 U24325 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21433), .B1(
        n21410), .B2(n21391), .ZN(n21392) );
  OAI211_X1 U24326 ( .C1(n21394), .C2(n21413), .A(n21393), .B(n21392), .ZN(
        P1_U3154) );
  AOI22_X1 U24327 ( .A1(n21430), .A2(n21396), .B1(n21428), .B2(n21395), .ZN(
        n21399) );
  AOI22_X1 U24328 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21433), .B1(
        n21432), .B2(n21397), .ZN(n21398) );
  OAI211_X1 U24329 ( .C1(n21400), .C2(n21436), .A(n21399), .B(n21398), .ZN(
        P1_U3155) );
  AOI22_X1 U24330 ( .A1(n21430), .A2(n21402), .B1(n21428), .B2(n21401), .ZN(
        n21405) );
  AOI22_X1 U24331 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21433), .B1(
        n21410), .B2(n21403), .ZN(n21404) );
  OAI211_X1 U24332 ( .C1(n21406), .C2(n21413), .A(n21405), .B(n21404), .ZN(
        P1_U3156) );
  AOI22_X1 U24333 ( .A1(n21430), .A2(n21408), .B1(n21428), .B2(n21407), .ZN(
        n21412) );
  AOI22_X1 U24334 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21433), .B1(
        n21410), .B2(n21409), .ZN(n21411) );
  OAI211_X1 U24335 ( .C1(n21414), .C2(n21413), .A(n21412), .B(n21411), .ZN(
        P1_U3157) );
  AOI22_X1 U24336 ( .A1(n21430), .A2(n21416), .B1(n21428), .B2(n21415), .ZN(
        n21419) );
  AOI22_X1 U24337 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21433), .B1(
        n21432), .B2(n21417), .ZN(n21418) );
  OAI211_X1 U24338 ( .C1(n21420), .C2(n21436), .A(n21419), .B(n21418), .ZN(
        P1_U3158) );
  AOI22_X1 U24339 ( .A1(n21430), .A2(n21422), .B1(n21428), .B2(n21421), .ZN(
        n21425) );
  AOI22_X1 U24340 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21433), .B1(
        n21432), .B2(n21423), .ZN(n21424) );
  OAI211_X1 U24341 ( .C1(n21426), .C2(n21436), .A(n21425), .B(n21424), .ZN(
        P1_U3159) );
  AOI22_X1 U24342 ( .A1(n21430), .A2(n21429), .B1(n21428), .B2(n21427), .ZN(
        n21435) );
  AOI22_X1 U24343 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21433), .B1(
        n21432), .B2(n21431), .ZN(n21434) );
  OAI211_X1 U24344 ( .C1(n21437), .C2(n21436), .A(n21435), .B(n21434), .ZN(
        P1_U3160) );
  AND2_X1 U24345 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21507), .ZN(
        P1_U3164) );
  NOR2_X1 U24346 ( .A1(n21510), .A2(n21613), .ZN(P1_U3165) );
  AND2_X1 U24347 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21507), .ZN(
        P1_U3166) );
  AND2_X1 U24348 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21507), .ZN(
        P1_U3167) );
  AND2_X1 U24349 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21507), .ZN(
        P1_U3168) );
  AND2_X1 U24350 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21507), .ZN(
        P1_U3169) );
  AND2_X1 U24351 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21507), .ZN(
        P1_U3170) );
  AND2_X1 U24352 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21507), .ZN(
        P1_U3171) );
  AND2_X1 U24353 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21507), .ZN(
        P1_U3172) );
  AND2_X1 U24354 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21507), .ZN(
        P1_U3173) );
  AND2_X1 U24355 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21507), .ZN(
        P1_U3174) );
  AND2_X1 U24356 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21507), .ZN(
        P1_U3175) );
  AND2_X1 U24357 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21507), .ZN(
        P1_U3176) );
  AND2_X1 U24358 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21507), .ZN(
        P1_U3177) );
  AND2_X1 U24359 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21507), .ZN(
        P1_U3178) );
  AND2_X1 U24360 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21507), .ZN(
        P1_U3179) );
  AND2_X1 U24361 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21507), .ZN(
        P1_U3180) );
  NOR2_X1 U24362 ( .A1(n21510), .A2(n21586), .ZN(P1_U3181) );
  AND2_X1 U24363 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21507), .ZN(
        P1_U3182) );
  AND2_X1 U24364 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21507), .ZN(
        P1_U3183) );
  AND2_X1 U24365 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21507), .ZN(
        P1_U3184) );
  INV_X1 U24366 ( .A(P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n21667) );
  NOR2_X1 U24367 ( .A1(n21510), .A2(n21667), .ZN(P1_U3185) );
  AND2_X1 U24368 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21507), .ZN(P1_U3186) );
  AND2_X1 U24369 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21507), .ZN(P1_U3187) );
  AND2_X1 U24370 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21507), .ZN(P1_U3188) );
  AND2_X1 U24371 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21507), .ZN(P1_U3189) );
  AND2_X1 U24372 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21507), .ZN(P1_U3190) );
  AND2_X1 U24373 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21507), .ZN(P1_U3191) );
  AND2_X1 U24374 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21507), .ZN(P1_U3192) );
  AND2_X1 U24375 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21507), .ZN(P1_U3193) );
  AOI21_X1 U24376 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21447), .A(n21442), 
        .ZN(n21451) );
  OAI21_X1 U24377 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(HOLD), .ZN(n21438) );
  OAI211_X1 U24378 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n21446), .A(n21438), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21439) );
  INV_X1 U24379 ( .A(n21439), .ZN(n21440) );
  OAI22_X1 U24380 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21451), .B1(n21531), 
        .B2(n21440), .ZN(P1_U3194) );
  OAI21_X1 U24381 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21446), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n21450) );
  AOI211_X1 U24382 ( .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(n21452), .A(
        n21442), .B(n21441), .ZN(n21445) );
  AOI21_X1 U24383 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21443), .A(n21445), 
        .ZN(n21449) );
  AOI22_X1 U24384 ( .A1(n21447), .A2(n21446), .B1(n21445), .B2(n21444), .ZN(
        n21448) );
  OAI22_X1 U24385 ( .A1(n21451), .A2(n21450), .B1(n21449), .B2(n21448), .ZN(
        P1_U3196) );
  NAND2_X1 U24386 ( .A1(n21531), .A2(n21452), .ZN(n21500) );
  INV_X1 U24387 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21453) );
  NAND2_X1 U24388 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21531), .ZN(n21497) );
  OAI222_X1 U24389 ( .A1(n21500), .A2(n14260), .B1(n21453), .B2(n21531), .C1(
        n15246), .C2(n21497), .ZN(P1_U3197) );
  INV_X1 U24390 ( .A(n21497), .ZN(n21502) );
  AOI222_X1 U24391 ( .A1(n21502), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21532), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21501), .ZN(n21454) );
  INV_X1 U24392 ( .A(n21454), .ZN(P1_U3198) );
  AOI222_X1 U24393 ( .A1(n21502), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n21532), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21501), .ZN(n21455) );
  INV_X1 U24394 ( .A(n21455), .ZN(P1_U3199) );
  AOI22_X1 U24395 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n21532), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n21501), .ZN(n21456) );
  OAI21_X1 U24396 ( .B1(n21457), .B2(n21497), .A(n21456), .ZN(P1_U3200) );
  AOI22_X1 U24397 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n21532), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n21501), .ZN(n21458) );
  OAI21_X1 U24398 ( .B1(n17520), .B2(n21497), .A(n21458), .ZN(P1_U3201) );
  INV_X1 U24399 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21460) );
  AOI22_X1 U24400 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n21532), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n21501), .ZN(n21459) );
  OAI21_X1 U24401 ( .B1(n21460), .B2(n21497), .A(n21459), .ZN(P1_U3202) );
  AOI22_X1 U24402 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21532), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n21502), .ZN(n21461) );
  OAI21_X1 U24403 ( .B1(n21623), .B2(n21500), .A(n21461), .ZN(P1_U3203) );
  INV_X1 U24404 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21462) );
  OAI222_X1 U24405 ( .A1(n21500), .A2(n21464), .B1(n21462), .B2(n21531), .C1(
        n21623), .C2(n21497), .ZN(P1_U3204) );
  INV_X1 U24406 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21463) );
  OAI222_X1 U24407 ( .A1(n21497), .A2(n21464), .B1(n21463), .B2(n21531), .C1(
        n15216), .C2(n21500), .ZN(P1_U3205) );
  INV_X1 U24408 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21465) );
  OAI222_X1 U24409 ( .A1(n21500), .A2(n21466), .B1(n21465), .B2(n21531), .C1(
        n15216), .C2(n21497), .ZN(P1_U3206) );
  AOI222_X1 U24410 ( .A1(n21502), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21532), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21501), .ZN(n21467) );
  INV_X1 U24411 ( .A(n21467), .ZN(P1_U3207) );
  AOI222_X1 U24412 ( .A1(n21502), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n21532), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n21501), .ZN(n21468) );
  INV_X1 U24413 ( .A(n21468), .ZN(P1_U3208) );
  INV_X1 U24414 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21469) );
  INV_X1 U24415 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21472) );
  OAI222_X1 U24416 ( .A1(n21497), .A2(n21470), .B1(n21469), .B2(n21531), .C1(
        n21472), .C2(n21500), .ZN(P1_U3209) );
  INV_X1 U24417 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21471) );
  INV_X1 U24418 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21473) );
  OAI222_X1 U24419 ( .A1(n21497), .A2(n21472), .B1(n21471), .B2(n21531), .C1(
        n21473), .C2(n21500), .ZN(P1_U3210) );
  INV_X1 U24420 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21474) );
  OAI222_X1 U24421 ( .A1(n21500), .A2(n21476), .B1(n21474), .B2(n21531), .C1(
        n21473), .C2(n21497), .ZN(P1_U3211) );
  AOI22_X1 U24422 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21532), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21501), .ZN(n21475) );
  OAI21_X1 U24423 ( .B1(n21476), .B2(n21497), .A(n21475), .ZN(P1_U3212) );
  AOI22_X1 U24424 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21532), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21502), .ZN(n21477) );
  OAI21_X1 U24425 ( .B1(n21479), .B2(n21500), .A(n21477), .ZN(P1_U3213) );
  INV_X1 U24426 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21478) );
  OAI222_X1 U24427 ( .A1(n21497), .A2(n21479), .B1(n21478), .B2(n21531), .C1(
        n21480), .C2(n21500), .ZN(P1_U3214) );
  INV_X1 U24428 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n21669) );
  INV_X1 U24429 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21482) );
  OAI222_X1 U24430 ( .A1(n21497), .A2(n21480), .B1(n21669), .B2(n21531), .C1(
        n21482), .C2(n21500), .ZN(P1_U3215) );
  INV_X1 U24431 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21481) );
  OAI222_X1 U24432 ( .A1(n21497), .A2(n21482), .B1(n21481), .B2(n21531), .C1(
        n21484), .C2(n21500), .ZN(P1_U3216) );
  INV_X1 U24433 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21483) );
  OAI222_X1 U24434 ( .A1(n21497), .A2(n21484), .B1(n21483), .B2(n21531), .C1(
        n21486), .C2(n21500), .ZN(P1_U3217) );
  AOI22_X1 U24435 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21532), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21501), .ZN(n21485) );
  OAI21_X1 U24436 ( .B1(n21486), .B2(n21497), .A(n21485), .ZN(P1_U3218) );
  AOI22_X1 U24437 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21532), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21502), .ZN(n21487) );
  OAI21_X1 U24438 ( .B1(n21489), .B2(n21500), .A(n21487), .ZN(P1_U3219) );
  INV_X1 U24439 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21488) );
  OAI222_X1 U24440 ( .A1(n21497), .A2(n21489), .B1(n21488), .B2(n21531), .C1(
        n21491), .C2(n21500), .ZN(P1_U3220) );
  INV_X1 U24441 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21490) );
  OAI222_X1 U24442 ( .A1(n21497), .A2(n21491), .B1(n21490), .B2(n21531), .C1(
        n21493), .C2(n21500), .ZN(P1_U3221) );
  INV_X1 U24443 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21492) );
  OAI222_X1 U24444 ( .A1(n21497), .A2(n21493), .B1(n21492), .B2(n21531), .C1(
        n21495), .C2(n21500), .ZN(P1_U3222) );
  AOI22_X1 U24445 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n21501), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21532), .ZN(n21494) );
  OAI21_X1 U24446 ( .B1(n21495), .B2(n21497), .A(n21494), .ZN(P1_U3223) );
  AOI22_X1 U24447 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n21502), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21532), .ZN(n21496) );
  OAI21_X1 U24448 ( .B1(n21498), .B2(n21500), .A(n21496), .ZN(P1_U3224) );
  INV_X1 U24449 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21499) );
  INV_X1 U24450 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n21656) );
  OAI222_X1 U24451 ( .A1(n21500), .A2(n21499), .B1(n21656), .B2(n21531), .C1(
        n21498), .C2(n21497), .ZN(P1_U3225) );
  AOI222_X1 U24452 ( .A1(n21502), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21532), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21501), .ZN(n21503) );
  INV_X1 U24453 ( .A(n21503), .ZN(P1_U3226) );
  INV_X1 U24454 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21504) );
  AOI22_X1 U24455 ( .A1(n21531), .A2(n21505), .B1(n21504), .B2(n21532), .ZN(
        P1_U3458) );
  MUX2_X1 U24456 ( .A(P1_BE_N_REG_2__SCAN_IN), .B(P1_BYTEENABLE_REG_2__SCAN_IN), .S(n21531), .Z(P1_U3459) );
  MUX2_X1 U24457 ( .A(P1_BE_N_REG_1__SCAN_IN), .B(P1_BYTEENABLE_REG_1__SCAN_IN), .S(n21531), .Z(P1_U3460) );
  MUX2_X1 U24458 ( .A(P1_BE_N_REG_0__SCAN_IN), .B(P1_BYTEENABLE_REG_0__SCAN_IN), .S(n21531), .Z(P1_U3461) );
  INV_X1 U24459 ( .A(n21508), .ZN(n21506) );
  AOI21_X1 U24460 ( .B1(n21515), .B2(n21507), .A(n21506), .ZN(P1_U3464) );
  OAI21_X1 U24461 ( .B1(n21510), .B2(n21509), .A(n21508), .ZN(P1_U3465) );
  NAND2_X1 U24462 ( .A1(n21511), .A2(n15246), .ZN(n21517) );
  AND2_X1 U24463 ( .A1(n21518), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n21512) );
  AOI22_X1 U24464 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(n21513), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n21512), .ZN(n21514) );
  OAI221_X1 U24465 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21516), .C1(n21515), .C2(n21517), .A(n21514), .ZN(P1_U3481) );
  OAI21_X1 U24466 ( .B1(n21518), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21517), 
        .ZN(n21519) );
  INV_X1 U24467 ( .A(n21519), .ZN(P1_U3482) );
  AOI22_X1 U24468 ( .A1(n21531), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21520), 
        .B2(n21532), .ZN(P1_U3483) );
  AOI211_X1 U24469 ( .C1(n21524), .C2(n21523), .A(n21522), .B(n21521), .ZN(
        n21530) );
  OAI211_X1 U24470 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n10084), .A(n21525), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21527) );
  AOI21_X1 U24471 ( .B1(n21527), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n21526), 
        .ZN(n21529) );
  NAND2_X1 U24472 ( .A1(n21530), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21528) );
  OAI21_X1 U24473 ( .B1(n21530), .B2(n21529), .A(n21528), .ZN(P1_U3485) );
  OAI22_X1 U24474 ( .A1(n21532), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n21531), .ZN(n21533) );
  INV_X1 U24475 ( .A(n21533), .ZN(P1_U3486) );
  NAND4_X1 U24476 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), 
        .A4(P3_UWORD_REG_2__SCAN_IN), .ZN(n21537) );
  NAND4_X1 U24477 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_EBX_REG_26__SCAN_IN), .A3(P3_ADDRESS_REG_29__SCAN_IN), .A4(n21674), 
        .ZN(n21536) );
  NAND4_X1 U24478 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(P1_DATAO_REG_24__SCAN_IN), .A4(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n21535) );
  NAND4_X1 U24479 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_EBX_REG_18__SCAN_IN), .A3(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A4(
        n21658), .ZN(n21534) );
  NOR4_X1 U24480 ( .A1(n21537), .A2(n21536), .A3(n21535), .A4(n21534), .ZN(
        n21687) );
  NAND3_X1 U24481 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n21557), .A3(n21558), 
        .ZN(n21555) );
  INV_X1 U24482 ( .A(n21538), .ZN(n21541) );
  NOR4_X1 U24483 ( .A1(P2_EBX_REG_3__SCAN_IN), .A2(P1_EAX_REG_27__SCAN_IN), 
        .A3(n21571), .A4(n21575), .ZN(n21540) );
  NOR4_X1 U24484 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(
        P1_EBX_REG_27__SCAN_IN), .A3(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n21539) );
  NAND4_X1 U24485 ( .A1(n21542), .A2(n21541), .A3(n21540), .A4(n21539), .ZN(
        n21554) );
  NOR4_X1 U24486 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(
        P1_LWORD_REG_13__SCAN_IN), .A3(P1_LWORD_REG_5__SCAN_IN), .A4(n21602), 
        .ZN(n21552) );
  INV_X1 U24487 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21577) );
  NAND4_X1 U24488 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(BUF1_REG_26__SCAN_IN), 
        .A3(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n21577), .ZN(n21545) );
  NAND3_X1 U24489 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_5__4__SCAN_IN), .A3(n21590), .ZN(n21544) );
  NAND4_X1 U24490 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_LWORD_REG_6__SCAN_IN), .A3(n21593), .A4(n21595), .ZN(n21543) );
  NOR4_X1 U24491 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21545), .A3(n21544), 
        .A4(n21543), .ZN(n21551) );
  NOR4_X1 U24492 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(P3_UWORD_REG_8__SCAN_IN), 
        .A3(n21646), .A4(n21645), .ZN(n21550) );
  INV_X1 U24493 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n21607) );
  NAND4_X1 U24494 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_30__SCAN_IN), .A3(P2_DATAO_REG_11__SCAN_IN), .A4(
        n21607), .ZN(n21548) );
  NAND3_X1 U24495 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_ADDRESS_REG_2__SCAN_IN), .A3(n21639), .ZN(n21547) );
  NAND4_X1 U24496 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_8__3__SCAN_IN), .A3(P3_PHYADDRPOINTER_REG_8__SCAN_IN), 
        .A4(n21623), .ZN(n21546) );
  NOR4_X1 U24497 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(n21548), .A3(n21547), 
        .A4(n21546), .ZN(n21549) );
  NAND4_X1 U24498 ( .A1(n21552), .A2(n21551), .A3(n21550), .A4(n21549), .ZN(
        n21553) );
  NOR4_X1 U24499 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n21555), .A3(n21554), 
        .A4(n21553), .ZN(n21686) );
  AOI22_X1 U24500 ( .A1(n21558), .A2(keyinput6), .B1(n21557), .B2(keyinput39), 
        .ZN(n21556) );
  OAI221_X1 U24501 ( .B1(n21558), .B2(keyinput6), .C1(n21557), .C2(keyinput39), 
        .A(n21556), .ZN(n21569) );
  AOI22_X1 U24502 ( .A1(n21561), .A2(keyinput23), .B1(keyinput46), .B2(n21560), 
        .ZN(n21559) );
  OAI221_X1 U24503 ( .B1(n21561), .B2(keyinput23), .C1(n21560), .C2(keyinput46), .A(n21559), .ZN(n21568) );
  AOI22_X1 U24504 ( .A1(n21563), .A2(keyinput33), .B1(n13448), .B2(keyinput20), 
        .ZN(n21562) );
  OAI221_X1 U24505 ( .B1(n21563), .B2(keyinput33), .C1(n13448), .C2(keyinput20), .A(n21562), .ZN(n21567) );
  AOI22_X1 U24506 ( .A1(n18257), .A2(keyinput49), .B1(n21565), .B2(keyinput14), 
        .ZN(n21564) );
  OAI221_X1 U24507 ( .B1(n18257), .B2(keyinput49), .C1(n21565), .C2(keyinput14), .A(n21564), .ZN(n21566) );
  NOR4_X1 U24508 ( .A1(n21569), .A2(n21568), .A3(n21567), .A4(n21566), .ZN(
        n21620) );
  AOI22_X1 U24509 ( .A1(n21572), .A2(keyinput56), .B1(n21571), .B2(keyinput12), 
        .ZN(n21570) );
  OAI221_X1 U24510 ( .B1(n21572), .B2(keyinput56), .C1(n21571), .C2(keyinput12), .A(n21570), .ZN(n21584) );
  AOI22_X1 U24511 ( .A1(n21575), .A2(keyinput51), .B1(n21574), .B2(keyinput13), 
        .ZN(n21573) );
  OAI221_X1 U24512 ( .B1(n21575), .B2(keyinput51), .C1(n21574), .C2(keyinput13), .A(n21573), .ZN(n21583) );
  AOI22_X1 U24513 ( .A1(n21577), .A2(keyinput57), .B1(keyinput40), .B2(n16706), 
        .ZN(n21576) );
  OAI221_X1 U24514 ( .B1(n21577), .B2(keyinput57), .C1(n16706), .C2(keyinput40), .A(n21576), .ZN(n21582) );
  AOI22_X1 U24515 ( .A1(n21580), .A2(keyinput59), .B1(keyinput24), .B2(n21579), 
        .ZN(n21578) );
  OAI221_X1 U24516 ( .B1(n21580), .B2(keyinput59), .C1(n21579), .C2(keyinput24), .A(n21578), .ZN(n21581) );
  NOR4_X1 U24517 ( .A1(n21584), .A2(n21583), .A3(n21582), .A4(n21581), .ZN(
        n21619) );
  AOI22_X1 U24518 ( .A1(n21587), .A2(keyinput19), .B1(keyinput30), .B2(n21586), 
        .ZN(n21585) );
  OAI221_X1 U24519 ( .B1(n21587), .B2(keyinput19), .C1(n21586), .C2(keyinput30), .A(n21585), .ZN(n21600) );
  INV_X1 U24520 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n21589) );
  AOI22_X1 U24521 ( .A1(n21590), .A2(keyinput15), .B1(n21589), .B2(keyinput10), 
        .ZN(n21588) );
  OAI221_X1 U24522 ( .B1(n21590), .B2(keyinput15), .C1(n21589), .C2(keyinput10), .A(n21588), .ZN(n21599) );
  AOI22_X1 U24523 ( .A1(n21593), .A2(keyinput28), .B1(keyinput16), .B2(n21592), 
        .ZN(n21591) );
  OAI221_X1 U24524 ( .B1(n21593), .B2(keyinput28), .C1(n21592), .C2(keyinput16), .A(n21591), .ZN(n21598) );
  AOI22_X1 U24525 ( .A1(n21596), .A2(keyinput25), .B1(n21595), .B2(keyinput4), 
        .ZN(n21594) );
  OAI221_X1 U24526 ( .B1(n21596), .B2(keyinput25), .C1(n21595), .C2(keyinput4), 
        .A(n21594), .ZN(n21597) );
  NOR4_X1 U24527 ( .A1(n21600), .A2(n21599), .A3(n21598), .A4(n21597), .ZN(
        n21618) );
  AOI22_X1 U24528 ( .A1(n21603), .A2(keyinput32), .B1(n21602), .B2(keyinput52), 
        .ZN(n21601) );
  OAI221_X1 U24529 ( .B1(n21603), .B2(keyinput32), .C1(n21602), .C2(keyinput52), .A(n21601), .ZN(n21616) );
  AOI22_X1 U24530 ( .A1(n21606), .A2(keyinput45), .B1(n21605), .B2(keyinput43), 
        .ZN(n21604) );
  OAI221_X1 U24531 ( .B1(n21606), .B2(keyinput45), .C1(n21605), .C2(keyinput43), .A(n21604), .ZN(n21610) );
  XNOR2_X1 U24532 ( .A(n21607), .B(keyinput41), .ZN(n21609) );
  XOR2_X1 U24533 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B(keyinput18), .Z(
        n21608) );
  OR3_X1 U24534 ( .A1(n21610), .A2(n21609), .A3(n21608), .ZN(n21615) );
  AOI22_X1 U24535 ( .A1(n21613), .A2(keyinput61), .B1(keyinput35), .B2(n21612), 
        .ZN(n21611) );
  OAI221_X1 U24536 ( .B1(n21613), .B2(keyinput61), .C1(n21612), .C2(keyinput35), .A(n21611), .ZN(n21614) );
  NOR3_X1 U24537 ( .A1(n21616), .A2(n21615), .A3(n21614), .ZN(n21617) );
  NAND4_X1 U24538 ( .A1(n21620), .A2(n21619), .A3(n21618), .A4(n21617), .ZN(
        n21685) );
  AOI22_X1 U24539 ( .A1(n21623), .A2(keyinput5), .B1(keyinput48), .B2(n21622), 
        .ZN(n21621) );
  OAI221_X1 U24540 ( .B1(n21623), .B2(keyinput5), .C1(n21622), .C2(keyinput48), 
        .A(n21621), .ZN(n21634) );
  AOI22_X1 U24541 ( .A1(n21626), .A2(keyinput11), .B1(n21625), .B2(keyinput7), 
        .ZN(n21624) );
  OAI221_X1 U24542 ( .B1(n21626), .B2(keyinput11), .C1(n21625), .C2(keyinput7), 
        .A(n21624), .ZN(n21633) );
  XNOR2_X1 U24543 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B(keyinput50), .ZN(
        n21629) );
  XNOR2_X1 U24544 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput54), 
        .ZN(n21628) );
  XNOR2_X1 U24545 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B(keyinput62), .ZN(
        n21627) );
  NAND3_X1 U24546 ( .A1(n21629), .A2(n21628), .A3(n21627), .ZN(n21632) );
  XNOR2_X1 U24547 ( .A(n21630), .B(keyinput3), .ZN(n21631) );
  NOR4_X1 U24548 ( .A1(n21634), .A2(n21633), .A3(n21632), .A4(n21631), .ZN(
        n21683) );
  AOI22_X1 U24549 ( .A1(n21637), .A2(keyinput26), .B1(n21636), .B2(keyinput2), 
        .ZN(n21635) );
  OAI221_X1 U24550 ( .B1(n21637), .B2(keyinput26), .C1(n21636), .C2(keyinput2), 
        .A(n21635), .ZN(n21650) );
  AOI22_X1 U24551 ( .A1(n21640), .A2(keyinput1), .B1(keyinput60), .B2(n21639), 
        .ZN(n21638) );
  OAI221_X1 U24552 ( .B1(n21640), .B2(keyinput1), .C1(n21639), .C2(keyinput60), 
        .A(n21638), .ZN(n21649) );
  AOI22_X1 U24553 ( .A1(n21643), .A2(keyinput21), .B1(n21642), .B2(keyinput37), 
        .ZN(n21641) );
  OAI221_X1 U24554 ( .B1(n21643), .B2(keyinput21), .C1(n21642), .C2(keyinput37), .A(n21641), .ZN(n21648) );
  AOI22_X1 U24555 ( .A1(n21646), .A2(keyinput38), .B1(keyinput36), .B2(n21645), 
        .ZN(n21644) );
  OAI221_X1 U24556 ( .B1(n21646), .B2(keyinput38), .C1(n21645), .C2(keyinput36), .A(n21644), .ZN(n21647) );
  NOR4_X1 U24557 ( .A1(n21650), .A2(n21649), .A3(n21648), .A4(n21647), .ZN(
        n21682) );
  AOI22_X1 U24558 ( .A1(n21653), .A2(keyinput8), .B1(n21652), .B2(keyinput44), 
        .ZN(n21651) );
  OAI221_X1 U24559 ( .B1(n21653), .B2(keyinput8), .C1(n21652), .C2(keyinput44), 
        .A(n21651), .ZN(n21664) );
  AOI22_X1 U24560 ( .A1(n21656), .A2(keyinput53), .B1(keyinput34), .B2(n21655), 
        .ZN(n21654) );
  OAI221_X1 U24561 ( .B1(n21656), .B2(keyinput53), .C1(n21655), .C2(keyinput34), .A(n21654), .ZN(n21663) );
  AOI22_X1 U24562 ( .A1(n11856), .A2(keyinput9), .B1(keyinput27), .B2(n21658), 
        .ZN(n21657) );
  OAI221_X1 U24563 ( .B1(n11856), .B2(keyinput9), .C1(n21658), .C2(keyinput27), 
        .A(n21657), .ZN(n21662) );
  AOI22_X1 U24564 ( .A1(n21660), .A2(keyinput17), .B1(n10967), .B2(keyinput29), 
        .ZN(n21659) );
  OAI221_X1 U24565 ( .B1(n21660), .B2(keyinput17), .C1(n10967), .C2(keyinput29), .A(n21659), .ZN(n21661) );
  NOR4_X1 U24566 ( .A1(n21664), .A2(n21663), .A3(n21662), .A4(n21661), .ZN(
        n21681) );
  AOI22_X1 U24567 ( .A1(n21667), .A2(keyinput22), .B1(n21666), .B2(keyinput58), 
        .ZN(n21665) );
  OAI221_X1 U24568 ( .B1(n21667), .B2(keyinput22), .C1(n21666), .C2(keyinput58), .A(n21665), .ZN(n21679) );
  AOI22_X1 U24569 ( .A1(n15322), .A2(keyinput47), .B1(keyinput63), .B2(n21669), 
        .ZN(n21668) );
  OAI221_X1 U24570 ( .B1(n15322), .B2(keyinput47), .C1(n21669), .C2(keyinput63), .A(n21668), .ZN(n21678) );
  AOI22_X1 U24571 ( .A1(n21672), .A2(keyinput55), .B1(keyinput0), .B2(n21671), 
        .ZN(n21670) );
  OAI221_X1 U24572 ( .B1(n21672), .B2(keyinput55), .C1(n21671), .C2(keyinput0), 
        .A(n21670), .ZN(n21677) );
  AOI22_X1 U24573 ( .A1(n21675), .A2(keyinput31), .B1(keyinput42), .B2(n21674), 
        .ZN(n21673) );
  OAI221_X1 U24574 ( .B1(n21675), .B2(keyinput31), .C1(n21674), .C2(keyinput42), .A(n21673), .ZN(n21676) );
  NOR4_X1 U24575 ( .A1(n21679), .A2(n21678), .A3(n21677), .A4(n21676), .ZN(
        n21680) );
  NAND4_X1 U24576 ( .A1(n21683), .A2(n21682), .A3(n21681), .A4(n21680), .ZN(
        n21684) );
  AOI211_X1 U24577 ( .C1(n21687), .C2(n21686), .A(n21685), .B(n21684), .ZN(
        n21698) );
  NOR2_X1 U24578 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20607), .ZN(
        n21694) );
  INV_X1 U24579 ( .A(n21688), .ZN(n21690) );
  OAI22_X1 U24580 ( .A1(n21692), .A2(n21691), .B1(n21690), .B2(n21689), .ZN(
        n21693) );
  NOR2_X1 U24581 ( .A1(n21694), .A2(n21693), .ZN(n21696) );
  MUX2_X1 U24582 ( .A(n20291), .B(n21696), .S(n21695), .Z(n21697) );
  XNOR2_X1 U24583 ( .A(n21698), .B(n21697), .ZN(P2_U3605) );
  BUF_X4 U11105 ( .A(n12263), .Z(n9552) );
  CLKBUF_X1 U11041 ( .A(n12953), .Z(n9583) );
  CLKBUF_X1 U11046 ( .A(n10623), .Z(n13299) );
  CLKBUF_X1 U11147 ( .A(n12112), .Z(n14446) );
  CLKBUF_X1 U12588 ( .A(n17632), .Z(n17638) );
  CLKBUF_X1 U12616 ( .A(n18633), .Z(n18639) );
endmodule

