

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9580, n9581, n9582, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
         n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
         n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
         n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574;

  INV_X1 U11024 ( .A(n18641), .ZN(n18728) );
  NOR2_X1 U11025 ( .A1(n20367), .A2(n20267), .ZN(n20311) );
  NAND2_X1 U11026 ( .A1(n16927), .A2(n16928), .ZN(n17026) );
  INV_X1 U11027 ( .A(n20610), .ZN(n16775) );
  BUF_X2 U11028 ( .A(n15292), .Z(n17366) );
  AND2_X1 U11029 ( .A1(n12629), .A2(n9606), .ZN(n14927) );
  NOR2_X1 U11030 ( .A1(n16008), .A2(n13186), .ZN(n13236) );
  NAND2_X2 U11031 ( .A1(n18978), .A2(n18991), .ZN(n19005) );
  AND2_X1 U11032 ( .A1(n17372), .A2(n17378), .ZN(n10496) );
  AND4_X1 U11033 ( .A1(n10866), .A2(n10867), .A3(n10868), .A4(n10864), .ZN(
        n9833) );
  OR2_X1 U11034 ( .A1(n13550), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17047) );
  CLKBUF_X2 U11036 ( .A(n13024), .Z(n19943) );
  OAI21_X2 U11037 ( .B1(n17445), .B2(n14157), .A(n13035), .ZN(n14704) );
  OAI21_X1 U11038 ( .B1(n14478), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12032), 
        .ZN(n9866) );
  CLKBUF_X2 U11039 ( .A(n12390), .Z(n14671) );
  INV_X1 U11040 ( .A(n14727), .ZN(n12525) );
  CLKBUF_X2 U11041 ( .A(n11931), .Z(n13692) );
  CLKBUF_X1 U11043 ( .A(n11874), .Z(n12911) );
  AND2_X1 U11044 ( .A1(n16746), .A2(n13133), .ZN(n10834) );
  AND2_X1 U11046 ( .A1(n12302), .A2(n14119), .ZN(n12450) );
  CLKBUF_X1 U11047 ( .A(n11954), .Z(n14275) );
  INV_X1 U11048 ( .A(n13514), .ZN(n18196) );
  NAND2_X1 U11049 ( .A1(n9942), .A2(n10739), .ZN(n10737) );
  CLKBUF_X1 U11050 ( .A(n11960), .Z(n14666) );
  NAND2_X1 U11051 ( .A1(n11895), .A2(n10610), .ZN(n11968) );
  CLKBUF_X3 U11053 ( .A(n9592), .Z(n9582) );
  AND2_X1 U11054 ( .A1(n11828), .A2(n11830), .ZN(n12098) );
  AND2_X1 U11055 ( .A1(n11830), .A2(n14087), .ZN(n11931) );
  AND2_X1 U11056 ( .A1(n11828), .A2(n14485), .ZN(n12117) );
  BUF_X1 U11057 ( .A(n12110), .Z(n9586) );
  AND2_X2 U11058 ( .A1(n11826), .A2(n11830), .ZN(n12116) );
  AND2_X2 U11059 ( .A1(n11826), .A2(n14481), .ZN(n11930) );
  AND2_X1 U11060 ( .A1(n11827), .A2(n11828), .ZN(n9592) );
  AND2_X2 U11061 ( .A1(n11819), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11826) );
  NAND3_X2 U11062 ( .A1(n10094), .A2(n10093), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10670) );
  AND2_X1 U11063 ( .A1(n11827), .A2(n11828), .ZN(n12110) );
  AND2_X1 U11066 ( .A1(n14087), .A2(n14485), .ZN(n12111) );
  NAND2_X1 U11067 ( .A1(n12047), .A2(n12046), .ZN(n12264) );
  AND4_X1 U11068 ( .A1(n10004), .A2(n10006), .A3(n10012), .A4(n10011), .ZN(
        n10003) );
  NAND2_X1 U11069 ( .A1(n12187), .A2(n12194), .ZN(n12620) );
  AND2_X1 U11070 ( .A1(n12133), .A2(n11897), .ZN(n12302) );
  OAI21_X1 U11071 ( .B1(n12620), .B2(n12275), .A(n12191), .ZN(n12192) );
  NAND2_X1 U11072 ( .A1(n10197), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12033) );
  AND2_X1 U11073 ( .A1(n10284), .A2(n12583), .ZN(n10283) );
  AND2_X1 U11074 ( .A1(n10807), .A2(n10591), .ZN(n10818) );
  BUF_X1 U11075 ( .A(n11961), .Z(n13652) );
  NAND2_X1 U11076 ( .A1(n14430), .A2(n12599), .ZN(n14410) );
  NAND3_X1 U11077 ( .A1(n12225), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n9972), .ZN(n12228) );
  NAND3_X1 U11078 ( .A1(n10064), .A2(n9960), .A3(n10568), .ZN(n12198) );
  XNOR2_X1 U11079 ( .A(n12192), .B(n21471), .ZN(n17378) );
  INV_X1 U11080 ( .A(n11118), .ZN(n11720) );
  INV_X1 U11081 ( .A(n11281), .ZN(n11426) );
  INV_X2 U11082 ( .A(n20006), .ZN(n13390) );
  OR2_X1 U11083 ( .A1(n10955), .A2(n10954), .ZN(n11076) );
  INV_X1 U11084 ( .A(n18202), .ZN(n17269) );
  AND2_X1 U11086 ( .A1(n17631), .A2(n17843), .ZN(n17617) );
  INV_X1 U11087 ( .A(n20750), .ZN(n20721) );
  BUF_X1 U11088 ( .A(n11968), .Z(n14207) );
  NAND2_X1 U11089 ( .A1(n12590), .A2(n12589), .ZN(n14186) );
  NAND2_X1 U11090 ( .A1(n14186), .A2(n14185), .ZN(n14430) );
  NAND2_X1 U11091 ( .A1(n15488), .A2(n15464), .ZN(n17401) );
  NAND2_X1 U11092 ( .A1(n12148), .A2(n12147), .ZN(n20889) );
  AND2_X1 U11094 ( .A1(n15663), .A2(n12530), .ZN(n13359) );
  INV_X1 U11095 ( .A(n20119), .ZN(n20467) );
  NOR2_X1 U11096 ( .A1(n20339), .A2(n20079), .ZN(n20325) );
  AND2_X1 U11097 ( .A1(n17573), .A2(n17843), .ZN(n17565) );
  INV_X1 U11098 ( .A(n18813), .ZN(n18780) );
  OR2_X1 U11099 ( .A1(n20797), .A2(n14275), .ZN(n14533) );
  NAND2_X1 U11100 ( .A1(n20405), .A2(n20404), .ZN(n20519) );
  INV_X1 U11101 ( .A(n17910), .ZN(n17918) );
  INV_X2 U11102 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14407) );
  OR2_X1 U11103 ( .A1(n13566), .A2(n18694), .ZN(n9580) );
  AND2_X1 U11104 ( .A1(n11830), .A2(n11829), .ZN(n11876) );
  AND2_X1 U11106 ( .A1(n11131), .A2(n9723), .ZN(n14601) );
  AND2_X2 U11107 ( .A1(n10046), .A2(n10084), .ZN(n9912) );
  AOI21_X2 U11108 ( .B1(n17309), .B2(n15968), .A(n17310), .ZN(n15734) );
  AOI21_X2 U11109 ( .B1(n11211), .B2(n11488), .A(n16268), .ZN(n11495) );
  AOI21_X2 U11110 ( .B1(n19538), .B2(n9682), .A(n14392), .ZN(n14388) );
  NAND2_X2 U11111 ( .A1(n18625), .A2(n18617), .ZN(n18614) );
  NOR2_X2 U11112 ( .A1(n11732), .A2(n11733), .ZN(n12554) );
  NAND2_X1 U11114 ( .A1(n12446), .A2(n14187), .ZN(n12361) );
  INV_X4 U11115 ( .A(n11598), .ZN(n9589) );
  NAND2_X4 U11116 ( .A1(n17144), .A2(n11536), .ZN(n11598) );
  XNOR2_X2 U11118 ( .A(n9916), .B(n9915), .ZN(n11182) );
  NOR3_X2 U11119 ( .A1(n19108), .A2(n13576), .A3(n13626), .ZN(n14385) );
  AND2_X4 U11120 ( .A1(n11533), .A2(n11532), .ZN(n18243) );
  BUF_X4 U11121 ( .A(n12110), .Z(n9587) );
  AND2_X2 U11122 ( .A1(n11821), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14481) );
  AND2_X1 U11123 ( .A1(n9913), .A2(n9914), .ZN(n11711) );
  INV_X1 U11124 ( .A(n18664), .ZN(n18684) );
  INV_X1 U11125 ( .A(n18808), .ZN(n18822) );
  INV_X1 U11126 ( .A(n18675), .ZN(n18686) );
  OR2_X1 U11127 ( .A1(n16799), .A2(n16797), .ZN(n20375) );
  OR2_X1 U11128 ( .A1(n16799), .A2(n16798), .ZN(n20465) );
  OR2_X1 U11129 ( .A1(n18817), .A2(n17098), .ZN(n18602) );
  AND3_X1 U11130 ( .A1(n15941), .A2(n16768), .A3(n10808), .ZN(n10889) );
  INV_X2 U11131 ( .A(n18810), .ZN(n18769) );
  OR2_X1 U11132 ( .A1(n10815), .A2(n13030), .ZN(n10812) );
  OAI21_X2 U11133 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19702), .A(n17547), 
        .ZN(n18810) );
  AND3_X1 U11134 ( .A1(n16768), .A2(n16733), .A3(n10817), .ZN(n20085) );
  NOR2_X1 U11135 ( .A1(n20829), .A2(n20959), .ZN(n21312) );
  INV_X1 U11136 ( .A(n10805), .ZN(n10807) );
  INV_X1 U11137 ( .A(n17445), .ZN(n10592) );
  CLKBUF_X2 U11138 ( .A(n13030), .Z(n19965) );
  NOR2_X2 U11139 ( .A1(n19580), .A2(n11678), .ZN(n17915) );
  OAI211_X1 U11140 ( .C1(n18431), .C2(n14392), .A(n14391), .B(n14390), .ZN(
        n19557) );
  OAI21_X1 U11141 ( .B1(n14388), .B2(n14146), .A(n19703), .ZN(n18293) );
  NAND2_X1 U11142 ( .A1(n14398), .A2(n10117), .ZN(n18973) );
  NOR2_X1 U11143 ( .A1(n9698), .A2(n10143), .ZN(n10142) );
  XNOR2_X1 U11144 ( .A(n13529), .B(n13527), .ZN(n18788) );
  AND2_X1 U11145 ( .A1(n11458), .A2(n10736), .ZN(n9594) );
  OR2_X1 U11146 ( .A1(n11963), .A2(n11947), .ZN(n13830) );
  OR2_X1 U11147 ( .A1(n11637), .A2(n11636), .ZN(n18494) );
  CLKBUF_X1 U11148 ( .A(n10719), .Z(n11464) );
  XNOR2_X1 U11149 ( .A(n13607), .B(n13609), .ZN(n13522) );
  NAND2_X1 U11150 ( .A1(n9807), .A2(n9806), .ZN(n11459) );
  AND2_X1 U11151 ( .A1(n11560), .A2(n11559), .ZN(n19131) );
  INV_X2 U11152 ( .A(n16856), .ZN(n11466) );
  NAND2_X1 U11153 ( .A1(n9921), .A2(n9920), .ZN(n10960) );
  NAND2_X1 U11154 ( .A1(n9809), .A2(n9808), .ZN(n10724) );
  NAND3_X1 U11155 ( .A1(n9907), .A2(n9906), .A3(n10695), .ZN(n9806) );
  NAND2_X2 U11156 ( .A1(n9830), .A2(n9828), .ZN(n16856) );
  BUF_X1 U11157 ( .A(n11967), .Z(n20842) );
  BUF_X1 U11158 ( .A(n11950), .Z(n11966) );
  INV_X2 U11159 ( .A(n10738), .ZN(n9588) );
  NOR2_X1 U11160 ( .A1(n10634), .A2(n10633), .ZN(n10747) );
  AND4_X1 U11161 ( .A1(n13425), .A2(n13430), .A3(n13426), .A4(n9710), .ZN(
        n10217) );
  AND2_X2 U11162 ( .A1(n13337), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10947) );
  INV_X4 U11163 ( .A(n18079), .ZN(n18192) );
  BUF_X2 U11164 ( .A(n11924), .Z(n12879) );
  INV_X4 U11165 ( .A(n18223), .ZN(n10450) );
  INV_X4 U11166 ( .A(n18196), .ZN(n18238) );
  INV_X1 U11167 ( .A(n13513), .ZN(n18200) );
  BUF_X2 U11168 ( .A(n11925), .Z(n12945) );
  AND2_X1 U11169 ( .A1(n11535), .A2(n14394), .ZN(n13511) );
  AND2_X1 U11170 ( .A1(n11535), .A2(n17144), .ZN(n13513) );
  CLKBUF_X2 U11171 ( .A(n11543), .Z(n17278) );
  CLKBUF_X3 U11172 ( .A(n13512), .Z(n18237) );
  BUF_X2 U11173 ( .A(n13672), .Z(n13693) );
  CLKBUF_X2 U11174 ( .A(n9585), .Z(n12118) );
  BUF_X2 U11175 ( .A(n12111), .Z(n9590) );
  AND2_X1 U11176 ( .A1(n17144), .A2(n11532), .ZN(n13512) );
  NOR2_X2 U11177 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13133) );
  AND2_X1 U11178 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14485) );
  AOI21_X1 U11179 ( .B1(n9643), .B2(n19946), .A(n9812), .ZN(n16495) );
  AOI21_X1 U11180 ( .B1(n9643), .B2(n16457), .A(n16232), .ZN(n16233) );
  AND2_X1 U11181 ( .A1(n10091), .A2(n9714), .ZN(n16562) );
  OR2_X1 U11182 ( .A1(n10335), .A2(n16208), .ZN(n10334) );
  NAND2_X1 U11183 ( .A1(n11082), .A2(n11757), .ZN(n16260) );
  NOR2_X1 U11184 ( .A1(n11706), .A2(n9900), .ZN(n9899) );
  XNOR2_X1 U11185 ( .A(n13771), .B(n13770), .ZN(n14740) );
  NAND2_X1 U11186 ( .A1(n11711), .A2(n9793), .ZN(n10336) );
  NAND2_X1 U11187 ( .A1(n9703), .A2(n9913), .ZN(n9834) );
  NAND2_X1 U11188 ( .A1(n11710), .A2(n10343), .ZN(n16280) );
  NAND2_X1 U11189 ( .A1(n11710), .A2(n10345), .ZN(n16354) );
  AND2_X1 U11190 ( .A1(n9932), .A2(n9930), .ZN(n16909) );
  AND2_X2 U11191 ( .A1(n9903), .A2(n9902), .ZN(n11710) );
  NAND2_X1 U11192 ( .A1(n9892), .A2(n10247), .ZN(n16225) );
  NAND2_X1 U11193 ( .A1(n16924), .A2(n9931), .ZN(n9930) );
  AND2_X1 U11194 ( .A1(n15201), .A2(n10323), .ZN(n9872) );
  AOI21_X1 U11195 ( .B1(n10340), .B2(n10339), .A(n9792), .ZN(n9914) );
  NAND2_X1 U11196 ( .A1(n10390), .A2(n11760), .ZN(n16251) );
  AND2_X1 U11197 ( .A1(n9580), .A2(n9937), .ZN(n9931) );
  XNOR2_X1 U11198 ( .A(n14729), .B(n14728), .ZN(n16069) );
  NAND2_X1 U11199 ( .A1(n9955), .A2(n15351), .ZN(n15201) );
  NAND2_X1 U11200 ( .A1(n13359), .A2(n13358), .ZN(n14729) );
  NAND2_X1 U11201 ( .A1(n16385), .A2(n10233), .ZN(n10307) );
  OR2_X1 U11202 ( .A1(n15210), .A2(n12226), .ZN(n15225) );
  AND2_X1 U11203 ( .A1(n10144), .A2(n16377), .ZN(n10389) );
  AND2_X1 U11204 ( .A1(n16386), .A2(n11018), .ZN(n10233) );
  AOI21_X1 U11205 ( .B1(n16417), .B2(n16418), .A(n9813), .ZN(n16385) );
  NAND2_X1 U11206 ( .A1(n10448), .A2(n10445), .ZN(n10446) );
  AND2_X1 U11207 ( .A1(n9965), .A2(n9717), .ZN(n10144) );
  CLKBUF_X1 U11208 ( .A(n11811), .Z(n15685) );
  INV_X1 U11209 ( .A(n14841), .ZN(n12878) );
  XNOR2_X1 U11210 ( .A(n9815), .B(n11472), .ZN(n16417) );
  AND2_X1 U11211 ( .A1(n18541), .A2(n18694), .ZN(n17101) );
  CLKBUF_X1 U11212 ( .A(n15728), .Z(n16125) );
  NAND2_X1 U11213 ( .A1(n10196), .A2(n15942), .ZN(n16432) );
  AND2_X1 U11214 ( .A1(n10311), .A2(n11204), .ZN(n11202) );
  NAND2_X1 U11215 ( .A1(n9816), .A2(n19791), .ZN(n9815) );
  NAND2_X1 U11216 ( .A1(n11196), .A2(n11195), .ZN(n16431) );
  AND2_X1 U11217 ( .A1(n10517), .A2(n10245), .ZN(n10244) );
  AND2_X1 U11218 ( .A1(n13564), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18541) );
  NAND2_X1 U11219 ( .A1(n10050), .A2(n11472), .ZN(n16420) );
  AOI21_X1 U11220 ( .B1(n10443), .B2(n10439), .A(n13562), .ZN(n13564) );
  NAND2_X1 U11221 ( .A1(n9881), .A2(n10342), .ZN(n11204) );
  OAI21_X1 U11222 ( .B1(n17120), .B2(n18575), .A(n18560), .ZN(n13562) );
  AOI21_X1 U11223 ( .B1(n10201), .B2(n12224), .A(n12223), .ZN(n10198) );
  NOR2_X2 U11224 ( .A1(n20116), .A2(n20375), .ZN(n20166) );
  INV_X1 U11225 ( .A(n10342), .ZN(n11198) );
  NOR2_X1 U11226 ( .A1(n18558), .A2(n10274), .ZN(n10439) );
  NOR2_X2 U11227 ( .A1(n20367), .A2(n20465), .ZN(n20515) );
  NAND2_X1 U11228 ( .A1(n14370), .A2(n10434), .ZN(n16024) );
  NAND2_X1 U11229 ( .A1(n10436), .A2(n9689), .ZN(n14370) );
  AND3_X1 U11230 ( .A1(n10002), .A2(n10010), .A3(n10819), .ZN(n10001) );
  AND2_X1 U11231 ( .A1(n10395), .A2(n16501), .ZN(n10394) );
  NAND2_X1 U11232 ( .A1(n9604), .A2(n9678), .ZN(n10146) );
  AND2_X1 U11233 ( .A1(n18570), .A2(n18575), .ZN(n18558) );
  AND2_X1 U11234 ( .A1(n9607), .A2(n9799), .ZN(n10038) );
  OAI21_X2 U11235 ( .B1(n18659), .B2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n18575), .ZN(n18625) );
  NAND2_X1 U11236 ( .A1(n10083), .A2(n10080), .ZN(n18659) );
  AND2_X1 U11237 ( .A1(n13023), .A2(n16177), .ZN(n14236) );
  NOR2_X2 U11238 ( .A1(n20930), .A2(n21232), .ZN(n20912) );
  OR2_X1 U11239 ( .A1(n13766), .A2(n11783), .ZN(n15694) );
  NAND2_X1 U11240 ( .A1(n12173), .A2(n12172), .ZN(n14463) );
  AOI21_X1 U11241 ( .B1(n10261), .B2(n10262), .A(n9880), .ZN(n9879) );
  NAND2_X1 U11242 ( .A1(n12604), .A2(n12603), .ZN(n14426) );
  AOI21_X1 U11243 ( .B1(n16828), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n13987), .ZN(n10012) );
  AND4_X1 U11244 ( .A1(n9820), .A2(n9819), .A3(n9818), .A4(n9817), .ZN(n10894)
         );
  NAND2_X1 U11245 ( .A1(n16799), .A2(n16797), .ZN(n20079) );
  NAND2_X1 U11246 ( .A1(n10263), .A2(n16768), .ZN(n19978) );
  AND3_X1 U11247 ( .A1(n15941), .A2(n16768), .A3(n10817), .ZN(n16828) );
  AND2_X1 U11248 ( .A1(n10816), .A2(n19965), .ZN(n10263) );
  NAND2_X1 U11249 ( .A1(n10818), .A2(n16768), .ZN(n10921) );
  OR2_X1 U11250 ( .A1(n12601), .A2(n12664), .ZN(n12604) );
  NOR2_X1 U11251 ( .A1(n18475), .A2(n18410), .ZN(n18413) );
  CLKBUF_X1 U11252 ( .A(n14667), .Z(n15166) );
  AND3_X1 U11253 ( .A1(n16768), .A2(n16733), .A3(n10808), .ZN(n20032) );
  NOR2_X1 U11254 ( .A1(n18480), .A2(n18417), .ZN(n18420) );
  NAND2_X1 U11255 ( .A1(n18740), .A2(n13549), .ZN(n13550) );
  NAND2_X2 U11256 ( .A1(n15151), .A2(n14209), .ZN(n15182) );
  OAI211_X1 U11257 ( .C1(n18751), .C2(n10069), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n10066), .ZN(n18740) );
  AOI21_X2 U11258 ( .B1(n11252), .B2(n11251), .A(n16888), .ZN(n11494) );
  OR2_X1 U11259 ( .A1(n14103), .A2(n12597), .ZN(n14104) );
  AND2_X1 U11260 ( .A1(n15037), .A2(n10463), .ZN(n14989) );
  NAND2_X1 U11261 ( .A1(n10325), .A2(n12059), .ZN(n10041) );
  NOR2_X1 U11262 ( .A1(n10813), .A2(n10592), .ZN(n10591) );
  NAND3_X1 U11263 ( .A1(n10139), .A2(n10138), .A3(n10267), .ZN(n10590) );
  CLKBUF_X1 U11264 ( .A(n14480), .Z(n21063) );
  NAND2_X1 U11265 ( .A1(n11745), .A2(n11746), .ZN(n11763) );
  NAND2_X2 U11266 ( .A1(n10272), .A2(n9938), .ZN(n18751) );
  AND2_X1 U11267 ( .A1(n11023), .A2(n10113), .ZN(n11745) );
  INV_X1 U11268 ( .A(n18877), .ZN(n18914) );
  NAND2_X1 U11269 ( .A1(n9984), .A2(n12284), .ZN(n14116) );
  NAND2_X1 U11270 ( .A1(n9898), .A2(n10800), .ZN(n10140) );
  NOR2_X1 U11271 ( .A1(n10072), .A2(n10068), .ZN(n10067) );
  NAND2_X1 U11272 ( .A1(n9895), .A2(n10765), .ZN(n10800) );
  NOR2_X1 U11273 ( .A1(n10465), .A2(n10464), .ZN(n10463) );
  NAND2_X1 U11274 ( .A1(n10142), .A2(n9896), .ZN(n10792) );
  NAND2_X1 U11275 ( .A1(n9941), .A2(n10735), .ZN(n10794) );
  AND2_X1 U11276 ( .A1(n10783), .A2(n10784), .ZN(n9896) );
  NAND2_X1 U11277 ( .A1(n10785), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9941) );
  AND3_X1 U11278 ( .A1(n10541), .A2(n10542), .A3(n10540), .ZN(n10795) );
  NOR2_X1 U11279 ( .A1(n10073), .A2(n13547), .ZN(n10072) );
  NAND2_X1 U11280 ( .A1(n9957), .A2(n20006), .ZN(n11033) );
  NAND2_X1 U11281 ( .A1(n10073), .A2(n13547), .ZN(n10071) );
  INV_X1 U11282 ( .A(n10466), .ZN(n10465) );
  NOR3_X1 U11283 ( .A1(n18494), .A2(n18493), .A3(n18492), .ZN(n18508) );
  NOR2_X1 U11284 ( .A1(n14385), .A2(n9600), .ZN(n19539) );
  CLKBUF_X1 U11285 ( .A(n11485), .Z(n16759) );
  XNOR2_X1 U11286 ( .A(n11508), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16910) );
  NOR2_X1 U11287 ( .A1(n10988), .A2(n10989), .ZN(n11001) );
  NAND2_X1 U11288 ( .A1(n11648), .A2(n13627), .ZN(n13626) );
  INV_X1 U11289 ( .A(n14987), .ZN(n10464) );
  INV_X2 U11290 ( .A(n13776), .ZN(n12555) );
  AND2_X2 U11291 ( .A1(n13545), .A2(n13502), .ZN(n18694) );
  NAND2_X2 U11292 ( .A1(n11458), .A2(n10347), .ZN(n13776) );
  NAND2_X1 U11293 ( .A1(n9894), .A2(n16856), .ZN(n16840) );
  CLKBUF_X1 U11294 ( .A(n11241), .Z(n14164) );
  AOI21_X1 U11295 ( .B1(n11086), .B2(n10524), .A(n10522), .ZN(n10989) );
  NOR2_X1 U11296 ( .A1(n10773), .A2(n10774), .ZN(n11445) );
  AND2_X1 U11297 ( .A1(n11948), .A2(n13830), .ZN(n12312) );
  INV_X1 U11298 ( .A(n9841), .ZN(n11458) );
  AND2_X1 U11299 ( .A1(n13536), .A2(n13475), .ZN(n13545) );
  OR2_X1 U11300 ( .A1(n13526), .A2(n13536), .ZN(n13527) );
  INV_X1 U11301 ( .A(n9824), .ZN(n11456) );
  INV_X2 U11302 ( .A(n12605), .ZN(n13787) );
  NAND2_X2 U11303 ( .A1(n11256), .A2(n11271), .ZN(n14727) );
  INV_X2 U11304 ( .A(n11294), .ZN(n14723) );
  CLKBUF_X2 U11305 ( .A(n11266), .Z(n12524) );
  INV_X2 U11306 ( .A(n11232), .ZN(n13987) );
  NAND2_X1 U11307 ( .A1(n9660), .A2(n9857), .ZN(n11289) );
  NAND2_X1 U11308 ( .A1(n11466), .A2(n9588), .ZN(n9824) );
  INV_X1 U11309 ( .A(n10719), .ZN(n19992) );
  NAND2_X1 U11310 ( .A1(n13986), .A2(n10960), .ZN(n13353) );
  INV_X1 U11311 ( .A(n11459), .ZN(n20002) );
  OR2_X1 U11312 ( .A1(n14208), .A2(n11972), .ZN(n15626) );
  AND2_X1 U11313 ( .A1(n16856), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14168) );
  AND2_X1 U11314 ( .A1(n11597), .A2(n11596), .ZN(n19117) );
  AND2_X1 U11315 ( .A1(n11540), .A2(n10300), .ZN(n19108) );
  NAND2_X2 U11316 ( .A1(n10738), .A2(n16856), .ZN(n11253) );
  AND2_X1 U11317 ( .A1(n13474), .A2(n13473), .ZN(n18418) );
  CLKBUF_X1 U11318 ( .A(n10724), .Z(n19997) );
  OR2_X1 U11319 ( .A1(n13501), .A2(n13500), .ZN(n13599) );
  BUF_X2 U11320 ( .A(n10720), .Z(n20015) );
  INV_X1 U11321 ( .A(n10724), .ZN(n11462) );
  OR2_X1 U11322 ( .A1(n10845), .A2(n10844), .ZN(n11272) );
  OR2_X1 U11323 ( .A1(n13458), .A2(n13457), .ZN(n13603) );
  OR2_X1 U11324 ( .A1(n10831), .A2(n10830), .ZN(n11186) );
  INV_X2 U11325 ( .A(n12149), .ZN(n10275) );
  OR2_X2 U11326 ( .A1(n13520), .A2(n13519), .ZN(n14215) );
  NAND3_X1 U11327 ( .A1(n9826), .A2(n9825), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9807) );
  NOR2_X2 U11328 ( .A1(n11613), .A2(n11612), .ZN(n19140) );
  AND2_X2 U11329 ( .A1(n11954), .A2(n13810), .ZN(n14187) );
  INV_X1 U11330 ( .A(n11954), .ZN(n20828) );
  CLKBUF_X1 U11331 ( .A(n11944), .Z(n12012) );
  NAND3_X1 U11332 ( .A1(n11843), .A2(n11842), .A3(n9637), .ZN(n12149) );
  AND2_X1 U11333 ( .A1(n9910), .A2(n9908), .ZN(n10738) );
  AND4_X1 U11334 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11560) );
  NAND3_X2 U11335 ( .A1(n10217), .A2(n13431), .A3(n13427), .ZN(n13609) );
  AND4_X1 U11336 ( .A1(n13462), .A2(n13461), .A3(n13460), .A4(n13459), .ZN(
        n13474) );
  INV_X2 U11337 ( .A(U214), .ZN(n17498) );
  NAND4_X2 U11338 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n13810) );
  NAND4_X1 U11339 ( .A1(n11873), .A2(n11872), .A3(n11871), .A4(n11870), .ZN(
        n11944) );
  NAND2_X1 U11340 ( .A1(n11886), .A2(n11885), .ZN(n11961) );
  NAND4_X2 U11341 ( .A1(n11918), .A2(n11917), .A3(n11916), .A4(n11915), .ZN(
        n11954) );
  AND4_X1 U11342 ( .A1(n11894), .A2(n11893), .A3(n11892), .A4(n11891), .ZN(
        n10610) );
  AND4_X1 U11343 ( .A1(n11884), .A2(n11883), .A3(n11882), .A4(n11881), .ZN(
        n11885) );
  BUF_X2 U11344 ( .A(n11902), .Z(n12931) );
  AND4_X1 U11345 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n11886) );
  AND4_X1 U11346 ( .A1(n11847), .A2(n11846), .A3(n11845), .A4(n11844), .ZN(
        n11853) );
  AND4_X1 U11347 ( .A1(n11851), .A2(n11850), .A3(n11849), .A4(n11848), .ZN(
        n11852) );
  AND4_X1 U11348 ( .A1(n11914), .A2(n11913), .A3(n11912), .A4(n11911), .ZN(
        n11915) );
  INV_X2 U11349 ( .A(n11603), .ZN(n18216) );
  AND4_X1 U11350 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11941) );
  AND4_X1 U11351 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11870) );
  AND4_X1 U11352 ( .A1(n11857), .A2(n11856), .A3(n11855), .A4(n11854), .ZN(
        n11873) );
  AND4_X1 U11353 ( .A1(n11861), .A2(n11860), .A3(n11859), .A4(n11858), .ZN(
        n11872) );
  AND4_X1 U11354 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11871) );
  OR2_X1 U11355 ( .A1(n10626), .A2(n10625), .ZN(n10634) );
  NAND2_X2 U11356 ( .A1(n20597), .A2(n20540), .ZN(n20599) );
  CLKBUF_X1 U11357 ( .A(n13132), .Z(n13335) );
  BUF_X4 U11358 ( .A(n11604), .Z(n18062) );
  INV_X2 U11359 ( .A(n11607), .ZN(n17954) );
  NAND2_X2 U11360 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21396), .ZN(n13891) );
  INV_X2 U11361 ( .A(n11598), .ZN(n18089) );
  NAND2_X2 U11362 ( .A1(n19682), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19678) );
  BUF_X2 U11363 ( .A(n11930), .Z(n12884) );
  BUF_X2 U11364 ( .A(n12712), .Z(n13691) );
  BUF_X2 U11365 ( .A(n12098), .Z(n12005) );
  INV_X2 U11366 ( .A(n18243), .ZN(n10303) );
  INV_X2 U11367 ( .A(n17535), .ZN(n17537) );
  AND2_X2 U11368 ( .A1(n10958), .A2(n16746), .ZN(n13132) );
  NOR2_X1 U11369 ( .A1(n19977), .A2(n20618), .ZN(n20511) );
  AND2_X2 U11370 ( .A1(n16745), .A2(n13133), .ZN(n10833) );
  AND2_X1 U11371 ( .A1(n11536), .A2(n14394), .ZN(n11524) );
  NOR2_X2 U11372 ( .A1(n15963), .A2(n15964), .ZN(n15966) );
  AND2_X2 U11373 ( .A1(n11827), .A2(n11829), .ZN(n12024) );
  AND2_X1 U11374 ( .A1(n14407), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11536) );
  AND2_X1 U11375 ( .A1(n9940), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11535) );
  AND2_X1 U11376 ( .A1(n14453), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11525) );
  AND2_X1 U11377 ( .A1(n11532), .A2(n14394), .ZN(n11543) );
  INV_X1 U11378 ( .A(n17162), .ZN(n14401) );
  AND3_X1 U11379 ( .A1(n17152), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11534) );
  AND2_X1 U11380 ( .A1(n17144), .A2(n11531), .ZN(n13514) );
  NAND2_X1 U11381 ( .A1(n10093), .A2(n16758), .ZN(n10628) );
  AND2_X2 U11382 ( .A1(n11829), .A2(n14485), .ZN(n13672) );
  AND2_X2 U11383 ( .A1(n11820), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11827) );
  AND2_X2 U11384 ( .A1(n10569), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11828) );
  INV_X1 U11385 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10569) );
  INV_X2 U11386 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n12586) );
  CLKBUF_X1 U11387 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15642) );
  INV_X4 U11388 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10093) );
  INV_X1 U11389 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10094) );
  INV_X2 U11390 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10958) );
  AND2_X1 U11391 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9905) );
  AND2_X1 U11392 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11531) );
  AND2_X1 U11393 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14394) );
  INV_X1 U11394 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17152) );
  NOR2_X2 U11395 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11532) );
  NOR2_X2 U11396 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17144) );
  NAND2_X1 U11397 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17162) );
  NOR2_X1 U11398 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11526) );
  INV_X1 U11399 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14453) );
  OAI211_X1 U11400 ( .C1(n13540), .C2(n13539), .A(1'b1), .B(n18748), .ZN(n9939) );
  AOI211_X2 U11402 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17916), .A(n17580), .B(
        n17579), .ZN(n17582) );
  INV_X4 U11403 ( .A(n17954), .ZN(n18174) );
  AND2_X4 U11404 ( .A1(n14394), .A2(n11531), .ZN(n17208) );
  NOR2_X2 U11405 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17669), .ZN(n17653) );
  AOI21_X2 U11406 ( .B1(n15735), .B2(n15968), .A(n16236), .ZN(n15705) );
  NAND2_X1 U11407 ( .A1(n18802), .A2(n13524), .ZN(n13529) );
  NOR2_X2 U11408 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17644), .ZN(n17630) );
  INV_X2 U11409 ( .A(n18202), .ZN(n9593) );
  NOR2_X2 U11410 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17622), .ZN(n17608) );
  NAND2_X2 U11411 ( .A1(n13550), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13637) );
  INV_X4 U11412 ( .A(n18198), .ZN(n17281) );
  NAND2_X1 U11413 ( .A1(n11525), .A2(n11535), .ZN(n18198) );
  NOR2_X2 U11414 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17602), .ZN(n17586) );
  NOR2_X2 U11415 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17834), .ZN(n17811) );
  NOR3_X4 U11416 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17896) );
  INV_X1 U11417 ( .A(n11946), .ZN(n9970) );
  NAND2_X1 U11418 ( .A1(n10960), .A2(n10720), .ZN(n10728) );
  NOR2_X1 U11419 ( .A1(n13810), .A2(n11954), .ZN(n11950) );
  NAND2_X1 U11420 ( .A1(n9912), .A2(n9608), .ZN(n9913) );
  NAND2_X1 U11421 ( .A1(n10253), .A2(n11766), .ZN(n10249) );
  NAND2_X1 U11422 ( .A1(n10252), .A2(n9696), .ZN(n10251) );
  INV_X1 U11423 ( .A(n11267), .ZN(n11294) );
  AND2_X1 U11424 ( .A1(n10736), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10347) );
  AND2_X1 U11425 ( .A1(n11445), .A2(n11464), .ZN(n11449) );
  NOR2_X1 U11426 ( .A1(n17445), .A2(n10804), .ZN(n10817) );
  NAND2_X1 U11427 ( .A1(n9835), .A2(n9919), .ZN(n10720) );
  AND2_X1 U11428 ( .A1(n10817), .A2(n13024), .ZN(n10809) );
  AND2_X1 U11429 ( .A1(n10121), .A2(n9674), .ZN(n9600) );
  NAND2_X1 U11430 ( .A1(n18751), .A2(n13544), .ZN(n13548) );
  NOR2_X1 U11431 ( .A1(n9834), .A2(n13730), .ZN(n13758) );
  NAND2_X1 U11432 ( .A1(n11710), .A2(n16234), .ZN(n16267) );
  BUF_X1 U11433 ( .A(n10797), .Z(n10796) );
  CLKBUF_X2 U11434 ( .A(n12024), .Z(n13667) );
  AND2_X1 U11435 ( .A1(n11969), .A2(n14207), .ZN(n12290) );
  AND3_X1 U11436 ( .A1(n12012), .A2(n14119), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12277) );
  NOR2_X1 U11437 ( .A1(n9642), .A2(n12015), .ZN(n10285) );
  NOR2_X1 U11438 ( .A1(n10533), .A2(n10116), .ZN(n10115) );
  NAND2_X1 U11439 ( .A1(n10534), .A2(n9666), .ZN(n10533) );
  INV_X1 U11440 ( .A(n10535), .ZN(n10534) );
  OR2_X1 U11441 ( .A1(n10536), .A2(n11050), .ZN(n10535) );
  NAND2_X2 U11442 ( .A1(n16745), .A2(n10958), .ZN(n13145) );
  NAND2_X2 U11443 ( .A1(n11107), .A2(n10093), .ZN(n13139) );
  AND2_X1 U11444 ( .A1(n10055), .A2(n10053), .ZN(n10342) );
  NAND2_X1 U11445 ( .A1(n13987), .A2(n10054), .ZN(n10053) );
  INV_X1 U11446 ( .A(n11309), .ZN(n10054) );
  NAND2_X1 U11447 ( .A1(n10729), .A2(n11459), .ZN(n11239) );
  NOR2_X1 U11448 ( .A1(n10293), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11533) );
  INV_X1 U11449 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U11451 ( .A1(n13003), .A2(n10210), .ZN(n10583) );
  INV_X1 U11452 ( .A(n13797), .ZN(n13683) );
  NOR2_X1 U11453 ( .A1(n10474), .A2(n14785), .ZN(n10472) );
  INV_X1 U11454 ( .A(n15210), .ZN(n9972) );
  NOR2_X1 U11455 ( .A1(n9692), .A2(n9609), .ZN(n10292) );
  NOR2_X1 U11456 ( .A1(n14954), .A2(n14955), .ZN(n14939) );
  OR2_X1 U11457 ( .A1(n9866), .A2(n20828), .ZN(n12137) );
  OR2_X1 U11458 ( .A1(n12319), .A2(n12390), .ZN(n14080) );
  INV_X1 U11459 ( .A(n11944), .ZN(n11956) );
  NAND2_X1 U11460 ( .A1(n11253), .A2(n11100), .ZN(n10968) );
  NAND2_X1 U11461 ( .A1(n11024), .A2(n11033), .ZN(n11023) );
  NAND2_X1 U11462 ( .A1(n10726), .A2(n9668), .ZN(n11241) );
  AND2_X1 U11463 ( .A1(n10094), .A2(n10093), .ZN(n10825) );
  NAND2_X1 U11464 ( .A1(n16024), .A2(n13185), .ZN(n10027) );
  AND2_X1 U11465 ( .A1(n16063), .A2(n15875), .ZN(n10557) );
  INV_X1 U11466 ( .A(n14602), .ZN(n10553) );
  AND2_X1 U11467 ( .A1(n12553), .A2(n10565), .ZN(n10564) );
  INV_X1 U11468 ( .A(n12559), .ZN(n10565) );
  OR2_X1 U11469 ( .A1(n10111), .A2(n9917), .ZN(n10105) );
  INV_X1 U11470 ( .A(n13385), .ZN(n9917) );
  NAND2_X1 U11471 ( .A1(n10102), .A2(n13385), .ZN(n10101) );
  NAND2_X1 U11472 ( .A1(n15731), .A2(n9754), .ZN(n11732) );
  NAND2_X1 U11473 ( .A1(n10112), .A2(n11076), .ZN(n11785) );
  INV_X1 U11474 ( .A(n15704), .ZN(n10112) );
  NOR2_X1 U11475 ( .A1(n9620), .A2(n10508), .ZN(n10507) );
  INV_X1 U11476 ( .A(n16123), .ZN(n10508) );
  OR2_X1 U11477 ( .A1(n14641), .A2(n15829), .ZN(n10515) );
  NAND2_X1 U11478 ( .A1(n9837), .A2(n9672), .ZN(n11045) );
  NAND2_X1 U11479 ( .A1(n10307), .A2(n9838), .ZN(n9837) );
  AND2_X1 U11480 ( .A1(n10389), .A2(n11741), .ZN(n9838) );
  OR3_X1 U11481 ( .A1(n14569), .A2(n14572), .A3(n10510), .ZN(n10509) );
  INV_X1 U11482 ( .A(n14579), .ZN(n10510) );
  NAND2_X1 U11483 ( .A1(n13987), .A2(n10588), .ZN(n10587) );
  INV_X1 U11484 ( .A(n11289), .ZN(n10588) );
  AND2_X1 U11485 ( .A1(n11255), .A2(n16814), .ZN(n11271) );
  NAND2_X1 U11486 ( .A1(n10772), .A2(n10771), .ZN(n10773) );
  NAND2_X1 U11487 ( .A1(n10770), .A2(n11462), .ZN(n10772) );
  AND2_X1 U11488 ( .A1(n10723), .A2(n10722), .ZN(n10726) );
  AND2_X1 U11489 ( .A1(n11459), .A2(n11255), .ZN(n10723) );
  AOI21_X1 U11490 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19571), .A(
        n11658), .ZN(n13575) );
  OR2_X1 U11491 ( .A1(n13572), .A2(n11666), .ZN(n13587) );
  INV_X1 U11492 ( .A(n13544), .ZN(n10073) );
  OR2_X1 U11493 ( .A1(n18694), .A2(n13546), .ZN(n13547) );
  NOR2_X1 U11494 ( .A1(n11651), .A2(n14142), .ZN(n10119) );
  INV_X1 U11495 ( .A(n19539), .ZN(n10120) );
  NAND2_X1 U11496 ( .A1(n11954), .A2(n12149), .ZN(n12390) );
  AND4_X1 U11497 ( .A1(n11929), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n11942) );
  AND4_X1 U11498 ( .A1(n11923), .A2(n11922), .A3(n11921), .A4(n11920), .ZN(
        n11943) );
  AND4_X1 U11499 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(
        n11940) );
  INV_X1 U11500 ( .A(n14187), .ZN(n13947) );
  OR2_X1 U11501 ( .A1(n13658), .A2(n14751), .ZN(n14753) );
  NAND2_X1 U11502 ( .A1(n12329), .A2(n12328), .ZN(n14089) );
  OR2_X1 U11503 ( .A1(n12330), .A2(n15614), .ZN(n14465) );
  NAND2_X1 U11504 ( .A1(n12362), .A2(n14671), .ZN(n14200) );
  NOR2_X1 U11505 ( .A1(n13853), .A2(n11958), .ZN(n11951) );
  NAND2_X1 U11506 ( .A1(n9987), .A2(n14115), .ZN(n12455) );
  NOR2_X1 U11507 ( .A1(n10286), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10282) );
  INV_X1 U11508 ( .A(n20640), .ZN(n14115) );
  NOR2_X2 U11509 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21265) );
  NAND2_X1 U11510 ( .A1(n11097), .A2(n11096), .ZN(n11228) );
  OR2_X1 U11511 ( .A1(n11095), .A2(n11094), .ZN(n11097) );
  NAND2_X1 U11512 ( .A1(n11788), .A2(n11780), .ZN(n13766) );
  NAND2_X1 U11513 ( .A1(n19728), .A2(n12545), .ZN(n19804) );
  OR2_X1 U11514 ( .A1(n13266), .A2(n13265), .ZN(n10428) );
  AOI21_X1 U11515 ( .B1(n16844), .B2(n14351), .A(n13350), .ZN(n14362) );
  AND3_X1 U11516 ( .A1(n16848), .A2(n13349), .A3(n15652), .ZN(n13350) );
  OR2_X1 U11517 ( .A1(n12511), .A2(n12514), .ZN(n12516) );
  NOR2_X1 U11518 ( .A1(n16194), .A2(n13768), .ZN(n16192) );
  AND3_X1 U11519 ( .A1(n11159), .A2(n11158), .A3(n11157), .ZN(n15822) );
  XNOR2_X1 U11520 ( .A(n10800), .B(n10799), .ZN(n10801) );
  AND2_X1 U11521 ( .A1(n10563), .A2(n10562), .ZN(n10560) );
  AND2_X1 U11522 ( .A1(n9793), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10549) );
  NAND2_X1 U11523 ( .A1(n16251), .A2(n10250), .ZN(n9892) );
  CLKBUF_X1 U11524 ( .A(n15819), .Z(n15820) );
  NAND2_X1 U11525 ( .A1(n10340), .A2(n10339), .ZN(n9902) );
  NOR2_X1 U11526 ( .A1(n10546), .A2(n9631), .ZN(n9901) );
  NAND2_X1 U11527 ( .A1(n14137), .A2(n14136), .ZN(n10019) );
  AND3_X1 U11528 ( .A1(n11292), .A2(n11291), .A3(n11290), .ZN(n15938) );
  NAND2_X1 U11529 ( .A1(n13015), .A2(n16814), .ZN(n13034) );
  NAND2_X1 U11530 ( .A1(n16775), .A2(n20622), .ZN(n20116) );
  NOR2_X1 U11531 ( .A1(n11649), .A2(n19117), .ZN(n10121) );
  NAND2_X1 U11532 ( .A1(n19709), .A2(n19108), .ZN(n14145) );
  INV_X1 U11533 ( .A(n17638), .ZN(n10371) );
  NAND2_X1 U11534 ( .A1(n19707), .A2(n18432), .ZN(n11678) );
  INV_X1 U11535 ( .A(n18694), .ZN(n18575) );
  NAND2_X1 U11536 ( .A1(n14116), .A2(n12574), .ZN(n20646) );
  NOR2_X1 U11537 ( .A1(n17335), .A2(n20640), .ZN(n12574) );
  INV_X1 U11538 ( .A(n17385), .ZN(n17370) );
  NAND2_X1 U11539 ( .A1(n17385), .A2(n14110), .ZN(n17377) );
  NAND2_X1 U11540 ( .A1(n19866), .A2(n20022), .ZN(n19855) );
  INV_X1 U11541 ( .A(n20622), .ZN(n16813) );
  AOI21_X1 U11542 ( .B1(n16505), .B2(n16443), .A(n16242), .ZN(n9950) );
  NAND2_X1 U11543 ( .A1(n16424), .A2(n14150), .ZN(n16455) );
  NAND2_X1 U11544 ( .A1(n16424), .A2(n13921), .ZN(n16441) );
  INV_X1 U11545 ( .A(n19964), .ZN(n19944) );
  NAND2_X2 U11546 ( .A1(n10796), .A2(n10793), .ZN(n17445) );
  NAND2_X1 U11547 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10240) );
  NAND2_X1 U11548 ( .A1(n20085), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n9817) );
  AND2_X1 U11549 ( .A1(n10518), .A2(n10396), .ZN(n10395) );
  OR2_X1 U11550 ( .A1(n11772), .A2(n16501), .ZN(n10396) );
  INV_X1 U11551 ( .A(n16239), .ZN(n10518) );
  INV_X1 U11552 ( .A(n10263), .ZN(n9880) );
  NAND2_X1 U11553 ( .A1(n19943), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10262) );
  NAND2_X1 U11554 ( .A1(n16768), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10261) );
  AND2_X1 U11555 ( .A1(n16733), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10188) );
  NAND2_X1 U11556 ( .A1(n15941), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10187) );
  NOR2_X1 U11557 ( .A1(n12764), .A2(n10574), .ZN(n10573) );
  INV_X1 U11558 ( .A(n10575), .ZN(n10574) );
  OR3_X1 U11559 ( .A1(n14953), .A2(n14952), .A3(n12763), .ZN(n12764) );
  BUF_X1 U11560 ( .A(n11919), .Z(n13698) );
  INV_X1 U11561 ( .A(n14625), .ZN(n10216) );
  INV_X1 U11562 ( .A(n12296), .ZN(n12279) );
  NAND2_X1 U11563 ( .A1(n12268), .A2(n12267), .ZN(n12280) );
  AOI21_X1 U11564 ( .B1(n15642), .B2(n21132), .A(n12274), .ZN(n12269) );
  NAND2_X1 U11565 ( .A1(n10326), .A2(n12059), .ZN(n10064) );
  INV_X1 U11566 ( .A(n14480), .ZN(n10326) );
  INV_X1 U11567 ( .A(n12193), .ZN(n10498) );
  OR2_X1 U11568 ( .A1(n12058), .A2(n12057), .ZN(n12168) );
  NAND2_X1 U11569 ( .A1(n11971), .A2(n14208), .ZN(n11973) );
  AOI21_X1 U11570 ( .B1(n10285), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9667), 
        .ZN(n10281) );
  NAND2_X1 U11571 ( .A1(n11955), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12046) );
  OR2_X1 U11572 ( .A1(n12012), .A2(n10287), .ZN(n12047) );
  NAND2_X1 U11573 ( .A1(n11978), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11990) );
  AND2_X1 U11574 ( .A1(n16259), .A2(n16377), .ZN(n9964) );
  NOR2_X1 U11575 ( .A1(n9676), .A2(n9836), .ZN(n10008) );
  AND2_X1 U11576 ( .A1(n16819), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9836) );
  AND2_X1 U11577 ( .A1(n11459), .A2(n10728), .ZN(n10205) );
  AND2_X1 U11578 ( .A1(n13361), .A2(n20015), .ZN(n9842) );
  INV_X1 U11579 ( .A(n14369), .ZN(n13263) );
  NAND2_X1 U11580 ( .A1(n9966), .A2(n9697), .ZN(n9856) );
  INV_X1 U11581 ( .A(n10664), .ZN(n9906) );
  INV_X1 U11582 ( .A(n10663), .ZN(n9907) );
  INV_X1 U11583 ( .A(n10676), .ZN(n9825) );
  NAND2_X1 U11584 ( .A1(n10701), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9920) );
  NAND2_X1 U11585 ( .A1(n10707), .A2(n10706), .ZN(n9921) );
  AOI21_X1 U11586 ( .B1(n19131), .B2(n11641), .A(n13582), .ZN(n11648) );
  NAND2_X1 U11587 ( .A1(n14215), .A2(n13609), .ZN(n13608) );
  NOR2_X1 U11588 ( .A1(n19140), .A2(n14145), .ZN(n11650) );
  AOI21_X1 U11589 ( .B1(n18174), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n10129), .ZN(n10128) );
  INV_X1 U11590 ( .A(n11581), .ZN(n10126) );
  OR2_X1 U11591 ( .A1(n10663), .A2(n10664), .ZN(n10752) );
  OR2_X1 U11592 ( .A1(n10675), .A2(n10676), .ZN(n10744) );
  NAND2_X1 U11593 ( .A1(n9588), .A2(n10739), .ZN(n10770) );
  NOR2_X1 U11594 ( .A1(n11253), .A2(n16902), .ZN(n10764) );
  AND4_X1 U11595 ( .A1(n11890), .A2(n11889), .A3(n11888), .A4(n11887), .ZN(
        n11895) );
  NAND2_X1 U11596 ( .A1(n11967), .A2(n11956), .ZN(n13651) );
  NOR2_X1 U11597 ( .A1(n14789), .A2(n14800), .ZN(n10211) );
  AND2_X1 U11598 ( .A1(n14813), .A2(n10571), .ZN(n10570) );
  NOR2_X1 U11599 ( .A1(n10577), .A2(n14914), .ZN(n10208) );
  NAND2_X1 U11600 ( .A1(n10578), .A2(n14863), .ZN(n10577) );
  INV_X1 U11601 ( .A(n10579), .ZN(n10578) );
  OR2_X1 U11602 ( .A1(n14947), .A2(n14948), .ZN(n14983) );
  INV_X1 U11603 ( .A(n14634), .ZN(n12628) );
  NOR2_X2 U11604 ( .A1(n13652), .A2(n12586), .ZN(n12756) );
  NAND2_X1 U11605 ( .A1(n12586), .A2(n21397), .ZN(n13797) );
  NAND2_X1 U11606 ( .A1(n15351), .A2(n10290), .ZN(n10289) );
  INV_X1 U11607 ( .A(n10291), .ZN(n10290) );
  INV_X1 U11608 ( .A(n14815), .ZN(n10475) );
  NAND2_X1 U11609 ( .A1(n12220), .A2(n10493), .ZN(n10201) );
  INV_X1 U11610 ( .A(n15300), .ZN(n12220) );
  NOR2_X1 U11611 ( .A1(n10482), .A2(n10481), .ZN(n10480) );
  INV_X1 U11612 ( .A(n14897), .ZN(n10482) );
  INV_X1 U11613 ( .A(n14915), .ZN(n10481) );
  NOR2_X1 U11614 ( .A1(n10467), .A2(n15007), .ZN(n10466) );
  INV_X1 U11615 ( .A(n9640), .ZN(n10467) );
  OR2_X1 U11616 ( .A1(n12104), .A2(n12103), .ZN(n12208) );
  INV_X1 U11617 ( .A(n9788), .ZN(n10461) );
  NAND2_X1 U11618 ( .A1(n14187), .A2(n14671), .ZN(n12440) );
  INV_X1 U11619 ( .A(n14446), .ZN(n10462) );
  OR2_X1 U11620 ( .A1(n14201), .A2(n13947), .ZN(n10456) );
  AND4_X1 U11621 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n10612) );
  AND3_X1 U11622 ( .A1(n11837), .A2(n11836), .A3(n11835), .ZN(n11842) );
  AOI22_X1 U11623 ( .A1(n11931), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13672), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11843) );
  INV_X1 U11624 ( .A(n20889), .ZN(n20866) );
  AND4_X1 U11625 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11918) );
  AND4_X1 U11626 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n11916) );
  AND4_X1 U11627 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11917) );
  NAND2_X1 U11628 ( .A1(n10527), .A2(n10526), .ZN(n11086) );
  NAND2_X1 U11629 ( .A1(n11253), .A2(n11222), .ZN(n10526) );
  NAND2_X1 U11630 ( .A1(n10959), .A2(n11225), .ZN(n10527) );
  NOR2_X1 U11631 ( .A1(n13382), .A2(n12536), .ZN(n13389) );
  AND2_X1 U11632 ( .A1(n10115), .A2(n11072), .ZN(n10114) );
  OR2_X1 U11633 ( .A1(n11041), .A2(n10535), .ZN(n11063) );
  NAND2_X1 U11634 ( .A1(n10537), .A2(n11049), .ZN(n10536) );
  INV_X1 U11635 ( .A(n11042), .ZN(n10537) );
  AND2_X1 U11636 ( .A1(n10530), .A2(n16066), .ZN(n10529) );
  INV_X1 U11637 ( .A(n12465), .ZN(n10399) );
  NOR2_X1 U11638 ( .A1(n15714), .A2(n15729), .ZN(n10505) );
  AND2_X1 U11639 ( .A1(n13056), .A2(n9756), .ZN(n10435) );
  AND2_X1 U11640 ( .A1(n13019), .A2(n13986), .ZN(n14369) );
  NOR2_X1 U11641 ( .A1(n13987), .A2(n16902), .ZN(n13019) );
  INV_X1 U11642 ( .A(n15789), .ZN(n10552) );
  INV_X1 U11643 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12492) );
  NAND2_X1 U11644 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10412) );
  INV_X1 U11645 ( .A(n14457), .ZN(n10555) );
  INV_X1 U11646 ( .A(n10959), .ZN(n11282) );
  INV_X1 U11647 ( .A(n10250), .ZN(n10246) );
  NAND2_X1 U11648 ( .A1(n13380), .A2(n16223), .ZN(n10100) );
  INV_X1 U11649 ( .A(n15700), .ZN(n10566) );
  NOR2_X1 U11650 ( .A1(n10394), .A2(n10254), .ZN(n10250) );
  NOR2_X1 U11651 ( .A1(n10181), .A2(n9684), .ZN(n10179) );
  NAND2_X1 U11652 ( .A1(n10356), .A2(n10357), .ZN(n10045) );
  AND2_X1 U11653 ( .A1(n9712), .A2(n10358), .ZN(n10357) );
  NAND2_X1 U11654 ( .A1(n10363), .A2(n10359), .ZN(n10358) );
  INV_X1 U11655 ( .A(n14608), .ZN(n10556) );
  AND2_X1 U11656 ( .A1(n10342), .A2(n11076), .ZN(n10206) );
  INV_X1 U11657 ( .A(n14418), .ZN(n11130) );
  INV_X1 U11658 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11472) );
  OR2_X1 U11659 ( .A1(n10888), .A2(n10887), .ZN(n11295) );
  NAND2_X1 U11660 ( .A1(n10268), .A2(n10799), .ZN(n10267) );
  NAND2_X1 U11661 ( .A1(n10088), .A2(n10140), .ZN(n10139) );
  INV_X1 U11662 ( .A(n10960), .ZN(n11254) );
  NAND2_X1 U11663 ( .A1(n10589), .A2(n10792), .ZN(n10797) );
  AND2_X1 U11664 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13029) );
  NOR2_X1 U11665 ( .A1(n9860), .A2(n9858), .ZN(n9857) );
  NAND2_X1 U11666 ( .A1(n11239), .A2(n10730), .ZN(n11452) );
  OAI21_X1 U11667 ( .B1(n16733), .B2(n14157), .A(n13018), .ZN(n13039) );
  OR2_X1 U11668 ( .A1(n13263), .A2(n20001), .ZN(n13021) );
  AND3_X1 U11669 ( .A1(n11247), .A2(n11246), .A3(n11245), .ZN(n14360) );
  AND2_X1 U11670 ( .A1(n13024), .A2(n10808), .ZN(n10810) );
  NOR2_X1 U11671 ( .A1(n17445), .A2(n10391), .ZN(n10808) );
  INV_X1 U11672 ( .A(n10804), .ZN(n10391) );
  NAND2_X1 U11673 ( .A1(n9811), .A2(n9810), .ZN(n10719) );
  INV_X1 U11674 ( .A(n10645), .ZN(n9877) );
  NAND2_X1 U11675 ( .A1(n10750), .A2(n10543), .ZN(n9809) );
  NAND2_X1 U11676 ( .A1(n10742), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9808) );
  NAND2_X2 U11677 ( .A1(n9805), .A2(n9804), .ZN(n11255) );
  INV_X1 U11678 ( .A(n10991), .ZN(n11103) );
  OR3_X1 U11679 ( .A1(n13576), .A2(n14399), .A3(n19135), .ZN(n14142) );
  INV_X1 U11680 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18195) );
  AND2_X1 U11681 ( .A1(n9650), .A2(n10378), .ZN(n10377) );
  INV_X1 U11682 ( .A(n18678), .ZN(n10378) );
  INV_X1 U11683 ( .A(n17866), .ZN(n10368) );
  NOR2_X1 U11684 ( .A1(n16955), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10445) );
  NAND2_X1 U11685 ( .A1(n11643), .A2(n10122), .ZN(n11649) );
  NOR2_X1 U11686 ( .A1(n14143), .A2(n10123), .ZN(n10122) );
  INV_X1 U11687 ( .A(n19140), .ZN(n10124) );
  INV_X1 U11688 ( .A(n19131), .ZN(n13576) );
  NOR2_X1 U11689 ( .A1(n18736), .A2(n13618), .ZN(n13619) );
  INV_X1 U11690 ( .A(n13622), .ZN(n9996) );
  NAND2_X1 U11691 ( .A1(n18757), .A2(n13614), .ZN(n13616) );
  AND2_X1 U11692 ( .A1(n13605), .A2(n13597), .ZN(n13604) );
  NAND2_X1 U11693 ( .A1(n13609), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10221) );
  NOR2_X1 U11694 ( .A1(n17162), .A2(n14407), .ZN(n14656) );
  INV_X1 U11695 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18107) );
  NAND2_X1 U11696 ( .A1(n11541), .A2(n10302), .ZN(n10301) );
  NAND2_X1 U11697 ( .A1(n11603), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10302) );
  OAI22_X1 U11698 ( .A1(n10450), .A2(n17207), .B1(n18113), .B2(n10303), .ZN(
        n11539) );
  INV_X1 U11699 ( .A(n13511), .ZN(n18079) );
  AND3_X1 U11700 ( .A1(n11618), .A2(n10454), .A3(n10161), .ZN(n11620) );
  AOI21_X1 U11701 ( .B1(n18089), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n10162), .ZN(n10161) );
  NOR2_X1 U11702 ( .A1(n13626), .A2(n14400), .ZN(n14389) );
  NOR2_X1 U11703 ( .A1(n11253), .A2(n19992), .ZN(n10736) );
  NOR2_X1 U11704 ( .A1(n12291), .A2(n12292), .ZN(n13950) );
  INV_X1 U11705 ( .A(n15071), .ZN(n20726) );
  AND2_X1 U11706 ( .A1(n12439), .A2(n12438), .ZN(n14785) );
  NAND2_X1 U11708 ( .A1(n20828), .A2(n13810), .ZN(n14273) );
  NAND2_X1 U11709 ( .A1(n12998), .A2(n9796), .ZN(n13791) );
  NAND2_X1 U11710 ( .A1(n13712), .A2(n13713), .ZN(n13790) );
  NAND2_X1 U11711 ( .A1(n12998), .A2(n9626), .ZN(n13686) );
  CLKBUF_X1 U11712 ( .A(n14775), .Z(n14776) );
  NOR3_X1 U11713 ( .A1(n12747), .A2(n12746), .A3(n12729), .ZN(n9886) );
  INV_X1 U11714 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12729) );
  INV_X1 U11715 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U11716 ( .A1(n12724), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12747) );
  NOR2_X1 U11717 ( .A1(n12615), .A2(n20701), .ZN(n12622) );
  NAND2_X1 U11718 ( .A1(n12228), .A2(n15201), .ZN(n15191) );
  NOR2_X1 U11719 ( .A1(n15456), .A2(n12339), .ZN(n15443) );
  NAND2_X1 U11720 ( .A1(n14942), .A2(n9749), .ZN(n14867) );
  INV_X1 U11721 ( .A(n14869), .ZN(n10477) );
  NAND2_X1 U11722 ( .A1(n14942), .A2(n10478), .ZN(n14892) );
  NAND2_X1 U11723 ( .A1(n14942), .A2(n10480), .ZN(n14899) );
  AND2_X1 U11724 ( .A1(n14942), .A2(n14915), .ZN(n14917) );
  AND2_X1 U11725 ( .A1(n9727), .A2(n10331), .ZN(n10330) );
  AND2_X1 U11726 ( .A1(n12411), .A2(n12410), .ZN(n14940) );
  XNOR2_X1 U11727 ( .A(n12183), .B(n12182), .ZN(n14526) );
  OR2_X1 U11728 ( .A1(n17401), .A2(n14469), .ZN(n17404) );
  OR2_X1 U11729 ( .A1(n12455), .A2(n17323), .ZN(n15488) );
  OR2_X1 U11730 ( .A1(n12455), .A2(n12327), .ZN(n15464) );
  INV_X1 U11731 ( .A(n15562), .ZN(n14469) );
  AND2_X1 U11732 ( .A1(n12585), .A2(n12584), .ZN(n14507) );
  NOR2_X1 U11733 ( .A1(n11999), .A2(n10317), .ZN(n10316) );
  INV_X1 U11734 ( .A(n11995), .ZN(n10317) );
  OAI21_X1 U11735 ( .B1(n14478), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12032), 
        .ZN(n10284) );
  NAND2_X1 U11736 ( .A1(n10491), .A2(n20951), .ZN(n21039) );
  NOR2_X1 U11737 ( .A1(n14508), .A2(n20866), .ZN(n21184) );
  OR2_X1 U11738 ( .A1(n14078), .A2(n21188), .ZN(n21270) );
  INV_X1 U11739 ( .A(n20855), .ZN(n20959) );
  NOR2_X1 U11740 ( .A1(n12601), .A2(n20951), .ZN(n21264) );
  INV_X1 U11741 ( .A(n14207), .ZN(n20851) );
  CLKBUF_X1 U11742 ( .A(n12450), .Z(n12451) );
  NOR2_X1 U11743 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15656) );
  XNOR2_X1 U11744 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U11745 ( .A1(n11777), .A2(n10528), .ZN(n11788) );
  NOR2_X1 U11746 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n10528) );
  NAND2_X1 U11747 ( .A1(n11777), .A2(n16006), .ZN(n11782) );
  OAI21_X1 U11748 ( .B1(n15705), .B2(n19815), .A(n16229), .ZN(n15706) );
  OAI21_X1 U11749 ( .B1(n15734), .B2(n19815), .A(n16246), .ZN(n15735) );
  NAND2_X1 U11750 ( .A1(n10516), .A2(n11761), .ZN(n11767) );
  NAND2_X1 U11751 ( .A1(n11763), .A2(n11780), .ZN(n10516) );
  OAI21_X1 U11752 ( .B1(n12502), .B2(n15763), .A(n16266), .ZN(n17309) );
  INV_X1 U11753 ( .A(n16847), .ZN(n13910) );
  OR2_X1 U11754 ( .A1(n10423), .A2(n10031), .ZN(n10426) );
  INV_X1 U11755 ( .A(n10428), .ZN(n10031) );
  NAND2_X1 U11756 ( .A1(n10023), .A2(n10022), .ZN(n16008) );
  NOR2_X1 U11757 ( .A1(n10026), .A2(n10429), .ZN(n10025) );
  NOR2_X1 U11758 ( .A1(n16016), .A2(n16015), .ZN(n16014) );
  NOR2_X1 U11759 ( .A1(n14562), .A2(n10503), .ZN(n10502) );
  NAND2_X1 U11760 ( .A1(n10504), .A2(n14575), .ZN(n10503) );
  INV_X1 U11761 ( .A(n14565), .ZN(n10504) );
  AND2_X1 U11762 ( .A1(n14237), .A2(n13038), .ZN(n10436) );
  NOR2_X1 U11763 ( .A1(n14165), .A2(n14164), .ZN(n14359) );
  INV_X1 U11764 ( .A(n13928), .ZN(n14048) );
  AND3_X1 U11765 ( .A1(n11714), .A2(n11713), .A3(n11712), .ZN(n15749) );
  AND2_X1 U11766 ( .A1(n11710), .A2(n10344), .ZN(n16297) );
  NAND2_X1 U11767 ( .A1(n11710), .A2(n10355), .ZN(n16569) );
  NOR2_X1 U11768 ( .A1(n16487), .A2(n11739), .ZN(n16463) );
  NAND2_X1 U11769 ( .A1(n13720), .A2(n13721), .ZN(n16465) );
  NOR2_X1 U11770 ( .A1(n16215), .A2(n9700), .ZN(n10193) );
  NOR2_X1 U11771 ( .A1(n16192), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10195) );
  OR2_X1 U11772 ( .A1(n16498), .A2(n11738), .ZN(n16487) );
  INV_X1 U11773 ( .A(n11711), .ZN(n16235) );
  AND3_X1 U11774 ( .A1(n11723), .A2(n11722), .A3(n11721), .ZN(n15719) );
  NOR2_X1 U11775 ( .A1(n10181), .A2(n10182), .ZN(n16528) );
  AND2_X1 U11776 ( .A1(n11794), .A2(n11793), .ZN(n15746) );
  NOR2_X1 U11777 ( .A1(n11441), .A2(n9620), .ZN(n15745) );
  CLKBUF_X1 U11778 ( .A(n9633), .Z(n15748) );
  OR2_X1 U11779 ( .A1(n10515), .A2(n10514), .ZN(n10513) );
  NAND2_X1 U11780 ( .A1(n15784), .A2(n15799), .ZN(n10514) );
  AND2_X1 U11781 ( .A1(n10344), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10343) );
  NAND2_X1 U11782 ( .A1(n9864), .A2(n11481), .ZN(n9863) );
  INV_X1 U11783 ( .A(n11480), .ZN(n9864) );
  NAND2_X1 U11784 ( .A1(n10314), .A2(n10360), .ZN(n10313) );
  INV_X1 U11785 ( .A(n16569), .ZN(n16310) );
  NAND2_X1 U11786 ( .A1(n11045), .A2(n9603), .ZN(n10365) );
  AND3_X1 U11787 ( .A1(n11153), .A2(n11152), .A3(n11151), .ZN(n14613) );
  NAND2_X1 U11788 ( .A1(n16665), .A2(n16295), .ZN(n16616) );
  NOR2_X1 U11789 ( .A1(n10182), .A2(n10180), .ZN(n16536) );
  INV_X1 U11790 ( .A(n11474), .ZN(n10180) );
  NAND2_X1 U11791 ( .A1(n10264), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10547) );
  INV_X1 U11792 ( .A(n16398), .ZN(n10264) );
  NAND2_X1 U11793 ( .A1(n16398), .A2(n11205), .ZN(n10548) );
  NAND2_X1 U11794 ( .A1(n10060), .A2(n9652), .ZN(n10340) );
  NAND2_X1 U11795 ( .A1(n10547), .A2(n10061), .ZN(n10060) );
  INV_X1 U11796 ( .A(n10548), .ZN(n10061) );
  INV_X1 U11797 ( .A(n9912), .ZN(n10338) );
  NAND2_X1 U11798 ( .A1(n9893), .A2(n11206), .ZN(n16398) );
  NAND2_X1 U11799 ( .A1(n11204), .A2(n13768), .ZN(n9893) );
  NAND2_X1 U11800 ( .A1(n9975), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10046) );
  AND2_X1 U11801 ( .A1(n11449), .A2(n11448), .ZN(n14351) );
  NAND2_X1 U11802 ( .A1(n13028), .A2(n10016), .ZN(n10018) );
  NOR2_X1 U11803 ( .A1(n13029), .A2(n10017), .ZN(n10016) );
  INV_X1 U11804 ( .A(n13027), .ZN(n10017) );
  NAND2_X1 U11805 ( .A1(n10021), .A2(n13029), .ZN(n10420) );
  NAND2_X1 U11806 ( .A1(n13028), .A2(n13027), .ZN(n10021) );
  AND2_X1 U11807 ( .A1(n11293), .A2(n11288), .ZN(n10500) );
  AND2_X1 U11808 ( .A1(n13033), .A2(n13032), .ZN(n14136) );
  XNOR2_X1 U11809 ( .A(n14704), .B(n13036), .ZN(n14137) );
  NAND2_X1 U11810 ( .A1(n11231), .A2(n11230), .ZN(n16844) );
  CLKBUF_X1 U11811 ( .A(n11107), .Z(n16757) );
  NAND2_X1 U11812 ( .A1(n10726), .A2(n10725), .ZN(n17298) );
  AND2_X1 U11813 ( .A1(n19992), .A2(n11462), .ZN(n10725) );
  AND2_X1 U11814 ( .A1(n14159), .A2(n14158), .ZN(n20119) );
  NAND2_X1 U11815 ( .A1(n16884), .A2(n14169), .ZN(n14158) );
  NAND2_X1 U11816 ( .A1(n16883), .A2(n16902), .ZN(n14159) );
  AND2_X1 U11817 ( .A1(n10810), .A2(n16733), .ZN(n20150) );
  NAND2_X1 U11818 ( .A1(n16775), .A2(n16813), .ZN(n20195) );
  NAND2_X1 U11819 ( .A1(n16799), .A2(n16798), .ZN(n20267) );
  INV_X1 U11820 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20335) );
  NAND2_X1 U11821 ( .A1(n20610), .A2(n16813), .ZN(n20367) );
  INV_X1 U11822 ( .A(n16733), .ZN(n10092) );
  NAND2_X1 U11823 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n14169) );
  INV_X1 U11824 ( .A(n19541), .ZN(n14140) );
  OR2_X1 U11825 ( .A1(n19541), .A2(n13588), .ZN(n19542) );
  AOI21_X1 U11826 ( .B1(n16908), .B2(n14141), .A(n19588), .ZN(n10134) );
  NAND2_X1 U11827 ( .A1(n11523), .A2(n11522), .ZN(n17573) );
  NAND2_X1 U11828 ( .A1(n17882), .A2(n11502), .ZN(n10380) );
  NAND2_X1 U11829 ( .A1(n18555), .A2(n11502), .ZN(n10381) );
  NAND2_X1 U11830 ( .A1(n11520), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U11831 ( .A1(n18289), .A2(n10156), .ZN(n18264) );
  AND2_X1 U11832 ( .A1(n18268), .A2(n9790), .ZN(n10156) );
  NOR2_X1 U11833 ( .A1(n18294), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n10297) );
  AND2_X1 U11834 ( .A1(n19140), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n10305) );
  AOI211_X1 U11835 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n11609), .B(n11608), .ZN(n11610) );
  INV_X1 U11836 ( .A(n10158), .ZN(n17180) );
  OAI21_X1 U11837 ( .B1(n9600), .B2(n14387), .A(n14386), .ZN(n18431) );
  XNOR2_X1 U11838 ( .A(n13616), .B(n10222), .ZN(n18747) );
  INV_X1 U11839 ( .A(n13615), .ZN(n10222) );
  NAND2_X1 U11840 ( .A1(n18747), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18746) );
  NAND2_X1 U11841 ( .A1(n17101), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16956) );
  NAND2_X1 U11842 ( .A1(n18540), .A2(n18575), .ZN(n10079) );
  AND2_X1 U11843 ( .A1(n18557), .A2(n17120), .ZN(n16959) );
  INV_X1 U11844 ( .A(n17157), .ZN(n17153) );
  NOR2_X1 U11845 ( .A1(n13628), .A2(n11649), .ZN(n13625) );
  INV_X1 U11846 ( .A(n19542), .ZN(n16907) );
  NAND2_X1 U11847 ( .A1(n17157), .A2(n10118), .ZN(n10117) );
  INV_X1 U11848 ( .A(n14399), .ZN(n10118) );
  INV_X1 U11849 ( .A(n10438), .ZN(n10437) );
  INV_X1 U11850 ( .A(n13637), .ZN(n18713) );
  NAND2_X1 U11851 ( .A1(n10438), .A2(n17047), .ZN(n18691) );
  NAND2_X1 U11852 ( .A1(n10071), .A2(n10074), .ZN(n10069) );
  NOR2_X1 U11853 ( .A1(n18775), .A2(n9994), .ZN(n18758) );
  AOI21_X1 U11854 ( .B1(n18776), .B2(n18777), .A(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U11855 ( .A1(n14389), .A2(n19721), .ZN(n19546) );
  NAND2_X1 U11856 ( .A1(n17157), .A2(n13625), .ZN(n19538) );
  INV_X2 U11857 ( .A(n18494), .ZN(n19709) );
  NAND2_X1 U11858 ( .A1(n18957), .A2(n19547), .ZN(n10133) );
  NAND2_X1 U11859 ( .A1(n9976), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10763) );
  OAI21_X1 U11860 ( .B1(n10737), .B2(n10760), .A(n10759), .ZN(n10761) );
  OR2_X1 U11861 ( .A1(n13943), .A2(n20640), .ZN(n13915) );
  NAND2_X1 U11862 ( .A1(n14278), .A2(n13915), .ZN(n21402) );
  INV_X1 U11863 ( .A(n20744), .ZN(n20723) );
  NAND2_X1 U11864 ( .A1(n14681), .A2(n14680), .ZN(n20750) );
  XNOR2_X1 U11865 ( .A(n14676), .B(n14675), .ZN(n15392) );
  INV_X1 U11866 ( .A(n14673), .ZN(n14676) );
  OR2_X1 U11867 ( .A1(n14764), .A2(n15114), .ZN(n13662) );
  OR3_X1 U11868 ( .A1(n14116), .A2(n20640), .A3(n14089), .ZN(n13656) );
  NAND2_X1 U11869 ( .A1(n15113), .A2(n20851), .ZN(n15114) );
  NAND2_X1 U11870 ( .A1(n14750), .A2(n14749), .ZN(n15189) );
  OR2_X1 U11871 ( .A1(n13685), .A2(n14748), .ZN(n14749) );
  AND2_X1 U11872 ( .A1(n13007), .A2(n13006), .ZN(n14763) );
  NAND2_X1 U11873 ( .A1(n13005), .A2(n13004), .ZN(n13006) );
  INV_X1 U11874 ( .A(n20811), .ZN(n17381) );
  NAND2_X1 U11875 ( .A1(n20646), .A2(n13010), .ZN(n17385) );
  NAND2_X1 U11876 ( .A1(n13008), .A2(n21265), .ZN(n20811) );
  AOI21_X1 U11877 ( .B1(n15392), .B2(n17424), .A(n15391), .ZN(n9980) );
  NOR3_X1 U11878 ( .A1(n15399), .A2(n15390), .A3(n9983), .ZN(n15388) );
  AND2_X1 U11879 ( .A1(n17404), .A2(n10324), .ZN(n9983) );
  NOR2_X1 U11880 ( .A1(n9982), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9981) );
  INV_X1 U11881 ( .A(n15389), .ZN(n9982) );
  XNOR2_X1 U11882 ( .A(n10487), .B(n15390), .ZN(n15387) );
  OAI21_X1 U11883 ( .B1(n13714), .B2(n10489), .A(n10202), .ZN(n10487) );
  NAND2_X1 U11884 ( .A1(n15351), .A2(n10324), .ZN(n10489) );
  NAND2_X1 U11885 ( .A1(n15191), .A2(n10203), .ZN(n10202) );
  XNOR2_X1 U11886 ( .A(n10278), .B(n10277), .ZN(n15394) );
  INV_X1 U11887 ( .A(n15187), .ZN(n10277) );
  MUX2_X1 U11888 ( .A(n12571), .B(n12570), .S(n12217), .Z(n12573) );
  NOR2_X1 U11889 ( .A1(n15439), .A2(n15424), .ZN(n15423) );
  INV_X1 U11890 ( .A(n17390), .ZN(n17424) );
  OR2_X1 U11891 ( .A1(n12455), .A2(n12314), .ZN(n17397) );
  CLKBUF_X1 U11892 ( .A(n14478), .Z(n21065) );
  INV_X1 U11894 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21397) );
  INV_X1 U11895 ( .A(n21265), .ZN(n21302) );
  NAND2_X1 U11896 ( .A1(n20917), .A2(n10491), .ZN(n10490) );
  INV_X1 U11897 ( .A(n12581), .ZN(n10492) );
  AOI21_X1 U11898 ( .B1(n14506), .B2(n14505), .A(n20855), .ZN(n20810) );
  INV_X1 U11899 ( .A(n21070), .ZN(n21090) );
  INV_X1 U11900 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21357) );
  NAND2_X1 U11901 ( .A1(n12532), .A2(n13910), .ZN(n13889) );
  NOR2_X1 U11902 ( .A1(n16840), .A2(n16888), .ZN(n12532) );
  NOR2_X1 U11903 ( .A1(n19815), .A2(n19838), .ZN(n15952) );
  OAI21_X1 U11904 ( .B1(n13742), .B2(n13743), .A(n19820), .ZN(n13746) );
  OAI21_X1 U11905 ( .B1(n13753), .B2(n19833), .A(n13752), .ZN(n13754) );
  INV_X1 U11906 ( .A(n19830), .ZN(n19773) );
  INV_X1 U11907 ( .A(n19776), .ZN(n19836) );
  INV_X1 U11908 ( .A(n19838), .ZN(n19820) );
  NAND2_X1 U11909 ( .A1(n19815), .A2(n19820), .ZN(n17314) );
  INV_X1 U11910 ( .A(n17314), .ZN(n19842) );
  AND2_X1 U11911 ( .A1(n19804), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19841) );
  AND2_X1 U11912 ( .A1(n19836), .A2(n10592), .ZN(n10392) );
  OR2_X1 U11913 ( .A1(n12561), .A2(n13773), .ZN(n16184) );
  NAND2_X1 U11914 ( .A1(n14370), .A2(n16175), .ZN(n16179) );
  AND2_X1 U11915 ( .A1(n13984), .A2(n16899), .ZN(n19866) );
  NAND2_X1 U11916 ( .A1(n14729), .A2(n13360), .ZN(n13753) );
  OR2_X1 U11917 ( .A1(n13359), .A2(n13358), .ZN(n13360) );
  OR2_X1 U11918 ( .A1(n13359), .A2(n12531), .ZN(n16080) );
  AOI211_X1 U11919 ( .C1(n12516), .C2(n12457), .A(n10404), .B(n10405), .ZN(
        n10403) );
  AND2_X1 U11920 ( .A1(n10406), .A2(n12457), .ZN(n10405) );
  NOR2_X1 U11921 ( .A1(n12516), .A2(n10407), .ZN(n10404) );
  OR2_X1 U11922 ( .A1(n13758), .A2(n10099), .ZN(n10098) );
  AOI21_X1 U11923 ( .B1(n16225), .B2(n10191), .A(n10598), .ZN(n11791) );
  NOR2_X1 U11924 ( .A1(n16215), .A2(n10194), .ZN(n10191) );
  AND2_X1 U11925 ( .A1(n10059), .A2(n13722), .ZN(n16208) );
  NAND2_X1 U11926 ( .A1(n10336), .A2(n16457), .ZN(n10335) );
  OAI21_X1 U11927 ( .B1(n16297), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16280), .ZN(n16551) );
  NAND2_X1 U11928 ( .A1(n16571), .A2(n16443), .ZN(n10258) );
  INV_X1 U11929 ( .A(n16298), .ZN(n10257) );
  NAND2_X1 U11930 ( .A1(n16564), .A2(n16577), .ZN(n10260) );
  NAND2_X1 U11931 ( .A1(n16310), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16564) );
  NOR2_X1 U11932 ( .A1(n16297), .A2(n16446), .ZN(n10259) );
  XNOR2_X1 U11933 ( .A(n16304), .B(n16303), .ZN(n16583) );
  NAND2_X1 U11934 ( .A1(n10362), .A2(n16306), .ZN(n16304) );
  NAND2_X1 U11935 ( .A1(n10365), .A2(n10363), .ZN(n10362) );
  INV_X1 U11936 ( .A(n16441), .ZN(n16452) );
  NAND2_X1 U11937 ( .A1(n13911), .A2(n11175), .ZN(n16424) );
  INV_X1 U11938 ( .A(n16455), .ZN(n16443) );
  NAND2_X1 U11939 ( .A1(n10110), .A2(n10107), .ZN(n13771) );
  NOR2_X1 U11940 ( .A1(n14720), .A2(n13768), .ZN(n13769) );
  OR2_X1 U11941 ( .A1(n10563), .A2(n10562), .ZN(n10558) );
  XNOR2_X1 U11942 ( .A(n13759), .B(n14733), .ZN(n14743) );
  XNOR2_X1 U11943 ( .A(n13395), .B(n13394), .ZN(n13733) );
  XNOR2_X1 U11944 ( .A(n13758), .B(n10539), .ZN(n10538) );
  INV_X1 U11945 ( .A(n10098), .ZN(n16190) );
  XNOR2_X1 U11946 ( .A(n13719), .B(n9658), .ZN(n10097) );
  NAND2_X1 U11947 ( .A1(n10106), .A2(n13385), .ZN(n13719) );
  NAND2_X1 U11948 ( .A1(n10111), .A2(n10244), .ZN(n10106) );
  NOR2_X1 U11949 ( .A1(n16208), .A2(n19963), .ZN(n10058) );
  AND2_X1 U11950 ( .A1(n15666), .A2(n11734), .ZN(n16210) );
  AND2_X1 U11951 ( .A1(n9989), .A2(n10059), .ZN(n16484) );
  NAND2_X1 U11952 ( .A1(n16225), .A2(n16223), .ZN(n16213) );
  XNOR2_X1 U11953 ( .A(n16241), .B(n16240), .ZN(n16506) );
  NAND2_X1 U11954 ( .A1(n10160), .A2(n11772), .ZN(n16241) );
  OAI21_X1 U11955 ( .B1(n16251), .B2(n11766), .A(n10253), .ZN(n10160) );
  AND2_X1 U11956 ( .A1(n16235), .A2(n9945), .ZN(n9944) );
  NAND2_X1 U11957 ( .A1(n9947), .A2(n16501), .ZN(n9945) );
  NAND2_X1 U11958 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U11959 ( .A1(n16267), .A2(n16501), .ZN(n9943) );
  OAI211_X1 U11960 ( .C1(n16267), .C2(n9803), .A(n10015), .B(n10014), .ZN(
        n16523) );
  NAND2_X1 U11961 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n10013), .ZN(
        n10015) );
  NAND2_X1 U11962 ( .A1(n10035), .A2(n16267), .ZN(n16547) );
  NAND2_X1 U11963 ( .A1(n10051), .A2(n16541), .ZN(n10035) );
  OAI21_X1 U11964 ( .B1(n11710), .B2(n10352), .A(n10349), .ZN(n9904) );
  AOI21_X1 U11965 ( .B1(n10351), .B2(n10350), .A(n9802), .ZN(n10349) );
  INV_X1 U11966 ( .A(n10353), .ZN(n10350) );
  AND2_X1 U11967 ( .A1(n10169), .A2(n16572), .ZN(n10168) );
  OR2_X1 U11968 ( .A1(n16573), .A2(n19949), .ZN(n10169) );
  INV_X1 U11969 ( .A(n16583), .ZN(n9844) );
  OAI21_X1 U11970 ( .B1(n16310), .B2(n10087), .A(n10085), .ZN(n16579) );
  INV_X1 U11971 ( .A(n10270), .ZN(n10087) );
  AOI21_X1 U11972 ( .B1(n10270), .B2(n16585), .A(n10086), .ZN(n10085) );
  NAND2_X1 U11973 ( .A1(n19963), .A2(n19956), .ZN(n10270) );
  NAND2_X1 U11974 ( .A1(n10348), .A2(n10351), .ZN(n16584) );
  NAND2_X1 U11975 ( .A1(n11710), .A2(n10353), .ZN(n10348) );
  NAND2_X1 U11976 ( .A1(n16581), .A2(n16582), .ZN(n9846) );
  CLKBUF_X3 U11977 ( .A(n10805), .Z(n16733) );
  NAND2_X1 U11978 ( .A1(n11494), .A2(n11487), .ZN(n19964) );
  INV_X1 U11979 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20627) );
  OR2_X1 U11980 ( .A1(n14704), .A2(n13989), .ZN(n20622) );
  INV_X1 U11981 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20619) );
  INV_X1 U11982 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20618) );
  NAND2_X1 U11983 ( .A1(n20619), .A2(n16814), .ZN(n20614) );
  NAND2_X1 U11984 ( .A1(n14366), .A2(n14365), .ZN(n17302) );
  AND2_X1 U11985 ( .A1(n20270), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20290) );
  INV_X1 U11986 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19582) );
  INV_X1 U11987 ( .A(n17569), .ZN(n10386) );
  NOR2_X1 U11988 ( .A1(n10385), .A2(n10384), .ZN(n10383) );
  NOR2_X1 U11989 ( .A1(n17918), .A2(n17572), .ZN(n10384) );
  INV_X1 U11990 ( .A(n17571), .ZN(n10385) );
  NAND2_X1 U11991 ( .A1(n17570), .A2(n17944), .ZN(n10387) );
  NOR2_X1 U11992 ( .A1(n17583), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n11684) );
  NAND2_X1 U11993 ( .A1(n17997), .A2(n9598), .ZN(n10153) );
  AND2_X1 U11994 ( .A1(n10153), .A2(n18270), .ZN(n17983) );
  AND2_X1 U11995 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n18000), .ZN(n17997) );
  NOR2_X1 U11996 ( .A1(n18277), .A2(n18069), .ZN(n18053) );
  NAND2_X1 U11997 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18088), .ZN(n18069) );
  NOR3_X1 U11998 ( .A1(n18120), .A2(n18123), .A3(n17710), .ZN(n18071) );
  NOR2_X1 U11999 ( .A1(n18157), .A2(n18153), .ZN(n18135) );
  AND2_X1 U12000 ( .A1(n10158), .A2(n10157), .ZN(n18289) );
  NOR2_X1 U12001 ( .A1(n17179), .A2(n19588), .ZN(n10157) );
  NAND2_X1 U12002 ( .A1(n18330), .A2(n19140), .ZN(n18324) );
  INV_X1 U12003 ( .A(n19140), .ZN(n18277) );
  NAND2_X1 U12004 ( .A1(n9936), .A2(n9933), .ZN(n9932) );
  AND2_X1 U12005 ( .A1(n13567), .A2(n9934), .ZN(n9933) );
  NAND2_X1 U12006 ( .A1(n9935), .A2(n13642), .ZN(n9934) );
  NAND2_X1 U12007 ( .A1(n17026), .A2(n10136), .ZN(n18588) );
  NOR2_X1 U12008 ( .A1(n18668), .A2(n10137), .ZN(n10136) );
  INV_X1 U12009 ( .A(n17096), .ZN(n10137) );
  OR2_X1 U12010 ( .A1(n18817), .A2(n18411), .ZN(n18641) );
  AND2_X1 U12011 ( .A1(n10440), .A2(n10443), .ZN(n16972) );
  NOR2_X1 U12012 ( .A1(n18558), .A2(n10441), .ZN(n10440) );
  AND2_X1 U12013 ( .A1(n9998), .A2(n18992), .ZN(n18901) );
  NAND2_X1 U12014 ( .A1(n18893), .A2(n9665), .ZN(n9998) );
  AND2_X1 U12015 ( .A1(n19086), .A2(n17098), .ZN(n18997) );
  AND2_X1 U12016 ( .A1(n18957), .A2(n19062), .ZN(n19057) );
  INV_X1 U12017 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19571) );
  INV_X1 U12018 ( .A(n17178), .ZN(n17174) );
  INV_X1 U12019 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U12020 ( .A1(n12264), .A2(n14275), .ZN(n12238) );
  OR2_X1 U12021 ( .A1(n12011), .A2(n12010), .ZN(n12013) );
  INV_X1 U12022 ( .A(n13776), .ZN(n10776) );
  NOR2_X1 U12023 ( .A1(n9959), .A2(n9701), .ZN(n9958) );
  NAND2_X1 U12024 ( .A1(n10915), .A2(n10916), .ZN(n9959) );
  NAND2_X1 U12025 ( .A1(n16828), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10239) );
  NOR2_X1 U12026 ( .A1(n10057), .A2(n10924), .ZN(n10056) );
  OR2_X1 U12027 ( .A1(n10925), .A2(n10926), .ZN(n10057) );
  NAND2_X1 U12028 ( .A1(n20150), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n9820) );
  NAND2_X1 U12029 ( .A1(n20032), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n9819) );
  NAND2_X1 U12030 ( .A1(n20197), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n9818) );
  AND2_X1 U12031 ( .A1(n10242), .A2(n10241), .ZN(n10893) );
  NAND2_X1 U12032 ( .A1(n16828), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10241) );
  NAND2_X1 U12033 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10242) );
  AND2_X1 U12034 ( .A1(n10737), .A2(n14168), .ZN(n10237) );
  AOI21_X1 U12035 ( .B1(n11232), .B2(n10171), .A(n9596), .ZN(n10170) );
  NOR2_X1 U12036 ( .A1(n14168), .A2(n11222), .ZN(n10171) );
  NAND2_X1 U12037 ( .A1(n9918), .A2(n10728), .ZN(n11235) );
  NOR2_X1 U12038 ( .A1(n18196), .A2(n10130), .ZN(n10129) );
  OR2_X1 U12039 ( .A1(n10645), .A2(n10646), .ZN(n10741) );
  AND2_X1 U12040 ( .A1(n12242), .A2(n12232), .ZN(n12256) );
  NOR2_X1 U12041 ( .A1(n15035), .A2(n10576), .ZN(n10575) );
  INV_X1 U12042 ( .A(n14650), .ZN(n10576) );
  INV_X1 U12043 ( .A(n12196), .ZN(n10333) );
  AND2_X1 U12044 ( .A1(n12175), .A2(n10328), .ZN(n10327) );
  NAND2_X1 U12045 ( .A1(n12059), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10328) );
  OR2_X1 U12046 ( .A1(n12081), .A2(n12080), .ZN(n12188) );
  AND2_X1 U12047 ( .A1(n12290), .A2(n12289), .ZN(n12315) );
  OR2_X1 U12048 ( .A1(n12030), .A2(n12029), .ZN(n12132) );
  NAND2_X1 U12049 ( .A1(n9832), .A2(n11976), .ZN(n11979) );
  NAND2_X1 U12050 ( .A1(n11975), .A2(n9622), .ZN(n9832) );
  AOI22_X1 U12051 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11931), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11832) );
  AOI21_X1 U12052 ( .B1(n11874), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n11875), .ZN(n11880) );
  AND2_X1 U12053 ( .A1(n10617), .A2(n10621), .ZN(n9911) );
  INV_X1 U12054 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10621) );
  AND3_X1 U12055 ( .A1(n9848), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n9847), .ZN(n9909) );
  NAND2_X1 U12056 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n9848) );
  NAND2_X1 U12057 ( .A1(n13327), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9847) );
  INV_X1 U12058 ( .A(n10978), .ZN(n9957) );
  CLKBUF_X1 U12059 ( .A(n10622), .Z(n13322) );
  CLKBUF_X1 U12060 ( .A(n13145), .Z(n13306) );
  OR2_X1 U12061 ( .A1(n10858), .A2(n10857), .ZN(n10959) );
  INV_X1 U12062 ( .A(n10395), .ZN(n10252) );
  INV_X1 U12063 ( .A(n16323), .ZN(n10359) );
  NAND2_X1 U12064 ( .A1(n11198), .A2(n10938), .ZN(n10311) );
  INV_X1 U12065 ( .A(n10938), .ZN(n9881) );
  AND2_X1 U12066 ( .A1(n10587), .A2(n11295), .ZN(n10586) );
  NAND2_X1 U12067 ( .A1(n13987), .A2(n9954), .ZN(n10145) );
  INV_X1 U12068 ( .A(n10800), .ZN(n10268) );
  AOI22_X1 U12069 ( .A1(n16819), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__3__SCAN_IN), .B2(n10890), .ZN(n10868) );
  NOR2_X1 U12070 ( .A1(n9879), .A2(n9878), .ZN(n9977) );
  OAI22_X1 U12071 ( .A1(n10860), .A2(n20344), .B1(n10921), .B2(n13221), .ZN(
        n9878) );
  NAND2_X1 U12072 ( .A1(n19983), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10011) );
  NAND2_X1 U12073 ( .A1(n20085), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10006) );
  NAND2_X1 U12074 ( .A1(n10889), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10004) );
  NAND2_X1 U12075 ( .A1(n10188), .A2(n10809), .ZN(n10184) );
  NAND2_X1 U12076 ( .A1(n20114), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10010) );
  NAND2_X1 U12077 ( .A1(n16803), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10005) );
  NAND2_X1 U12078 ( .A1(n20226), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10009) );
  NAND2_X1 U12079 ( .A1(n20032), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10007) );
  NOR2_X1 U12080 ( .A1(n9588), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11267) );
  INV_X1 U12081 ( .A(n10876), .ZN(n9860) );
  AOI21_X1 U12082 ( .B1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B2(n10881), .A(n9695), .ZN(n9859) );
  INV_X1 U12083 ( .A(n10820), .ZN(n13138) );
  AND2_X1 U12084 ( .A1(n10719), .A2(n10724), .ZN(n11242) );
  NAND2_X1 U12085 ( .A1(n10805), .A2(n17445), .ZN(n10815) );
  NAND2_X1 U12086 ( .A1(n10263), .A2(n19943), .ZN(n10919) );
  INV_X1 U12087 ( .A(n10646), .ZN(n9876) );
  AOI22_X1 U12088 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13339), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10654) );
  NAND2_X1 U12089 ( .A1(n10696), .A2(n10695), .ZN(n9919) );
  INV_X1 U12090 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10695) );
  AND2_X1 U12091 ( .A1(n20627), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10991) );
  XNOR2_X1 U12092 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10969) );
  INV_X1 U12093 ( .A(n14215), .ZN(n9993) );
  NOR2_X1 U12094 ( .A1(n18196), .A2(n10163), .ZN(n10162) );
  INV_X1 U12095 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10163) );
  NOR2_X1 U12096 ( .A1(n14824), .A2(n10572), .ZN(n10571) );
  NOR2_X1 U12097 ( .A1(n12831), .A2(n12830), .ZN(n9891) );
  INV_X1 U12098 ( .A(n13709), .ZN(n13679) );
  NAND2_X1 U12099 ( .A1(n10580), .A2(n14901), .ZN(n10579) );
  INV_X1 U12100 ( .A(n14880), .ZN(n10580) );
  NOR2_X1 U12101 ( .A1(n12781), .A2(n12780), .ZN(n9889) );
  INV_X1 U12102 ( .A(n9775), .ZN(n10213) );
  INV_X1 U12103 ( .A(n11953), .ZN(n12309) );
  AND2_X1 U12104 ( .A1(n12311), .A2(n12315), .ZN(n12310) );
  OAI21_X1 U12105 ( .B1(n12280), .B2(n12278), .A(n12277), .ZN(n9986) );
  NOR2_X1 U12106 ( .A1(n9601), .A2(n9755), .ZN(n9985) );
  NAND2_X1 U12107 ( .A1(n10040), .A2(n10041), .ZN(n12176) );
  NOR2_X1 U12108 ( .A1(n12567), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10291) );
  NOR2_X1 U12109 ( .A1(n14894), .A2(n10479), .ZN(n10478) );
  INV_X1 U12110 ( .A(n10480), .ZN(n10479) );
  AND4_X1 U12111 ( .A1(n12109), .A2(n15309), .A3(n15298), .A4(n15302), .ZN(
        n10331) );
  INV_X1 U12112 ( .A(n15036), .ZN(n10468) );
  INV_X1 U12113 ( .A(n17371), .ZN(n10497) );
  NOR2_X1 U12114 ( .A1(n13651), .A2(n11896), .ZN(n11897) );
  AND2_X1 U12115 ( .A1(n12321), .A2(n12320), .ZN(n12328) );
  NAND2_X1 U12116 ( .A1(n9868), .A2(n12156), .ZN(n12164) );
  NAND2_X1 U12117 ( .A1(n14190), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9868) );
  OR2_X1 U12118 ( .A1(n12124), .A2(n12123), .ZN(n12150) );
  INV_X1 U12119 ( .A(n12015), .ZN(n10286) );
  AND2_X1 U12120 ( .A1(n12000), .A2(n10281), .ZN(n9923) );
  NAND2_X1 U12121 ( .A1(n10281), .A2(n9969), .ZN(n9925) );
  INV_X1 U12122 ( .A(n10285), .ZN(n9969) );
  NAND2_X1 U12123 ( .A1(n11994), .A2(n11993), .ZN(n11995) );
  INV_X1 U12124 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21064) );
  INV_X1 U12125 ( .A(n11960), .ZN(n11967) );
  AOI21_X1 U12126 ( .B1(n21399), .B2(n14504), .A(n17358), .ZN(n20814) );
  INV_X1 U12127 ( .A(n10728), .ZN(n10722) );
  AND2_X1 U12128 ( .A1(n19772), .A2(n10531), .ZN(n10530) );
  NAND2_X1 U12129 ( .A1(n11021), .A2(n19772), .ZN(n11031) );
  OAI21_X1 U12130 ( .B1(n13390), .B2(n9954), .A(n9953), .ZN(n9952) );
  NAND2_X1 U12131 ( .A1(n13390), .A2(n14376), .ZN(n9953) );
  INV_X1 U12132 ( .A(n10525), .ZN(n10524) );
  NAND2_X1 U12133 ( .A1(n10962), .A2(n10961), .ZN(n10523) );
  CLKBUF_X1 U12134 ( .A(n13139), .Z(n13331) );
  NAND2_X1 U12135 ( .A1(n13332), .A2(n9791), .ZN(n13324) );
  CLKBUF_X1 U12136 ( .A(n10690), .Z(n13279) );
  INV_X1 U12137 ( .A(n15802), .ZN(n11163) );
  INV_X1 U12138 ( .A(n15986), .ZN(n10424) );
  INV_X1 U12139 ( .A(n15990), .ZN(n10427) );
  INV_X1 U12140 ( .A(n10029), .ZN(n10026) );
  NAND2_X1 U12141 ( .A1(n10431), .A2(n10430), .ZN(n10429) );
  INV_X1 U12142 ( .A(n16015), .ZN(n10430) );
  NOR2_X1 U12143 ( .A1(n13185), .A2(n16009), .ZN(n10028) );
  NAND2_X1 U12144 ( .A1(n13185), .A2(n16022), .ZN(n10029) );
  NAND2_X1 U12145 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10408) );
  NOR2_X1 U12146 ( .A1(n12506), .A2(n10402), .ZN(n12512) );
  AND2_X1 U12147 ( .A1(n12498), .A2(n9762), .ZN(n12503) );
  NOR2_X1 U12148 ( .A1(n11177), .A2(n10401), .ZN(n10400) );
  INV_X1 U12149 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10401) );
  NOR2_X1 U12150 ( .A1(n16403), .A2(n10417), .ZN(n10416) );
  INV_X1 U12151 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10417) );
  INV_X1 U12152 ( .A(n12473), .ZN(n10415) );
  AND2_X1 U12153 ( .A1(n9669), .A2(n14590), .ZN(n10554) );
  INV_X1 U12154 ( .A(n9898), .ZN(n10799) );
  NOR2_X1 U12155 ( .A1(n16217), .A2(n16227), .ZN(n10550) );
  OR2_X1 U12156 ( .A1(n11766), .A2(n16253), .ZN(n10584) );
  INV_X1 U12157 ( .A(n15719), .ZN(n10567) );
  NAND2_X1 U12158 ( .A1(n11474), .A2(n9686), .ZN(n10181) );
  AND2_X1 U12159 ( .A1(n11752), .A2(n9708), .ZN(n9963) );
  NOR2_X1 U12160 ( .A1(n16555), .A2(n10346), .ZN(n10344) );
  NOR2_X1 U12161 ( .A1(n16303), .A2(n10361), .ZN(n10360) );
  INV_X1 U12162 ( .A(n16306), .ZN(n10361) );
  AND2_X1 U12163 ( .A1(n16296), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10355) );
  NAND2_X1 U12164 ( .A1(n11015), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16386) );
  NAND2_X1 U12165 ( .A1(n10310), .A2(n10976), .ZN(n11015) );
  OR2_X1 U12166 ( .A1(n10937), .A2(n10936), .ZN(n11309) );
  INV_X1 U12167 ( .A(n11202), .ZN(n10255) );
  NAND2_X1 U12168 ( .A1(n11182), .A2(n13768), .ZN(n9816) );
  AND2_X1 U12169 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10432) );
  AND2_X1 U12170 ( .A1(n9841), .A2(n10236), .ZN(n10781) );
  INV_X1 U12171 ( .A(n10782), .ZN(n10143) );
  NAND2_X1 U12172 ( .A1(n9588), .A2(n9681), .ZN(n11281) );
  OR2_X1 U12173 ( .A1(n13263), .A2(n13164), .ZN(n13036) );
  CLKBUF_X1 U12174 ( .A(n13138), .Z(n16755) );
  NAND2_X1 U12175 ( .A1(n9854), .A2(n9853), .ZN(n11231) );
  NAND2_X1 U12176 ( .A1(n16902), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9853) );
  NAND2_X1 U12177 ( .A1(n9855), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U12178 ( .A1(n9856), .A2(n11228), .ZN(n9855) );
  NAND2_X1 U12179 ( .A1(n15941), .A2(n10810), .ZN(n20371) );
  INV_X1 U12180 ( .A(n10675), .ZN(n9826) );
  NAND2_X1 U12181 ( .A1(n16787), .A2(n20467), .ZN(n16789) );
  INV_X1 U12182 ( .A(n16786), .ZN(n16787) );
  AND2_X1 U12183 ( .A1(n9823), .A2(n9821), .ZN(n16855) );
  INV_X1 U12184 ( .A(n17297), .ZN(n9821) );
  AOI21_X1 U12185 ( .B1(n18223), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(n9694), .ZN(n10453) );
  NOR2_X1 U12186 ( .A1(n18672), .A2(n18769), .ZN(n16914) );
  OR2_X1 U12187 ( .A1(n10441), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10274) );
  INV_X1 U12188 ( .A(n10071), .ZN(n10068) );
  NAND2_X1 U12189 ( .A1(n9661), .A2(n10125), .ZN(n11638) );
  NOR2_X1 U12190 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  NAND2_X1 U12191 ( .A1(n10733), .A2(n11241), .ZN(n9976) );
  INV_X1 U12192 ( .A(n10770), .ZN(n10758) );
  NAND2_X1 U12193 ( .A1(n12357), .A2(n12356), .ZN(n12360) );
  INV_X1 U12194 ( .A(n20738), .ZN(n20718) );
  OR3_X1 U12195 ( .A1(n21402), .A2(n17416), .A3(n13798), .ZN(n15059) );
  INV_X1 U12196 ( .A(n14427), .ZN(n13786) );
  MUX2_X1 U12197 ( .A(n14686), .B(n13711), .S(n13797), .Z(n13713) );
  NAND2_X1 U12198 ( .A1(n10582), .A2(n14748), .ZN(n10581) );
  INV_X1 U12199 ( .A(n10583), .ZN(n10582) );
  AND2_X1 U12200 ( .A1(n10211), .A2(n10210), .ZN(n10209) );
  NOR2_X1 U12201 ( .A1(n12959), .A2(n15217), .ZN(n12960) );
  NAND2_X1 U12202 ( .A1(n12960), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12997) );
  NAND2_X1 U12203 ( .A1(n9890), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12907) );
  OR2_X1 U12204 ( .A1(n12907), .A2(n12906), .ZN(n12959) );
  CLKBUF_X1 U12205 ( .A(n14797), .Z(n14798) );
  NAND2_X1 U12206 ( .A1(n9891), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12862) );
  AND2_X1 U12207 ( .A1(n10208), .A2(n14854), .ZN(n10207) );
  NAND2_X1 U12208 ( .A1(n9888), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12831) );
  INV_X1 U12209 ( .A(n9891), .ZN(n12860) );
  NAND2_X1 U12210 ( .A1(n9889), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12813) );
  INV_X1 U12211 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14903) );
  CLKBUF_X1 U12212 ( .A(n14911), .Z(n14912) );
  NAND2_X1 U12213 ( .A1(n12779), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12781) );
  INV_X1 U12214 ( .A(n12778), .ZN(n12779) );
  INV_X1 U12215 ( .A(n9889), .ZN(n12812) );
  NAND2_X1 U12216 ( .A1(n9886), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12778) );
  CLKBUF_X1 U12217 ( .A(n14927), .Z(n14928) );
  NOR2_X1 U12218 ( .A1(n12680), .A2(n12679), .ZN(n12724) );
  NAND2_X1 U12219 ( .A1(n9885), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12680) );
  INV_X1 U12220 ( .A(n12665), .ZN(n9885) );
  NAND2_X1 U12221 ( .A1(n12659), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12665) );
  INV_X1 U12222 ( .A(n10215), .ZN(n10214) );
  NOR2_X1 U12223 ( .A1(n10215), .A2(n9775), .ZN(n10212) );
  AND2_X1 U12224 ( .A1(n12630), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12659) );
  AND2_X1 U12225 ( .A1(n12622), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12630) );
  OAI21_X1 U12226 ( .B1(n12620), .B2(n12664), .A(n12619), .ZN(n14553) );
  AND2_X1 U12227 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12576) );
  AND2_X1 U12228 ( .A1(n12576), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12611) );
  AND2_X1 U12229 ( .A1(n12229), .A2(n10319), .ZN(n10318) );
  NAND2_X1 U12230 ( .A1(n10320), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10319) );
  AND2_X1 U12231 ( .A1(n10488), .A2(n15395), .ZN(n10203) );
  NOR2_X1 U12232 ( .A1(n15351), .A2(n10324), .ZN(n10488) );
  NAND2_X1 U12233 ( .A1(n10062), .A2(n12228), .ZN(n10322) );
  INV_X1 U12234 ( .A(n10288), .ZN(n10062) );
  OAI21_X1 U12235 ( .B1(n12227), .B2(n12217), .A(n9759), .ZN(n10288) );
  NAND2_X1 U12236 ( .A1(n9872), .A2(n12228), .ZN(n13714) );
  INV_X1 U12237 ( .A(n15404), .ZN(n10323) );
  NAND2_X1 U12238 ( .A1(n12217), .A2(n15425), .ZN(n9929) );
  NOR2_X1 U12239 ( .A1(n10471), .A2(n10476), .ZN(n10470) );
  INV_X1 U12240 ( .A(n14774), .ZN(n10476) );
  INV_X1 U12241 ( .A(n10472), .ZN(n10471) );
  NAND2_X1 U12242 ( .A1(n14835), .A2(n10473), .ZN(n14808) );
  NAND2_X1 U12243 ( .A1(n14835), .A2(n14815), .ZN(n14814) );
  INV_X1 U12244 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15469) );
  NOR2_X2 U12245 ( .A1(n14867), .A2(n14856), .ZN(n14855) );
  AND2_X1 U12246 ( .A1(n12423), .A2(n12422), .ZN(n14869) );
  NOR2_X1 U12247 ( .A1(n9974), .A2(n9962), .ZN(n9961) );
  INV_X1 U12248 ( .A(n15310), .ZN(n9962) );
  NAND2_X1 U12249 ( .A1(n10329), .A2(n10200), .ZN(n15239) );
  INV_X1 U12250 ( .A(n10201), .ZN(n10200) );
  AND2_X1 U12251 ( .A1(n12417), .A2(n12416), .ZN(n14915) );
  INV_X1 U12252 ( .A(n14940), .ZN(n12412) );
  NAND2_X1 U12253 ( .A1(n9973), .A2(n15310), .ZN(n15300) );
  AND2_X1 U12254 ( .A1(n15330), .A2(n12108), .ZN(n15320) );
  AND2_X1 U12255 ( .A1(n15037), .A2(n10466), .ZN(n15009) );
  AND3_X1 U12256 ( .A1(n12105), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n12243), 
        .ZN(n12106) );
  NAND2_X1 U12257 ( .A1(n10065), .A2(n12211), .ZN(n17364) );
  NAND2_X1 U12258 ( .A1(n12634), .A2(n12243), .ZN(n10065) );
  NOR2_X1 U12259 ( .A1(n10461), .A2(n9785), .ZN(n10460) );
  NOR2_X1 U12260 ( .A1(n14447), .A2(n10461), .ZN(n10458) );
  NAND2_X1 U12261 ( .A1(n10459), .A2(n10462), .ZN(n14527) );
  NAND2_X1 U12262 ( .A1(n12581), .A2(n12243), .ZN(n12173) );
  AND2_X1 U12263 ( .A1(n17401), .A2(n14191), .ZN(n15565) );
  OR2_X1 U12264 ( .A1(n12601), .A2(n12275), .ZN(n12163) );
  XNOR2_X1 U12265 ( .A(n12164), .B(n14262), .ZN(n14252) );
  AND3_X1 U12266 ( .A1(n11985), .A2(n11984), .A3(n12325), .ZN(n11988) );
  INV_X1 U12267 ( .A(n11830), .ZN(n14487) );
  CLKBUF_X1 U12268 ( .A(n13830), .Z(n13831) );
  OR3_X1 U12269 ( .A1(n13974), .A2(n13973), .A3(n13972), .ZN(n17324) );
  OR2_X1 U12270 ( .A1(n12581), .A2(n10491), .ZN(n20930) );
  OR2_X1 U12271 ( .A1(n21039), .A2(n21262), .ZN(n21014) );
  NAND2_X1 U12272 ( .A1(n12581), .A2(n12601), .ZN(n21161) );
  NOR2_X1 U12273 ( .A1(n20819), .A2(n12586), .ZN(n21190) );
  INV_X1 U12274 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21234) );
  NAND2_X1 U12275 ( .A1(n20867), .A2(n20866), .ZN(n21232) );
  INV_X1 U12276 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21432) );
  NAND2_X1 U12277 ( .A1(n20889), .A2(n14508), .ZN(n21262) );
  NAND2_X1 U12278 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21296) );
  NAND2_X1 U12279 ( .A1(n14508), .A2(n20866), .ZN(n21155) );
  AOI21_X1 U12280 ( .B1(n21234), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20959), 
        .ZN(n21306) );
  NOR2_X2 U12281 ( .A1(n20811), .A2(n13852), .ZN(n20849) );
  NOR2_X2 U12282 ( .A1(n20812), .A2(n20811), .ZN(n20850) );
  INV_X1 U12283 ( .A(n14116), .ZN(n14096) );
  NAND2_X1 U12284 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n14504) );
  INV_X1 U12285 ( .A(n21404), .ZN(n17352) );
  NAND2_X1 U12286 ( .A1(n9824), .A2(n11253), .ZN(n11455) );
  AND2_X1 U12287 ( .A1(n11092), .A2(n11091), .ZN(n11226) );
  OAI21_X1 U12288 ( .B1(n20633), .B2(n11493), .A(n11112), .ZN(n11250) );
  CLKBUF_X1 U12289 ( .A(n15678), .Z(n15688) );
  AND2_X1 U12290 ( .A1(n10114), .A2(n16035), .ZN(n10113) );
  NOR2_X1 U12291 ( .A1(n12496), .A2(n16285), .ZN(n12498) );
  AND2_X1 U12292 ( .A1(n11068), .A2(n11071), .ZN(n15794) );
  NAND2_X1 U12293 ( .A1(n10411), .A2(n10410), .ZN(n10409) );
  INV_X1 U12294 ( .A(n10412), .ZN(n10411) );
  NOR2_X1 U12295 ( .A1(n10413), .A2(n12492), .ZN(n10410) );
  INV_X1 U12296 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12494) );
  OR2_X1 U12297 ( .A1(n9632), .A2(n12494), .ZN(n12496) );
  OR2_X1 U12298 ( .A1(n11041), .A2(n10536), .ZN(n11051) );
  INV_X1 U12299 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12480) );
  NAND2_X1 U12300 ( .A1(n12459), .A2(n12458), .ZN(n12502) );
  NAND2_X1 U12301 ( .A1(n14733), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12458) );
  NOR2_X1 U12302 ( .A1(n12464), .A2(n10398), .ZN(n10397) );
  NAND2_X1 U12303 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U12304 ( .A1(n11012), .A2(n9651), .ZN(n10981) );
  INV_X1 U12305 ( .A(n9952), .ZN(n11013) );
  INV_X1 U12306 ( .A(n19804), .ZN(n19827) );
  AND3_X1 U12307 ( .A1(n12558), .A2(n12557), .A3(n12556), .ZN(n12559) );
  AND3_X1 U12308 ( .A1(n11166), .A2(n11165), .A3(n11164), .ZN(n15789) );
  AND2_X1 U12309 ( .A1(n12527), .A2(n12526), .ZN(n15660) );
  NOR2_X2 U12310 ( .A1(n15661), .A2(n15660), .ZN(n15663) );
  AND2_X1 U12311 ( .A1(n11804), .A2(n11803), .ZN(n15714) );
  NAND2_X1 U12312 ( .A1(n11802), .A2(n11801), .ZN(n15713) );
  AND2_X1 U12313 ( .A1(n10435), .A2(n16025), .ZN(n10434) );
  AND2_X1 U12314 ( .A1(n14370), .A2(n10435), .ZN(n16031) );
  OR2_X1 U12315 ( .A1(n10515), .A2(n10512), .ZN(n10511) );
  INV_X1 U12316 ( .A(n15799), .ZN(n10512) );
  AND2_X1 U12317 ( .A1(n11432), .A2(n11431), .ZN(n15829) );
  OR2_X1 U12318 ( .A1(n14585), .A2(n14641), .ZN(n15830) );
  INV_X1 U12319 ( .A(n14575), .ZN(n10501) );
  OR2_X1 U12320 ( .A1(n19898), .A2(n13373), .ZN(n16160) );
  OR2_X1 U12321 ( .A1(n19898), .A2(n13362), .ZN(n14269) );
  AND2_X2 U12322 ( .A1(n13372), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n16790)
         );
  OR3_X1 U12323 ( .A1(n12518), .A2(n12457), .A3(n10408), .ZN(n10407) );
  OR2_X1 U12324 ( .A1(n12518), .A2(n10408), .ZN(n10406) );
  NOR3_X1 U12325 ( .A1(n12516), .A2(n12518), .A3(n16200), .ZN(n13734) );
  INV_X1 U12326 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13730) );
  INV_X1 U12327 ( .A(n16223), .ZN(n10194) );
  INV_X1 U12328 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U12329 ( .A1(n12498), .A2(n10400), .ZN(n12500) );
  INV_X1 U12330 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16285) );
  INV_X1 U12331 ( .A(n16322), .ZN(n10364) );
  NOR3_X1 U12332 ( .A1(n9629), .A2(n10413), .A3(n12486), .ZN(n12490) );
  NOR2_X1 U12333 ( .A1(n9629), .A2(n12486), .ZN(n12488) );
  AND3_X1 U12334 ( .A1(n11150), .A2(n11149), .A3(n11148), .ZN(n14608) );
  NOR2_X1 U12335 ( .A1(n12473), .A2(n10414), .ZN(n12482) );
  NAND2_X1 U12336 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n9602), .ZN(
        n10414) );
  AND3_X1 U12337 ( .A1(n11142), .A2(n11141), .A3(n11140), .ZN(n15889) );
  AND3_X1 U12338 ( .A1(n11139), .A2(n11138), .A3(n11137), .ZN(n14602) );
  NAND2_X1 U12339 ( .A1(n10415), .A2(n10416), .ZN(n12477) );
  AND3_X1 U12340 ( .A1(n11134), .A2(n11133), .A3(n11132), .ZN(n14457) );
  OR2_X1 U12341 ( .A1(n12471), .A2(n21556), .ZN(n12473) );
  INV_X1 U12342 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16403) );
  NOR2_X1 U12343 ( .A1(n12473), .A2(n16403), .ZN(n12475) );
  AND3_X1 U12344 ( .A1(n11124), .A2(n11123), .A3(n11122), .ZN(n14374) );
  NAND2_X1 U12345 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12465) );
  NAND2_X1 U12346 ( .A1(n16677), .A2(n9679), .ZN(n16475) );
  NOR2_X1 U12347 ( .A1(n13762), .A2(n10104), .ZN(n10103) );
  INV_X1 U12348 ( .A(n13718), .ZN(n10104) );
  NOR2_X1 U12349 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  INV_X1 U12350 ( .A(n13760), .ZN(n10108) );
  INV_X1 U12351 ( .A(n13761), .ZN(n10109) );
  AND2_X1 U12352 ( .A1(n11254), .A2(n9588), .ZN(n11256) );
  AND2_X1 U12353 ( .A1(n10564), .A2(n13772), .ZN(n10563) );
  INV_X1 U12354 ( .A(n13779), .ZN(n10562) );
  OR3_X1 U12355 ( .A1(n13750), .A2(n13768), .A3(n10539), .ZN(n13761) );
  NAND2_X1 U12356 ( .A1(n10390), .A2(n9827), .ZN(n10111) );
  AND2_X1 U12357 ( .A1(n10247), .A2(n11760), .ZN(n9827) );
  NOR2_X1 U12358 ( .A1(n10100), .A2(n9691), .ZN(n10517) );
  NAND2_X1 U12359 ( .A1(n10246), .A2(n10247), .ZN(n10245) );
  INV_X1 U12360 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16217) );
  AND3_X1 U12361 ( .A1(n11726), .A2(n11725), .A3(n11724), .ZN(n15700) );
  OR2_X1 U12362 ( .A1(n15741), .A2(n11771), .ZN(n11772) );
  NAND2_X1 U12363 ( .A1(n15731), .A2(n9736), .ZN(n15717) );
  NAND2_X1 U12364 ( .A1(n10044), .A2(n9750), .ZN(n11082) );
  NAND2_X1 U12365 ( .A1(n10045), .A2(n9747), .ZN(n10044) );
  CLKBUF_X1 U12366 ( .A(n11441), .Z(n11703) );
  OR2_X1 U12367 ( .A1(n16605), .A2(n10269), .ZN(n10086) );
  NOR2_X1 U12368 ( .A1(n19954), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10269) );
  NOR2_X1 U12369 ( .A1(n19963), .A2(n10354), .ZN(n10353) );
  INV_X1 U12370 ( .A(n10355), .ZN(n10354) );
  INV_X1 U12371 ( .A(n14613), .ZN(n11154) );
  NAND2_X1 U12372 ( .A1(n11045), .A2(n16330), .ZN(n16324) );
  NAND2_X1 U12373 ( .A1(n11710), .A2(n16296), .ZN(n16317) );
  NOR2_X1 U12374 ( .A1(n16724), .A2(n9798), .ZN(n11477) );
  AND3_X1 U12375 ( .A1(n11129), .A2(n11128), .A3(n11127), .ZN(n14418) );
  NAND2_X1 U12377 ( .A1(n16432), .A2(n11006), .ZN(n9814) );
  CLKBUF_X1 U12378 ( .A(n16169), .Z(n16170) );
  INV_X1 U12379 ( .A(n11295), .ZN(n11183) );
  AND2_X1 U12380 ( .A1(n10178), .A2(n10174), .ZN(n16737) );
  NAND2_X1 U12381 ( .A1(n16565), .A2(n19940), .ZN(n10178) );
  INV_X1 U12382 ( .A(n10175), .ZN(n10174) );
  OAI21_X1 U12383 ( .B1(n19954), .B2(n19939), .A(n19941), .ZN(n10175) );
  NAND2_X1 U12384 ( .A1(n10785), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9897) );
  INV_X1 U12385 ( .A(n10720), .ZN(n13986) );
  NAND2_X1 U12386 ( .A1(n14152), .A2(n14151), .ZN(n14154) );
  INV_X1 U12387 ( .A(n12502), .ZN(n15968) );
  AND2_X2 U12388 ( .A1(n10613), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16745) );
  NOR2_X2 U12389 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16758) );
  INV_X1 U12390 ( .A(n9905), .ZN(n14348) );
  INV_X1 U12391 ( .A(n13039), .ZN(n13020) );
  NAND2_X1 U12392 ( .A1(n14364), .A2(n14363), .ZN(n16863) );
  OR2_X1 U12393 ( .A1(n20034), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19982) );
  NOR2_X1 U12394 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20080) );
  INV_X1 U12395 ( .A(n16791), .ZN(n20013) );
  INV_X1 U12396 ( .A(n20339), .ZN(n20405) );
  INV_X1 U12397 ( .A(n20465), .ZN(n20404) );
  NOR2_X2 U12398 ( .A1(n16788), .A2(n16789), .ZN(n20021) );
  NOR2_X2 U12399 ( .A1(n16790), .A2(n16789), .ZN(n16791) );
  AND2_X1 U12400 ( .A1(n20467), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20023) );
  INV_X1 U12401 ( .A(n16899), .ZN(n16888) );
  OAI21_X1 U12402 ( .B1(n11223), .B2(n11104), .A(n11228), .ZN(n16847) );
  OR2_X1 U12403 ( .A1(n13587), .A2(n11668), .ZN(n11669) );
  NOR2_X1 U12404 ( .A1(n11500), .A2(n10375), .ZN(n11520) );
  OR3_X1 U12405 ( .A1(n17577), .A2(n16963), .A3(n18821), .ZN(n10375) );
  NAND2_X1 U12406 ( .A1(n10374), .A2(n17843), .ZN(n11523) );
  AND2_X1 U12407 ( .A1(n17596), .A2(n17843), .ZN(n17588) );
  OR2_X1 U12408 ( .A1(n17588), .A2(n17589), .ZN(n10374) );
  OR2_X1 U12409 ( .A1(n17617), .A2(n17618), .ZN(n10382) );
  OR2_X1 U12410 ( .A1(n17674), .A2(n18639), .ZN(n10372) );
  NOR2_X1 U12411 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17709), .ZN(n17700) );
  NOR2_X1 U12412 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17737), .ZN(n17721) );
  NOR2_X1 U12413 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17790), .ZN(n17773) );
  NOR2_X1 U12414 ( .A1(n17915), .A2(n17924), .ZN(n17650) );
  NOR2_X1 U12415 ( .A1(n10150), .A2(n17645), .ZN(n10147) );
  INV_X1 U12416 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n10150) );
  NOR2_X1 U12417 ( .A1(n18037), .A2(n10149), .ZN(n10148) );
  OR2_X1 U12418 ( .A1(n14144), .A2(n10159), .ZN(n10158) );
  AND2_X1 U12419 ( .A1(n14389), .A2(n19547), .ZN(n10159) );
  NAND2_X1 U12420 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18429), .ZN(n18417) );
  OR2_X1 U12421 ( .A1(n13444), .A2(n13443), .ZN(n13597) );
  NOR2_X1 U12422 ( .A1(n11638), .A2(n19131), .ZN(n14450) );
  INV_X1 U12423 ( .A(n13636), .ZN(n9935) );
  INV_X1 U12424 ( .A(n10446), .ZN(n13566) );
  NOR2_X1 U12425 ( .A1(n13563), .A2(n16960), .ZN(n10444) );
  NOR3_X1 U12426 ( .A1(n11500), .A2(n17577), .A3(n16963), .ZN(n16916) );
  OR2_X1 U12427 ( .A1(n18844), .A2(n18854), .ZN(n18550) );
  AND2_X1 U12428 ( .A1(n9728), .A2(n17743), .ZN(n18630) );
  INV_X1 U12429 ( .A(n18642), .ZN(n10376) );
  AND2_X1 U12430 ( .A1(n17743), .A2(n10377), .ZN(n18656) );
  NAND2_X1 U12431 ( .A1(n17743), .A2(n9650), .ZN(n18671) );
  NOR2_X1 U12432 ( .A1(n18783), .A2(n17846), .ZN(n10367) );
  INV_X1 U12433 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17846) );
  NOR2_X1 U12434 ( .A1(n17866), .A2(n18783), .ZN(n18762) );
  NOR2_X1 U12435 ( .A1(n10369), .A2(n18783), .ZN(n10366) );
  NOR2_X1 U12436 ( .A1(n19592), .A2(n21509), .ZN(n18790) );
  NAND2_X1 U12437 ( .A1(n10449), .A2(n10446), .ZN(n16925) );
  INV_X1 U12438 ( .A(n16959), .ZN(n17118) );
  OR2_X1 U12439 ( .A1(n17135), .A2(n17120), .ZN(n10231) );
  AND2_X1 U12440 ( .A1(n18694), .A2(n10442), .ZN(n10441) );
  NAND2_X1 U12441 ( .A1(n13561), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10443) );
  OR3_X1 U12442 ( .A1(n13637), .A2(n18668), .A3(n18571), .ZN(n18844) );
  AND2_X1 U12443 ( .A1(n17121), .A2(n10225), .ZN(n10224) );
  INV_X1 U12444 ( .A(n10226), .ZN(n10225) );
  AND2_X1 U12445 ( .A1(n13555), .A2(n17131), .ZN(n17096) );
  NOR2_X1 U12446 ( .A1(n18867), .A2(n10000), .ZN(n18871) );
  OR2_X1 U12447 ( .A1(n18869), .A2(n18868), .ZN(n10000) );
  NOR2_X1 U12448 ( .A1(n18883), .A2(n19082), .ZN(n18893) );
  AOI21_X1 U12449 ( .B1(n13553), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10081), .ZN(n10080) );
  AND2_X1 U12450 ( .A1(n18694), .A2(n10082), .ZN(n10081) );
  AND2_X1 U12451 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17131) );
  OAI21_X1 U12452 ( .B1(n19545), .B2(n18937), .A(n18930), .ZN(n18867) );
  INV_X1 U12453 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18912) );
  NAND2_X1 U12454 ( .A1(n10227), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10226) );
  NOR2_X1 U12455 ( .A1(n18912), .A2(n10228), .ZN(n10227) );
  AND2_X1 U12456 ( .A1(n19543), .A2(n18411), .ZN(n18971) );
  NOR2_X1 U12457 ( .A1(n18956), .A2(n18940), .ZN(n18701) );
  NAND2_X1 U12458 ( .A1(n18701), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18700) );
  INV_X1 U12459 ( .A(n16994), .ZN(n18939) );
  NAND2_X1 U12460 ( .A1(n13623), .A2(n17049), .ZN(n18972) );
  NAND2_X1 U12461 ( .A1(n13620), .A2(n9995), .ZN(n17050) );
  AOI21_X1 U12462 ( .B1(n13619), .B2(n9996), .A(n9662), .ZN(n9995) );
  INV_X1 U12463 ( .A(n13619), .ZN(n13621) );
  NAND2_X1 U12464 ( .A1(n17050), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17049) );
  NAND2_X1 U12465 ( .A1(n18746), .A2(n13617), .ZN(n18737) );
  NAND2_X1 U12466 ( .A1(n18758), .A2(n18759), .ZN(n18757) );
  NAND2_X1 U12467 ( .A1(n18784), .A2(n13613), .ZN(n18776) );
  NOR2_X1 U12468 ( .A1(n18776), .A2(n18777), .ZN(n18775) );
  XNOR2_X1 U12469 ( .A(n13611), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18800) );
  OAI21_X1 U12470 ( .B1(n14215), .B2(n10219), .A(n10218), .ZN(n13610) );
  NAND2_X1 U12471 ( .A1(n14215), .A2(n13609), .ZN(n10218) );
  NAND2_X1 U12472 ( .A1(n10221), .A2(n10220), .ZN(n10219) );
  NOR2_X1 U12473 ( .A1(n11542), .A2(n10301), .ZN(n10300) );
  AND4_X1 U12474 ( .A1(n11587), .A2(n11586), .A3(n11585), .A4(n11584), .ZN(
        n11597) );
  NOR2_X1 U12475 ( .A1(n11623), .A2(n11622), .ZN(n19122) );
  INV_X1 U12476 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11621) );
  INV_X1 U12477 ( .A(n11638), .ZN(n19135) );
  NAND2_X1 U12478 ( .A1(n19591), .A2(n19106), .ZN(n19252) );
  INV_X1 U12479 ( .A(n14273), .ZN(n21398) );
  INV_X1 U12480 ( .A(n20702), .ZN(n20736) );
  AND2_X1 U12481 ( .A1(n21402), .A2(n13799), .ZN(n20735) );
  XNOR2_X1 U12482 ( .A(n14201), .B(n12360), .ZN(n10457) );
  AND2_X1 U12483 ( .A1(n21402), .A2(n13801), .ZN(n15071) );
  NOR2_X1 U12484 ( .A1(n9887), .A2(n9751), .ZN(n20744) );
  AND2_X1 U12485 ( .A1(n15059), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20738) );
  INV_X1 U12486 ( .A(n15114), .ZN(n15104) );
  INV_X1 U12487 ( .A(n15108), .ZN(n15111) );
  INV_X1 U12488 ( .A(n14763), .ZN(n15121) );
  NAND2_X1 U12489 ( .A1(n15151), .A2(n13854), .ZN(n15153) );
  CLKBUF_X1 U12490 ( .A(n13850), .Z(n15165) );
  INV_X1 U12491 ( .A(n15153), .ZN(n15164) );
  INV_X1 U12492 ( .A(n15151), .ZN(n15179) );
  NOR2_X1 U12493 ( .A1(n15179), .A2(n14209), .ZN(n15180) );
  NAND2_X1 U12494 ( .A1(n13837), .A2(n13836), .ZN(n15151) );
  OR2_X1 U12495 ( .A1(n13835), .A2(n13948), .ZN(n13836) );
  NAND2_X1 U12496 ( .A1(n13973), .A2(n14115), .ZN(n13837) );
  INV_X1 U12497 ( .A(n15180), .ZN(n14639) );
  AND2_X1 U12498 ( .A1(n14118), .A2(n17346), .ZN(n20766) );
  INV_X1 U12499 ( .A(n20766), .ZN(n20786) );
  INV_X2 U12500 ( .A(n20772), .ZN(n20783) );
  INV_X1 U12501 ( .A(n14536), .ZN(n20797) );
  INV_X1 U12502 ( .A(n14533), .ZN(n20805) );
  INV_X1 U12503 ( .A(n20804), .ZN(n14536) );
  XNOR2_X1 U12504 ( .A(n13793), .B(n13813), .ZN(n14681) );
  INV_X1 U12505 ( .A(n13791), .ZN(n13792) );
  OAI21_X1 U12506 ( .B1(n13712), .B2(n13713), .A(n13790), .ZN(n14689) );
  AOI21_X1 U12507 ( .B1(n14789), .B2(n14787), .A(n14788), .ZN(n15203) );
  INV_X1 U12508 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15217) );
  INV_X1 U12509 ( .A(n9886), .ZN(n12697) );
  AND2_X1 U12510 ( .A1(n14969), .A2(n14968), .ZN(n15328) );
  INV_X1 U12511 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20701) );
  XNOR2_X1 U12512 ( .A(n9869), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13825) );
  NAND2_X1 U12513 ( .A1(n9871), .A2(n9870), .ZN(n9869) );
  AND2_X1 U12514 ( .A1(n10321), .A2(n10318), .ZN(n9870) );
  NAND3_X1 U12515 ( .A1(n13714), .A2(n10322), .A3(n9753), .ZN(n9871) );
  XNOR2_X1 U12516 ( .A(n12449), .B(n12448), .ZN(n15084) );
  MUX2_X1 U12517 ( .A(n14674), .B(n14671), .S(n14753), .Z(n12449) );
  INV_X1 U12518 ( .A(n15396), .ZN(n15417) );
  INV_X1 U12519 ( .A(n15190), .ZN(n9971) );
  NAND2_X1 U12520 ( .A1(n15443), .A2(n12340), .ZN(n15439) );
  NAND2_X1 U12521 ( .A1(n12227), .A2(n12226), .ZN(n15212) );
  NAND2_X1 U12522 ( .A1(n15472), .A2(n12338), .ZN(n15456) );
  AND2_X1 U12523 ( .A1(n12336), .A2(n12335), .ZN(n15502) );
  NAND2_X1 U12524 ( .A1(n10499), .A2(n12193), .ZN(n17374) );
  INV_X1 U12525 ( .A(n17378), .ZN(n10036) );
  NAND2_X1 U12526 ( .A1(n10486), .A2(n10485), .ZN(n10484) );
  OR2_X1 U12527 ( .A1(n12455), .A2(n14089), .ZN(n15562) );
  NAND2_X1 U12528 ( .A1(n12455), .A2(n20716), .ZN(n14196) );
  OR2_X1 U12529 ( .A1(n12455), .A2(n12454), .ZN(n17390) );
  INV_X1 U12530 ( .A(n17397), .ZN(n17429) );
  INV_X1 U12531 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12593) );
  INV_X1 U12532 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14101) );
  NOR2_X1 U12533 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15629) );
  OAI21_X1 U12534 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21197), .A(n13978), 
        .ZN(n15640) );
  OAI211_X1 U12535 ( .C1(n20825), .C2(n20822), .A(n20820), .B(n21134), .ZN(
        n20857) );
  NOR2_X2 U12536 ( .A1(n20930), .A2(n21262), .ZN(n20946) );
  OAI21_X1 U12537 ( .B1(n10603), .B2(n20960), .A(n21276), .ZN(n20977) );
  OAI21_X1 U12538 ( .B1(n21267), .B2(n20955), .A(n20954), .ZN(n20975) );
  OAI211_X1 U12539 ( .C1(n10593), .C2(n21197), .A(n21134), .B(n21074), .ZN(
        n21091) );
  NOR2_X2 U12540 ( .A1(n21161), .A2(n21232), .ZN(n21150) );
  OAI211_X1 U12541 ( .C1(n10602), .C2(n21197), .A(n21276), .B(n21196), .ZN(
        n21227) );
  AOI22_X1 U12542 ( .A1(n21195), .A2(n21192), .B1(n21190), .B2(n21189), .ZN(
        n21231) );
  OAI211_X1 U12543 ( .C1(n21410), .C2(n21277), .A(n21276), .B(n21275), .ZN(
        n21421) );
  AND2_X1 U12544 ( .A1(n20855), .A2(n20821), .ZN(n21300) );
  AND2_X1 U12545 ( .A1(n20855), .A2(n20833), .ZN(n21318) );
  AND2_X1 U12546 ( .A1(n20855), .A2(n20836), .ZN(n21323) );
  AND2_X1 U12547 ( .A1(n20855), .A2(n20839), .ZN(n21329) );
  AND2_X1 U12548 ( .A1(n20855), .A2(n20843), .ZN(n21335) );
  AND2_X1 U12549 ( .A1(n20855), .A2(n20846), .ZN(n21341) );
  INV_X1 U12550 ( .A(n21415), .ZN(n21351) );
  NOR2_X1 U12551 ( .A1(n14096), .A2(n21197), .ZN(n17358) );
  NAND2_X1 U12552 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21404) );
  INV_X1 U12553 ( .A(n17359), .ZN(n21399) );
  AOI221_X1 U12554 ( .B1(n10287), .B2(n21357), .C1(n17350), .C2(n21357), .A(
        n17435), .ZN(n17439) );
  INV_X1 U12555 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n13869) );
  CLKBUF_X1 U12556 ( .A(n11455), .Z(n15652) );
  NAND2_X1 U12557 ( .A1(n14157), .A2(n14156), .ZN(n16884) );
  INV_X1 U12558 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20408) );
  INV_X1 U12559 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19748) );
  NAND2_X1 U12560 ( .A1(n13765), .A2(n13398), .ZN(n13767) );
  OAI211_X1 U12561 ( .C1(n11777), .C2(n9786), .A(n11782), .B(n11780), .ZN(
        n15704) );
  INV_X1 U12562 ( .A(n11777), .ZN(n11779) );
  NAND2_X1 U12564 ( .A1(n14717), .A2(n12541), .ZN(n19830) );
  OR2_X1 U12565 ( .A1(n11425), .A2(n11424), .ZN(n19847) );
  OR2_X1 U12566 ( .A1(n11397), .A2(n11396), .ZN(n14616) );
  OR2_X1 U12567 ( .A1(n11370), .A2(n11369), .ZN(n16062) );
  OR2_X1 U12568 ( .A1(n11356), .A2(n11355), .ZN(n19854) );
  OR2_X1 U12569 ( .A1(n11327), .A2(n11326), .ZN(n14595) );
  INV_X2 U12570 ( .A(n19866), .ZN(n16065) );
  NAND2_X1 U12571 ( .A1(n10425), .A2(n15986), .ZN(n15982) );
  NAND2_X1 U12572 ( .A1(n13269), .A2(n10426), .ZN(n10425) );
  NAND2_X1 U12573 ( .A1(n15991), .A2(n15990), .ZN(n10030) );
  AND2_X1 U12574 ( .A1(n9649), .A2(n13158), .ZN(n10596) );
  INV_X1 U12575 ( .A(n16160), .ZN(n19868) );
  NAND2_X1 U12576 ( .A1(n10436), .A2(n9752), .ZN(n16178) );
  NAND2_X1 U12577 ( .A1(n14362), .A2(n13351), .ZN(n13352) );
  AND2_X1 U12578 ( .A1(n14167), .A2(n20526), .ZN(n19928) );
  OR2_X1 U12579 ( .A1(n14048), .A2(n13926), .ZN(n13993) );
  OR2_X1 U12580 ( .A1(n13889), .A2(n12562), .ZN(n13928) );
  INV_X1 U12581 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21556) );
  OAI21_X1 U12582 ( .B1(n16466), .B2(n19964), .A(n16464), .ZN(n9968) );
  NAND2_X1 U12583 ( .A1(n10336), .A2(n16462), .ZN(n16191) );
  NAND2_X1 U12584 ( .A1(n16461), .A2(n19960), .ZN(n16468) );
  XNOR2_X1 U12585 ( .A(n16199), .B(n16198), .ZN(n16460) );
  NAND2_X1 U12586 ( .A1(n10192), .A2(n10599), .ZN(n16199) );
  NAND2_X1 U12587 ( .A1(n9946), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16250) );
  INV_X1 U12588 ( .A(n10051), .ZN(n16268) );
  OR2_X1 U12589 ( .A1(n16605), .A2(n9862), .ZN(n9861) );
  OR2_X1 U12590 ( .A1(n9865), .A2(n9863), .ZN(n9862) );
  INV_X1 U12591 ( .A(n11695), .ZN(n9865) );
  OR2_X1 U12592 ( .A1(n16605), .A2(n9863), .ZN(n11698) );
  NOR2_X1 U12593 ( .A1(n16605), .A2(n11480), .ZN(n16554) );
  OR2_X1 U12594 ( .A1(n16559), .A2(n16561), .ZN(n10090) );
  NAND2_X1 U12595 ( .A1(n10365), .A2(n16322), .ZN(n16308) );
  AND2_X1 U12596 ( .A1(n16536), .A2(n11476), .ZN(n16633) );
  INV_X1 U12597 ( .A(n11710), .ZN(n16379) );
  NAND2_X1 U12598 ( .A1(n10544), .A2(n10547), .ZN(n16391) );
  NAND2_X1 U12599 ( .A1(n10338), .A2(n10548), .ZN(n10544) );
  INV_X1 U12600 ( .A(n10340), .ZN(n10545) );
  NAND2_X1 U12601 ( .A1(n11477), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16695) );
  XNOR2_X1 U12602 ( .A(n9912), .B(n9655), .ZN(n16699) );
  NAND2_X1 U12603 ( .A1(n16737), .A2(n9851), .ZN(n16727) );
  NAND2_X1 U12604 ( .A1(n9852), .A2(n16736), .ZN(n9851) );
  INV_X1 U12605 ( .A(n16449), .ZN(n10164) );
  NAND2_X1 U12606 ( .A1(n10177), .A2(n10176), .ZN(n19941) );
  INV_X1 U12607 ( .A(n11494), .ZN(n10177) );
  INV_X1 U12608 ( .A(n16797), .ZN(n16798) );
  INV_X1 U12609 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16860) );
  AND2_X1 U12610 ( .A1(n10019), .A2(n9671), .ZN(n14223) );
  NAND2_X1 U12611 ( .A1(n14442), .A2(n11288), .ZN(n15939) );
  INV_X1 U12612 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17363) );
  AOI21_X1 U12613 ( .B1(n10592), .B2(n14702), .A(n14701), .ZN(n16868) );
  XNOR2_X1 U12614 ( .A(n14137), .B(n14136), .ZN(n16797) );
  AND2_X1 U12615 ( .A1(n16844), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16883) );
  NOR2_X2 U12616 ( .A1(n20267), .A2(n20116), .ZN(n20020) );
  OAI21_X1 U12617 ( .B1(n19986), .B2(n19985), .A(n19984), .ZN(n20027) );
  AND2_X1 U12618 ( .A1(n19981), .A2(n20467), .ZN(n20025) );
  OAI21_X1 U12619 ( .B1(n20088), .B2(n20087), .A(n20086), .ZN(n20105) );
  OAI21_X1 U12620 ( .B1(n20138), .B2(n16814), .A(n20122), .ZN(n20140) );
  OAI21_X1 U12621 ( .B1(n20153), .B2(n20152), .A(n20151), .ZN(n20170) );
  NOR2_X1 U12622 ( .A1(n20195), .A2(n20375), .ZN(n20177) );
  INV_X1 U12623 ( .A(n20191), .ZN(n20180) );
  NOR2_X1 U12624 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20200), .ZN(
        n20189) );
  AND2_X1 U12625 ( .A1(n16809), .A2(n16808), .ZN(n20190) );
  AND2_X1 U12626 ( .A1(n20270), .A2(n20627), .ZN(n20236) );
  NAND2_X1 U12627 ( .A1(n20233), .A2(n20232), .ZN(n20260) );
  INV_X1 U12628 ( .A(n10889), .ZN(n20268) );
  OAI21_X1 U12629 ( .B1(n10889), .B2(n20290), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20271) );
  AND2_X1 U12630 ( .A1(n16831), .A2(n16817), .ZN(n20309) );
  OAI21_X1 U12631 ( .B1(n16818), .B2(n20309), .A(n20467), .ZN(n20312) );
  OAI21_X1 U12632 ( .B1(n16826), .B2(n16821), .A(n16820), .ZN(n20310) );
  NOR2_X1 U12633 ( .A1(n20367), .A2(n20079), .ZN(n20340) );
  OAI21_X1 U12634 ( .B1(n20342), .B2(n20338), .A(n20337), .ZN(n20362) );
  INV_X1 U12635 ( .A(n20497), .ZN(n20391) );
  AOI22_X1 U12636 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16791), .ZN(n20439) );
  OAI22_X1 U12637 ( .A1(n21495), .A2(n20013), .B1(n16076), .B2(n20011), .ZN(
        n20440) );
  OAI22_X1 U12638 ( .A1(n20014), .A2(n20013), .B1(n20012), .B2(n20011), .ZN(
        n20446) );
  AOI22_X1 U12639 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n16791), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n20021), .ZN(n20473) );
  INV_X1 U12640 ( .A(n20419), .ZN(n20470) );
  AND2_X1 U12641 ( .A1(n20023), .A2(n16856), .ZN(n20461) );
  AOI22_X1 U12642 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n16791), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n20021), .ZN(n20479) );
  INV_X1 U12643 ( .A(n20421), .ZN(n20476) );
  AND2_X1 U12644 ( .A1(n20023), .A2(n11232), .ZN(n20474) );
  AND2_X1 U12645 ( .A1(n20467), .A2(n19989), .ZN(n20475) );
  AOI22_X1 U12646 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16791), .ZN(n20485) );
  INV_X1 U12647 ( .A(n20426), .ZN(n20482) );
  AND2_X1 U12648 ( .A1(n20023), .A2(n19992), .ZN(n20480) );
  AND2_X1 U12649 ( .A1(n20467), .A2(n19993), .ZN(n20481) );
  INV_X1 U12650 ( .A(n20434), .ZN(n20488) );
  AND2_X1 U12651 ( .A1(n20023), .A2(n19997), .ZN(n20486) );
  AND2_X1 U12652 ( .A1(n20467), .A2(n19998), .ZN(n20487) );
  AOI22_X1 U12653 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16791), .ZN(n20497) );
  INV_X1 U12654 ( .A(n20439), .ZN(n20494) );
  AND2_X1 U12655 ( .A1(n20467), .A2(n20003), .ZN(n20493) );
  INV_X1 U12656 ( .A(n20443), .ZN(n20500) );
  AND2_X1 U12657 ( .A1(n20023), .A2(n20006), .ZN(n20498) );
  AND2_X1 U12658 ( .A1(n20467), .A2(n20007), .ZN(n20499) );
  INV_X1 U12659 ( .A(n20440), .ZN(n20503) );
  INV_X1 U12660 ( .A(n20449), .ZN(n20506) );
  AND2_X1 U12661 ( .A1(n20023), .A2(n20015), .ZN(n20504) );
  AND2_X1 U12662 ( .A1(n20467), .A2(n20016), .ZN(n20505) );
  INV_X1 U12663 ( .A(n20446), .ZN(n20509) );
  INV_X1 U12664 ( .A(n20458), .ZN(n20514) );
  AND2_X1 U12665 ( .A1(n20467), .A2(n20026), .ZN(n20512) );
  INV_X1 U12666 ( .A(n20463), .ZN(n20459) );
  OR2_X1 U12667 ( .A1(n12461), .A2(n12460), .ZN(n19838) );
  NAND2_X1 U12668 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n16887) );
  AND2_X1 U12669 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13867), .ZN(n16904) );
  NOR3_X1 U12670 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20533), .A3(n19734), 
        .ZN(n20526) );
  INV_X1 U12671 ( .A(n19707), .ZN(n19720) );
  INV_X1 U12672 ( .A(n14385), .ZN(n18493) );
  INV_X1 U12673 ( .A(n10121), .ZN(n17546) );
  INV_X1 U12674 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19591) );
  NAND2_X1 U12675 ( .A1(n19703), .A2(n14140), .ZN(n18492) );
  AOI21_X1 U12676 ( .B1(n19005), .B2(n16908), .A(n10132), .ZN(n10131) );
  OAI21_X1 U12677 ( .B1(n10135), .B2(n19709), .A(n10134), .ZN(n10132) );
  AND2_X1 U12678 ( .A1(n10379), .A2(n9766), .ZN(n17598) );
  NOR2_X1 U12679 ( .A1(n17632), .A2(n10370), .ZN(n17633) );
  NOR2_X1 U12680 ( .A1(n18579), .A2(n17639), .ZN(n17638) );
  AND2_X1 U12681 ( .A1(n17654), .A2(n17843), .ZN(n17639) );
  NOR2_X1 U12682 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17684), .ZN(n17672) );
  NOR2_X1 U12683 ( .A1(n17664), .A2(n17665), .ZN(n17663) );
  AND2_X1 U12684 ( .A1(n10372), .A2(n17843), .ZN(n17664) );
  NOR2_X1 U12685 ( .A1(n17882), .A2(n10373), .ZN(n17674) );
  AND2_X1 U12686 ( .A1(n18593), .A2(n17719), .ZN(n10373) );
  INV_X1 U12687 ( .A(n10372), .ZN(n17673) );
  NOR2_X1 U12688 ( .A1(n17906), .A2(n17651), .ZN(n17726) );
  NOR2_X1 U12689 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17760), .ZN(n17747) );
  NOR2_X1 U12690 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17798), .ZN(n17797) );
  INV_X1 U12691 ( .A(n17887), .ZN(n17928) );
  INV_X1 U12692 ( .A(n17916), .ZN(n17929) );
  INV_X1 U12693 ( .A(n17650), .ZN(n17930) );
  NAND2_X1 U12694 ( .A1(n17997), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17989) );
  AND2_X1 U12695 ( .A1(n18053), .A2(n9628), .ZN(n18000) );
  NOR2_X1 U12696 ( .A1(n18120), .A2(n10154), .ZN(n18088) );
  NOR2_X1 U12697 ( .A1(n18264), .A2(n10155), .ZN(n18173) );
  NAND2_X1 U12698 ( .A1(n9783), .A2(n9624), .ZN(n10155) );
  NOR2_X1 U12699 ( .A1(n18231), .A2(n18230), .ZN(n18234) );
  NOR2_X1 U12700 ( .A1(n18308), .A2(n10296), .ZN(n10294) );
  OR2_X1 U12701 ( .A1(n10297), .A2(n10299), .ZN(n10296) );
  INV_X1 U12702 ( .A(n10297), .ZN(n10295) );
  NOR2_X1 U12703 ( .A1(n18438), .A2(n18316), .ZN(n18311) );
  NAND2_X1 U12704 ( .A1(n18330), .A2(n10304), .ZN(n18316) );
  AND2_X1 U12705 ( .A1(n9625), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U12706 ( .A1(n18330), .A2(n10305), .ZN(n18325) );
  OAI211_X1 U12707 ( .C1(n18216), .C2(n17962), .A(n11611), .B(n11610), .ZN(
        n11612) );
  INV_X1 U12708 ( .A(n18368), .ZN(n18337) );
  INV_X1 U12709 ( .A(n18374), .ZN(n18362) );
  INV_X1 U12710 ( .A(n13603), .ZN(n18421) );
  INV_X1 U12711 ( .A(n13597), .ZN(n18426) );
  INV_X1 U12712 ( .A(n18382), .ZN(n18427) );
  AND2_X1 U12713 ( .A1(n14450), .A2(n14241), .ZN(n18382) );
  INV_X1 U12714 ( .A(n18398), .ZN(n18430) );
  NAND2_X1 U12715 ( .A1(n18460), .A2(n18432), .ZN(n18457) );
  NOR2_X1 U12716 ( .A1(n18492), .A2(n18431), .ZN(n18460) );
  INV_X1 U12717 ( .A(n18460), .ZN(n18490) );
  AOI211_X1 U12718 ( .C1(n19705), .C2(n18494), .A(n18493), .B(n18492), .ZN(
        n18532) );
  INV_X1 U12719 ( .A(n18508), .ZN(n18536) );
  NOR2_X1 U12720 ( .A1(n18533), .A2(n19709), .ZN(n18534) );
  AOI21_X1 U12721 ( .B1(n18540), .B2(n10447), .A(n18641), .ZN(n10075) );
  NOR2_X1 U12722 ( .A1(n18597), .A2(n18599), .ZN(n18581) );
  AND2_X1 U12723 ( .A1(n17026), .A2(n13551), .ZN(n18664) );
  INV_X1 U12724 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18783) );
  INV_X1 U12725 ( .A(n16915), .ZN(n19206) );
  INV_X1 U12726 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19592) );
  NAND2_X1 U12727 ( .A1(n10448), .A2(n10447), .ZN(n16939) );
  OAI21_X1 U12728 ( .B1(n10077), .B2(n18411), .A(n10076), .ZN(n17102) );
  NAND2_X1 U12729 ( .A1(n17099), .A2(n18411), .ZN(n10076) );
  AND2_X1 U12730 ( .A1(n10232), .A2(n10229), .ZN(n18825) );
  AOI211_X1 U12731 ( .C1(n17117), .C2(n18971), .A(n18833), .B(n10230), .ZN(
        n10229) );
  OR2_X1 U12732 ( .A1(n16959), .A2(n19545), .ZN(n10232) );
  NAND2_X1 U12733 ( .A1(n10231), .A2(n17119), .ZN(n10230) );
  OR2_X1 U12734 ( .A1(n19082), .A2(n18867), .ZN(n18920) );
  AND2_X1 U12735 ( .A1(n13593), .A2(n19703), .ZN(n19062) );
  INV_X1 U12736 ( .A(n18973), .ZN(n18991) );
  NAND2_X1 U12737 ( .A1(n10437), .A2(n17047), .ZN(n17043) );
  NAND2_X1 U12738 ( .A1(n18751), .A2(n10072), .ZN(n10070) );
  INV_X1 U12739 ( .A(n19062), .ZN(n19082) );
  NOR2_X1 U12740 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n17540) );
  NOR2_X1 U12741 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19690), .ZN(
        n19578) );
  AOI211_X1 U12742 ( .C1(n19703), .C2(n19557), .A(n19107), .B(n14393), .ZN(
        n17178) );
  NOR2_X1 U12743 ( .A1(n19709), .A2(n19139), .ZN(n19425) );
  NOR2_X1 U12744 ( .A1(n19117), .A2(n19139), .ZN(n19497) );
  NAND2_X1 U12745 ( .A1(n10133), .A2(n16908), .ZN(n19577) );
  NAND2_X1 U12746 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19710) );
  INV_X1 U12747 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19690) );
  INV_X1 U12748 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21395) );
  NOR2_X1 U12749 ( .A1(n16788), .A2(n13863), .ZN(n17455) );
  NOR2_X2 U12750 ( .A1(n17498), .A2(n17455), .ZN(n17499) );
  INV_X1 U12751 ( .A(U212), .ZN(n17501) );
  NAND2_X1 U12752 ( .A1(n13774), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10542) );
  NAND2_X1 U12753 ( .A1(n14763), .A2(n15108), .ZN(n13664) );
  NAND2_X1 U12754 ( .A1(n15394), .A2(n17382), .ZN(n10276) );
  OAI21_X1 U12755 ( .B1(n15189), .B2(n20811), .A(n15188), .ZN(n10280) );
  AOI21_X1 U12756 ( .B1(n14763), .B2(n17381), .A(n13013), .ZN(n13014) );
  OAI21_X1 U12757 ( .B1(n15393), .B2(n17397), .A(n9978), .ZN(P1_U3001) );
  INV_X1 U12758 ( .A(n9979), .ZN(n9978) );
  OAI21_X1 U12759 ( .B1(n15388), .B2(n9981), .A(n9980), .ZN(n9979) );
  XNOR2_X1 U12760 ( .A(n21160), .B(n12601), .ZN(n14690) );
  NAND2_X1 U12761 ( .A1(n10492), .A2(n10490), .ZN(n14695) );
  INV_X1 U12762 ( .A(n13754), .ZN(n13756) );
  NAND2_X1 U12763 ( .A1(n12563), .A2(n19836), .ZN(n12564) );
  INV_X1 U12764 ( .A(n12523), .ZN(n12566) );
  AOI21_X1 U12765 ( .B1(n12549), .B2(n19812), .A(n12548), .ZN(n12565) );
  NOR2_X1 U12766 ( .A1(n19835), .A2(n10392), .ZN(n19845) );
  NAND2_X1 U12767 ( .A1(n19866), .A2(n10592), .ZN(n13990) );
  NOR2_X1 U12768 ( .A1(n13783), .A2(n13782), .ZN(n13784) );
  NOR2_X1 U12769 ( .A1(n13738), .A2(n13737), .ZN(n13739) );
  NAND2_X1 U12770 ( .A1(n10538), .A2(n16457), .ZN(n13740) );
  NAND2_X1 U12771 ( .A1(n13733), .A2(n16435), .ZN(n13741) );
  OAI21_X1 U12772 ( .B1(n10098), .B2(n16446), .A(n10095), .ZN(P2_U2985) );
  AOI21_X1 U12773 ( .B1(n10097), .B2(n16435), .A(n10096), .ZN(n10095) );
  OR2_X1 U12774 ( .A1(n16189), .A2(n16188), .ZN(n10096) );
  OAI211_X1 U12775 ( .C1(n16211), .C2(n16459), .A(n10337), .B(n10334), .ZN(
        P2_U2987) );
  AOI21_X1 U12776 ( .B1(n16210), .B2(n16443), .A(n16209), .ZN(n10337) );
  INV_X1 U12777 ( .A(n9949), .ZN(n9948) );
  OAI21_X1 U12778 ( .B1(n16506), .B2(n16459), .A(n9950), .ZN(n9949) );
  NAND2_X1 U12779 ( .A1(n16523), .A2(n16457), .ZN(n16249) );
  INV_X1 U12780 ( .A(n10265), .ZN(n16271) );
  OAI21_X1 U12781 ( .B1(n16547), .B2(n16446), .A(n10266), .ZN(n10265) );
  AOI21_X1 U12782 ( .B1(n16270), .B2(n16443), .A(n16269), .ZN(n10266) );
  INV_X1 U12783 ( .A(n10309), .ZN(n10308) );
  OAI21_X1 U12784 ( .B1(n16551), .B2(n16446), .A(n16289), .ZN(n10309) );
  AOI21_X1 U12785 ( .B1(n10260), .B2(n10259), .A(n10256), .ZN(n16299) );
  NAND2_X1 U12786 ( .A1(n10258), .A2(n10257), .ZN(n10256) );
  OAI211_X1 U12787 ( .C1(n16583), .C2(n16459), .A(n10235), .B(n10234), .ZN(
        P2_U2998) );
  AOI21_X1 U12788 ( .B1(n19851), .B2(n16443), .A(n16305), .ZN(n10234) );
  NAND2_X1 U12789 ( .A1(n9670), .A2(n16457), .ZN(n10235) );
  NOR2_X1 U12790 ( .A1(n13920), .A2(n10393), .ZN(n13923) );
  AND2_X1 U12791 ( .A1(n16443), .A2(n10592), .ZN(n10393) );
  NAND2_X1 U12792 ( .A1(n10538), .A2(n19946), .ZN(n13405) );
  NOR2_X1 U12793 ( .A1(n13729), .A2(n13728), .ZN(n13732) );
  NAND2_X1 U12794 ( .A1(n10058), .A2(n10336), .ZN(n11818) );
  OAI21_X1 U12795 ( .B1(n16485), .B2(n19974), .A(n9849), .ZN(P2_U3020) );
  AOI21_X1 U12796 ( .B1(n16484), .B2(n19946), .A(n9850), .ZN(n9849) );
  OR2_X1 U12797 ( .A1(n16482), .A2(n16483), .ZN(n9850) );
  OR2_X1 U12798 ( .A1(n16493), .A2(n16494), .ZN(n9812) );
  NAND2_X1 U12799 ( .A1(n9944), .A2(n9943), .ZN(n16509) );
  AOI21_X1 U12800 ( .B1(n16523), .B2(n19946), .A(n16522), .ZN(n16524) );
  OAI21_X1 U12801 ( .B1(n16547), .B2(n19963), .A(n16548), .ZN(n10043) );
  NAND2_X1 U12802 ( .A1(n9904), .A2(n10168), .ZN(n16574) );
  OAI211_X1 U12803 ( .C1(n16586), .C2(n16585), .A(n9845), .B(n9843), .ZN(
        P2_U3030) );
  AOI21_X1 U12804 ( .B1(n16584), .B2(n16585), .A(n9846), .ZN(n9845) );
  NAND2_X1 U12805 ( .A1(n9844), .A2(n17444), .ZN(n9843) );
  AND2_X1 U12806 ( .A1(n9823), .A2(n9822), .ZN(n17299) );
  NOR2_X1 U12807 ( .A1(n17297), .A2(n17296), .ZN(n9822) );
  NAND2_X1 U12808 ( .A1(n10388), .A2(n9677), .ZN(P3_U2640) );
  OR2_X1 U12809 ( .A1(n17565), .A2(n9789), .ZN(n10388) );
  NOR4_X1 U12810 ( .A1(n11684), .A2(n17567), .A3(n11683), .A4(n11682), .ZN(
        n11685) );
  AOI22_X1 U12811 ( .A1(n17983), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n10152), 
        .B2(n17982), .ZN(n17984) );
  INV_X1 U12812 ( .A(n10153), .ZN(n10152) );
  NAND2_X1 U12813 ( .A1(n18053), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n18038) );
  NOR2_X1 U12814 ( .A1(n18120), .A2(n18123), .ZN(n18104) );
  NOR4_X1 U12815 ( .A1(n18588), .A2(n18856), .A3(n10442), .A4(n18854), .ZN(
        n16980) );
  OAI21_X1 U12816 ( .B1(n16923), .B2(n19095), .A(n13647), .ZN(n13648) );
  NAND2_X1 U12817 ( .A1(n9704), .A2(n9997), .ZN(P3_U2842) );
  OAI21_X1 U12818 ( .B1(n18901), .B2(n18897), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9997) );
  OAI21_X1 U12819 ( .B1(n18899), .B2(n19012), .A(n18898), .ZN(n9999) );
  NAND2_X1 U12820 ( .A1(n17455), .A2(U214), .ZN(U212) );
  INV_X1 U12821 ( .A(n10795), .ZN(n10769) );
  AND2_X2 U12822 ( .A1(n13336), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10839) );
  INV_X1 U12823 ( .A(n17208), .ZN(n11548) );
  INV_X2 U12825 ( .A(n14659), .ZN(n18244) );
  NAND2_X1 U12826 ( .A1(n12878), .A2(n12877), .ZN(n14823) );
  AND2_X1 U12827 ( .A1(n14576), .A2(n10502), .ZN(n14548) );
  OR2_X1 U12828 ( .A1(n14549), .A2(n14569), .ZN(n14568) );
  AND4_X1 U12829 ( .A1(n10331), .A2(n15296), .A3(n9733), .A4(n15320), .ZN(
        n9595) );
  AND2_X1 U12830 ( .A1(n11225), .A2(n11222), .ZN(n9596) );
  AND2_X1 U12831 ( .A1(n9605), .A2(n11693), .ZN(n9597) );
  INV_X2 U12832 ( .A(n16910), .ZN(n17882) );
  AND3_X1 U12833 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_26__SCAN_IN), .ZN(n9598) );
  AND2_X2 U12834 ( .A1(n13334), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10832) );
  INV_X1 U12835 ( .A(n11524), .ZN(n18202) );
  NAND2_X1 U12836 ( .A1(n17743), .A2(n9641), .ZN(n11504) );
  NAND2_X1 U12837 ( .A1(n10216), .A2(n12628), .ZN(n10215) );
  AND2_X2 U12838 ( .A1(n13338), .A2(n10635), .ZN(n10882) );
  INV_X1 U12839 ( .A(n18251), .ZN(n11603) );
  NAND2_X1 U12840 ( .A1(n14913), .A2(n14901), .ZN(n14879) );
  AND2_X1 U12841 ( .A1(n11802), .A2(n9738), .ZN(n15684) );
  AND2_X1 U12842 ( .A1(n10212), .A2(n12629), .ZN(n14646) );
  AND2_X1 U12843 ( .A1(n12878), .A2(n10571), .ZN(n14812) );
  NAND2_X1 U12844 ( .A1(n15888), .A2(n10557), .ZN(n14607) );
  NOR3_X1 U12845 ( .A1(n14549), .A2(n14569), .A3(n14572), .ZN(n9599) );
  NAND2_X1 U12846 ( .A1(n12629), .A2(n12628), .ZN(n14624) );
  NOR2_X1 U12847 ( .A1(n14549), .A2(n10509), .ZN(n14578) );
  NAND2_X2 U12848 ( .A1(n9894), .A2(n10764), .ZN(n11118) );
  AND2_X1 U12849 ( .A1(n12297), .A2(n12264), .ZN(n9601) );
  AND2_X1 U12850 ( .A1(n10416), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9602) );
  AND2_X1 U12851 ( .A1(n16323), .A2(n16330), .ZN(n9603) );
  INV_X1 U12852 ( .A(n9631), .ZN(n10339) );
  AND4_X1 U12853 ( .A1(n10894), .A2(n10893), .A3(n10892), .A4(n10891), .ZN(
        n9604) );
  AND2_X1 U12854 ( .A1(n11163), .A2(n10552), .ZN(n9605) );
  AND3_X1 U12855 ( .A1(n10216), .A2(n12628), .A3(n9765), .ZN(n9606) );
  INV_X1 U12856 ( .A(n13547), .ZN(n10074) );
  AND2_X1 U12857 ( .A1(n9961), .A2(n9683), .ZN(n9607) );
  OAI21_X1 U12858 ( .B1(n17047), .B2(n9784), .A(n18575), .ZN(n10083) );
  AND2_X1 U12859 ( .A1(n10547), .A2(n10339), .ZN(n9608) );
  AND2_X1 U12860 ( .A1(n15379), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9609) );
  OR2_X1 U12861 ( .A1(n12306), .A2(n11946), .ZN(n9610) );
  AND2_X1 U12862 ( .A1(n9861), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9611) );
  AND2_X1 U12863 ( .A1(n13776), .A2(n10775), .ZN(n9612) );
  AND2_X1 U12864 ( .A1(n9725), .A2(n10727), .ZN(n9613) );
  AND2_X1 U12865 ( .A1(n10985), .A2(n10976), .ZN(n9614) );
  AND2_X1 U12866 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n9615) );
  AND2_X1 U12867 ( .A1(n9597), .A2(n9787), .ZN(n9616) );
  INV_X2 U12868 ( .A(n11076), .ZN(n13768) );
  OR3_X1 U12869 ( .A1(n14562), .A2(n11315), .A3(n10501), .ZN(n9617) );
  AND2_X1 U12870 ( .A1(n10525), .A2(n10519), .ZN(n9618) );
  OR2_X1 U12871 ( .A1(n10532), .A2(n11013), .ZN(n9619) );
  OR2_X1 U12872 ( .A1(n11444), .A2(n15746), .ZN(n9620) );
  NOR2_X1 U12873 ( .A1(n15981), .A2(n10424), .ZN(n9621) );
  AND2_X1 U12874 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n9622) );
  INV_X1 U12875 ( .A(n11033), .ZN(n11778) );
  INV_X2 U12876 ( .A(n12217), .ZN(n15351) );
  AND2_X1 U12877 ( .A1(n9736), .A2(n10566), .ZN(n9623) );
  AND4_X1 U12878 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_9__SCAN_IN), .ZN(n9624) );
  AND2_X1 U12879 ( .A1(n10305), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n9625) );
  AND2_X1 U12880 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9626) );
  AND2_X1 U12881 ( .A1(n10148), .A2(n10147), .ZN(n9627) );
  AND2_X1 U12882 ( .A1(n9627), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n9628) );
  OR2_X1 U12883 ( .A1(n12484), .A2(n12480), .ZN(n9629) );
  AND2_X2 U12884 ( .A1(n13132), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10846) );
  OAI21_X2 U12885 ( .B1(n12582), .B2(n10568), .A(n12167), .ZN(n12601) );
  INV_X1 U12886 ( .A(n9887), .ZN(n15058) );
  INV_X1 U12887 ( .A(n9852), .ZN(n19970) );
  NAND2_X1 U12888 ( .A1(n19956), .A2(n19954), .ZN(n9852) );
  AND4_X1 U12889 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n12322), .ZN(
        n9630) );
  INV_X1 U12890 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10543) );
  AND2_X1 U12891 ( .A1(n11207), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9631) );
  AND2_X2 U12892 ( .A1(n13334), .A2(n10543), .ZN(n10852) );
  INV_X2 U12893 ( .A(n9588), .ZN(n11232) );
  NAND2_X1 U12894 ( .A1(n14646), .A2(n10575), .ZN(n14947) );
  INV_X2 U12895 ( .A(n13810), .ZN(n11955) );
  NAND2_X1 U12896 ( .A1(n14370), .A2(n13056), .ZN(n16028) );
  OR2_X1 U12897 ( .A1(n9629), .A2(n10409), .ZN(n9632) );
  NAND2_X1 U12898 ( .A1(n15801), .A2(n9616), .ZN(n9633) );
  NAND2_X1 U12899 ( .A1(n11023), .A2(n10114), .ZN(n9634) );
  NOR2_X1 U12900 ( .A1(n14585), .A2(n10515), .ZN(n9635) );
  AND2_X1 U12901 ( .A1(n14855), .A2(n14840), .ZN(n14832) );
  NOR2_X1 U12902 ( .A1(n9633), .A2(n15749), .ZN(n15747) );
  NAND2_X1 U12903 ( .A1(n14646), .A2(n14650), .ZN(n14649) );
  NOR2_X1 U12904 ( .A1(n14900), .A2(n10579), .ZN(n14864) );
  NOR2_X1 U12905 ( .A1(n19005), .A2(n18494), .ZN(n18957) );
  AND2_X1 U12906 ( .A1(n12799), .A2(n10208), .ZN(n14853) );
  NAND3_X1 U12907 ( .A1(n10561), .A2(n10559), .A3(n10558), .ZN(n14738) );
  NAND2_X1 U12908 ( .A1(n15801), .A2(n9597), .ZN(n11173) );
  AND2_X1 U12909 ( .A1(n11534), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11549) );
  NAND2_X1 U12910 ( .A1(n11021), .A2(n10529), .ZN(n11024) );
  NAND2_X1 U12911 ( .A1(n10307), .A2(n10389), .ZN(n9636) );
  AND4_X1 U12912 ( .A1(n11841), .A2(n11840), .A3(n11839), .A4(n11838), .ZN(
        n9637) );
  INV_X1 U12913 ( .A(n10182), .ZN(n16677) );
  NAND2_X1 U12914 ( .A1(n16701), .A2(n16705), .ZN(n10182) );
  AND2_X1 U12915 ( .A1(n11023), .A2(n10115), .ZN(n9638) );
  INV_X1 U12916 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17577) );
  AND2_X1 U12917 ( .A1(n18330), .A2(n9625), .ZN(n9639) );
  NOR2_X1 U12918 ( .A1(n15023), .A2(n10468), .ZN(n9640) );
  NOR2_X1 U12919 ( .A1(n14408), .A2(n14542), .ZN(n14541) );
  AND2_X1 U12920 ( .A1(n10377), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9641) );
  NOR2_X1 U12921 ( .A1(n12465), .A2(n12464), .ZN(n12463) );
  NOR2_X1 U12922 ( .A1(n12158), .A2(n12047), .ZN(n9642) );
  INV_X1 U12923 ( .A(n10041), .ZN(n20951) );
  AND2_X1 U12924 ( .A1(n16228), .A2(n16216), .ZN(n9643) );
  AND2_X1 U12925 ( .A1(n12629), .A2(n10214), .ZN(n14626) );
  NAND2_X1 U12926 ( .A1(n15731), .A2(n15732), .ZN(n15716) );
  AND2_X1 U12927 ( .A1(n11802), .A2(n10505), .ZN(n9644) );
  OR3_X1 U12928 ( .A1(n9629), .A2(n10412), .A3(n10413), .ZN(n9645) );
  NAND2_X1 U12929 ( .A1(n11710), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16353) );
  INV_X1 U12930 ( .A(n9918), .ZN(n10739) );
  AND2_X1 U12931 ( .A1(n15731), .A2(n9623), .ZN(n9646) );
  AND2_X1 U12932 ( .A1(n14835), .A2(n10472), .ZN(n9647) );
  NAND2_X1 U12933 ( .A1(n10415), .A2(n9602), .ZN(n9648) );
  AND2_X1 U12934 ( .A1(n13118), .A2(n13117), .ZN(n9649) );
  AND2_X1 U12935 ( .A1(n18703), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9650) );
  AND2_X1 U12936 ( .A1(n10973), .A2(n9952), .ZN(n9651) );
  XOR2_X1 U12937 ( .A(n11206), .B(n11330), .Z(n9652) );
  AND2_X1 U12938 ( .A1(n15801), .A2(n9605), .ZN(n9653) );
  NOR2_X1 U12939 ( .A1(n14585), .A2(n10511), .ZN(n15783) );
  AND2_X1 U12940 ( .A1(n10557), .A2(n10556), .ZN(n9654) );
  NAND2_X1 U12941 ( .A1(n15801), .A2(n11163), .ZN(n15788) );
  XOR2_X1 U12942 ( .A(n16398), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(n9655) );
  OR2_X1 U12943 ( .A1(n11041), .A2(n11042), .ZN(n9656) );
  XNOR2_X1 U12944 ( .A(n10791), .B(n11115), .ZN(n9657) );
  NAND2_X1 U12945 ( .A1(n13760), .A2(n13718), .ZN(n9658) );
  XOR2_X1 U12946 ( .A(n17566), .B(n17565), .Z(n9659) );
  AND4_X1 U12947 ( .A1(n10872), .A2(n10871), .A3(n10870), .A4(n10869), .ZN(
        n9660) );
  AND4_X1 U12948 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n9661) );
  NOR2_X1 U12949 ( .A1(n14775), .A2(n10581), .ZN(n13712) );
  NAND2_X1 U12950 ( .A1(n10506), .A2(n11442), .ZN(n11795) );
  AND2_X1 U12951 ( .A1(n18738), .A2(n18737), .ZN(n9662) );
  OAI21_X1 U12952 ( .B1(n10338), .B2(n10546), .A(n10545), .ZN(n16392) );
  AND3_X1 U12953 ( .A1(n10865), .A2(n9977), .A3(n10863), .ZN(n9663) );
  AND2_X1 U12954 ( .A1(n12942), .A2(n10209), .ZN(n13002) );
  NAND2_X1 U12955 ( .A1(n11023), .A2(n11025), .ZN(n11041) );
  INV_X1 U12956 ( .A(n16267), .ZN(n9946) );
  INV_X1 U12957 ( .A(n11253), .ZN(n11225) );
  OR2_X1 U12958 ( .A1(n15084), .A2(n17390), .ZN(n9664) );
  OR2_X1 U12959 ( .A1(n18975), .A2(n18892), .ZN(n9665) );
  OR2_X1 U12960 ( .A1(n20006), .A2(n11062), .ZN(n9666) );
  AND2_X1 U12961 ( .A1(n9642), .A2(n12015), .ZN(n9667) );
  AND3_X1 U12962 ( .A1(n19992), .A2(n11462), .A3(n11466), .ZN(n9668) );
  AND2_X1 U12963 ( .A1(n11130), .A2(n10555), .ZN(n9669) );
  XNOR2_X1 U12964 ( .A(n10794), .B(n10795), .ZN(n10806) );
  XOR2_X1 U12965 ( .A(n16569), .B(n16585), .Z(n9670) );
  NAND2_X1 U12966 ( .A1(n15320), .A2(n12109), .ZN(n15299) );
  AND2_X2 U12967 ( .A1(n13339), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10948) );
  OR2_X1 U12968 ( .A1(n14704), .A2(n13037), .ZN(n9671) );
  INV_X1 U12969 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16902) );
  INV_X1 U12970 ( .A(n10448), .ZN(n18540) );
  AND2_X1 U12971 ( .A1(n13565), .A2(n18830), .ZN(n10448) );
  AND3_X1 U12972 ( .A1(n16331), .A2(n16345), .A3(n16342), .ZN(n9672) );
  OR2_X1 U12973 ( .A1(n15995), .A2(n15998), .ZN(n9673) );
  AND2_X1 U12974 ( .A1(n18494), .A2(n19108), .ZN(n9674) );
  AND2_X1 U12975 ( .A1(n10332), .A2(n10330), .ZN(n9675) );
  AND2_X1 U12976 ( .A1(n10890), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9676) );
  AND3_X1 U12977 ( .A1(n10387), .A2(n10386), .A3(n10383), .ZN(n9677) );
  AND3_X1 U12978 ( .A1(n10903), .A2(n10902), .A3(n10901), .ZN(n9678) );
  AND2_X1 U12979 ( .A1(n11474), .A2(n19970), .ZN(n9679) );
  NAND2_X1 U12980 ( .A1(n11033), .A2(n9956), .ZN(n11021) );
  NOR2_X1 U12981 ( .A1(n10596), .A2(n16014), .ZN(n9680) );
  AND2_X1 U12982 ( .A1(n10960), .A2(n16814), .ZN(n9681) );
  OR2_X1 U12983 ( .A1(n18493), .A2(n19709), .ZN(n9682) );
  OR2_X1 U12984 ( .A1(n13419), .A2(n13418), .ZN(n13607) );
  NAND2_X1 U12985 ( .A1(n10329), .A2(n9607), .ZN(n15258) );
  AND2_X1 U12986 ( .A1(n10493), .A2(n12221), .ZN(n9683) );
  NOR2_X1 U12987 ( .A1(n19970), .A2(n16510), .ZN(n9684) );
  AND2_X1 U12988 ( .A1(n12185), .A2(n10333), .ZN(n9685) );
  INV_X1 U12989 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10714) );
  OR2_X1 U12990 ( .A1(n19970), .A2(n16234), .ZN(n9686) );
  AND2_X1 U12991 ( .A1(n12300), .A2(n15644), .ZN(n9687) );
  AND2_X1 U12992 ( .A1(n10426), .A2(n10030), .ZN(n9688) );
  NAND2_X1 U12993 ( .A1(n13039), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9689) );
  AND3_X1 U12994 ( .A1(n16463), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16462), .ZN(n9690) );
  NOR2_X1 U12995 ( .A1(n16192), .A2(n13399), .ZN(n9691) );
  NAND2_X1 U12996 ( .A1(n15297), .A2(n12214), .ZN(n9692) );
  OR2_X1 U12997 ( .A1(n14585), .A2(n10513), .ZN(n11700) );
  NAND2_X1 U12998 ( .A1(n11021), .A2(n10530), .ZN(n9693) );
  INV_X1 U12999 ( .A(n14143), .ZN(n19127) );
  OR2_X1 U13000 ( .A1(n11573), .A2(n11572), .ZN(n14143) );
  AND2_X1 U13001 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n9694) );
  AND2_X1 U13002 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n9695) );
  NAND2_X1 U13003 ( .A1(n11772), .A2(n16501), .ZN(n9696) );
  OR2_X1 U13004 ( .A1(n11226), .A2(n11225), .ZN(n9697) );
  AND2_X1 U13005 ( .A1(n9594), .A2(n10432), .ZN(n9698) );
  OR2_X1 U13006 ( .A1(n10298), .A2(n18370), .ZN(n9699) );
  INV_X1 U13007 ( .A(n11775), .ZN(n11773) );
  NOR2_X1 U13008 ( .A1(n11767), .A2(n11768), .ZN(n11775) );
  OR2_X1 U13009 ( .A1(n10194), .A2(n10195), .ZN(n9700) );
  INV_X1 U13010 ( .A(n14800), .ZN(n12941) );
  NAND2_X1 U13011 ( .A1(n10240), .A2(n10239), .ZN(n9701) );
  INV_X1 U13012 ( .A(n10352), .ZN(n10351) );
  NOR2_X1 U13013 ( .A1(n16592), .A2(n16568), .ZN(n10352) );
  INV_X1 U13014 ( .A(n10254), .ZN(n10253) );
  NAND2_X1 U13015 ( .A1(n10585), .A2(n10584), .ZN(n10254) );
  NAND2_X1 U13016 ( .A1(n12799), .A2(n12798), .ZN(n14900) );
  NAND2_X1 U13017 ( .A1(n12998), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9702) );
  INV_X1 U13018 ( .A(n9928), .ZN(n12569) );
  AND2_X1 U13019 ( .A1(n9914), .A2(n10549), .ZN(n9703) );
  OR2_X1 U13020 ( .A1(n12217), .A2(n15544), .ZN(n15310) );
  NOR2_X1 U13021 ( .A1(n18896), .A2(n9999), .ZN(n9704) );
  AND3_X1 U13022 ( .A1(n13433), .A2(n13432), .A3(n10451), .ZN(n9705) );
  NAND2_X1 U13023 ( .A1(n10097), .A2(n17444), .ZN(n9706) );
  AND3_X1 U13024 ( .A1(n10005), .A2(n10009), .A3(n10007), .ZN(n9707) );
  AND2_X1 U13025 ( .A1(n14835), .A2(n10470), .ZN(n13657) );
  AND3_X1 U13026 ( .A1(n11751), .A2(n16261), .A3(n9964), .ZN(n9708) );
  INV_X1 U13027 ( .A(n10547), .ZN(n10546) );
  NOR2_X1 U13028 ( .A1(n19131), .A2(n19135), .ZN(n11643) );
  AND2_X1 U13029 ( .A1(n13491), .A2(n10453), .ZN(n9709) );
  INV_X1 U13030 ( .A(n9890), .ZN(n12905) );
  NOR2_X1 U13031 ( .A1(n12862), .A2(n12861), .ZN(n9890) );
  INV_X1 U13032 ( .A(n9888), .ZN(n12829) );
  NOR2_X1 U13033 ( .A1(n12813), .A2(n14903), .ZN(n9888) );
  AND3_X1 U13034 ( .A1(n13428), .A2(n13429), .A3(n13424), .ZN(n9710) );
  AND2_X1 U13035 ( .A1(n10307), .A2(n10144), .ZN(n9711) );
  INV_X1 U13036 ( .A(n14777), .ZN(n10210) );
  AND2_X1 U13037 ( .A1(n10360), .A2(n11742), .ZN(n9712) );
  AND2_X1 U13038 ( .A1(n10018), .A2(n10420), .ZN(n9713) );
  NOR2_X1 U13039 ( .A1(n10364), .A2(n11055), .ZN(n10363) );
  INV_X1 U13040 ( .A(n10363), .ZN(n10314) );
  AND3_X1 U13041 ( .A1(n11373), .A2(n11372), .A3(n11371), .ZN(n14569) );
  NOR2_X1 U13042 ( .A1(n16560), .A2(n10090), .ZN(n9714) );
  AND2_X1 U13043 ( .A1(n11462), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9715) );
  AND2_X1 U13044 ( .A1(n9914), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9716) );
  AND2_X1 U13045 ( .A1(n16387), .A2(n16399), .ZN(n9717) );
  AND2_X1 U13046 ( .A1(n9603), .A2(n10360), .ZN(n9718) );
  AND2_X1 U13047 ( .A1(n15190), .A2(n10291), .ZN(n9719) );
  AND2_X1 U13048 ( .A1(n12225), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9720) );
  AND2_X1 U13049 ( .A1(n11466), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9721) );
  AND2_X1 U13050 ( .A1(n10205), .A2(n9842), .ZN(n9722) );
  AND2_X1 U13051 ( .A1(n10554), .A2(n10553), .ZN(n9723) );
  AND2_X1 U13052 ( .A1(n10382), .A2(n17843), .ZN(n9724) );
  AND2_X1 U13053 ( .A1(n17298), .A2(n11466), .ZN(n9725) );
  AND2_X1 U13054 ( .A1(n11182), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11200) );
  INV_X1 U13055 ( .A(n11200), .ZN(n10243) );
  AND2_X1 U13056 ( .A1(n9654), .A2(n11154), .ZN(n9726) );
  AND2_X1 U13057 ( .A1(n15296), .A2(n15320), .ZN(n9727) );
  AND2_X1 U13058 ( .A1(n9641), .A2(n10376), .ZN(n9728) );
  AND2_X1 U13059 ( .A1(n13403), .A2(n10606), .ZN(n9729) );
  AND2_X1 U13060 ( .A1(n10144), .A2(n9963), .ZN(n9730) );
  INV_X1 U13061 ( .A(n10248), .ZN(n10247) );
  OAI21_X1 U13062 ( .B1(n10394), .B2(n10249), .A(n10251), .ZN(n10248) );
  OR2_X1 U13063 ( .A1(n10670), .A2(n10659), .ZN(n9731) );
  NAND2_X1 U13064 ( .A1(n11449), .A2(n9715), .ZN(n9732) );
  INV_X1 U13065 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12464) );
  NAND2_X1 U13066 ( .A1(n17101), .A2(n10444), .ZN(n10449) );
  NAND2_X1 U13067 ( .A1(n12217), .A2(n15522), .ZN(n9733) );
  AND2_X1 U13068 ( .A1(n10327), .A2(n9685), .ZN(n9734) );
  INV_X1 U13069 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18821) );
  INV_X1 U13070 ( .A(n19963), .ZN(n19946) );
  AND2_X1 U13071 ( .A1(n11114), .A2(n11232), .ZN(n16435) );
  INV_X1 U13072 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n16814) );
  NAND2_X1 U13073 ( .A1(n13637), .A2(n18694), .ZN(n10438) );
  NAND2_X1 U13074 ( .A1(n18277), .A2(n14241), .ZN(n18425) );
  INV_X1 U13075 ( .A(n18425), .ZN(n18370) );
  INV_X1 U13076 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10418) );
  INV_X1 U13077 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12518) );
  NOR2_X1 U13078 ( .A1(n15050), .A2(n15049), .ZN(n14651) );
  AND2_X1 U13079 ( .A1(n14601), .A2(n11143), .ZN(n15888) );
  NAND2_X1 U13080 ( .A1(n14576), .A2(n14575), .ZN(n14561) );
  NAND2_X1 U13081 ( .A1(n15037), .A2(n15036), .ZN(n15022) );
  AND2_X1 U13082 ( .A1(n18053), .A2(n9627), .ZN(n9735) );
  NAND2_X1 U13083 ( .A1(n11449), .A2(n11462), .ZN(n11484) );
  NAND2_X1 U13084 ( .A1(n18053), .A2(n10148), .ZN(n10151) );
  AND2_X1 U13085 ( .A1(n10567), .A2(n15732), .ZN(n9736) );
  NAND2_X1 U13086 ( .A1(n11131), .A2(n10554), .ZN(n14591) );
  AND2_X1 U13087 ( .A1(n15888), .A2(n16063), .ZN(n15874) );
  NAND2_X1 U13088 ( .A1(n12498), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11176) );
  NAND2_X1 U13089 ( .A1(n11131), .A2(n11130), .ZN(n14417) );
  AND2_X1 U13090 ( .A1(n14666), .A2(n14275), .ZN(n12243) );
  INV_X1 U13091 ( .A(n19974), .ZN(n17444) );
  OR2_X1 U13092 ( .A1(n12516), .A2(n16200), .ZN(n9737) );
  OAI21_X1 U13093 ( .B1(n14727), .B2(n19748), .A(n11261), .ZN(n14267) );
  AND2_X1 U13094 ( .A1(n10505), .A2(n15699), .ZN(n9738) );
  AND2_X1 U13095 ( .A1(n10859), .A2(n10586), .ZN(n9739) );
  AND2_X1 U13096 ( .A1(n15888), .A2(n9726), .ZN(n14614) );
  AND2_X1 U13097 ( .A1(n11131), .A2(n9669), .ZN(n14458) );
  OR2_X1 U13098 ( .A1(n15351), .A2(n15395), .ZN(n9740) );
  INV_X1 U13099 ( .A(n11025), .ZN(n10116) );
  OR2_X1 U13100 ( .A1(n10167), .A2(n13164), .ZN(n9741) );
  OR2_X1 U13101 ( .A1(n10167), .A2(n13171), .ZN(n9742) );
  OR2_X1 U13102 ( .A1(n10167), .A2(n13189), .ZN(n9743) );
  OR2_X1 U13103 ( .A1(n10167), .A2(n19996), .ZN(n9744) );
  OR2_X1 U13104 ( .A1(n10167), .A2(n20001), .ZN(n9745) );
  NAND2_X1 U13105 ( .A1(n11494), .A2(n20630), .ZN(n19974) );
  NAND2_X1 U13106 ( .A1(n15888), .A2(n9654), .ZN(n9746) );
  NOR3_X1 U13107 ( .A1(n12506), .A2(n16238), .A3(n12505), .ZN(n12508) );
  INV_X1 U13108 ( .A(n12877), .ZN(n10572) );
  INV_X1 U13109 ( .A(n11303), .ZN(n9954) );
  NAND2_X1 U13110 ( .A1(n18972), .A2(n18939), .ZN(n18956) );
  AND3_X1 U13111 ( .A1(n11758), .A2(n11756), .A3(n11754), .ZN(n9747) );
  INV_X1 U13112 ( .A(n16908), .ZN(n10135) );
  AND2_X1 U13113 ( .A1(n13560), .A2(n18625), .ZN(n9748) );
  INV_X1 U13114 ( .A(n11315), .ZN(n14576) );
  NAND2_X1 U13115 ( .A1(n15037), .A2(n9640), .ZN(n10469) );
  AND2_X1 U13116 ( .A1(n10478), .A2(n10477), .ZN(n9749) );
  AND2_X1 U13117 ( .A1(n16282), .A2(n11743), .ZN(n9750) );
  INV_X1 U13118 ( .A(n19956), .ZN(n16565) );
  NAND2_X1 U13119 ( .A1(n16902), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14157) );
  INV_X1 U13120 ( .A(n14157), .ZN(n10020) );
  AND2_X1 U13121 ( .A1(n21402), .A2(n11966), .ZN(n9751) );
  AND2_X1 U13122 ( .A1(n16177), .A2(n16176), .ZN(n9752) );
  INV_X1 U13123 ( .A(n11946), .ZN(n20832) );
  AND2_X1 U13124 ( .A1(n9740), .A2(n15390), .ZN(n9753) );
  AND2_X1 U13125 ( .A1(n9623), .A2(n15687), .ZN(n9754) );
  INV_X1 U13126 ( .A(n11444), .ZN(n11442) );
  AND2_X1 U13127 ( .A1(n10287), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9755) );
  AND4_X1 U13128 ( .A1(n16030), .A2(n16029), .A3(n16042), .A4(n16033), .ZN(
        n9756) );
  AND2_X1 U13129 ( .A1(n11001), .A2(n11002), .ZN(n11012) );
  INV_X1 U13130 ( .A(n11012), .ZN(n10532) );
  INV_X1 U13131 ( .A(n16009), .ZN(n10431) );
  AND3_X1 U13132 ( .A1(n12678), .A2(n12677), .A3(n12676), .ZN(n15035) );
  INV_X1 U13133 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15755) );
  OR2_X1 U13134 ( .A1(n15319), .A2(n12219), .ZN(n9974) );
  INV_X1 U13135 ( .A(n10474), .ZN(n10473) );
  OR2_X1 U13136 ( .A1(n10475), .A2(n14806), .ZN(n10474) );
  AND2_X1 U13137 ( .A1(n10521), .A2(n10520), .ZN(n9757) );
  NAND2_X1 U13138 ( .A1(n10709), .A2(n10737), .ZN(n9758) );
  AND2_X1 U13139 ( .A1(n12217), .A2(n10289), .ZN(n9759) );
  OR2_X1 U13140 ( .A1(n12506), .A2(n12505), .ZN(n9760) );
  INV_X1 U13141 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10287) );
  INV_X1 U13142 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12486) );
  AND2_X1 U13143 ( .A1(n12166), .A2(n12165), .ZN(n9761) );
  AND2_X1 U13144 ( .A1(n10400), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9762) );
  AND2_X1 U13145 ( .A1(n9738), .A2(n15686), .ZN(n9763) );
  NOR2_X1 U13146 ( .A1(n13185), .A2(n16022), .ZN(n9764) );
  AND2_X1 U13147 ( .A1(n10573), .A2(n10213), .ZN(n9765) );
  AND2_X1 U13148 ( .A1(n10380), .A2(n17843), .ZN(n9766) );
  AND2_X1 U13149 ( .A1(n18370), .A2(n10295), .ZN(n9767) );
  OR2_X1 U13150 ( .A1(n10670), .A2(n13135), .ZN(n9768) );
  OR2_X1 U13151 ( .A1(n10670), .A2(n13149), .ZN(n9769) );
  AND2_X1 U13152 ( .A1(n9621), .A2(n10427), .ZN(n9770) );
  AND2_X1 U13153 ( .A1(n9739), .A2(n10145), .ZN(n9771) );
  AND2_X1 U13154 ( .A1(n10859), .A2(n10587), .ZN(n9772) );
  AND2_X1 U13155 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n9773) );
  INV_X1 U13156 ( .A(n16423), .ZN(n10176) );
  NOR2_X1 U13157 ( .A1(n19594), .A2(n19582), .ZN(n19703) );
  INV_X1 U13158 ( .A(n19703), .ZN(n19588) );
  OR2_X1 U13159 ( .A1(n19728), .A2(n12535), .ZN(n19833) );
  OR2_X1 U13160 ( .A1(n13911), .A2(n11232), .ZN(n16446) );
  INV_X1 U13161 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U13162 ( .A1(n10458), .A2(n10462), .ZN(n9774) );
  INV_X1 U13163 ( .A(n18411), .ZN(n17098) );
  INV_X1 U13164 ( .A(n16446), .ZN(n16457) );
  AND4_X1 U13165 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n9775) );
  OR2_X1 U13166 ( .A1(n10167), .A2(n13221), .ZN(n9776) );
  OR2_X1 U13167 ( .A1(n10167), .A2(n13244), .ZN(n9777) );
  OR2_X1 U13168 ( .A1(n10167), .A2(n13251), .ZN(n9778) );
  OR2_X1 U13169 ( .A1(n10167), .A2(n20010), .ZN(n9779) );
  OR2_X1 U13170 ( .A1(n10167), .A2(n13280), .ZN(n9780) );
  OR2_X1 U13171 ( .A1(n10167), .A2(n20019), .ZN(n9781) );
  OR2_X1 U13172 ( .A1(n10167), .A2(n13304), .ZN(n9782) );
  AND4_X1 U13173 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(P3_EBX_REG_5__SCAN_IN), .ZN(n9783) );
  OR3_X1 U13174 ( .A1(n13552), .A2(n16991), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U13175 ( .A1(n12376), .A2(n12375), .ZN(n9785) );
  OR2_X1 U13176 ( .A1(n20006), .A2(n16006), .ZN(n9786) );
  INV_X1 U13177 ( .A(n16955), .ZN(n10447) );
  INV_X1 U13178 ( .A(n14141), .ZN(n19547) );
  NAND3_X1 U13179 ( .A1(n11172), .A2(n11171), .A3(n11170), .ZN(n9787) );
  NAND3_X1 U13180 ( .A1(n12372), .A2(n12386), .A3(n12371), .ZN(n9788) );
  OR2_X1 U13181 ( .A1(n17919), .A2(n17566), .ZN(n9789) );
  AND2_X1 U13182 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .ZN(n9790) );
  INV_X1 U13183 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12505) );
  AND3_X1 U13184 ( .A1(n10367), .A2(n10368), .A3(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17016) );
  OR2_X1 U13185 ( .A1(n10167), .A2(n13323), .ZN(n9791) );
  OR2_X1 U13186 ( .A1(n11735), .A2(n11738), .ZN(n9792) );
  NAND2_X1 U13187 ( .A1(n10366), .A2(n10368), .ZN(n17020) );
  AND2_X1 U13188 ( .A1(n10550), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9793) );
  AND3_X1 U13189 ( .A1(n18128), .A2(n18129), .A3(n10455), .ZN(n9794) );
  AND3_X1 U13190 ( .A1(n18246), .A2(n18245), .A3(n10452), .ZN(n9795) );
  INV_X1 U13191 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16725) );
  AND2_X1 U13192 ( .A1(n9626), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9796) );
  INV_X1 U13193 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16736) );
  INV_X1 U13194 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10130) );
  OR2_X1 U13195 ( .A1(n11500), .A2(n16963), .ZN(n9797) );
  OR2_X1 U13196 ( .A1(n16725), .A2(n11472), .ZN(n9798) );
  INV_X1 U13197 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16006) );
  INV_X1 U13198 ( .A(n10346), .ZN(n10345) );
  NAND2_X1 U13199 ( .A1(n9801), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10346) );
  AND3_X1 U13200 ( .A1(n15501), .A2(n15240), .A3(n15491), .ZN(n9799) );
  OR2_X1 U13201 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9800) );
  AND2_X1 U13202 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n9801) );
  INV_X1 U13203 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16568) );
  INV_X1 U13204 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10204) );
  INV_X1 U13205 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10442) );
  INV_X1 U13206 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10228) );
  INV_X1 U13207 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10149) );
  INV_X1 U13208 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10082) );
  INV_X1 U13209 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10531) );
  INV_X1 U13210 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10013) );
  INV_X1 U13211 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10324) );
  INV_X1 U13212 ( .A(n15395), .ZN(n10320) );
  INV_X1 U13213 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10273) );
  INV_X1 U13214 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n10299) );
  INV_X1 U13215 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10306) );
  INV_X1 U13216 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10539) );
  INV_X1 U13217 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10413) );
  INV_X1 U13218 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10369) );
  NAND2_X1 U13219 ( .A1(n16577), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9802) );
  OR2_X1 U13220 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n10013), .ZN(
        n9803) );
  NOR2_X2 U13221 ( .A1(n20852), .A2(n10275), .ZN(n21322) );
  OR3_X1 U13222 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20814), .A3(n21197), 
        .ZN(n20852) );
  AND4_X2 U13223 ( .A1(n10719), .A2(n10724), .A3(n11459), .A4(n11255), .ZN(
        n9942) );
  NAND2_X1 U13224 ( .A1(n10743), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9804) );
  NAND2_X1 U13225 ( .A1(n10751), .A2(n10706), .ZN(n9805) );
  NAND3_X1 U13226 ( .A1(n9877), .A2(n9876), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9810) );
  NAND2_X1 U13227 ( .A1(n10747), .A2(n10635), .ZN(n9811) );
  AND2_X1 U13228 ( .A1(n9815), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9813) );
  NAND2_X1 U13229 ( .A1(n9814), .A2(n11011), .ZN(n16418) );
  AND2_X1 U13230 ( .A1(n10809), .A2(n16733), .ZN(n20197) );
  NOR2_X1 U13231 ( .A1(n17298), .A2(n9824), .ZN(n9823) );
  NAND2_X1 U13232 ( .A1(n9829), .A2(n10714), .ZN(n9828) );
  NAND4_X1 U13233 ( .A1(n10710), .A2(n10712), .A3(n10711), .A4(n10713), .ZN(
        n9829) );
  NAND2_X1 U13234 ( .A1(n9831), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9830) );
  NAND4_X1 U13235 ( .A1(n10715), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n9831) );
  AND2_X2 U13236 ( .A1(n11975), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10197) );
  INV_X1 U13237 ( .A(n10197), .ZN(n11996) );
  AND2_X2 U13238 ( .A1(n10166), .A2(n10587), .ZN(n10987) );
  NAND2_X2 U13239 ( .A1(n9833), .A2(n9663), .ZN(n10166) );
  AND2_X1 U13240 ( .A1(n9834), .A2(n13730), .ZN(n10099) );
  NAND2_X1 U13241 ( .A1(n16191), .A2(n9834), .ZN(n16469) );
  NAND2_X2 U13242 ( .A1(n9595), .A2(n10332), .ZN(n10329) );
  NAND3_X1 U13243 ( .A1(n9595), .A2(n12224), .A3(n10332), .ZN(n10199) );
  NAND2_X2 U13244 ( .A1(n10612), .A2(n10611), .ZN(n11946) );
  NAND2_X1 U13245 ( .A1(n10275), .A2(n20832), .ZN(n11958) );
  AND3_X1 U13246 ( .A1(n12583), .A2(n9734), .A3(n9866), .ZN(n9960) );
  NAND3_X1 U13247 ( .A1(n13714), .A2(n9740), .A3(n10322), .ZN(n10278) );
  NAND4_X1 U13248 ( .A1(n9921), .A2(n9919), .A3(n9920), .A4(n9835), .ZN(n9918)
         );
  NAND2_X1 U13249 ( .A1(n10689), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9835) );
  INV_X1 U13250 ( .A(n11182), .ZN(n10050) );
  NOR2_X2 U13251 ( .A1(n10803), .A2(n19943), .ZN(n16819) );
  NAND2_X1 U13252 ( .A1(n10205), .A2(n9839), .ZN(n10089) );
  INV_X1 U13253 ( .A(n9840), .ZN(n9839) );
  NAND3_X1 U13254 ( .A1(n20015), .A2(n13361), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9840) );
  NAND3_X1 U13255 ( .A1(n10205), .A2(n9842), .A3(n11462), .ZN(n9841) );
  NAND2_X1 U13256 ( .A1(n9913), .A2(n9716), .ZN(n16216) );
  AND2_X2 U13257 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11107) );
  INV_X2 U13258 ( .A(n13139), .ZN(n13327) );
  AND2_X2 U13259 ( .A1(n13327), .A2(n10714), .ZN(n10847) );
  NAND3_X1 U13260 ( .A1(n10875), .A2(n10874), .A3(n9859), .ZN(n9858) );
  AND2_X1 U13261 ( .A1(n12583), .A2(n9866), .ZN(n12582) );
  OR2_X1 U13262 ( .A1(n12583), .A2(n9866), .ZN(n12584) );
  NAND2_X1 U13263 ( .A1(n9867), .A2(n10496), .ZN(n10495) );
  NAND2_X1 U13264 ( .A1(n9867), .A2(n17378), .ZN(n10499) );
  XNOR2_X1 U13265 ( .A(n9867), .B(n10036), .ZN(n17430) );
  NAND2_X2 U13266 ( .A1(n9922), .A2(n12184), .ZN(n9867) );
  XNOR2_X1 U13267 ( .A(n12155), .B(n12154), .ZN(n14190) );
  NAND2_X1 U13268 ( .A1(n9873), .A2(n10243), .ZN(n9875) );
  NAND2_X1 U13269 ( .A1(n10034), .A2(n10032), .ZN(n9873) );
  NAND3_X1 U13270 ( .A1(n9875), .A2(n11199), .A3(n9874), .ZN(n9975) );
  NAND3_X1 U13271 ( .A1(n16419), .A2(n16420), .A3(n10255), .ZN(n9874) );
  NAND2_X2 U13272 ( .A1(n10047), .A2(n11197), .ZN(n16419) );
  NAND2_X2 U13273 ( .A1(n10818), .A2(n19943), .ZN(n20344) );
  NAND2_X1 U13274 ( .A1(n10206), .A2(n9881), .ZN(n11206) );
  NAND2_X2 U13275 ( .A1(n10782), .A2(n10238), .ZN(n10785) );
  AND3_X2 U13276 ( .A1(n9884), .A2(n9883), .A3(n9882), .ZN(n10782) );
  NAND3_X1 U13277 ( .A1(n10727), .A2(n17298), .A3(n9721), .ZN(n9882) );
  NAND2_X1 U13278 ( .A1(n10777), .A2(n11466), .ZN(n9883) );
  NAND2_X1 U13279 ( .A1(n10237), .A2(n10709), .ZN(n9884) );
  NOR2_X2 U13280 ( .A1(n14681), .A2(n14679), .ZN(n9887) );
  INV_X2 U13281 ( .A(n11118), .ZN(n13774) );
  INV_X2 U13282 ( .A(n10737), .ZN(n9894) );
  NAND2_X1 U13283 ( .A1(n10785), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9895) );
  NAND3_X1 U13284 ( .A1(n10767), .A2(n10766), .A3(n10768), .ZN(n9898) );
  NAND3_X1 U13285 ( .A1(n9732), .A2(n9612), .A3(n9897), .ZN(n10589) );
  NAND3_X1 U13286 ( .A1(n10141), .A2(n10140), .A3(n10797), .ZN(n10138) );
  NAND2_X1 U13287 ( .A1(n9899), .A2(n19946), .ZN(n11708) );
  AOI21_X1 U13288 ( .B1(n9899), .B2(n16457), .A(n16277), .ZN(n16278) );
  AND2_X1 U13289 ( .A1(n16280), .A2(n11707), .ZN(n9900) );
  NAND3_X1 U13290 ( .A1(n10046), .A2(n10084), .A3(n9901), .ZN(n9903) );
  AND2_X4 U13291 ( .A1(n9905), .A2(n10958), .ZN(n13336) );
  AND2_X1 U13292 ( .A1(n13133), .A2(n9905), .ZN(n13119) );
  NAND4_X1 U13293 ( .A1(n10616), .A2(n10614), .A3(n10615), .A4(n9909), .ZN(
        n9908) );
  NAND4_X1 U13294 ( .A1(n10619), .A2(n9911), .A3(n10618), .A4(n10620), .ZN(
        n9910) );
  NAND3_X1 U13295 ( .A1(n13404), .A2(n13405), .A3(n9729), .ZN(P2_U3016) );
  NAND2_X1 U13296 ( .A1(n10146), .A2(n10145), .ZN(n9915) );
  NAND4_X2 U13297 ( .A1(n9707), .A2(n10001), .A3(n10003), .A4(n10008), .ZN(
        n10341) );
  AND3_X2 U13298 ( .A1(n10166), .A2(n9739), .A3(n10341), .ZN(n9916) );
  NAND3_X1 U13299 ( .A1(n10486), .A2(n14526), .A3(n10485), .ZN(n9922) );
  NAND2_X1 U13300 ( .A1(n12174), .A2(n14471), .ZN(n10485) );
  NAND2_X1 U13301 ( .A1(n9923), .A2(n13976), .ZN(n9924) );
  NAND2_X1 U13302 ( .A1(n9924), .A2(n9925), .ZN(n9927) );
  NAND2_X2 U13303 ( .A1(n10283), .A2(n10568), .ZN(n12167) );
  NAND2_X2 U13304 ( .A1(n9927), .A2(n9926), .ZN(n10568) );
  NAND3_X1 U13305 ( .A1(n13976), .A2(n10282), .A3(n12000), .ZN(n9926) );
  NAND2_X1 U13306 ( .A1(n15231), .A2(n9929), .ZN(n9928) );
  NAND2_X2 U13307 ( .A1(n15241), .A2(n15190), .ZN(n15231) );
  NAND3_X1 U13308 ( .A1(n13560), .A2(n18625), .A3(n18854), .ZN(n18570) );
  NAND3_X1 U13309 ( .A1(n18577), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n18570), .ZN(n13561) );
  NAND3_X1 U13310 ( .A1(n9932), .A2(n18728), .A3(n9930), .ZN(n16922) );
  NAND2_X1 U13311 ( .A1(n16925), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16924) );
  NAND3_X1 U13312 ( .A1(n10449), .A2(n13642), .A3(n9580), .ZN(n9936) );
  INV_X1 U13313 ( .A(n13567), .ZN(n9937) );
  NAND2_X1 U13314 ( .A1(n13540), .A2(n13539), .ZN(n13541) );
  XNOR2_X1 U13315 ( .A(n13540), .B(n13538), .ZN(n18760) );
  INV_X1 U13316 ( .A(n9939), .ZN(n9938) );
  NAND2_X1 U13317 ( .A1(n10067), .A2(n18751), .ZN(n10066) );
  INV_X1 U13318 ( .A(n10794), .ZN(n10052) );
  NAND2_X1 U13319 ( .A1(n10722), .A2(n9942), .ZN(n11099) );
  NOR2_X4 U13320 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11830) );
  NAND3_X1 U13321 ( .A1(n12309), .A2(n11946), .A3(n11950), .ZN(n11947) );
  OAI21_X1 U13322 ( .B1(n13853), .B2(n14119), .A(n11946), .ZN(n12316) );
  NOR2_X1 U13323 ( .A1(n13969), .A2(n11946), .ZN(n13970) );
  MUX2_X1 U13324 ( .A(n11962), .B(n12309), .S(n11946), .Z(n11965) );
  NAND3_X1 U13325 ( .A1(n9944), .A2(n9943), .A3(n16457), .ZN(n9951) );
  NAND2_X1 U13326 ( .A1(n9951), .A2(n9948), .ZN(P2_U2990) );
  NAND2_X1 U13327 ( .A1(n9719), .A2(n15241), .ZN(n9955) );
  INV_X1 U13328 ( .A(n15231), .ZN(n12227) );
  NAND2_X1 U13329 ( .A1(n9957), .A2(n15902), .ZN(n9956) );
  NAND4_X1 U13330 ( .A1(n10056), .A2(n10917), .A3(n10918), .A4(n9958), .ZN(
        n10055) );
  NAND2_X4 U13331 ( .A1(n12198), .A2(n12106), .ZN(n12217) );
  NAND2_X1 U13332 ( .A1(n10310), .A2(n9614), .ZN(n9965) );
  INV_X1 U13333 ( .A(n11015), .ZN(n16384) );
  NAND2_X1 U13334 ( .A1(n15351), .A2(n9800), .ZN(n10493) );
  NAND2_X1 U13335 ( .A1(n9967), .A2(n11224), .ZN(n9966) );
  NAND2_X1 U13336 ( .A1(n10172), .A2(n10170), .ZN(n9967) );
  AOI211_X2 U13337 ( .C1(n16465), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n9690), .B(n9968), .ZN(n16467) );
  NAND2_X2 U13339 ( .A1(n10315), .A2(n11999), .ZN(n13976) );
  AND2_X2 U13340 ( .A1(n9970), .A2(n12149), .ZN(n12133) );
  NAND2_X1 U13341 ( .A1(n9720), .A2(n9971), .ZN(n15192) );
  INV_X1 U13342 ( .A(n9974), .ZN(n9973) );
  OAI21_X1 U13343 ( .B1(n9975), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10046), .ZN(n16711) );
  INV_X1 U13344 ( .A(n9976), .ZN(n10734) );
  NAND3_X1 U13345 ( .A1(n12281), .A2(n9986), .A3(n9985), .ZN(n9984) );
  NAND3_X1 U13346 ( .A1(n12308), .A2(n9988), .A3(n9610), .ZN(n9987) );
  OR2_X1 U13347 ( .A1(n12307), .A2(n20832), .ZN(n9988) );
  NAND2_X1 U13348 ( .A1(n16216), .A2(n16217), .ZN(n9989) );
  INV_X2 U13349 ( .A(n11955), .ZN(n14119) );
  NAND3_X1 U13350 ( .A1(n9992), .A2(n9991), .A3(n9990), .ZN(n13611) );
  NAND2_X1 U13351 ( .A1(n13607), .A2(n14206), .ZN(n9990) );
  NAND3_X1 U13352 ( .A1(n14243), .A2(n14215), .A3(n13609), .ZN(n9991) );
  NAND2_X1 U13353 ( .A1(n9993), .A2(n13607), .ZN(n9992) );
  NOR2_X2 U13354 ( .A1(n18956), .A2(n10226), .ZN(n18937) );
  INV_X1 U13355 ( .A(n10183), .ZN(n10002) );
  NAND2_X1 U13356 ( .A1(n16267), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10014) );
  NAND4_X1 U13357 ( .A1(n10420), .A2(n9671), .A3(n10019), .A4(n10018), .ZN(
        n10419) );
  NAND3_X1 U13358 ( .A1(n10027), .A2(n10025), .A3(n10024), .ZN(n10022) );
  NAND2_X1 U13359 ( .A1(n13118), .A2(n9764), .ZN(n10024) );
  NAND2_X1 U13360 ( .A1(n9649), .A2(n10028), .ZN(n10023) );
  NAND3_X1 U13361 ( .A1(n10027), .A2(n10029), .A3(n10024), .ZN(n16016) );
  NAND2_X1 U13362 ( .A1(n10033), .A2(n11202), .ZN(n10032) );
  INV_X1 U13363 ( .A(n16420), .ZN(n10033) );
  NAND3_X1 U13364 ( .A1(n10047), .A2(n11202), .A3(n11197), .ZN(n10034) );
  NAND3_X1 U13365 ( .A1(n12166), .A2(n12165), .A3(n10037), .ZN(n10486) );
  NAND2_X1 U13366 ( .A1(n14463), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10037) );
  NAND2_X1 U13367 ( .A1(n10329), .A2(n10038), .ZN(n10039) );
  NAND2_X1 U13368 ( .A1(n10039), .A2(n15351), .ZN(n15241) );
  NAND2_X1 U13369 ( .A1(n15231), .A2(n15425), .ZN(n12225) );
  INV_X1 U13370 ( .A(n12167), .ZN(n10040) );
  XNOR2_X2 U13371 ( .A(n10041), .B(n12167), .ZN(n12581) );
  OAI21_X1 U13372 ( .B1(n16549), .B2(n19974), .A(n10042), .ZN(P2_U3025) );
  INV_X1 U13373 ( .A(n10043), .ZN(n10042) );
  INV_X1 U13374 ( .A(n16429), .ZN(n10049) );
  NAND2_X1 U13375 ( .A1(n10048), .A2(n16431), .ZN(n10047) );
  NAND2_X1 U13376 ( .A1(n10049), .A2(n16725), .ZN(n10048) );
  NAND2_X1 U13377 ( .A1(n11710), .A2(n16538), .ZN(n10051) );
  NAND2_X1 U13378 ( .A1(n10052), .A2(n10795), .ZN(n10551) );
  NAND2_X1 U13379 ( .A1(n11711), .A2(n10550), .ZN(n10059) );
  XNOR2_X1 U13380 ( .A(n11979), .B(n11990), .ZN(n12016) );
  INV_X1 U13381 ( .A(n12016), .ZN(n20919) );
  NAND2_X1 U13382 ( .A1(n12018), .A2(n20919), .ZN(n20860) );
  AND2_X1 U13383 ( .A1(n10568), .A2(n10327), .ZN(n10063) );
  AND3_X2 U13384 ( .A1(n10064), .A2(n12582), .A3(n10063), .ZN(n12186) );
  INV_X1 U13385 ( .A(n12198), .ZN(n12207) );
  OAI211_X1 U13386 ( .C1(n18751), .C2(n10074), .A(n10071), .B(n10070), .ZN(
        n18741) );
  AND2_X1 U13387 ( .A1(n10077), .A2(n10075), .ZN(n16957) );
  NAND2_X1 U13388 ( .A1(n10079), .A2(n10078), .ZN(n10077) );
  NOR2_X1 U13389 ( .A1(n18541), .A2(n17108), .ZN(n10078) );
  NAND2_X1 U13390 ( .A1(n11203), .A2(n11202), .ZN(n10084) );
  INV_X1 U13391 ( .A(n11201), .ZN(n16422) );
  NAND2_X1 U13392 ( .A1(n16419), .A2(n16420), .ZN(n11201) );
  NAND4_X1 U13393 ( .A1(n10684), .A2(n10682), .A3(n10681), .A4(n10683), .ZN(
        n10751) );
  NAND4_X1 U13394 ( .A1(n10677), .A2(n10680), .A3(n10679), .A4(n10678), .ZN(
        n10743) );
  INV_X1 U13395 ( .A(n10551), .ZN(n10088) );
  OAI21_X2 U13396 ( .B1(n11461), .B2(n16902), .A(n10089), .ZN(n10777) );
  OR2_X1 U13397 ( .A1(n16551), .A2(n19963), .ZN(n10091) );
  NAND2_X2 U13398 ( .A1(n10092), .A2(n10809), .ZN(n20463) );
  INV_X4 U13399 ( .A(n10670), .ZN(n13334) );
  NAND4_X1 U13400 ( .A1(n9651), .A2(n11001), .A3(n11002), .A4(n10980), .ZN(
        n10978) );
  INV_X1 U13401 ( .A(n10244), .ZN(n10102) );
  NAND3_X1 U13402 ( .A1(n10105), .A2(n13718), .A3(n10101), .ZN(n13763) );
  NAND3_X1 U13403 ( .A1(n10105), .A2(n10103), .A3(n10101), .ZN(n10110) );
  AOI21_X2 U13404 ( .B1(n17157), .B2(n13629), .A(n13628), .ZN(n14398) );
  NOR2_X2 U13405 ( .A1(n10120), .A2(n10119), .ZN(n17157) );
  NAND3_X1 U13406 ( .A1(n19108), .A2(n19122), .A3(n10124), .ZN(n10123) );
  NAND3_X1 U13407 ( .A1(n11582), .A2(n11583), .A3(n10128), .ZN(n10127) );
  INV_X1 U13408 ( .A(n10131), .ZN(n17547) );
  NAND2_X1 U13409 ( .A1(n10769), .A2(n10794), .ZN(n10141) );
  NAND4_X1 U13410 ( .A1(n10146), .A2(n10341), .A3(n9771), .A4(n10166), .ZN(
        n10938) );
  INV_X1 U13411 ( .A(n10151), .ZN(n18005) );
  NAND3_X1 U13412 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_18__SCAN_IN), 
        .A3(P3_EBX_REG_17__SCAN_IN), .ZN(n10154) );
  INV_X1 U13413 ( .A(n18071), .ZN(n18103) );
  XNOR2_X2 U13414 ( .A(n10987), .B(n10986), .ZN(n10165) );
  NAND2_X1 U13415 ( .A1(n10165), .A2(n16449), .ZN(n11196) );
  NAND2_X1 U13416 ( .A1(n10165), .A2(n13768), .ZN(n10196) );
  XNOR2_X1 U13417 ( .A(n10165), .B(n10164), .ZN(n16740) );
  AND3_X1 U13418 ( .A1(n10341), .A2(n9772), .A3(n10166), .ZN(n11184) );
  CLKBUF_X1 U13419 ( .A(n10670), .Z(n10167) );
  MUX2_X1 U13420 ( .A(n11255), .B(n20015), .S(n11459), .Z(n10721) );
  NAND3_X1 U13421 ( .A1(n10173), .A2(n11221), .A3(n11220), .ZN(n10172) );
  NAND3_X1 U13422 ( .A1(n11216), .A2(n11215), .A3(n11466), .ZN(n10173) );
  NAND2_X1 U13423 ( .A1(n16677), .A2(n10179), .ZN(n16474) );
  NAND2_X1 U13424 ( .A1(n16733), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10186) );
  OAI211_X1 U13425 ( .C1(n20463), .C2(n10190), .A(n10185), .B(n10184), .ZN(
        n10183) );
  NAND2_X1 U13426 ( .A1(n10189), .A2(n10810), .ZN(n10185) );
  NAND2_X1 U13427 ( .A1(n10187), .A2(n10186), .ZN(n10189) );
  INV_X1 U13428 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U13429 ( .A1(n16225), .A2(n10193), .ZN(n10192) );
  NAND2_X1 U13430 ( .A1(n10197), .A2(n15642), .ZN(n12045) );
  NAND2_X1 U13431 ( .A1(n12137), .A2(n12136), .ZN(n12155) );
  NAND2_X1 U13432 ( .A1(n14107), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12154) );
  AND2_X2 U13433 ( .A1(n10199), .A2(n10198), .ZN(n15190) );
  NAND2_X2 U13434 ( .A1(n10292), .A2(n12215), .ZN(n10332) );
  NAND2_X1 U13435 ( .A1(n20921), .A2(n10287), .ZN(n12148) );
  XNOR2_X2 U13436 ( .A(n12035), .B(n9630), .ZN(n20921) );
  NAND3_X1 U13437 ( .A1(n12148), .A2(n12147), .A3(n12243), .ZN(n12153) );
  NOR2_X2 U13438 ( .A1(n10204), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16746) );
  XNOR2_X2 U13439 ( .A(n10590), .B(n9657), .ZN(n10805) );
  NAND2_X1 U13440 ( .A1(n13976), .A2(n12000), .ZN(n14078) );
  NAND2_X1 U13441 ( .A1(n12799), .A2(n10207), .ZN(n14841) );
  NAND2_X1 U13442 ( .A1(n12942), .A2(n10211), .ZN(n14775) );
  NAND2_X1 U13443 ( .A1(n12942), .A2(n12941), .ZN(n14787) );
  NAND2_X1 U13444 ( .A1(n15387), .A2(n17382), .ZN(n13717) );
  NAND2_X1 U13445 ( .A1(n14480), .A2(n10287), .ZN(n10325) );
  INV_X1 U13446 ( .A(n10280), .ZN(n10279) );
  AOI21_X1 U13447 ( .B1(n9594), .B2(n9615), .A(n9773), .ZN(n10540) );
  NAND2_X1 U13448 ( .A1(n14927), .A2(n14929), .ZN(n14911) );
  NAND2_X1 U13449 ( .A1(n10279), .A2(n10276), .ZN(P1_U2970) );
  INV_X1 U13450 ( .A(n12582), .ZN(n12585) );
  NOR2_X1 U13451 ( .A1(n14409), .A2(n12600), .ZN(n12607) );
  INV_X1 U13452 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10220) );
  INV_X1 U13453 ( .A(n18956), .ZN(n10223) );
  NAND2_X1 U13454 ( .A1(n10223), .A2(n10224), .ZN(n18845) );
  NAND3_X1 U13455 ( .A1(n9841), .A2(n10764), .A3(n10236), .ZN(n10238) );
  NAND3_X1 U13456 ( .A1(n11239), .A2(n10730), .A3(n10724), .ZN(n10236) );
  NAND2_X1 U13457 ( .A1(n10271), .A2(n13541), .ZN(n18749) );
  NAND2_X1 U13458 ( .A1(n18760), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10271) );
  NAND2_X1 U13459 ( .A1(n13541), .A2(n10273), .ZN(n10272) );
  AND2_X2 U13460 ( .A1(n11535), .A2(n11533), .ZN(n11604) );
  NAND2_X1 U13461 ( .A1(n10275), .A2(n13810), .ZN(n12362) );
  AND3_X1 U13462 ( .A1(n11830), .A2(n14087), .A3(
        P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U13463 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11931), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U13464 ( .A1(n20860), .A2(n12019), .ZN(n14478) );
  INV_X1 U13465 ( .A(n12601), .ZN(n10491) );
  NOR2_X1 U13466 ( .A1(n18308), .A2(n10299), .ZN(n10298) );
  NOR2_X1 U13467 ( .A1(n10294), .A2(n9767), .ZN(n18295) );
  INV_X1 U13468 ( .A(n18308), .ZN(n18303) );
  INV_X1 U13469 ( .A(n10298), .ZN(n18302) );
  OAI22_X1 U13470 ( .A1(n10450), .A2(n11606), .B1(n17226), .B2(n10303), .ZN(
        n11609) );
  OAI22_X1 U13471 ( .A1(n10450), .A2(n17220), .B1(n17221), .B2(n10303), .ZN(
        n17223) );
  OAI22_X1 U13472 ( .A1(n10450), .A2(n17206), .B1(n17207), .B2(n10303), .ZN(
        n17211) );
  OAI22_X1 U13473 ( .A1(n10450), .A2(n18201), .B1(n17233), .B2(n10303), .ZN(
        n17236) );
  OAI22_X1 U13474 ( .A1(n10450), .A2(n17246), .B1(n17247), .B2(n10303), .ZN(
        n17251) );
  OAI22_X1 U13475 ( .A1(n10450), .A2(n17262), .B1(n17263), .B2(n10303), .ZN(
        n17266) );
  OAI22_X1 U13476 ( .A1(n10450), .A2(n17950), .B1(n17951), .B2(n10303), .ZN(
        n17953) );
  OAI22_X1 U13477 ( .A1(n10450), .A2(n18010), .B1(n18011), .B2(n10303), .ZN(
        n18015) );
  OAI22_X1 U13478 ( .A1(n10450), .A2(n18021), .B1(n18022), .B2(n10303), .ZN(
        n18026) );
  OAI22_X1 U13479 ( .A1(n10450), .A2(n18106), .B1(n18107), .B2(n10303), .ZN(
        n18110) );
  OAI22_X1 U13480 ( .A1(n10450), .A2(n18138), .B1(n18139), .B2(n10303), .ZN(
        n18143) );
  OAI22_X1 U13481 ( .A1(n10450), .A2(n18076), .B1(n18077), .B2(n10303), .ZN(
        n18081) );
  NAND2_X1 U13482 ( .A1(n9730), .A2(n10307), .ZN(n10390) );
  NAND2_X1 U13483 ( .A1(n16290), .A2(n10308), .ZN(P2_U2996) );
  NAND3_X1 U13484 ( .A1(n11204), .A2(n13768), .A3(n10311), .ZN(n10310) );
  NAND2_X1 U13485 ( .A1(n11045), .A2(n9718), .ZN(n10312) );
  NAND2_X1 U13486 ( .A1(n10312), .A2(n10313), .ZN(n11688) );
  NAND2_X1 U13487 ( .A1(n12019), .A2(n11995), .ZN(n10315) );
  NAND2_X1 U13488 ( .A1(n12019), .A2(n10316), .ZN(n12000) );
  NAND3_X1 U13489 ( .A1(n12228), .A2(n15201), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U13490 ( .A1(n12186), .A2(n12185), .ZN(n12194) );
  NAND2_X1 U13491 ( .A1(n10341), .A2(n10859), .ZN(n10986) );
  NAND2_X1 U13492 ( .A1(n16324), .A2(n10363), .ZN(n10356) );
  INV_X1 U13493 ( .A(n9594), .ZN(n11470) );
  NAND2_X1 U13494 ( .A1(n17017), .A2(n17016), .ZN(n17783) );
  OAI21_X1 U13495 ( .B1(n11515), .B2(n11514), .A(n19598), .ZN(n10370) );
  NAND2_X1 U13496 ( .A1(n10371), .A2(n17843), .ZN(n11515) );
  INV_X1 U13497 ( .A(n10374), .ZN(n17587) );
  INV_X1 U13498 ( .A(n11523), .ZN(n17575) );
  NAND2_X1 U13499 ( .A1(n10379), .A2(n10380), .ZN(n17609) );
  OR2_X2 U13500 ( .A1(n17617), .A2(n10381), .ZN(n10379) );
  INV_X1 U13501 ( .A(n10382), .ZN(n17616) );
  NAND2_X1 U13502 ( .A1(n10399), .A2(n10397), .ZN(n12471) );
  NAND3_X1 U13503 ( .A1(n10399), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12469) );
  NAND3_X1 U13504 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10402) );
  INV_X1 U13505 ( .A(n10403), .ZN(n13781) );
  NAND2_X1 U13506 ( .A1(n10419), .A2(n10420), .ZN(n14235) );
  NAND2_X1 U13507 ( .A1(n10422), .A2(n10421), .ZN(n15980) );
  NAND3_X1 U13508 ( .A1(n10428), .A2(n13269), .A3(n9770), .ZN(n10421) );
  NAND2_X1 U13509 ( .A1(n13292), .A2(n9621), .ZN(n10422) );
  NAND2_X1 U13510 ( .A1(n13269), .A2(n10427), .ZN(n10423) );
  NAND2_X1 U13511 ( .A1(n10428), .A2(n13269), .ZN(n15991) );
  INV_X2 U13513 ( .A(n13024), .ZN(n16768) );
  XNOR2_X2 U13514 ( .A(n10802), .B(n10801), .ZN(n13024) );
  NAND3_X1 U13515 ( .A1(n10438), .A2(n13551), .A3(n17047), .ZN(n13553) );
  NAND2_X1 U13516 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11552) );
  NAND2_X1 U13517 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11590) );
  NAND2_X1 U13518 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13466) );
  NAND2_X1 U13519 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13482) );
  NAND2_X1 U13520 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10451) );
  NAND2_X1 U13521 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10452) );
  NAND2_X1 U13522 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10454) );
  NAND2_X1 U13523 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10455) );
  AND2_X4 U13524 ( .A1(n11534), .A2(n14407), .ZN(n18223) );
  NAND2_X1 U13525 ( .A1(n10456), .A2(n12360), .ZN(n14255) );
  XNOR2_X1 U13526 ( .A(n10457), .B(n14187), .ZN(n14193) );
  OAI21_X1 U13527 ( .B1(n15079), .B2(n10457), .A(n15072), .ZN(n15077) );
  NAND2_X1 U13528 ( .A1(n12369), .A2(n12368), .ZN(n14447) );
  INV_X1 U13529 ( .A(n14447), .ZN(n10459) );
  NAND3_X1 U13530 ( .A1(n10460), .A2(n10459), .A3(n10462), .ZN(n14555) );
  XNOR2_X1 U13531 ( .A(n10484), .B(n10483), .ZN(n14546) );
  INV_X1 U13532 ( .A(n14526), .ZN(n10483) );
  NAND2_X1 U13533 ( .A1(n10495), .A2(n10494), .ZN(n15292) );
  AOI21_X1 U13534 ( .B1(n10498), .B2(n17372), .A(n10497), .ZN(n10494) );
  NAND2_X1 U13535 ( .A1(n14442), .A2(n10500), .ZN(n15937) );
  NAND2_X2 U13536 ( .A1(n14440), .A2(n14439), .ZN(n14442) );
  NAND2_X1 U13537 ( .A1(n11802), .A2(n9763), .ZN(n11811) );
  INV_X1 U13538 ( .A(n11441), .ZN(n10506) );
  NAND2_X1 U13539 ( .A1(n10506), .A2(n10507), .ZN(n15728) );
  NAND2_X1 U13540 ( .A1(n13390), .A2(n10962), .ZN(n10519) );
  NAND2_X1 U13541 ( .A1(n13390), .A2(n10961), .ZN(n10520) );
  NAND2_X1 U13542 ( .A1(n11086), .A2(n20006), .ZN(n10521) );
  NOR2_X1 U13543 ( .A1(n20006), .A2(n10523), .ZN(n10522) );
  NAND2_X1 U13544 ( .A1(n11272), .A2(n20006), .ZN(n10525) );
  NAND2_X1 U13545 ( .A1(n11117), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10541) );
  NAND2_X1 U13546 ( .A1(n10798), .A2(n10551), .ZN(n10802) );
  AND2_X1 U13547 ( .A1(n12554), .A2(n10564), .ZN(n13773) );
  NAND2_X1 U13548 ( .A1(n12554), .A2(n10560), .ZN(n10559) );
  NAND2_X1 U13549 ( .A1(n12554), .A2(n12553), .ZN(n12560) );
  OR2_X1 U13550 ( .A1(n12554), .A2(n10562), .ZN(n10561) );
  NAND2_X1 U13551 ( .A1(n12878), .A2(n10570), .ZN(n14797) );
  INV_X1 U13552 ( .A(n14797), .ZN(n12942) );
  NOR2_X1 U13553 ( .A1(n14775), .A2(n10583), .ZN(n13685) );
  INV_X1 U13554 ( .A(n16244), .ZN(n10585) );
  AOI21_X1 U13555 ( .B1(n16251), .B2(n16253), .A(n11766), .ZN(n16243) );
  OR2_X1 U13556 ( .A1(n10589), .A2(n10792), .ZN(n10793) );
  NOR2_X1 U13557 ( .A1(n10590), .A2(n11116), .ZN(n16437) );
  NAND2_X1 U13558 ( .A1(n10807), .A2(n17445), .ZN(n10814) );
  NAND2_X1 U13559 ( .A1(n13266), .A2(n13265), .ZN(n13269) );
  NAND2_X1 U13560 ( .A1(n13240), .A2(n9673), .ZN(n13266) );
  INV_X1 U13561 ( .A(n15801), .ZN(n15821) );
  AND2_X1 U13562 ( .A1(n14238), .A2(n14237), .ZN(n20610) );
  OAI211_X1 U13563 ( .C1(n16469), .C2(n19963), .A(n16468), .B(n16467), .ZN(
        n16470) );
  INV_X1 U13564 ( .A(n13685), .ZN(n13007) );
  NAND2_X1 U13565 ( .A1(n14629), .A2(n10597), .ZN(n15050) );
  NAND2_X2 U13566 ( .A1(n12560), .A2(n15667), .ZN(n16466) );
  NAND2_X1 U13567 ( .A1(n12217), .A2(n12129), .ZN(n15379) );
  XNOR2_X1 U13568 ( .A(n12217), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15330) );
  INV_X1 U13569 ( .A(n15392), .ZN(n14677) );
  OAI21_X1 U13570 ( .B1(n15084), .B2(n15079), .A(n13818), .ZN(n13819) );
  NAND2_X1 U13571 ( .A1(n11792), .A2(n17444), .ZN(n11816) );
  INV_X1 U13572 ( .A(n14255), .ZN(n12369) );
  NOR2_X2 U13573 ( .A1(n16280), .A2(n11707), .ZN(n11706) );
  INV_X1 U13574 ( .A(n16211), .ZN(n11792) );
  NAND2_X1 U13575 ( .A1(n13758), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13759) );
  AOI21_X1 U13576 ( .B1(n13825), .B2(n17382), .A(n13824), .ZN(n13826) );
  NAND2_X1 U13577 ( .A1(n16190), .A2(n19946), .ZN(n13731) );
  CLKBUF_X1 U13578 ( .A(n16385), .Z(n16411) );
  AOI21_X1 U13579 ( .B1(n16069), .B2(n19960), .A(n14739), .ZN(n14742) );
  INV_X1 U13580 ( .A(n11549), .ZN(n14659) );
  NOR2_X1 U13581 ( .A1(n21191), .A2(n21156), .ZN(n10593) );
  NOR2_X1 U13582 ( .A1(n13378), .A2(n10604), .ZN(n10594) );
  AND2_X1 U13583 ( .A1(n12206), .A2(n12205), .ZN(n10595) );
  AND2_X1 U13584 ( .A1(n14635), .A2(n14628), .ZN(n10597) );
  OR2_X1 U13585 ( .A1(n18917), .A2(n18912), .ZN(n18668) );
  OR2_X1 U13586 ( .A1(n16193), .A2(n16212), .ZN(n10598) );
  INV_X1 U13587 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12468) );
  AND2_X2 U13588 ( .A1(n13849), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20812)
         );
  OR2_X1 U13589 ( .A1(n16195), .A2(n16194), .ZN(n10599) );
  AND2_X1 U13590 ( .A1(n11426), .A2(n11076), .ZN(n10600) );
  AND3_X1 U13591 ( .A1(n12761), .A2(n12760), .A3(n12759), .ZN(n10601) );
  OR2_X1 U13592 ( .A1(n19607), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19717) );
  INV_X2 U13593 ( .A(n19717), .ZN(n19682) );
  INV_X1 U13594 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12226) );
  INV_X2 U13595 ( .A(n18532), .ZN(n18533) );
  INV_X1 U13596 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18724) );
  INV_X1 U13597 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11774) );
  INV_X1 U13598 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13164) );
  NOR3_X1 U13599 ( .A1(n12350), .A2(n12349), .A3(n12348), .ZN(n12351) );
  INV_X1 U13600 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14733) );
  INV_X1 U13601 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11653) );
  INV_X1 U13602 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n19000) );
  INV_X2 U13603 ( .A(n19704), .ZN(n18488) );
  INV_X2 U13604 ( .A(n18534), .ZN(n18529) );
  INV_X1 U13605 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17301) );
  NOR2_X1 U13606 ( .A1(n21191), .A2(n21295), .ZN(n10602) );
  NOR2_X1 U13607 ( .A1(n21191), .A2(n21007), .ZN(n10603) );
  NAND2_X1 U13608 ( .A1(n15650), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n13907) );
  INV_X1 U13609 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12221) );
  OR2_X2 U13610 ( .A1(n13889), .A2(n11232), .ZN(n14077) );
  OR2_X1 U13611 ( .A1(n19898), .A2(n13353), .ZN(n16164) );
  INV_X1 U13612 ( .A(n13633), .ZN(n18992) );
  INV_X1 U13613 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21197) );
  OR2_X2 U13614 ( .A1(n13009), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20716) );
  INV_X1 U13615 ( .A(n20716), .ZN(n17416) );
  AND2_X1 U13616 ( .A1(n19870), .A2(BUF2_REG_30__SCAN_IN), .ZN(n10604) );
  NOR2_X1 U13617 ( .A1(n14207), .A2(n12586), .ZN(n12621) );
  INV_X1 U13618 ( .A(n12621), .ZN(n12605) );
  AND2_X1 U13619 ( .A1(n9737), .A2(n12517), .ZN(n10605) );
  NAND2_X1 U13620 ( .A1(n13656), .A2(n13655), .ZN(n15113) );
  INV_X1 U13621 ( .A(n15113), .ZN(n13660) );
  INV_X1 U13622 ( .A(n20646), .ZN(n17382) );
  AND2_X1 U13623 ( .A1(n18277), .A2(n18289), .ZN(n18286) );
  INV_X2 U13624 ( .A(n18286), .ZN(n18270) );
  NAND2_X2 U13625 ( .A1(n13352), .A2(n16899), .ZN(n19898) );
  OR2_X1 U13626 ( .A1(n13753), .A2(n19949), .ZN(n10606) );
  OR2_X1 U13627 ( .A1(n13753), .A2(n16168), .ZN(n10607) );
  AND3_X1 U13628 ( .A1(n14737), .A2(n14736), .A3(n14735), .ZN(n10608) );
  INV_X1 U13629 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16877) );
  BUF_X1 U13630 ( .A(n10807), .Z(n15941) );
  AND2_X1 U13631 ( .A1(n11426), .A2(n11309), .ZN(n10609) );
  INV_X1 U13632 ( .A(n12554), .ZN(n15666) );
  INV_X1 U13633 ( .A(n16400), .ZN(n11016) );
  AND4_X1 U13634 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n10611) );
  INV_X1 U13635 ( .A(n12256), .ZN(n12235) );
  AOI22_X1 U13636 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11883) );
  OR2_X1 U13637 ( .A1(n12955), .A2(n12954), .ZN(n12964) );
  OR2_X1 U13638 ( .A1(n12093), .A2(n12092), .ZN(n12199) );
  INV_X1 U13639 ( .A(n12294), .ZN(n12265) );
  INV_X1 U13640 ( .A(n12133), .ZN(n12288) );
  INV_X1 U13641 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12230) );
  INV_X1 U13642 ( .A(n11048), .ZN(n11049) );
  AOI22_X1 U13643 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13326), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10619) );
  INV_X1 U13644 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10635) );
  INV_X1 U13645 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11652) );
  OR2_X1 U13646 ( .A1(n12240), .A2(n12244), .ZN(n12242) );
  INV_X1 U13647 ( .A(n14914), .ZN(n12798) );
  AND2_X1 U13648 ( .A1(n12272), .A2(n12271), .ZN(n12274) );
  OR2_X1 U13649 ( .A1(n12069), .A2(n12068), .ZN(n12177) );
  INV_X1 U13650 ( .A(n12013), .ZN(n12158) );
  AND2_X1 U13651 ( .A1(n17324), .A2(n21357), .ZN(n14500) );
  NOR2_X1 U13652 ( .A1(n17301), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11094) );
  OR2_X1 U13653 ( .A1(n10914), .A2(n10913), .ZN(n11303) );
  OR2_X1 U13654 ( .A1(n10953), .A2(n10952), .ZN(n10954) );
  NOR2_X1 U13655 ( .A1(n11017), .A2(n11016), .ZN(n11018) );
  INV_X1 U13656 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10706) );
  AND2_X1 U13657 ( .A1(n11653), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13569) );
  INV_X1 U13658 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17207) );
  INV_X1 U13659 ( .A(n18668), .ZN(n13551) );
  OR2_X1 U13660 ( .A1(n12274), .A2(n12273), .ZN(n12296) );
  INV_X1 U13661 ( .A(n12440), .ZN(n12413) );
  INV_X1 U13662 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12830) );
  INV_X1 U13663 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12780) );
  INV_X1 U13664 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12130) );
  INV_X1 U13665 ( .A(n12243), .ZN(n12275) );
  INV_X1 U13666 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n21552) );
  OR3_X1 U13667 ( .A1(n11095), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n17363), .ZN(n11102) );
  INV_X1 U13668 ( .A(n15729), .ZN(n11801) );
  INV_X1 U13669 ( .A(n16172), .ZN(n11301) );
  INV_X1 U13670 ( .A(n13383), .ZN(n13384) );
  AND2_X1 U13671 ( .A1(n11103), .A2(n10992), .ZN(n11218) );
  INV_X1 U13672 ( .A(n19117), .ZN(n13582) );
  INV_X1 U13673 ( .A(n18564), .ZN(n11514) );
  INV_X1 U13674 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18057) );
  NAND2_X1 U13675 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12270), .ZN(
        n12298) );
  INV_X1 U13676 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12861) );
  INV_X1 U13677 ( .A(n14254), .ZN(n12368) );
  NAND2_X1 U13678 ( .A1(n12765), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13709) );
  INV_X1 U13679 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12679) );
  NAND2_X1 U13680 ( .A1(n12131), .A2(n12130), .ZN(n15296) );
  NAND2_X1 U13681 ( .A1(n12045), .A2(n12044), .ZN(n20953) );
  INV_X1 U13682 ( .A(n12534), .ZN(n14358) );
  INV_X1 U13683 ( .A(n11778), .ZN(n11780) );
  INV_X1 U13684 ( .A(n15665), .ZN(n12553) );
  AND2_X1 U13685 ( .A1(n13209), .A2(n13208), .ZN(n13233) );
  OR2_X1 U13686 ( .A1(n13106), .A2(n13105), .ZN(n16025) );
  INV_X1 U13687 ( .A(n11701), .ZN(n11439) );
  NOR2_X1 U13688 ( .A1(n10598), .A2(n13384), .ZN(n13385) );
  AND3_X1 U13689 ( .A1(n11162), .A2(n11161), .A3(n11160), .ZN(n15802) );
  AND3_X1 U13690 ( .A1(n11731), .A2(n11730), .A3(n11729), .ZN(n11733) );
  INV_X1 U13691 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16227) );
  AND2_X1 U13692 ( .A1(n16357), .A2(n16359), .ZN(n16342) );
  INV_X1 U13693 ( .A(n11312), .ZN(n14582) );
  INV_X1 U13694 ( .A(n11186), .ZN(n11265) );
  OR2_X1 U13695 ( .A1(n13030), .A2(n14157), .ZN(n13033) );
  NOR2_X2 U13696 ( .A1(n10812), .A2(n16768), .ZN(n16803) );
  INV_X1 U13697 ( .A(n20614), .ZN(n20266) );
  AND3_X1 U13698 ( .A1(n20335), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20372) );
  OR3_X1 U13699 ( .A1(n13573), .A2(n13572), .A3(n13586), .ZN(n13574) );
  INV_X1 U13700 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17226) );
  INV_X1 U13701 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18113) );
  AND2_X1 U13702 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17120) );
  AND2_X1 U13703 ( .A1(n17034), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17017) );
  NOR2_X1 U13704 ( .A1(n18411), .A2(n18414), .ZN(n13502) );
  INV_X1 U13705 ( .A(n19546), .ZN(n18916) );
  NAND2_X1 U13706 ( .A1(n15629), .A2(n10287), .ZN(n13009) );
  AND2_X1 U13707 ( .A1(n20708), .A2(n14883), .ZN(n15053) );
  INV_X1 U13708 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13813) );
  AND2_X1 U13709 ( .A1(n12405), .A2(n12404), .ZN(n14987) );
  NAND2_X1 U13710 ( .A1(n13834), .A2(n13833), .ZN(n13973) );
  AND2_X1 U13711 ( .A1(n14273), .A2(n17352), .ZN(n14274) );
  AOI21_X1 U13712 ( .B1(n14983), .B2(n14951), .A(n14950), .ZN(n14985) );
  INV_X1 U13713 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20665) );
  OR3_X1 U13714 ( .A1(n15452), .A2(n15425), .A3(n15424), .ZN(n15396) );
  AND2_X1 U13715 ( .A1(n12432), .A2(n12431), .ZN(n14833) );
  INV_X1 U13716 ( .A(n14465), .ZN(n15590) );
  INV_X1 U13717 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14261) );
  OR2_X1 U13718 ( .A1(n21063), .A2(n20817), .ZN(n20891) );
  OR2_X1 U13719 ( .A1(n21039), .A2(n21232), .ZN(n21004) );
  NOR2_X1 U13720 ( .A1(n21190), .A2(n20959), .ZN(n21134) );
  INV_X1 U13721 ( .A(n21065), .ZN(n21273) );
  NOR2_X1 U13722 ( .A1(n21126), .A2(n20959), .ZN(n21276) );
  NAND2_X1 U13723 ( .A1(n21357), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17355) );
  NAND2_X1 U13724 ( .A1(n12540), .A2(n12538), .ZN(n19809) );
  OR2_X1 U13725 ( .A1(n11342), .A2(n11341), .ZN(n14600) );
  OR2_X1 U13726 ( .A1(n14236), .A2(n14235), .ZN(n14238) );
  AND2_X1 U13727 ( .A1(n11438), .A2(n11437), .ZN(n11701) );
  INV_X1 U13728 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16238) );
  AND2_X1 U13729 ( .A1(n11258), .A2(n11257), .ZN(n11444) );
  INV_X1 U13730 ( .A(n19960), .ZN(n19949) );
  NOR2_X1 U13731 ( .A1(n11250), .A2(n11249), .ZN(n11251) );
  OR2_X1 U13732 ( .A1(n20032), .A2(n20031), .ZN(n20037) );
  AND2_X1 U13733 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20078) );
  OR2_X1 U13734 ( .A1(n16803), .A2(n16802), .ZN(n16809) );
  AND2_X1 U13735 ( .A1(n16831), .A2(n20335), .ZN(n20270) );
  OR2_X1 U13736 ( .A1(n16828), .A2(n16827), .ZN(n16834) );
  NAND2_X1 U13737 ( .A1(n20610), .A2(n20622), .ZN(n20339) );
  AND2_X1 U13738 ( .A1(n16877), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12543) );
  NAND2_X1 U13739 ( .A1(n13575), .A2(n11669), .ZN(n19541) );
  INV_X1 U13740 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17764) );
  INV_X1 U13741 ( .A(n17915), .ZN(n17906) );
  INV_X1 U13742 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18255) );
  INV_X1 U13743 ( .A(n18293), .ZN(n14241) );
  INV_X1 U13744 ( .A(n16914), .ZN(n18595) );
  INV_X1 U13745 ( .A(n17744), .ZN(n18703) );
  INV_X1 U13746 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17035) );
  NAND2_X1 U13747 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17866) );
  NAND2_X1 U13748 ( .A1(n19591), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18672) );
  INV_X1 U13749 ( .A(n19075), .ZN(n17135) );
  AND2_X1 U13750 ( .A1(n18976), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18977) );
  AND2_X1 U13751 ( .A1(n13596), .A2(n13595), .ZN(n19543) );
  INV_X1 U13752 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21541) );
  NAND2_X1 U13753 ( .A1(n19570), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19229) );
  AND2_X1 U13754 ( .A1(n12451), .A2(n14115), .ZN(n13794) );
  OR2_X1 U13755 ( .A1(n17355), .A2(n10287), .ZN(n20640) );
  AND2_X1 U13756 ( .A1(n15071), .A2(n14825), .ZN(n20672) );
  NAND2_X1 U13757 ( .A1(n15059), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14679) );
  INV_X1 U13758 ( .A(n15101), .ZN(n15108) );
  INV_X1 U13759 ( .A(n14383), .ZN(n20807) );
  OR2_X1 U13760 ( .A1(n14278), .A2(n14274), .ZN(n20804) );
  INV_X1 U13761 ( .A(n14949), .ZN(n15019) );
  INV_X1 U13762 ( .A(n17377), .ZN(n17379) );
  INV_X1 U13763 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14194) );
  NOR2_X1 U13764 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20814), .ZN(n20855) );
  OAI22_X1 U13765 ( .A1(n20825), .A2(n20824), .B1(n21069), .B2(n20955), .ZN(
        n20856) );
  INV_X1 U13766 ( .A(n20930), .ZN(n20918) );
  INV_X1 U13767 ( .A(n20929), .ZN(n20947) );
  NOR2_X2 U13768 ( .A1(n20930), .A2(n21155), .ZN(n20976) );
  INV_X1 U13769 ( .A(n21004), .ZN(n21030) );
  INV_X1 U13770 ( .A(n21014), .ZN(n21058) );
  OAI21_X1 U13771 ( .B1(n21097), .B2(n21096), .A(n21306), .ZN(n21119) );
  INV_X1 U13772 ( .A(n21128), .ZN(n21149) );
  NOR2_X2 U13773 ( .A1(n21161), .A2(n21262), .ZN(n21180) );
  INV_X1 U13774 ( .A(n21198), .ZN(n21226) );
  AND2_X1 U13775 ( .A1(n21264), .A2(n21184), .ZN(n21258) );
  INV_X1 U13776 ( .A(n21417), .ZN(n21292) );
  INV_X1 U13777 ( .A(n21355), .ZN(n21308) );
  AND2_X1 U13778 ( .A1(n20855), .A2(n20854), .ZN(n21349) );
  NOR2_X1 U13779 ( .A1(n13907), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n13878) );
  CLKBUF_X1 U13780 ( .A(n13878), .Z(n13905) );
  INV_X1 U13781 ( .A(n16080), .ZN(n12549) );
  INV_X1 U13782 ( .A(n19809), .ZN(n19829) );
  INV_X1 U13783 ( .A(n19833), .ZN(n19812) );
  INV_X1 U13784 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16001) );
  OR2_X1 U13785 ( .A1(n11411), .A2(n11410), .ZN(n14620) );
  INV_X1 U13786 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n16066) );
  OR2_X1 U13787 ( .A1(n16179), .A2(n14415), .ZN(n14594) );
  INV_X1 U13788 ( .A(n19855), .ZN(n19863) );
  AND2_X1 U13789 ( .A1(n13291), .A2(n13290), .ZN(n15986) );
  NOR2_X1 U13790 ( .A1(n14269), .A2(n16788), .ZN(n19869) );
  INV_X1 U13791 ( .A(n16164), .ZN(n19903) );
  AND2_X1 U13792 ( .A1(n14644), .A2(n13361), .ZN(n19899) );
  INV_X1 U13793 ( .A(n19908), .ZN(n19989) );
  INV_X1 U13794 ( .A(n19897), .ZN(n19993) );
  INV_X2 U13795 ( .A(n13993), .ZN(n14073) );
  INV_X1 U13796 ( .A(n14077), .ZN(n13926) );
  AND2_X1 U13797 ( .A1(n15788), .A2(n15803), .ZN(n16571) );
  AND2_X1 U13798 ( .A1(n14592), .A2(n14591), .ZN(n16678) );
  AND2_X1 U13799 ( .A1(n14371), .A2(n14375), .ZN(n19800) );
  INV_X1 U13800 ( .A(n16424), .ZN(n16450) );
  INV_X1 U13801 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16632) );
  OR2_X1 U13802 ( .A1(n14702), .A2(n9594), .ZN(n11471) );
  AND2_X1 U13803 ( .A1(n11494), .A2(n11447), .ZN(n19960) );
  INV_X1 U13804 ( .A(n20035), .ZN(n20053) );
  INV_X1 U13805 ( .A(n16793), .ZN(n20071) );
  AND2_X1 U13806 ( .A1(n20080), .A2(n20078), .ZN(n20104) );
  NOR2_X1 U13807 ( .A1(n20195), .A2(n20079), .ZN(n20131) );
  NAND2_X1 U13808 ( .A1(n16806), .A2(n16805), .ZN(n20191) );
  NOR2_X2 U13809 ( .A1(n20465), .A2(n20116), .ZN(n20218) );
  OAI21_X1 U13810 ( .B1(n20273), .B2(n20272), .A(n20271), .ZN(n20291) );
  AND2_X1 U13811 ( .A1(n16834), .A2(n16833), .ZN(n20329) );
  INV_X1 U13812 ( .A(n20343), .ZN(n20361) );
  NOR2_X2 U13813 ( .A1(n20339), .A2(n20375), .ZN(n20400) );
  NAND2_X1 U13814 ( .A1(n20416), .A2(n20415), .ZN(n20454) );
  AND2_X1 U13815 ( .A1(n20467), .A2(n19867), .ZN(n20462) );
  AND2_X1 U13816 ( .A1(n20023), .A2(n20002), .ZN(n20492) );
  AND2_X1 U13817 ( .A1(n20023), .A2(n20022), .ZN(n20510) );
  AND2_X1 U13818 ( .A1(n12543), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16899) );
  NOR2_X1 U13819 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19734) );
  INV_X1 U13820 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20540) );
  AOI21_X1 U13821 ( .B1(n19539), .B2(n19538), .A(n18492), .ZN(n19707) );
  NOR2_X2 U13822 ( .A1(n19690), .A2(n17924), .ZN(n17910) );
  AND2_X1 U13823 ( .A1(n19720), .A2(n11675), .ZN(n17924) );
  NAND2_X1 U13824 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n18135), .ZN(n18120) );
  INV_X1 U13825 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18231) );
  INV_X1 U13826 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18269) );
  NOR2_X2 U13827 ( .A1(n18425), .A2(n19135), .ZN(n18368) );
  AND4_X1 U13828 ( .A1(n13479), .A2(n13478), .A3(n13477), .A4(n13476), .ZN(
        n13490) );
  INV_X1 U13829 ( .A(n19108), .ZN(n18432) );
  INV_X1 U13830 ( .A(n18536), .ZN(n18530) );
  AND2_X1 U13831 ( .A1(n17096), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17121) );
  INV_X1 U13832 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18940) );
  AND2_X1 U13833 ( .A1(n17540), .A2(n11672), .ZN(n13633) );
  INV_X1 U13834 ( .A(n19090), .ZN(n19066) );
  AND2_X1 U13835 ( .A1(n19062), .A2(n19543), .ZN(n19086) );
  NAND2_X1 U13836 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19096) );
  NOR2_X1 U13837 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19690), .ZN(n19107) );
  INV_X1 U13838 ( .A(n19205), .ZN(n19198) );
  INV_X1 U13839 ( .A(n19223), .ZN(n19225) );
  INV_X1 U13840 ( .A(n19250), .ZN(n19243) );
  NOR2_X1 U13841 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19185) );
  INV_X1 U13842 ( .A(n19340), .ZN(n19328) );
  INV_X1 U13843 ( .A(n19362), .ZN(n19355) );
  INV_X1 U13844 ( .A(n19407), .ZN(n19414) );
  INV_X1 U13845 ( .A(n19500), .ZN(n19458) );
  INV_X1 U13846 ( .A(n19710), .ZN(n19705) );
  INV_X1 U13847 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19618) );
  INV_X1 U13848 ( .A(n16790), .ZN(n16788) );
  NAND2_X1 U13849 ( .A1(n14116), .A2(n13794), .ZN(n14278) );
  INV_X1 U13850 ( .A(n21396), .ZN(n21407) );
  INV_X1 U13851 ( .A(n13819), .ZN(n13820) );
  INV_X1 U13852 ( .A(n20735), .ZN(n15079) );
  AND2_X1 U13853 ( .A1(n13662), .A2(n13661), .ZN(n13663) );
  NAND2_X1 U13854 ( .A1(n15113), .A2(n14207), .ZN(n15101) );
  INV_X1 U13855 ( .A(n15328), .ZN(n15174) );
  NAND2_X1 U13856 ( .A1(n20766), .A2(n14119), .ZN(n14135) );
  NAND2_X1 U13857 ( .A1(n20786), .A2(n20774), .ZN(n20772) );
  OR2_X1 U13858 ( .A1(n14278), .A2(n14277), .ZN(n14383) );
  INV_X1 U13859 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21471) );
  INV_X1 U13860 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21132) );
  INV_X1 U13861 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13981) );
  NAND2_X1 U13862 ( .A1(n20918), .A2(n21184), .ZN(n20887) );
  AOI22_X1 U13863 ( .A1(n20895), .A2(n20892), .B1(n21006), .B2(n21126), .ZN(
        n20916) );
  AOI22_X1 U13864 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20925), .B1(n20927), 
        .B2(n20924), .ZN(n20950) );
  OR2_X1 U13865 ( .A1(n21039), .A2(n20952), .ZN(n21003) );
  AOI22_X1 U13866 ( .A1(n21011), .A2(n21008), .B1(n21006), .B2(n21190), .ZN(
        n21034) );
  OR2_X1 U13867 ( .A1(n21039), .A2(n21155), .ZN(n21070) );
  NAND2_X1 U13868 ( .A1(n21062), .A2(n21184), .ZN(n21122) );
  AOI22_X1 U13869 ( .A1(n21130), .A2(n21127), .B1(n21126), .B2(n21266), .ZN(
        n21154) );
  OR2_X1 U13870 ( .A1(n21161), .A2(n21155), .ZN(n21198) );
  INV_X1 U13871 ( .A(n21300), .ZN(n21201) );
  INV_X1 U13872 ( .A(n21335), .ZN(n21220) );
  NAND2_X1 U13873 ( .A1(n21264), .A2(n21233), .ZN(n21417) );
  NAND2_X1 U13874 ( .A1(n21264), .A2(n21263), .ZN(n21415) );
  NAND2_X1 U13875 ( .A1(n21264), .A2(n20813), .ZN(n21355) );
  INV_X1 U13876 ( .A(n21385), .ZN(n21361) );
  INV_X1 U13877 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n15650) );
  INV_X1 U13878 ( .A(n13907), .ZN(n21396) );
  INV_X1 U13879 ( .A(n13878), .ZN(n21376) );
  AND2_X1 U13880 ( .A1(n13889), .A2(n19837), .ZN(n19728) );
  NAND2_X1 U13881 ( .A1(n11250), .A2(n11113), .ZN(n13911) );
  OR2_X1 U13882 ( .A1(n15976), .A2(n19776), .ZN(n13755) );
  NAND2_X1 U13883 ( .A1(n14048), .A2(n20408), .ZN(n19776) );
  INV_X1 U13884 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19788) );
  XNOR2_X1 U13885 ( .A(n9713), .B(n14223), .ZN(n16799) );
  INV_X1 U13886 ( .A(n19869), .ZN(n16154) );
  INV_X1 U13887 ( .A(n16518), .ZN(n16122) );
  INV_X1 U13888 ( .A(n19899), .ZN(n16168) );
  INV_X1 U13889 ( .A(n19898), .ZN(n14644) );
  NOR2_X1 U13890 ( .A1(n19903), .A2(n19899), .ZN(n16183) );
  AND2_X1 U13891 ( .A1(n16160), .A2(n14269), .ZN(n19907) );
  NAND2_X1 U13892 ( .A1(n19928), .A2(n14168), .ZN(n19910) );
  INV_X1 U13893 ( .A(n14475), .ZN(n19930) );
  INV_X1 U13894 ( .A(n19928), .ZN(n19938) );
  INV_X1 U13895 ( .A(n16435), .ZN(n16459) );
  INV_X1 U13896 ( .A(n13402), .ZN(n13403) );
  NOR2_X1 U13897 ( .A1(n11705), .A2(n11704), .ZN(n11709) );
  NAND2_X1 U13898 ( .A1(n11494), .A2(n20632), .ZN(n19963) );
  INV_X1 U13899 ( .A(n17302), .ZN(n16773) );
  INV_X1 U13900 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20001) );
  INV_X1 U13901 ( .A(n20020), .ZN(n20058) );
  AOI211_X2 U13902 ( .C1(n16793), .C2(n16781), .A(n20119), .B(n16780), .ZN(
        n20077) );
  INV_X1 U13903 ( .A(n20097), .ZN(n20109) );
  INV_X1 U13904 ( .A(n20131), .ZN(n20143) );
  INV_X1 U13905 ( .A(n20166), .ZN(n20174) );
  INV_X1 U13906 ( .A(n20177), .ZN(n20194) );
  OR2_X1 U13907 ( .A1(n20195), .A2(n20465), .ZN(n20258) );
  NAND2_X1 U13908 ( .A1(n20405), .A2(n20222), .ZN(n20295) );
  INV_X1 U13909 ( .A(n20311), .ZN(n20308) );
  INV_X1 U13910 ( .A(n20325), .ZN(n20333) );
  INV_X1 U13911 ( .A(n20340), .ZN(n20366) );
  NAND2_X1 U13912 ( .A1(n20369), .A2(n20368), .ZN(n20452) );
  AOI22_X1 U13913 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16791), .ZN(n20458) );
  INV_X1 U13914 ( .A(n20606), .ZN(n20521) );
  INV_X1 U13915 ( .A(HOLD), .ZN(n21363) );
  INV_X1 U13916 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21509) );
  NAND2_X1 U13917 ( .A1(n9659), .A2(n19598), .ZN(n11686) );
  INV_X1 U13918 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17793) );
  NAND2_X1 U13919 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19601), .ZN(n17879) );
  INV_X1 U13920 ( .A(n17884), .ZN(n19723) );
  INV_X1 U13921 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18288) );
  INV_X1 U13922 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19125) );
  NOR2_X1 U13923 ( .A1(n18465), .A2(n18391), .ZN(n18394) );
  AND2_X1 U13924 ( .A1(n13490), .A2(n13489), .ZN(n18411) );
  AND2_X1 U13925 ( .A1(n18380), .A2(n18379), .ZN(n18429) );
  INV_X1 U13926 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18441) );
  INV_X1 U13927 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21491) );
  NAND2_X1 U13928 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18552), .ZN(n19704) );
  INV_X1 U13929 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18480) );
  INV_X1 U13930 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19105) );
  INV_X1 U13931 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18895) );
  INV_X1 U13932 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18830) );
  INV_X1 U13933 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18854) );
  INV_X1 U13934 ( .A(n18997), .ZN(n19012) );
  INV_X1 U13935 ( .A(n13633), .ZN(n18988) );
  OR2_X1 U13936 ( .A1(n19062), .A2(n18905), .ZN(n19090) );
  INV_X1 U13937 ( .A(n19057), .ZN(n19095) );
  INV_X1 U13938 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19568) );
  INV_X1 U13939 ( .A(n19289), .ZN(n19296) );
  INV_X1 U13940 ( .A(n19508), .ZN(n19377) );
  INV_X1 U13941 ( .A(n19522), .ZN(n19412) );
  INV_X1 U13942 ( .A(n19497), .ZN(n19461) );
  INV_X1 U13943 ( .A(n19452), .ZN(n19487) );
  INV_X1 U13944 ( .A(n19404), .ZN(n19519) );
  INV_X1 U13945 ( .A(n17879), .ZN(n19598) );
  INV_X1 U13946 ( .A(n19687), .ZN(n19602) );
  INV_X1 U13947 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19615) );
  INV_X1 U13948 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19628) );
  INV_X1 U13949 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19658) );
  INV_X1 U13950 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19134) );
  INV_X1 U13951 ( .A(n17499), .ZN(n17503) );
  INV_X1 U13952 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20544) );
  NAND2_X1 U13953 ( .A1(n13664), .A2(n13663), .ZN(P1_U2844) );
  OAI211_X1 U13954 ( .C1(n16279), .C2(n19974), .A(n11709), .B(n11708), .ZN(
        P2_U3027) );
  NAND2_X1 U13955 ( .A1(n11686), .A2(n11685), .ZN(P3_U2641) );
  NAND4_X1 U13956 ( .A1(n20812), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13862), .A4(
        n13861), .ZN(U214) );
  INV_X1 U13957 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10613) );
  NAND2_X2 U13958 ( .A1(n16745), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10622) );
  INV_X4 U13959 ( .A(n10622), .ZN(n13337) );
  INV_X2 U13960 ( .A(n13145), .ZN(n13326) );
  AOI22_X1 U13961 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13326), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10616) );
  INV_X2 U13962 ( .A(n10628), .ZN(n10690) );
  AOI22_X1 U13963 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13964 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10614) );
  AND2_X4 U13965 ( .A1(n11107), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10820) );
  AOI22_X1 U13966 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13967 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13968 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10617) );
  INV_X1 U13969 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13199) );
  INV_X1 U13970 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10623) );
  OAI22_X1 U13971 ( .A1(n10622), .A2(n13199), .B1(n13138), .B2(n10623), .ZN(
        n10626) );
  INV_X1 U13972 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13202) );
  INV_X1 U13973 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10624) );
  OAI22_X1 U13974 ( .A1(n13145), .A2(n13202), .B1(n13139), .B2(n10624), .ZN(
        n10625) );
  NAND2_X1 U13975 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10632) );
  INV_X1 U13976 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10627) );
  OR2_X1 U13977 ( .A1(n10670), .A2(n10627), .ZN(n10631) );
  OR2_X1 U13978 ( .A1(n10628), .A2(n19996), .ZN(n10630) );
  NAND2_X1 U13979 ( .A1(n13336), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10629) );
  NAND4_X1 U13980 ( .A1(n10632), .A2(n10631), .A3(n10630), .A4(n10629), .ZN(
        n10633) );
  NAND2_X1 U13981 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10639) );
  INV_X2 U13982 ( .A(n13145), .ZN(n13339) );
  NAND2_X1 U13983 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10638) );
  NAND2_X1 U13984 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10637) );
  NAND2_X1 U13985 ( .A1(n13327), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10636) );
  NAND4_X1 U13986 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10646) );
  NAND2_X1 U13987 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10644) );
  INV_X1 U13988 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10640) );
  OR2_X1 U13989 ( .A1(n10670), .A2(n10640), .ZN(n10643) );
  INV_X1 U13990 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13189) );
  OR2_X1 U13991 ( .A1(n10628), .A2(n13189), .ZN(n10642) );
  NAND2_X1 U13992 ( .A1(n13336), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10641) );
  NAND4_X1 U13993 ( .A1(n10644), .A2(n10643), .A3(n10642), .A4(n10641), .ZN(
        n10645) );
  NOR2_X1 U13994 ( .A1(n9588), .A2(n19992), .ZN(n10708) );
  AOI22_X1 U13995 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13339), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13996 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13997 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13998 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10647) );
  NAND4_X1 U13999 ( .A1(n10650), .A2(n10649), .A3(n10648), .A4(n10647), .ZN(
        n10750) );
  AOI22_X1 U14000 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U14001 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U14002 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10651) );
  NAND4_X1 U14003 ( .A1(n10654), .A2(n10653), .A3(n10652), .A4(n10651), .ZN(
        n10742) );
  NAND2_X1 U14004 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10658) );
  NAND2_X1 U14005 ( .A1(n13326), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10657) );
  NAND2_X1 U14006 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10656) );
  NAND2_X1 U14007 ( .A1(n13327), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10655) );
  NAND4_X1 U14008 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10664) );
  INV_X1 U14009 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10659) );
  NAND2_X1 U14010 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10662) );
  INV_X1 U14011 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13244) );
  OR2_X1 U14012 ( .A1(n10628), .A2(n13244), .ZN(n10661) );
  NAND2_X1 U14013 ( .A1(n13336), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10660) );
  NAND4_X1 U14014 ( .A1(n9731), .A2(n10662), .A3(n10661), .A4(n10660), .ZN(
        n10663) );
  NAND2_X1 U14015 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10668) );
  NAND2_X1 U14016 ( .A1(n13326), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10667) );
  NAND2_X1 U14017 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10666) );
  NAND2_X1 U14018 ( .A1(n13327), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10665) );
  NAND4_X1 U14019 ( .A1(n10668), .A2(n10667), .A3(n10666), .A4(n10665), .ZN(
        n10676) );
  INV_X1 U14020 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10669) );
  OR2_X1 U14021 ( .A1(n10670), .A2(n10669), .ZN(n10674) );
  NAND2_X1 U14022 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10673) );
  INV_X1 U14023 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13251) );
  OR2_X1 U14024 ( .A1(n10628), .A2(n13251), .ZN(n10672) );
  NAND2_X1 U14025 ( .A1(n13336), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10671) );
  NAND4_X1 U14026 ( .A1(n10674), .A2(n10673), .A3(n10672), .A4(n10671), .ZN(
        n10675) );
  AOI22_X1 U14027 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U14028 ( .A1(n13327), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U14029 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U14030 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13339), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U14031 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13339), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U14032 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U14033 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U14034 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U14035 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13326), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U14036 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U14037 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U14038 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10685) );
  NAND4_X1 U14039 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        n10689) );
  AOI22_X1 U14040 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13326), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U14041 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U14042 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U14043 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10691) );
  NAND4_X1 U14044 ( .A1(n10694), .A2(n10693), .A3(n10692), .A4(n10691), .ZN(
        n10696) );
  AOI22_X1 U14045 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13339), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U14046 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U14047 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U14048 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10697) );
  NAND4_X1 U14049 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n10701) );
  AOI22_X1 U14050 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13339), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U14051 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U14052 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U14053 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10702) );
  NAND4_X1 U14054 ( .A1(n10705), .A2(n10704), .A3(n10703), .A4(n10702), .ZN(
        n10707) );
  NAND2_X1 U14055 ( .A1(n10708), .A2(n11099), .ZN(n10709) );
  AOI22_X1 U14056 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U14057 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10820), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U14058 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U14059 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U14060 ( .A1(n13132), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U14061 ( .A1(n10820), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U14062 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U14063 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13326), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10715) );
  NAND2_X1 U14064 ( .A1(n13353), .A2(n19997), .ZN(n10771) );
  NAND4_X1 U14065 ( .A1(n10721), .A2(n11464), .A3(n10728), .A4(n10771), .ZN(
        n10727) );
  AND2_X1 U14066 ( .A1(n13353), .A2(n9588), .ZN(n11461) );
  INV_X1 U14067 ( .A(n11235), .ZN(n10729) );
  NAND2_X1 U14068 ( .A1(n13353), .A2(n20002), .ZN(n11243) );
  AND2_X1 U14069 ( .A1(n11243), .A2(n20022), .ZN(n10730) );
  NOR2_X1 U14070 ( .A1(n19997), .A2(n19992), .ZN(n10732) );
  AND2_X1 U14071 ( .A1(n11254), .A2(n20015), .ZN(n10731) );
  NAND4_X1 U14072 ( .A1(n11456), .A2(n10732), .A3(n10731), .A4(n20022), .ZN(
        n10733) );
  NAND2_X1 U14073 ( .A1(n10734), .A2(n16840), .ZN(n11485) );
  AOI22_X1 U14074 ( .A1(n11485), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n15656), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10735) );
  NAND2_X1 U14075 ( .A1(n14168), .A2(n9588), .ZN(n10760) );
  NAND2_X1 U14076 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10740) );
  NOR2_X1 U14077 ( .A1(n10741), .A2(n10740), .ZN(n10746) );
  INV_X1 U14078 ( .A(n10742), .ZN(n10745) );
  NAND4_X1 U14079 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n10756) );
  INV_X1 U14080 ( .A(n10747), .ZN(n10749) );
  NAND2_X1 U14081 ( .A1(n10543), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10748) );
  NOR2_X1 U14082 ( .A1(n10749), .A2(n10748), .ZN(n10754) );
  INV_X1 U14083 ( .A(n10750), .ZN(n10753) );
  NAND4_X1 U14084 ( .A1(n10754), .A2(n10753), .A3(n10752), .A4(n10751), .ZN(
        n10755) );
  NAND2_X1 U14085 ( .A1(n10756), .A2(n10755), .ZN(n10757) );
  NAND3_X1 U14086 ( .A1(n10758), .A2(n11455), .A3(n10757), .ZN(n10759) );
  INV_X1 U14087 ( .A(n10761), .ZN(n10762) );
  NAND2_X2 U14088 ( .A1(n10763), .A2(n10762), .ZN(n11117) );
  AOI21_X1 U14089 ( .B1(n16902), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10765) );
  NAND2_X1 U14090 ( .A1(n11117), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10768) );
  NAND2_X1 U14091 ( .A1(n10776), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U14092 ( .A1(n13774), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10766) );
  NAND3_X1 U14093 ( .A1(n11455), .A2(n20002), .A3(n20022), .ZN(n10774) );
  NAND2_X1 U14094 ( .A1(n15656), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10775) );
  INV_X1 U14095 ( .A(n15656), .ZN(n10779) );
  NAND2_X1 U14096 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10778) );
  OAI211_X1 U14097 ( .C1(n11118), .C2(n19748), .A(n10779), .B(n10778), .ZN(
        n10780) );
  AOI21_X1 U14098 ( .B1(n10781), .B2(n10777), .A(n10780), .ZN(n10784) );
  NAND2_X1 U14099 ( .A1(n11117), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10783) );
  NAND2_X1 U14100 ( .A1(n10785), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10787) );
  NAND2_X1 U14101 ( .A1(n15656), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10786) );
  NAND2_X1 U14102 ( .A1(n10787), .A2(n10786), .ZN(n10791) );
  INV_X1 U14103 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10790) );
  NAND2_X1 U14104 ( .A1(n11117), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10789) );
  AOI22_X1 U14105 ( .A1(n13774), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10788) );
  OAI211_X1 U14106 ( .C1(n13776), .C2(n10790), .A(n10789), .B(n10788), .ZN(
        n11115) );
  INV_X1 U14107 ( .A(n10806), .ZN(n10804) );
  XNOR2_X2 U14108 ( .A(n10804), .B(n10796), .ZN(n13030) );
  OR2_X2 U14109 ( .A1(n10814), .A2(n19965), .ZN(n10803) );
  NAND2_X1 U14110 ( .A1(n10806), .A2(n10797), .ZN(n10798) );
  NOR2_X2 U14111 ( .A1(n10803), .A2(n16768), .ZN(n10890) );
  INV_X1 U14112 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10811) );
  NOR2_X4 U14113 ( .A1(n10812), .A2(n19943), .ZN(n16782) );
  INV_X1 U14114 ( .A(n13030), .ZN(n10813) );
  INV_X1 U14115 ( .A(n20344), .ZN(n20336) );
  AOI22_X1 U14116 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n16782), .B1(
        n20336), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10819) );
  INV_X1 U14117 ( .A(n10815), .ZN(n10816) );
  INV_X1 U14118 ( .A(n19978), .ZN(n19983) );
  INV_X1 U14119 ( .A(n10919), .ZN(n20114) );
  INV_X1 U14120 ( .A(n10921), .ZN(n20226) );
  AOI22_X1 U14122 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10824) );
  AND2_X2 U14123 ( .A1(n13327), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10931) );
  AOI22_X1 U14124 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10823) );
  AND2_X2 U14125 ( .A1(n13337), .A2(n10635), .ZN(n10873) );
  AOI22_X1 U14126 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10822) );
  CLKBUF_X3 U14127 ( .A(n10820), .Z(n13338) );
  AND2_X2 U14128 ( .A1(n13338), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10908) );
  AOI22_X1 U14129 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10821) );
  NAND4_X1 U14130 ( .A1(n10824), .A2(n10823), .A3(n10822), .A4(n10821), .ZN(
        n10831) );
  AOI22_X1 U14131 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U14132 ( .A1(n10948), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U14134 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n13119), .B1(
        n13120), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U14135 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10826) );
  NAND4_X1 U14136 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10830) );
  AND2_X1 U14137 ( .A1(n11186), .A2(n13987), .ZN(n13917) );
  AOI22_X1 U14138 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10873), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U14139 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U14140 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13119), .B1(
        n13120), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U14141 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10835) );
  NAND4_X1 U14142 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(
        n10845) );
  AOI22_X1 U14143 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U14144 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10908), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U14145 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10847), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U14146 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10882), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10840) );
  NAND4_X1 U14147 ( .A1(n10843), .A2(n10842), .A3(n10841), .A4(n10840), .ZN(
        n10844) );
  NAND2_X1 U14148 ( .A1(n13917), .A2(n11272), .ZN(n11190) );
  AOI22_X1 U14149 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U14150 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U14151 ( .A1(n10948), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U14152 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10908), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10848) );
  NAND4_X1 U14153 ( .A1(n10851), .A2(n10850), .A3(n10849), .A4(n10848), .ZN(
        n10858) );
  AOI22_X1 U14154 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U14155 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U14156 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13119), .B1(
        n13120), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U14157 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10853) );
  NAND4_X1 U14158 ( .A1(n10856), .A2(n10855), .A3(n10854), .A4(n10853), .ZN(
        n10857) );
  NAND2_X1 U14159 ( .A1(n11190), .A2(n11282), .ZN(n10859) );
  INV_X1 U14160 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10860) );
  INV_X1 U14161 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13221) );
  INV_X1 U14162 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10861) );
  INV_X1 U14163 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13222) );
  OAI22_X1 U14164 ( .A1(n10861), .A2(n20463), .B1(n20371), .B2(n13222), .ZN(
        n10862) );
  INV_X1 U14165 ( .A(n10862), .ZN(n10863) );
  AOI22_X1 U14166 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n16828), .B1(
        n10889), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U14167 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20197), .B1(
        n20150), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U14168 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n16782), .B1(
        n16803), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U14169 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20085), .B1(
        n20032), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U14170 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U14171 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U14172 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13119), .B1(
        n13120), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U14173 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U14174 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U14175 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10882), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U14176 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U14177 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U14178 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U14179 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13119), .B1(
        n13120), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U14180 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10877) );
  NAND4_X1 U14181 ( .A1(n10880), .A2(n10879), .A3(n10878), .A4(n10877), .ZN(
        n10888) );
  AOI22_X1 U14182 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U14183 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10885) );
  AOI22_X1 U14184 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10884) );
  AOI22_X1 U14185 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10882), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10883) );
  NAND4_X1 U14186 ( .A1(n10886), .A2(n10885), .A3(n10884), .A4(n10883), .ZN(
        n10887) );
  AOI22_X1 U14187 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n16803), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U14188 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n16782), .B1(
        n16819), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10891) );
  INV_X1 U14189 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10895) );
  INV_X1 U14190 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20010) );
  OAI22_X1 U14191 ( .A1(n10895), .A2(n10919), .B1(n19978), .B2(n20010), .ZN(
        n10896) );
  INV_X1 U14192 ( .A(n10896), .ZN(n10903) );
  INV_X1 U14193 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10897) );
  INV_X1 U14194 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13280) );
  OAI22_X1 U14195 ( .A1(n10897), .A2(n20344), .B1(n10921), .B2(n13280), .ZN(
        n10898) );
  INV_X1 U14196 ( .A(n10898), .ZN(n10902) );
  INV_X1 U14197 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10899) );
  INV_X1 U14198 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13281) );
  OAI22_X1 U14199 ( .A1(n10899), .A2(n20463), .B1(n20371), .B2(n13281), .ZN(
        n10900) );
  INV_X1 U14200 ( .A(n10900), .ZN(n10901) );
  AOI22_X1 U14201 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U14202 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U14203 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n13119), .B1(
        n13120), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U14204 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10904) );
  NAND4_X1 U14205 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n10914) );
  AOI22_X1 U14206 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U14207 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U14208 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U14209 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n10882), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10909) );
  NAND4_X1 U14210 ( .A1(n10912), .A2(n10911), .A3(n10910), .A4(n10909), .ZN(
        n10913) );
  AOI22_X1 U14211 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n16782), .B1(
        n16819), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U14212 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n16803), .B1(
        n10890), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U14213 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20085), .B1(
        n20032), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U14214 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20197), .B1(
        n20150), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10916) );
  INV_X1 U14215 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10920) );
  INV_X1 U14216 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20019) );
  OAI22_X1 U14217 ( .A1(n10920), .A2(n10919), .B1(n19978), .B2(n20019), .ZN(
        n10926) );
  INV_X1 U14218 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10922) );
  INV_X1 U14219 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13304) );
  OAI22_X1 U14220 ( .A1(n10922), .A2(n20344), .B1(n10921), .B2(n13304), .ZN(
        n10925) );
  INV_X1 U14221 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10923) );
  INV_X1 U14222 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13305) );
  OAI22_X1 U14223 ( .A1(n10923), .A2(n20463), .B1(n20371), .B2(n13305), .ZN(
        n10924) );
  AOI22_X1 U14224 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U14225 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U14226 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13119), .B1(
        n13120), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U14227 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10927) );
  NAND4_X1 U14228 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n10937) );
  AOI22_X1 U14229 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U14230 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U14231 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U14232 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10882), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10932) );
  NAND4_X1 U14233 ( .A1(n10935), .A2(n10934), .A3(n10933), .A4(n10932), .ZN(
        n10936) );
  AOI22_X1 U14234 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U14235 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14236 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14237 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10882), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10939) );
  NAND4_X1 U14238 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10955) );
  AOI22_X1 U14239 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U14240 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13119), .B1(
        n13120), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10945) );
  NAND2_X1 U14241 ( .A1(n10852), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10944) );
  NAND2_X1 U14242 ( .A1(n10832), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10943) );
  NAND4_X1 U14243 ( .A1(n10946), .A2(n10945), .A3(n10944), .A4(n10943), .ZN(
        n10953) );
  INV_X1 U14244 ( .A(n10947), .ZN(n11108) );
  INV_X1 U14245 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10951) );
  INV_X1 U14246 ( .A(n10948), .ZN(n10950) );
  INV_X1 U14247 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10949) );
  OAI22_X1 U14248 ( .A1(n11108), .A2(n10951), .B1(n10950), .B2(n10949), .ZN(
        n10952) );
  NAND2_X1 U14249 ( .A1(n11217), .A2(n10991), .ZN(n10957) );
  NAND2_X1 U14250 ( .A1(n20335), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10956) );
  NAND2_X1 U14251 ( .A1(n10957), .A2(n10956), .ZN(n10965) );
  XNOR2_X1 U14252 ( .A(n10958), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10963) );
  XNOR2_X1 U14253 ( .A(n10965), .B(n10963), .ZN(n11222) );
  INV_X1 U14254 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10961) );
  CLKBUF_X3 U14255 ( .A(n10960), .Z(n20006) );
  NOR2_X1 U14256 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10962) );
  INV_X1 U14257 ( .A(n10963), .ZN(n10964) );
  NAND2_X1 U14258 ( .A1(n10965), .A2(n10964), .ZN(n10967) );
  NAND2_X1 U14259 ( .A1(n16860), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10966) );
  NAND2_X1 U14260 ( .A1(n10967), .A2(n10966), .ZN(n10970) );
  XNOR2_X1 U14261 ( .A(n10970), .B(n10969), .ZN(n11100) );
  OAI21_X1 U14262 ( .B1(n11289), .B2(n11253), .A(n10968), .ZN(n11090) );
  MUX2_X1 U14263 ( .A(n11090), .B(P2_EBX_REG_3__SCAN_IN), .S(n13390), .Z(
        n10988) );
  NAND2_X1 U14264 ( .A1(n10970), .A2(n10969), .ZN(n10972) );
  NAND2_X1 U14265 ( .A1(n20618), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10971) );
  NAND2_X1 U14266 ( .A1(n10972), .A2(n10971), .ZN(n11095) );
  MUX2_X1 U14267 ( .A(n11295), .B(n11102), .S(n11253), .Z(n11091) );
  INV_X1 U14268 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11121) );
  MUX2_X1 U14269 ( .A(n11091), .B(n11121), .S(n13390), .Z(n11002) );
  INV_X1 U14270 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14376) );
  INV_X1 U14271 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n14420) );
  MUX2_X1 U14272 ( .A(n11309), .B(n14420), .S(n13390), .Z(n10973) );
  INV_X1 U14273 ( .A(n10973), .ZN(n10974) );
  NAND2_X1 U14274 ( .A1(n9619), .A2(n10974), .ZN(n10975) );
  AND2_X1 U14275 ( .A1(n10981), .A2(n10975), .ZN(n15929) );
  INV_X1 U14276 ( .A(n15929), .ZN(n10976) );
  INV_X1 U14277 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14460) );
  MUX2_X1 U14278 ( .A(n14460), .B(n11076), .S(n20006), .Z(n10980) );
  INV_X1 U14279 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n15902) );
  NOR2_X1 U14280 ( .A1(n20006), .A2(n15902), .ZN(n10977) );
  AND2_X1 U14281 ( .A1(n10978), .A2(n10977), .ZN(n10979) );
  OR2_X1 U14282 ( .A1(n11021), .A2(n10979), .ZN(n15905) );
  NOR2_X1 U14283 ( .A1(n15905), .A2(n13768), .ZN(n10982) );
  NAND2_X1 U14284 ( .A1(n10982), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16388) );
  INV_X1 U14285 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16704) );
  XNOR2_X1 U14286 ( .A(n10981), .B(n10980), .ZN(n10984) );
  NAND2_X1 U14287 ( .A1(n10984), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16400) );
  AND3_X1 U14288 ( .A1(n16388), .A2(n16704), .A3(n16400), .ZN(n10985) );
  INV_X1 U14289 ( .A(n10982), .ZN(n10983) );
  INV_X1 U14290 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U14291 ( .A1(n10983), .A2(n11330), .ZN(n16387) );
  INV_X1 U14292 ( .A(n10984), .ZN(n15917) );
  NAND2_X1 U14293 ( .A1(n15917), .A2(n11205), .ZN(n16399) );
  XNOR2_X1 U14294 ( .A(n10989), .B(n10988), .ZN(n15942) );
  NAND2_X1 U14295 ( .A1(n9757), .A2(n9618), .ZN(n10990) );
  NAND2_X1 U14296 ( .A1(n10990), .A2(n10989), .ZN(n15958) );
  XNOR2_X1 U14297 ( .A(n15958), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13961) );
  NAND2_X1 U14298 ( .A1(n10093), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10992) );
  MUX2_X1 U14299 ( .A(n11186), .B(n11218), .S(n11253), .Z(n11085) );
  MUX2_X1 U14300 ( .A(P2_EBX_REG_0__SCAN_IN), .B(n11085), .S(n20006), .Z(
        n19828) );
  NAND2_X1 U14301 ( .A1(n19828), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13935) );
  INV_X1 U14302 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13933) );
  INV_X1 U14303 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13992) );
  NAND3_X1 U14304 ( .A1(n11254), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10993) );
  NAND2_X1 U14305 ( .A1(n9618), .A2(n10993), .ZN(n15969) );
  AOI21_X1 U14306 ( .B1(n13935), .B2(n13933), .A(n15969), .ZN(n10994) );
  INV_X1 U14307 ( .A(n10994), .ZN(n10997) );
  INV_X1 U14308 ( .A(n13935), .ZN(n10995) );
  NAND2_X1 U14309 ( .A1(n10995), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10996) );
  NAND2_X1 U14310 ( .A1(n10997), .A2(n10996), .ZN(n13960) );
  NAND2_X1 U14311 ( .A1(n13961), .A2(n13960), .ZN(n11000) );
  INV_X1 U14312 ( .A(n15958), .ZN(n10998) );
  NAND2_X1 U14313 ( .A1(n10998), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10999) );
  NAND2_X1 U14314 ( .A1(n11000), .A2(n10999), .ZN(n16447) );
  INV_X1 U14315 ( .A(n11001), .ZN(n11004) );
  INV_X1 U14316 ( .A(n11002), .ZN(n11003) );
  XNOR2_X1 U14317 ( .A(n11004), .B(n11003), .ZN(n19808) );
  NAND2_X1 U14318 ( .A1(n19808), .A2(n16725), .ZN(n11007) );
  OAI21_X1 U14319 ( .B1(n16447), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11007), .ZN(n11005) );
  INV_X1 U14320 ( .A(n11005), .ZN(n11006) );
  NAND3_X1 U14321 ( .A1(n11007), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n16447), .ZN(n11010) );
  INV_X1 U14322 ( .A(n19808), .ZN(n11008) );
  NAND2_X1 U14323 ( .A1(n11008), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11009) );
  AND2_X1 U14324 ( .A1(n11010), .A2(n11009), .ZN(n11011) );
  NAND2_X1 U14325 ( .A1(n10532), .A2(n11013), .ZN(n11014) );
  NAND2_X1 U14326 ( .A1(n9619), .A2(n11014), .ZN(n19791) );
  INV_X1 U14327 ( .A(n16388), .ZN(n11017) );
  INV_X1 U14328 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n19772) );
  NOR2_X1 U14329 ( .A1(n11021), .A2(n19772), .ZN(n11019) );
  MUX2_X1 U14330 ( .A(n11021), .B(n11019), .S(n13390), .Z(n11020) );
  INV_X1 U14331 ( .A(n11020), .ZN(n11022) );
  NAND2_X1 U14332 ( .A1(n11022), .A2(n11031), .ZN(n11038) );
  INV_X1 U14333 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16638) );
  OAI21_X1 U14334 ( .B1(n11038), .B2(n13768), .A(n16638), .ZN(n16377) );
  NAND2_X1 U14335 ( .A1(n13390), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U14336 ( .A1(n11024), .A2(n10116), .ZN(n11026) );
  NAND2_X1 U14337 ( .A1(n11041), .A2(n11026), .ZN(n15878) );
  OR2_X1 U14338 ( .A1(n15878), .A2(n13768), .ZN(n11027) );
  NAND2_X1 U14339 ( .A1(n11027), .A2(n16632), .ZN(n16344) );
  NOR2_X1 U14340 ( .A1(n20006), .A2(n16066), .ZN(n11028) );
  AOI21_X1 U14341 ( .B1(n9693), .B2(n11028), .A(n11778), .ZN(n11029) );
  NAND2_X1 U14342 ( .A1(n11024), .A2(n11029), .ZN(n19757) );
  OR2_X1 U14343 ( .A1(n19757), .A2(n13768), .ZN(n11030) );
  INV_X1 U14344 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16640) );
  NAND2_X1 U14345 ( .A1(n11030), .A2(n16640), .ZN(n16360) );
  NAND2_X1 U14346 ( .A1(n13390), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11032) );
  MUX2_X1 U14347 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n11032), .S(n11031), .Z(
        n11034) );
  AND2_X1 U14348 ( .A1(n11034), .A2(n11033), .ZN(n15892) );
  AND2_X1 U14349 ( .A1(n15892), .A2(n11076), .ZN(n11037) );
  INV_X1 U14350 ( .A(n11037), .ZN(n11035) );
  INV_X1 U14351 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16658) );
  NAND2_X1 U14352 ( .A1(n11035), .A2(n16658), .ZN(n16369) );
  AND2_X1 U14353 ( .A1(n16360), .A2(n16369), .ZN(n11036) );
  AND2_X1 U14354 ( .A1(n16344), .A2(n11036), .ZN(n11741) );
  NAND2_X1 U14355 ( .A1(n11037), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16370) );
  INV_X1 U14356 ( .A(n11038), .ZN(n19775) );
  AND2_X1 U14357 ( .A1(n11076), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11039) );
  NAND2_X1 U14358 ( .A1(n19775), .A2(n11039), .ZN(n16376) );
  AND2_X1 U14359 ( .A1(n16370), .A2(n16376), .ZN(n16357) );
  NAND2_X1 U14360 ( .A1(n11076), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11040) );
  OR2_X1 U14361 ( .A1(n19757), .A2(n11040), .ZN(n16359) );
  INV_X1 U14362 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n15862) );
  NOR2_X1 U14363 ( .A1(n20006), .A2(n15862), .ZN(n11042) );
  NAND2_X1 U14364 ( .A1(n11041), .A2(n11042), .ZN(n11043) );
  NAND2_X1 U14365 ( .A1(n9656), .A2(n11043), .ZN(n15865) );
  OR2_X1 U14366 ( .A1(n15865), .A2(n13768), .ZN(n11044) );
  INV_X1 U14367 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16618) );
  OR2_X1 U14368 ( .A1(n11044), .A2(n16618), .ZN(n16331) );
  OR3_X1 U14369 ( .A1(n15878), .A2(n13768), .A3(n16632), .ZN(n16345) );
  NAND2_X1 U14370 ( .A1(n11044), .A2(n16618), .ZN(n16330) );
  INV_X1 U14371 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n15853) );
  NOR2_X1 U14372 ( .A1(n20006), .A2(n15853), .ZN(n11048) );
  XNOR2_X1 U14373 ( .A(n9656), .B(n11048), .ZN(n15856) );
  INV_X1 U14374 ( .A(n15856), .ZN(n11046) );
  NAND2_X1 U14375 ( .A1(n11046), .A2(n11076), .ZN(n11047) );
  INV_X1 U14376 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16598) );
  NAND2_X1 U14377 ( .A1(n11047), .A2(n16598), .ZN(n16323) );
  OR3_X1 U14378 ( .A1(n15856), .A2(n13768), .A3(n16598), .ZN(n16322) );
  INV_X1 U14379 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n15838) );
  NOR2_X1 U14380 ( .A1(n20006), .A2(n15838), .ZN(n11050) );
  NAND2_X1 U14381 ( .A1(n11051), .A2(n11050), .ZN(n11052) );
  NAND2_X1 U14382 ( .A1(n11063), .A2(n11052), .ZN(n15839) );
  NOR2_X1 U14383 ( .A1(n15839), .A2(n13768), .ZN(n11053) );
  NAND2_X1 U14384 ( .A1(n11053), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16307) );
  INV_X1 U14385 ( .A(n16307), .ZN(n11055) );
  INV_X1 U14386 ( .A(n11053), .ZN(n11054) );
  NAND2_X1 U14387 ( .A1(n11054), .A2(n16568), .ZN(n16306) );
  INV_X1 U14388 ( .A(n11063), .ZN(n11056) );
  INV_X1 U14389 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n15824) );
  NAND2_X1 U14390 ( .A1(n11056), .A2(n15824), .ZN(n11061) );
  NOR2_X1 U14391 ( .A1(n20006), .A2(n15824), .ZN(n11057) );
  AOI21_X1 U14392 ( .B1(n11063), .B2(n11057), .A(n11778), .ZN(n11058) );
  NAND2_X1 U14393 ( .A1(n11061), .A2(n11058), .ZN(n15827) );
  NOR2_X1 U14394 ( .A1(n15827), .A2(n13768), .ZN(n11075) );
  INV_X1 U14395 ( .A(n11075), .ZN(n11059) );
  XNOR2_X1 U14396 ( .A(n11059), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11751) );
  INV_X1 U14397 ( .A(n11751), .ZN(n16303) );
  INV_X1 U14398 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n15808) );
  NOR2_X1 U14399 ( .A1(n20006), .A2(n15808), .ZN(n11060) );
  NAND2_X1 U14400 ( .A1(n11061), .A2(n11060), .ZN(n11064) );
  NOR2_X1 U14401 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n11062) );
  INV_X1 U14402 ( .A(n9638), .ZN(n11066) );
  NAND2_X1 U14403 ( .A1(n11064), .A2(n11066), .ZN(n15809) );
  NOR2_X1 U14404 ( .A1(n15809), .A2(n13768), .ZN(n11074) );
  INV_X1 U14405 ( .A(n11074), .ZN(n11065) );
  INV_X1 U14406 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16577) );
  NAND2_X1 U14407 ( .A1(n11065), .A2(n16577), .ZN(n11742) );
  NAND2_X1 U14408 ( .A1(n13390), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11067) );
  MUX2_X1 U14409 ( .A(n13390), .B(n11067), .S(n11066), .Z(n11068) );
  INV_X1 U14410 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n16043) );
  NAND2_X1 U14411 ( .A1(n9638), .A2(n16043), .ZN(n11071) );
  AND2_X1 U14412 ( .A1(n11076), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11069) );
  NAND2_X1 U14413 ( .A1(n15794), .A2(n11069), .ZN(n16281) );
  INV_X1 U14414 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11169) );
  NOR2_X1 U14415 ( .A1(n20006), .A2(n11169), .ZN(n11070) );
  NAND2_X1 U14416 ( .A1(n11071), .A2(n11070), .ZN(n11073) );
  OAI21_X1 U14417 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n13390), .ZN(n11072) );
  NAND2_X1 U14418 ( .A1(n11073), .A2(n9634), .ZN(n15774) );
  INV_X1 U14419 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11707) );
  OR3_X1 U14420 ( .A1(n15774), .A2(n13768), .A3(n11707), .ZN(n11690) );
  AND2_X1 U14421 ( .A1(n16281), .A2(n11690), .ZN(n11758) );
  NAND2_X1 U14422 ( .A1(n11074), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11756) );
  NAND2_X1 U14423 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11754) );
  NAND2_X1 U14424 ( .A1(n15794), .A2(n11076), .ZN(n11077) );
  INV_X1 U14425 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16553) );
  NAND2_X1 U14426 ( .A1(n11077), .A2(n16553), .ZN(n16282) );
  OR2_X1 U14427 ( .A1(n15774), .A2(n13768), .ZN(n11078) );
  NAND2_X1 U14428 ( .A1(n11078), .A2(n11707), .ZN(n11743) );
  NAND2_X1 U14429 ( .A1(n13390), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11079) );
  XNOR2_X1 U14430 ( .A(n9634), .B(n11079), .ZN(n15768) );
  AND2_X1 U14431 ( .A1(n11076), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11080) );
  NAND2_X1 U14432 ( .A1(n15768), .A2(n11080), .ZN(n11757) );
  INV_X1 U14433 ( .A(n16260), .ZN(n11084) );
  NAND2_X1 U14434 ( .A1(n15768), .A2(n11076), .ZN(n11081) );
  INV_X1 U14435 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11488) );
  NAND2_X1 U14436 ( .A1(n11081), .A2(n11488), .ZN(n16259) );
  AOI21_X1 U14437 ( .B1(n16259), .B2(n11757), .A(n11082), .ZN(n11083) );
  AOI21_X1 U14438 ( .B1(n11084), .B2(n16259), .A(n11083), .ZN(n11498) );
  INV_X1 U14439 ( .A(n11085), .ZN(n11089) );
  INV_X1 U14440 ( .A(n11217), .ZN(n11088) );
  INV_X1 U14441 ( .A(n11086), .ZN(n11087) );
  OAI21_X1 U14442 ( .B1(n11089), .B2(n11088), .A(n11087), .ZN(n11093) );
  INV_X1 U14443 ( .A(n11090), .ZN(n11092) );
  NAND2_X1 U14444 ( .A1(n11093), .A2(n11226), .ZN(n11098) );
  NAND2_X1 U14445 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17301), .ZN(
        n11096) );
  NAND2_X1 U14446 ( .A1(n11098), .A2(n11228), .ZN(n20633) );
  INV_X1 U14447 ( .A(n11099), .ZN(n16857) );
  AND2_X1 U14448 ( .A1(n13987), .A2(n16856), .ZN(n11236) );
  NAND2_X1 U14449 ( .A1(n16857), .A2(n11236), .ZN(n11493) );
  INV_X1 U14450 ( .A(n11100), .ZN(n11101) );
  NAND2_X1 U14451 ( .A1(n11102), .A2(n11101), .ZN(n11223) );
  XNOR2_X1 U14452 ( .A(n11217), .B(n11103), .ZN(n11215) );
  NAND2_X1 U14453 ( .A1(n11222), .A2(n11215), .ZN(n11104) );
  NAND2_X1 U14454 ( .A1(n11222), .A2(n11218), .ZN(n11105) );
  OAI21_X1 U14455 ( .B1(n11223), .B2(n11105), .A(n16877), .ZN(n11106) );
  OR2_X1 U14456 ( .A1(n16847), .A2(n11106), .ZN(n11111) );
  AOI21_X1 U14457 ( .B1(n16757), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17297) );
  NAND2_X1 U14458 ( .A1(n11108), .A2(n17297), .ZN(n11109) );
  INV_X1 U14459 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n16853) );
  NAND2_X1 U14460 ( .A1(n11109), .A2(n16853), .ZN(n11110) );
  NAND2_X1 U14461 ( .A1(n11110), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20620) );
  NAND2_X1 U14462 ( .A1(n11111), .A2(n20620), .ZN(n20629) );
  NAND3_X1 U14463 ( .A1(n16857), .A2(n11232), .A3(n20629), .ZN(n11112) );
  AND2_X1 U14464 ( .A1(n16856), .A2(n16899), .ZN(n11113) );
  INV_X1 U14465 ( .A(n13911), .ZN(n11114) );
  INV_X1 U14466 ( .A(n11115), .ZN(n11116) );
  NAND2_X1 U14468 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11120) );
  AOI22_X1 U14469 ( .A1(n11720), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11119) );
  OAI211_X1 U14470 ( .C1(n11121), .C2(n13776), .A(n11120), .B(n11119), .ZN(
        n16436) );
  NAND2_X1 U14471 ( .A1(n16437), .A2(n16436), .ZN(n14373) );
  INV_X1 U14472 ( .A(n14373), .ZN(n11126) );
  NAND2_X1 U14473 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14474 ( .A1(n12555), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11123) );
  AOI22_X1 U14475 ( .A1(n11720), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11122) );
  INV_X1 U14476 ( .A(n14374), .ZN(n11125) );
  NAND2_X1 U14477 ( .A1(n11126), .A2(n11125), .ZN(n14371) );
  INV_X2 U14478 ( .A(n14371), .ZN(n11131) );
  NAND2_X1 U14479 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11129) );
  NAND2_X1 U14480 ( .A1(n12555), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U14481 ( .A1(n11720), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11127) );
  NAND2_X1 U14482 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14483 ( .A1(n12555), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U14484 ( .A1(n11720), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14485 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11136) );
  AOI22_X1 U14486 ( .A1(n11720), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11135) );
  OAI211_X1 U14487 ( .C1(n15902), .C2(n13776), .A(n11136), .B(n11135), .ZN(
        n14590) );
  NAND2_X1 U14488 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11139) );
  NAND2_X1 U14489 ( .A1(n12555), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11138) );
  AOI22_X1 U14490 ( .A1(n11720), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11137) );
  NAND2_X1 U14491 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11142) );
  NAND2_X1 U14492 ( .A1(n12555), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11141) );
  AOI22_X1 U14493 ( .A1(n11720), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11140) );
  INV_X1 U14494 ( .A(n15889), .ZN(n11143) );
  NAND2_X1 U14495 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11145) );
  AOI22_X1 U14496 ( .A1(n13774), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11144) );
  OAI211_X1 U14497 ( .C1(n16066), .C2(n13776), .A(n11145), .B(n11144), .ZN(
        n16063) );
  INV_X1 U14498 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n15877) );
  NAND2_X1 U14499 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11147) );
  AOI22_X1 U14500 ( .A1(n13774), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11146) );
  OAI211_X1 U14501 ( .C1(n15877), .C2(n13776), .A(n11147), .B(n11146), .ZN(
        n15875) );
  NAND2_X1 U14502 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11150) );
  NAND2_X1 U14503 ( .A1(n12555), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14504 ( .A1(n11720), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11148) );
  NAND2_X1 U14505 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11153) );
  NAND2_X1 U14506 ( .A1(n12555), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11152) );
  AOI22_X1 U14507 ( .A1(n11720), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11151) );
  NAND2_X1 U14508 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11156) );
  AOI22_X1 U14509 ( .A1(n11720), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11155) );
  OAI211_X1 U14510 ( .C1(n15838), .C2(n13776), .A(n11156), .B(n11155), .ZN(
        n15835) );
  NAND2_X1 U14511 ( .A1(n14614), .A2(n15835), .ZN(n15819) );
  NAND2_X1 U14512 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11159) );
  NAND2_X1 U14513 ( .A1(n12555), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11158) );
  AOI22_X1 U14514 ( .A1(n11720), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11157) );
  NOR2_X4 U14515 ( .A1(n15819), .A2(n15822), .ZN(n15801) );
  NAND2_X1 U14516 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11162) );
  NAND2_X1 U14517 ( .A1(n12555), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11161) );
  AOI22_X1 U14518 ( .A1(n11720), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11160) );
  NAND2_X1 U14519 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11166) );
  NAND2_X1 U14520 ( .A1(n12555), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U14521 ( .A1(n11720), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11164) );
  NAND2_X1 U14522 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11168) );
  AOI22_X1 U14523 ( .A1(n11720), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11167) );
  OAI211_X1 U14524 ( .C1(n11169), .C2(n13776), .A(n11168), .B(n11167), .ZN(
        n11693) );
  INV_X1 U14525 ( .A(n11173), .ZN(n11174) );
  NAND2_X1 U14526 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11172) );
  NAND2_X1 U14527 ( .A1(n12555), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14528 ( .A1(n11720), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11170) );
  OAI21_X1 U14529 ( .B1(n11174), .B2(n9787), .A(n15748), .ZN(n16034) );
  INV_X1 U14530 ( .A(n16034), .ZN(n11181) );
  NOR2_X1 U14531 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19730) );
  INV_X1 U14532 ( .A(n19730), .ZN(n17296) );
  NAND2_X1 U14533 ( .A1(n20614), .A2(n17296), .ZN(n14437) );
  NAND2_X1 U14534 ( .A1(n14437), .A2(n16902), .ZN(n11175) );
  AND2_X1 U14535 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n14150) );
  NAND2_X1 U14536 ( .A1(n12482), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12484) );
  NAND2_X1 U14537 ( .A1(n11176), .A2(n11177), .ZN(n11178) );
  NAND2_X1 U14538 ( .A1(n12500), .A2(n11178), .ZN(n15761) );
  NAND2_X1 U14539 ( .A1(n20408), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12461) );
  NAND2_X1 U14540 ( .A1(n14157), .A2(n12461), .ZN(n13921) );
  AND2_X2 U14541 ( .A1(n15656), .A2(n20266), .ZN(n16423) );
  NAND2_X1 U14542 ( .A1(n16423), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11491) );
  NAND2_X1 U14543 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11179) );
  OAI211_X1 U14544 ( .C1(n15761), .C2(n16441), .A(n11491), .B(n11179), .ZN(
        n11180) );
  AOI21_X1 U14545 ( .B1(n11181), .B2(n16443), .A(n11180), .ZN(n11213) );
  XNOR2_X2 U14546 ( .A(n11184), .B(n11183), .ZN(n16429) );
  INV_X1 U14547 ( .A(n13917), .ZN(n11185) );
  NAND2_X1 U14548 ( .A1(n11185), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13919) );
  INV_X1 U14549 ( .A(n13919), .ZN(n11187) );
  XNOR2_X1 U14550 ( .A(n11265), .B(n11272), .ZN(n11188) );
  NAND2_X1 U14551 ( .A1(n11187), .A2(n11188), .ZN(n11189) );
  XNOR2_X1 U14552 ( .A(n13919), .B(n11188), .ZN(n13930) );
  NAND2_X1 U14553 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13930), .ZN(
        n13931) );
  NAND2_X1 U14554 ( .A1(n11189), .A2(n13931), .ZN(n11191) );
  XOR2_X1 U14555 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11191), .Z(
        n13958) );
  XNOR2_X1 U14556 ( .A(n11190), .B(n11282), .ZN(n13959) );
  NAND2_X1 U14557 ( .A1(n13958), .A2(n13959), .ZN(n11193) );
  NAND2_X1 U14558 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11191), .ZN(
        n11192) );
  NAND2_X1 U14559 ( .A1(n11193), .A2(n11192), .ZN(n11194) );
  XNOR2_X1 U14560 ( .A(n11194), .B(n16736), .ZN(n16449) );
  NAND2_X1 U14561 ( .A1(n11194), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11195) );
  NAND2_X1 U14562 ( .A1(n16429), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11197) );
  NAND2_X1 U14563 ( .A1(n11200), .A2(n11198), .ZN(n11199) );
  NAND2_X1 U14564 ( .A1(n11201), .A2(n10243), .ZN(n11203) );
  INV_X1 U14565 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11205) );
  INV_X1 U14566 ( .A(n11206), .ZN(n11207) );
  NAND4_X1 U14567 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U14568 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16615) );
  NOR2_X1 U14569 ( .A1(n11208), .A2(n16615), .ZN(n11482) );
  INV_X1 U14570 ( .A(n11482), .ZN(n16555) );
  INV_X1 U14571 ( .A(n11706), .ZN(n11211) );
  AND2_X1 U14572 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11209) );
  AND2_X1 U14573 ( .A1(n11482), .A2(n11209), .ZN(n11489) );
  AND2_X1 U14574 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16641) );
  NAND2_X1 U14575 ( .A1(n16641), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11475) );
  NOR2_X1 U14576 ( .A1(n11475), .A2(n11488), .ZN(n11210) );
  NAND2_X1 U14577 ( .A1(n11489), .A2(n11210), .ZN(n16537) );
  NAND2_X1 U14578 ( .A1(n11495), .A2(n16457), .ZN(n11212) );
  OAI211_X1 U14579 ( .C1(n11498), .C2(n16459), .A(n11213), .B(n11212), .ZN(
        P2_U2994) );
  INV_X1 U14580 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19726) );
  NOR2_X1 U14581 ( .A1(n19726), .A2(n20540), .ZN(n20533) );
  NAND2_X1 U14582 ( .A1(n16887), .A2(n20526), .ZN(n12534) );
  NAND2_X1 U14583 ( .A1(n19992), .A2(n14358), .ZN(n11234) );
  NAND2_X1 U14584 ( .A1(n11456), .A2(n11222), .ZN(n11221) );
  INV_X1 U14585 ( .A(n11218), .ZN(n11214) );
  NAND2_X1 U14586 ( .A1(n13987), .A2(n11214), .ZN(n11216) );
  NAND2_X1 U14587 ( .A1(n11218), .A2(n11217), .ZN(n11219) );
  NAND2_X1 U14588 ( .A1(n11225), .A2(n11219), .ZN(n11220) );
  INV_X1 U14589 ( .A(n11223), .ZN(n11224) );
  NAND2_X1 U14590 ( .A1(n11231), .A2(n11466), .ZN(n11227) );
  NAND2_X1 U14591 ( .A1(n11227), .A2(n20002), .ZN(n11233) );
  INV_X1 U14592 ( .A(n11228), .ZN(n11229) );
  NAND2_X1 U14593 ( .A1(n14168), .A2(n11229), .ZN(n11230) );
  NAND2_X1 U14594 ( .A1(n16844), .A2(n11232), .ZN(n14165) );
  MUX2_X1 U14595 ( .A(n11234), .B(n11233), .S(n14165), .Z(n11252) );
  MUX2_X1 U14596 ( .A(n10737), .B(n11464), .S(n13987), .Z(n11248) );
  INV_X1 U14597 ( .A(n16887), .ZN(n20532) );
  OR2_X1 U14598 ( .A1(n16847), .A2(n20532), .ZN(n13348) );
  NAND3_X1 U14599 ( .A1(n9894), .A2(n13910), .A3(n14358), .ZN(n11247) );
  NAND2_X1 U14600 ( .A1(n11235), .A2(n20022), .ZN(n11237) );
  NAND2_X1 U14601 ( .A1(n11237), .A2(n11236), .ZN(n11453) );
  AOI21_X1 U14602 ( .B1(n20002), .B2(n13987), .A(n16856), .ZN(n11238) );
  OAI21_X1 U14603 ( .B1(n11238), .B2(n13361), .A(n11464), .ZN(n11240) );
  AND3_X1 U14604 ( .A1(n11453), .A2(n11240), .A3(n11239), .ZN(n11246) );
  NAND2_X1 U14605 ( .A1(n11243), .A2(n11242), .ZN(n11244) );
  NAND2_X1 U14606 ( .A1(n14164), .A2(n11244), .ZN(n11245) );
  OAI21_X1 U14607 ( .B1(n11248), .B2(n13348), .A(n14360), .ZN(n11249) );
  NOR2_X1 U14608 ( .A1(n11099), .A2(n11253), .ZN(n20630) );
  NOR2_X1 U14609 ( .A1(n11255), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14610 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U14611 ( .A1(n12525), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11257) );
  INV_X1 U14612 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17446) );
  NAND2_X1 U14613 ( .A1(n13361), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11259) );
  OAI211_X1 U14614 ( .C1(n9588), .C2(n17446), .A(n11259), .B(n16814), .ZN(
        n11260) );
  INV_X1 U14615 ( .A(n11260), .ZN(n11261) );
  INV_X1 U14616 ( .A(n13353), .ZN(n11262) );
  NAND2_X1 U14617 ( .A1(n11267), .A2(n11262), .ZN(n11280) );
  INV_X1 U14618 ( .A(n11271), .ZN(n11263) );
  OAI21_X1 U14619 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n16814), .A(
        n11263), .ZN(n11264) );
  OAI211_X2 U14620 ( .C1(n11265), .C2(n11281), .A(n11280), .B(n11264), .ZN(
        n14268) );
  NAND2_X1 U14621 ( .A1(n14267), .A2(n14268), .ZN(n11276) );
  INV_X1 U14622 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20542) );
  NAND2_X1 U14623 ( .A1(n11266), .A2(P2_EAX_REG_1__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U14624 ( .A1(n11267), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11268) );
  OAI211_X1 U14625 ( .C1(n14727), .C2(n20542), .A(n11269), .B(n11268), .ZN(
        n11275) );
  XNOR2_X1 U14626 ( .A(n11276), .B(n11275), .ZN(n14152) );
  AND2_X1 U14627 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11270) );
  AOI21_X1 U14628 ( .B1(n11271), .B2(n13353), .A(n11270), .ZN(n11274) );
  NAND2_X1 U14629 ( .A1(n11426), .A2(n11272), .ZN(n11273) );
  AND2_X1 U14630 ( .A1(n11274), .A2(n11273), .ZN(n14151) );
  INV_X1 U14631 ( .A(n11275), .ZN(n11277) );
  NAND2_X1 U14632 ( .A1(n11277), .A2(n11276), .ZN(n11278) );
  NAND2_X1 U14633 ( .A1(n14154), .A2(n11278), .ZN(n11287) );
  NAND2_X1 U14634 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11279) );
  OAI211_X1 U14635 ( .C1(n11282), .C2(n11281), .A(n11280), .B(n11279), .ZN(
        n11285) );
  XNOR2_X1 U14636 ( .A(n11287), .B(n11285), .ZN(n14440) );
  AOI22_X1 U14637 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n11284) );
  NAND2_X1 U14638 ( .A1(n12525), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11283) );
  AND2_X1 U14639 ( .A1(n11284), .A2(n11283), .ZN(n14439) );
  INV_X1 U14640 ( .A(n11285), .ZN(n11286) );
  NAND2_X1 U14641 ( .A1(n11287), .A2(n11286), .ZN(n11288) );
  AOI22_X1 U14642 ( .A1(n11426), .A2(n11289), .B1(n12524), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14643 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11291) );
  NAND2_X1 U14644 ( .A1(n12525), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11290) );
  INV_X1 U14645 ( .A(n15938), .ZN(n11293) );
  INV_X1 U14646 ( .A(n15937), .ZN(n11302) );
  NAND2_X1 U14647 ( .A1(n11426), .A2(n11295), .ZN(n11297) );
  NAND2_X1 U14648 ( .A1(n12524), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n11296) );
  OAI211_X1 U14649 ( .C1(n11294), .C2(n16725), .A(n11297), .B(n11296), .ZN(
        n11298) );
  INV_X1 U14650 ( .A(n11298), .ZN(n11300) );
  NAND2_X1 U14651 ( .A1(n12525), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11299) );
  AND2_X1 U14652 ( .A1(n11300), .A2(n11299), .ZN(n16172) );
  NAND2_X1 U14653 ( .A1(n11302), .A2(n11301), .ZN(n16169) );
  INV_X1 U14654 ( .A(n16169), .ZN(n11311) );
  NAND2_X1 U14655 ( .A1(n11426), .A2(n11303), .ZN(n11305) );
  NAND2_X1 U14656 ( .A1(n12524), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n11304) );
  OAI211_X1 U14657 ( .C1(n11294), .C2(n11472), .A(n11305), .B(n11304), .ZN(
        n11306) );
  INV_X1 U14658 ( .A(n11306), .ZN(n11308) );
  NAND2_X1 U14659 ( .A1(n12525), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11307) );
  AND2_X1 U14660 ( .A1(n11308), .A2(n11307), .ZN(n16171) );
  INV_X1 U14661 ( .A(n16171), .ZN(n11310) );
  AOI21_X1 U14662 ( .B1(n11311), .B2(n11310), .A(n10609), .ZN(n11312) );
  INV_X1 U14663 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20550) );
  NAND2_X1 U14664 ( .A1(n12524), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U14665 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11313) );
  OAI211_X1 U14666 ( .C1(n14727), .C2(n20550), .A(n11314), .B(n11313), .ZN(
        n14583) );
  AOI21_X1 U14667 ( .B1(n14582), .B2(n14583), .A(n10600), .ZN(n11315) );
  INV_X1 U14668 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20552) );
  NAND2_X1 U14669 ( .A1(n12524), .A2(P2_EAX_REG_7__SCAN_IN), .ZN(n11317) );
  NAND2_X1 U14670 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11316) );
  OAI211_X1 U14671 ( .C1(n14727), .C2(n20552), .A(n11317), .B(n11316), .ZN(
        n14575) );
  INV_X1 U14672 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20554) );
  NOR2_X1 U14673 ( .A1(n14727), .A2(n20554), .ZN(n11332) );
  AOI22_X1 U14674 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14675 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14676 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14677 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11318) );
  NAND4_X1 U14678 ( .A1(n11321), .A2(n11320), .A3(n11319), .A4(n11318), .ZN(
        n11327) );
  AOI22_X1 U14679 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14680 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14681 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14682 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n10908), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11322) );
  NAND4_X1 U14683 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11326) );
  NAND2_X1 U14684 ( .A1(n11426), .A2(n14595), .ZN(n11329) );
  NAND2_X1 U14685 ( .A1(n12524), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n11328) );
  OAI211_X1 U14686 ( .C1(n11294), .C2(n11330), .A(n11329), .B(n11328), .ZN(
        n11331) );
  NOR2_X1 U14687 ( .A1(n11332), .A2(n11331), .ZN(n14562) );
  INV_X1 U14688 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20556) );
  NOR2_X1 U14689 ( .A1(n14727), .A2(n20556), .ZN(n11346) );
  AOI22_X1 U14690 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10948), .B1(
        n10947), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14691 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14692 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14693 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11333) );
  NAND4_X1 U14694 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(
        n11342) );
  AOI22_X1 U14695 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14696 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11339) );
  INV_X1 U14697 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n21485) );
  AOI22_X1 U14698 ( .A1(n10908), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14699 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11337) );
  NAND4_X1 U14700 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n11341) );
  NAND2_X1 U14701 ( .A1(n11426), .A2(n14600), .ZN(n11344) );
  NAND2_X1 U14702 ( .A1(n12524), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n11343) );
  OAI211_X1 U14703 ( .C1(n11294), .C2(n16638), .A(n11344), .B(n11343), .ZN(
        n11345) );
  NOR2_X1 U14704 ( .A1(n11346), .A2(n11345), .ZN(n14565) );
  NAND2_X1 U14705 ( .A1(n12525), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14706 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10873), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14707 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14708 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14709 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11347) );
  NAND4_X1 U14710 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n11356) );
  AOI22_X1 U14711 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14712 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10908), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14713 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10882), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14714 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10931), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11351) );
  NAND4_X1 U14715 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11355) );
  NAND2_X1 U14716 ( .A1(n11426), .A2(n19854), .ZN(n11359) );
  NAND2_X1 U14717 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11358) );
  NAND2_X1 U14718 ( .A1(n12524), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n11357) );
  NAND4_X1 U14719 ( .A1(n11360), .A2(n11359), .A3(n11358), .A4(n11357), .ZN(
        n14550) );
  NAND2_X1 U14720 ( .A1(n14548), .A2(n14550), .ZN(n14549) );
  AOI22_X1 U14721 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U14722 ( .A1(n12525), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14723 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14724 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14725 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14726 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11361) );
  NAND4_X1 U14727 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11370) );
  AOI22_X1 U14728 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14729 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14730 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14731 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11365) );
  NAND4_X1 U14732 ( .A1(n11368), .A2(n11367), .A3(n11366), .A4(n11365), .ZN(
        n11369) );
  NAND2_X1 U14733 ( .A1(n11426), .A2(n16062), .ZN(n11371) );
  INV_X1 U14734 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20562) );
  NOR2_X1 U14735 ( .A1(n14727), .A2(n20562), .ZN(n11387) );
  AOI22_X1 U14736 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10873), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14737 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14738 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14739 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11374) );
  NAND4_X1 U14740 ( .A1(n11377), .A2(n11376), .A3(n11375), .A4(n11374), .ZN(
        n11383) );
  AOI22_X1 U14741 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14742 ( .A1(n10948), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14743 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10931), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14744 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10908), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11378) );
  NAND4_X1 U14745 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n11382) );
  OR2_X1 U14746 ( .A1(n11383), .A2(n11382), .ZN(n16058) );
  NAND2_X1 U14747 ( .A1(n11426), .A2(n16058), .ZN(n11385) );
  NAND2_X1 U14748 ( .A1(n12524), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n11384) );
  OAI211_X1 U14749 ( .C1(n11294), .C2(n16632), .A(n11385), .B(n11384), .ZN(
        n11386) );
  NOR2_X1 U14750 ( .A1(n11387), .A2(n11386), .ZN(n14572) );
  NAND2_X1 U14751 ( .A1(n12525), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14752 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14753 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14754 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14755 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11388) );
  NAND4_X1 U14756 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n11397) );
  AOI22_X1 U14757 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14758 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14759 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14760 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11392) );
  NAND4_X1 U14761 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(
        n11396) );
  NAND2_X1 U14762 ( .A1(n11426), .A2(n14616), .ZN(n11400) );
  NAND2_X1 U14763 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11399) );
  NAND2_X1 U14764 ( .A1(n12524), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U14765 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n14579) );
  NAND2_X1 U14766 ( .A1(n12525), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14767 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10948), .B1(
        n10846), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14768 ( .A1(n10881), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14769 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10908), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14770 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10847), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11402) );
  NAND4_X1 U14771 ( .A1(n11405), .A2(n11404), .A3(n11403), .A4(n11402), .ZN(
        n11411) );
  AOI22_X1 U14772 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14773 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14774 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14775 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11406) );
  NAND4_X1 U14776 ( .A1(n11409), .A2(n11408), .A3(n11407), .A4(n11406), .ZN(
        n11410) );
  NAND2_X1 U14777 ( .A1(n11426), .A2(n14620), .ZN(n11414) );
  NAND2_X1 U14778 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11413) );
  NAND2_X1 U14779 ( .A1(n12524), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n11412) );
  NAND4_X1 U14780 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11412), .ZN(
        n14586) );
  NAND2_X1 U14781 ( .A1(n14578), .A2(n14586), .ZN(n14585) );
  INV_X1 U14782 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20568) );
  NOR2_X1 U14783 ( .A1(n14727), .A2(n20568), .ZN(n11430) );
  AOI22_X1 U14784 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14785 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14786 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14787 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11416) );
  NAND4_X1 U14788 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n11425) );
  AOI22_X1 U14789 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14790 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14791 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14792 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11420) );
  NAND4_X1 U14793 ( .A1(n11423), .A2(n11422), .A3(n11421), .A4(n11420), .ZN(
        n11424) );
  NAND2_X1 U14794 ( .A1(n11426), .A2(n19847), .ZN(n11428) );
  NAND2_X1 U14795 ( .A1(n12524), .A2(P2_EAX_REG_15__SCAN_IN), .ZN(n11427) );
  OAI211_X1 U14796 ( .C1(n11294), .C2(n16568), .A(n11428), .B(n11427), .ZN(
        n11429) );
  NOR2_X1 U14797 ( .A1(n11430), .A2(n11429), .ZN(n14641) );
  AOI22_X1 U14798 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n11432) );
  NAND2_X1 U14799 ( .A1(n12525), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11431) );
  INV_X1 U14800 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20572) );
  NAND2_X1 U14801 ( .A1(n12524), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n11434) );
  NAND2_X1 U14802 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11433) );
  OAI211_X1 U14803 ( .C1(n14727), .C2(n20572), .A(n11434), .B(n11433), .ZN(
        n15799) );
  INV_X1 U14804 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20573) );
  NAND2_X1 U14805 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11436) );
  NAND2_X1 U14806 ( .A1(n12524), .A2(P2_EAX_REG_18__SCAN_IN), .ZN(n11435) );
  OAI211_X1 U14807 ( .C1(n14727), .C2(n20573), .A(n11436), .B(n11435), .ZN(
        n15784) );
  INV_X1 U14808 ( .A(n11700), .ZN(n11440) );
  AOI22_X1 U14809 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U14810 ( .A1(n12525), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11437) );
  NAND2_X1 U14811 ( .A1(n11440), .A2(n11439), .ZN(n11441) );
  INV_X1 U14812 ( .A(n11795), .ZN(n11443) );
  AOI21_X1 U14813 ( .B1(n11444), .B2(n11703), .A(n11443), .ZN(n16139) );
  NAND2_X1 U14814 ( .A1(n9758), .A2(n11445), .ZN(n16845) );
  NAND2_X1 U14815 ( .A1(n16840), .A2(n14164), .ZN(n16848) );
  NAND2_X1 U14816 ( .A1(n16848), .A2(n11232), .ZN(n11446) );
  NAND2_X1 U14817 ( .A1(n16845), .A2(n11446), .ZN(n11447) );
  AND2_X1 U14818 ( .A1(n13987), .A2(n20006), .ZN(n11448) );
  NAND2_X1 U14819 ( .A1(n11494), .A2(n14351), .ZN(n19956) );
  NAND2_X1 U14820 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19958) );
  INV_X1 U14821 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11450) );
  AND2_X1 U14822 ( .A1(n19958), .A2(n11450), .ZN(n19940) );
  INV_X1 U14823 ( .A(n19940), .ZN(n11451) );
  NOR2_X1 U14824 ( .A1(n19958), .A2(n11450), .ZN(n19939) );
  AOI21_X1 U14825 ( .B1(n16565), .B2(n11451), .A(n19939), .ZN(n16735) );
  NOR2_X1 U14826 ( .A1(n16735), .A2(n16736), .ZN(n16713) );
  NAND2_X1 U14827 ( .A1(n11452), .A2(n11232), .ZN(n14699) );
  NAND2_X1 U14828 ( .A1(n14699), .A2(n11453), .ZN(n11454) );
  NAND2_X1 U14829 ( .A1(n11454), .A2(n19997), .ZN(n11469) );
  AND2_X1 U14830 ( .A1(n11456), .A2(n11464), .ZN(n11457) );
  NAND2_X1 U14831 ( .A1(n11458), .A2(n11457), .ZN(n13351) );
  OAI21_X1 U14832 ( .B1(n11459), .B2(n15652), .A(n13351), .ZN(n11460) );
  NOR2_X1 U14833 ( .A1(n11460), .A2(n9613), .ZN(n11468) );
  OAI21_X1 U14834 ( .B1(n9722), .B2(n11461), .A(n15652), .ZN(n11463) );
  NAND2_X1 U14835 ( .A1(n11463), .A2(n11462), .ZN(n11465) );
  MUX2_X1 U14836 ( .A(n11466), .B(n11465), .S(n11464), .Z(n11467) );
  NAND3_X1 U14837 ( .A1(n11469), .A2(n11468), .A3(n11467), .ZN(n14702) );
  NAND2_X1 U14838 ( .A1(n11494), .A2(n11471), .ZN(n19954) );
  NAND2_X1 U14839 ( .A1(n16713), .A2(n9852), .ZN(n16724) );
  NAND2_X1 U14840 ( .A1(n11477), .A2(n16704), .ZN(n16701) );
  AOI21_X1 U14841 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n19970), .ZN(n16714) );
  NOR2_X1 U14842 ( .A1(n16714), .A2(n16727), .ZN(n16705) );
  NAND2_X1 U14843 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16682) );
  INV_X1 U14844 ( .A(n16682), .ZN(n11473) );
  OR2_X1 U14845 ( .A1(n19970), .A2(n11473), .ZN(n11474) );
  INV_X1 U14846 ( .A(n11475), .ZN(n16295) );
  OR2_X1 U14847 ( .A1(n19970), .A2(n16295), .ZN(n11476) );
  NOR2_X1 U14848 ( .A1(n16615), .A2(n16598), .ZN(n16566) );
  OR2_X1 U14849 ( .A1(n16616), .A2(n16566), .ZN(n11478) );
  NAND2_X1 U14850 ( .A1(n16633), .A2(n11478), .ZN(n16605) );
  INV_X1 U14851 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16585) );
  NOR3_X1 U14852 ( .A1(n16568), .A2(n16585), .A3(n16577), .ZN(n11479) );
  NOR2_X1 U14853 ( .A1(n19970), .A2(n11479), .ZN(n11480) );
  OR2_X1 U14854 ( .A1(n19970), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11481) );
  NAND3_X1 U14855 ( .A1(n11482), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n11707), .ZN(n11483) );
  OR2_X1 U14856 ( .A1(n16616), .A2(n11483), .ZN(n11695) );
  NAND2_X1 U14857 ( .A1(n16759), .A2(n13987), .ZN(n11486) );
  NAND2_X1 U14858 ( .A1(n11484), .A2(n11486), .ZN(n11487) );
  INV_X1 U14859 ( .A(n16616), .ZN(n16629) );
  NAND3_X1 U14860 ( .A1(n16629), .A2(n11489), .A3(n11488), .ZN(n11490) );
  OAI211_X1 U14861 ( .C1(n16034), .C2(n19964), .A(n11491), .B(n11490), .ZN(
        n11492) );
  AOI211_X1 U14862 ( .C1(n16139), .C2(n19960), .A(n9611), .B(n11492), .ZN(
        n11497) );
  INV_X1 U14863 ( .A(n11493), .ZN(n20632) );
  NAND2_X1 U14864 ( .A1(n11495), .A2(n19946), .ZN(n11496) );
  OAI211_X1 U14865 ( .C1(n11498), .C2(n19974), .A(n11497), .B(n11496), .ZN(
        P2_U3026) );
  NAND2_X1 U14866 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17033) );
  NOR2_X1 U14867 ( .A1(n17033), .A2(n17035), .ZN(n17034) );
  NOR2_X2 U14868 ( .A1(n17793), .A2(n17783), .ZN(n17743) );
  NAND2_X1 U14869 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17744) );
  NAND2_X1 U14870 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18678) );
  NAND2_X1 U14871 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18642) );
  NAND2_X1 U14872 ( .A1(n18630), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18597) );
  NAND2_X1 U14873 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18599) );
  NAND2_X1 U14874 ( .A1(n18581), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11501) );
  NAND2_X1 U14875 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18553) );
  NOR2_X2 U14876 ( .A1(n11501), .A2(n18553), .ZN(n16973) );
  NAND2_X1 U14877 ( .A1(n16973), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14878 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16963) );
  INV_X1 U14879 ( .A(n11520), .ZN(n11499) );
  XNOR2_X1 U14880 ( .A(n11499), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17566) );
  INV_X1 U14881 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18543) );
  OR2_X1 U14882 ( .A1(n18821), .A2(n11500), .ZN(n11517) );
  NOR2_X1 U14883 ( .A1(n18543), .A2(n11517), .ZN(n11516) );
  NOR2_X1 U14884 ( .A1(n16963), .A2(n11517), .ZN(n16917) );
  INV_X1 U14885 ( .A(n16917), .ZN(n11521) );
  OAI21_X1 U14886 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11516), .A(
        n11521), .ZN(n16966) );
  INV_X1 U14887 ( .A(n16966), .ZN(n17589) );
  NOR2_X1 U14888 ( .A1(n18821), .A2(n11501), .ZN(n11505) );
  INV_X1 U14889 ( .A(n11505), .ZN(n11513) );
  NOR2_X1 U14890 ( .A1(n18553), .A2(n11513), .ZN(n11503) );
  OAI21_X1 U14891 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n11503), .A(
        n11517), .ZN(n11502) );
  INV_X1 U14892 ( .A(n11502), .ZN(n17610) );
  INV_X1 U14893 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18568) );
  NOR2_X1 U14894 ( .A1(n18568), .A2(n11513), .ZN(n11512) );
  INV_X1 U14895 ( .A(n11503), .ZN(n16961) );
  OAI21_X1 U14896 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n11512), .A(
        n16961), .ZN(n18555) );
  INV_X1 U14897 ( .A(n18555), .ZN(n17618) );
  INV_X1 U14898 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18583) );
  INV_X1 U14899 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17662) );
  INV_X1 U14900 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11507) );
  NOR2_X1 U14901 ( .A1(n18821), .A2(n11504), .ZN(n16984) );
  INV_X1 U14902 ( .A(n16984), .ZN(n17707) );
  NOR2_X1 U14903 ( .A1(n18642), .A2(n17707), .ZN(n18593) );
  INV_X1 U14904 ( .A(n18593), .ZN(n17690) );
  NOR2_X1 U14905 ( .A1(n11507), .A2(n17690), .ZN(n11506) );
  NAND2_X1 U14906 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11506), .ZN(
        n11510) );
  NOR2_X1 U14907 ( .A1(n17662), .A2(n11510), .ZN(n11509) );
  INV_X1 U14908 ( .A(n11509), .ZN(n18551) );
  AOI21_X1 U14909 ( .B1(n18583), .B2(n18551), .A(n11505), .ZN(n18579) );
  OAI21_X1 U14910 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11506), .A(
        n11510), .ZN(n18609) );
  INV_X1 U14911 ( .A(n18609), .ZN(n17665) );
  AOI21_X1 U14912 ( .B1(n11507), .B2(n17690), .A(n11506), .ZN(n18639) );
  NOR2_X1 U14913 ( .A1(n18821), .A2(n18671), .ZN(n18673) );
  NAND2_X1 U14914 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18673), .ZN(
        n17731) );
  NOR2_X1 U14915 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17731), .ZN(
        n17719) );
  NOR2_X1 U14916 ( .A1(n17663), .A2(n17882), .ZN(n17656) );
  INV_X1 U14917 ( .A(n17656), .ZN(n11511) );
  AOI21_X1 U14918 ( .B1(n17662), .B2(n11510), .A(n11509), .ZN(n18596) );
  NAND2_X1 U14919 ( .A1(n11511), .A2(n18601), .ZN(n17654) );
  AOI21_X1 U14920 ( .B1(n18568), .B2(n11513), .A(n11512), .ZN(n18564) );
  NAND2_X1 U14921 ( .A1(n11515), .A2(n11514), .ZN(n17631) );
  INV_X1 U14922 ( .A(n17598), .ZN(n11519) );
  AOI21_X1 U14923 ( .B1(n18543), .B2(n11517), .A(n11516), .ZN(n18538) );
  INV_X1 U14924 ( .A(n18538), .ZN(n11518) );
  NAND2_X1 U14925 ( .A1(n11519), .A2(n11518), .ZN(n17596) );
  AOI21_X1 U14926 ( .B1(n17577), .B2(n11521), .A(n11520), .ZN(n17576) );
  INV_X1 U14927 ( .A(n17576), .ZN(n11522) );
  NOR3_X1 U14928 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n19601) );
  AOI22_X1 U14929 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11530) );
  INV_X2 U14930 ( .A(n18200), .ZN(n18235) );
  AOI22_X1 U14931 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11529) );
  INV_X2 U14932 ( .A(n18198), .ZN(n18248) );
  AOI22_X1 U14933 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17281), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11528) );
  AND2_X2 U14934 ( .A1(n11525), .A2(n11532), .ZN(n11607) );
  AND2_X2 U14935 ( .A1(n14401), .A2(n11526), .ZN(n11605) );
  AOI22_X1 U14936 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11527) );
  NAND4_X1 U14937 ( .A1(n11530), .A2(n11529), .A3(n11528), .A4(n11527), .ZN(
        n11542) );
  NAND2_X2 U14938 ( .A1(n14656), .A2(n14453), .ZN(n18251) );
  AOI22_X1 U14939 ( .A1(n11604), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11541) );
  INV_X1 U14940 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11537) );
  OAI22_X1 U14941 ( .A1(n18079), .A2(n11537), .B1(n11598), .B2(n18107), .ZN(
        n11538) );
  AOI211_X1 U14942 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n11539), .B(n11538), .ZN(n11540) );
  AOI22_X1 U14943 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11547) );
  BUF_X4 U14944 ( .A(n11543), .Z(n18236) );
  AOI22_X1 U14945 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14946 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14947 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14948 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11553) );
  INV_X1 U14949 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17263) );
  NAND2_X1 U14950 ( .A1(n18243), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11551) );
  NAND2_X1 U14951 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11550) );
  NAND4_X1 U14952 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11558) );
  INV_X1 U14953 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U14954 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11555) );
  NAND2_X1 U14955 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11554) );
  OAI211_X1 U14956 ( .C1(n18216), .C2(n11556), .A(n11555), .B(n11554), .ZN(
        n11557) );
  NOR2_X1 U14957 ( .A1(n11558), .A2(n11557), .ZN(n11559) );
  INV_X1 U14958 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18161) );
  NAND2_X1 U14959 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11562) );
  NAND2_X1 U14960 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11561) );
  OAI211_X1 U14961 ( .C1(n18216), .C2(n18161), .A(n11562), .B(n11561), .ZN(
        n11563) );
  INV_X1 U14962 ( .A(n11563), .ZN(n11567) );
  AOI22_X1 U14963 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11566) );
  INV_X2 U14964 ( .A(n18200), .ZN(n18219) );
  AOI22_X1 U14965 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18219), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11565) );
  NAND2_X1 U14966 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11564) );
  NAND4_X1 U14967 ( .A1(n11567), .A2(n11566), .A3(n11565), .A4(n11564), .ZN(
        n11573) );
  AOI22_X1 U14968 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14969 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14970 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14971 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11568) );
  NAND4_X1 U14972 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11572) );
  INV_X1 U14973 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18013) );
  NAND2_X1 U14974 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11575) );
  NAND2_X1 U14975 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11574) );
  OAI211_X1 U14976 ( .C1(n18216), .C2(n18013), .A(n11575), .B(n11574), .ZN(
        n11576) );
  INV_X1 U14977 ( .A(n11576), .ZN(n11580) );
  AOI22_X1 U14978 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14979 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U14980 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11577) );
  AOI22_X1 U14981 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14982 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14983 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14984 ( .A1(n19127), .A2(n19135), .ZN(n11641) );
  AOI22_X1 U14985 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14986 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14987 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14988 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14989 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11591) );
  INV_X1 U14990 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17233) );
  NAND2_X1 U14991 ( .A1(n18243), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11589) );
  NAND2_X1 U14992 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11588) );
  NAND4_X1 U14993 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n11595) );
  NAND2_X1 U14994 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11593) );
  NAND2_X1 U14995 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11592) );
  OAI211_X1 U14996 ( .C1(n18216), .C2(n18195), .A(n11593), .B(n11592), .ZN(
        n11594) );
  NOR2_X1 U14997 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  AOI22_X1 U14998 ( .A1(n17208), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9589), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14999 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U15000 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18219), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U15001 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17281), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11599) );
  NAND4_X1 U15002 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11613) );
  INV_X1 U15003 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17962) );
  AOI22_X1 U15004 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11611) );
  INV_X1 U15005 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11606) );
  INV_X1 U15006 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17961) );
  INV_X1 U15007 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17963) );
  OAI22_X1 U15008 ( .A1(n17954), .A2(n17961), .B1(n18196), .B2(n17963), .ZN(
        n11608) );
  AOI22_X1 U15009 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n17281), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U15010 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U15011 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U15012 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11614) );
  NAND4_X1 U15013 ( .A1(n11617), .A2(n11616), .A3(n11615), .A4(n11614), .ZN(
        n11623) );
  AOI22_X1 U15014 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U15015 ( .A1(n11604), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11619) );
  OAI211_X1 U15016 ( .C1(n18216), .C2(n11621), .A(n11620), .B(n11619), .ZN(
        n11622) );
  NOR2_X1 U15017 ( .A1(n19140), .A2(n19122), .ZN(n13627) );
  INV_X1 U15018 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11626) );
  NAND2_X1 U15019 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11625) );
  NAND2_X1 U15020 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11624) );
  OAI211_X1 U15021 ( .C1(n18251), .C2(n11626), .A(n11625), .B(n11624), .ZN(
        n11627) );
  INV_X1 U15022 ( .A(n11627), .ZN(n11631) );
  AOI22_X1 U15023 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U15024 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11629) );
  NAND2_X1 U15025 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11628) );
  NAND4_X1 U15026 ( .A1(n11631), .A2(n11630), .A3(n11629), .A4(n11628), .ZN(
        n11637) );
  AOI22_X1 U15027 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U15028 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U15029 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U15030 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11632) );
  NAND4_X1 U15031 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11636) );
  INV_X1 U15032 ( .A(n11643), .ZN(n11640) );
  OR2_X1 U15033 ( .A1(n19140), .A2(n14450), .ZN(n14147) );
  NAND3_X1 U15034 ( .A1(n19709), .A2(n18432), .A3(n14147), .ZN(n13578) );
  NOR2_X1 U15035 ( .A1(n9674), .A2(n11650), .ZN(n11647) );
  AOI21_X1 U15036 ( .B1(n19117), .B2(n19108), .A(n14450), .ZN(n11639) );
  AOI21_X1 U15037 ( .B1(n11641), .B2(n11640), .A(n11639), .ZN(n11646) );
  NOR2_X1 U15038 ( .A1(n19140), .A2(n11643), .ZN(n11644) );
  NOR2_X1 U15039 ( .A1(n9674), .A2(n13582), .ZN(n11642) );
  OAI22_X1 U15040 ( .A1(n19127), .A2(n11644), .B1(n11643), .B2(n11642), .ZN(
        n11645) );
  AOI211_X1 U15041 ( .C1(n11647), .C2(n19122), .A(n11646), .B(n11645), .ZN(
        n13577) );
  OAI211_X1 U15042 ( .C1(n19122), .C2(n11648), .A(n13578), .B(n13577), .ZN(
        n13628) );
  INV_X1 U15043 ( .A(n11650), .ZN(n11651) );
  NAND2_X1 U15044 ( .A1(n19117), .A2(n19122), .ZN(n14399) );
  NAND2_X1 U15045 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19592), .ZN(n19594) );
  MUX2_X1 U15046 ( .A(n11652), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13568) );
  NAND2_X1 U15047 ( .A1(n13568), .A2(n13569), .ZN(n11667) );
  NAND2_X1 U15048 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n11652), .ZN(
        n11654) );
  NAND2_X1 U15049 ( .A1(n11667), .A2(n11654), .ZN(n11665) );
  MUX2_X1 U15050 ( .A(n19568), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11664) );
  NAND2_X1 U15051 ( .A1(n11665), .A2(n11664), .ZN(n11656) );
  NAND2_X1 U15052 ( .A1(n19568), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11655) );
  NAND2_X1 U15053 ( .A1(n11656), .A2(n11655), .ZN(n11657) );
  NAND2_X1 U15054 ( .A1(n11657), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11661) );
  OAI22_X1 U15055 ( .A1(n11657), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19571), .ZN(n11659) );
  AOI21_X1 U15056 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11661), .A(
        n11659), .ZN(n11658) );
  NAND2_X1 U15057 ( .A1(n11659), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11663) );
  NOR2_X1 U15058 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19571), .ZN(
        n11660) );
  NAND2_X1 U15059 ( .A1(n11661), .A2(n11660), .ZN(n11662) );
  NAND2_X1 U15060 ( .A1(n11663), .A2(n11662), .ZN(n13572) );
  XNOR2_X1 U15061 ( .A(n11665), .B(n11664), .ZN(n11666) );
  OAI21_X1 U15062 ( .B1(n13569), .B2(n13568), .A(n11667), .ZN(n11668) );
  NAND2_X1 U15063 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18494), .ZN(n11670) );
  AOI211_X4 U15064 ( .C1(n21509), .C2(n19710), .A(n11678), .B(n11670), .ZN(
        n17887) );
  NAND2_X1 U15065 ( .A1(n17896), .A2(n18269), .ZN(n17886) );
  NOR2_X1 U15066 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17886), .ZN(n17873) );
  INV_X1 U15067 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18158) );
  NAND2_X1 U15068 ( .A1(n17873), .A2(n18158), .ZN(n17863) );
  NOR2_X1 U15069 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17863), .ZN(n17844) );
  NAND2_X1 U15070 ( .A1(n17844), .A2(n18255), .ZN(n17834) );
  NAND2_X1 U15071 ( .A1(n17811), .A2(n18231), .ZN(n17798) );
  INV_X1 U15072 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n18188) );
  NAND2_X1 U15073 ( .A1(n17797), .A2(n18188), .ZN(n17790) );
  NAND2_X1 U15074 ( .A1(n17773), .A2(n17764), .ZN(n17760) );
  INV_X1 U15075 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17738) );
  NAND2_X1 U15076 ( .A1(n17747), .A2(n17738), .ZN(n17737) );
  INV_X1 U15077 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17710) );
  NAND2_X1 U15078 ( .A1(n17721), .A2(n17710), .ZN(n17709) );
  INV_X1 U15079 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17686) );
  NAND2_X1 U15080 ( .A1(n17700), .A2(n17686), .ZN(n17684) );
  INV_X1 U15081 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18037) );
  NAND2_X1 U15082 ( .A1(n17672), .A2(n18037), .ZN(n17669) );
  INV_X1 U15083 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17645) );
  NAND2_X1 U15084 ( .A1(n17653), .A2(n17645), .ZN(n17644) );
  INV_X1 U15085 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17623) );
  NAND2_X1 U15086 ( .A1(n17630), .A2(n17623), .ZN(n17622) );
  INV_X1 U15087 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17936) );
  NAND2_X1 U15088 ( .A1(n17608), .A2(n17936), .ZN(n17602) );
  INV_X1 U15089 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17982) );
  NAND2_X1 U15090 ( .A1(n17586), .A2(n17982), .ZN(n11680) );
  NAND2_X1 U15091 ( .A1(n17887), .A2(n11680), .ZN(n17583) );
  INV_X1 U15092 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19670) );
  INV_X1 U15093 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19666) );
  INV_X1 U15094 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19607) );
  NOR2_X1 U15095 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n17544) );
  INV_X1 U15096 ( .A(n17544), .ZN(n11671) );
  NAND3_X1 U15097 ( .A1(n19615), .A2(n19678), .A3(n11671), .ZN(n19708) );
  AOI211_X1 U15098 ( .C1(n19708), .C2(n19709), .A(n19705), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n11679) );
  INV_X1 U15099 ( .A(n11679), .ZN(n19580) );
  INV_X1 U15100 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19663) );
  INV_X1 U15101 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19640) );
  INV_X1 U15102 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19633) );
  INV_X1 U15103 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19624) );
  NAND3_X1 U15104 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17892) );
  NOR2_X1 U15105 ( .A1(n19624), .A2(n17892), .ZN(n17871) );
  NAND2_X1 U15106 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17871), .ZN(n17833) );
  NOR2_X1 U15107 ( .A1(n19628), .A2(n17833), .ZN(n17839) );
  NAND2_X1 U15108 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17839), .ZN(n17824) );
  NOR2_X1 U15109 ( .A1(n19633), .A2(n17824), .ZN(n17781) );
  NAND4_X1 U15110 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17781), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n17775) );
  NOR2_X1 U15111 ( .A1(n19640), .A2(n17775), .ZN(n17763) );
  NAND3_X1 U15112 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17763), .ZN(n17651) );
  INV_X1 U15113 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19654) );
  INV_X1 U15114 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19652) );
  INV_X1 U15115 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19650) );
  INV_X1 U15116 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19648) );
  INV_X1 U15117 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19646) );
  NOR3_X1 U15118 ( .A1(n19650), .A2(n19648), .A3(n19646), .ZN(n17695) );
  INV_X1 U15119 ( .A(n17695), .ZN(n17683) );
  NOR3_X1 U15120 ( .A1(n19654), .A2(n19652), .A3(n17683), .ZN(n17678) );
  NAND2_X1 U15121 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17678), .ZN(n17652) );
  NOR3_X1 U15122 ( .A1(n19658), .A2(n17651), .A3(n17652), .ZN(n17649) );
  NAND2_X1 U15123 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17649), .ZN(n17637) );
  NOR2_X1 U15124 ( .A1(n19663), .A2(n17637), .ZN(n17628) );
  NAND3_X1 U15125 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17915), .A3(n17628), 
        .ZN(n17619) );
  NOR2_X1 U15126 ( .A1(n19666), .A2(n17619), .ZN(n17607) );
  NAND2_X1 U15127 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n17607), .ZN(n17605) );
  NOR2_X1 U15128 ( .A1(n19670), .A2(n17605), .ZN(n17585) );
  NAND3_X1 U15129 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n17585), .ZN(n17563) );
  NOR2_X1 U15130 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17563), .ZN(n17567) );
  NAND2_X1 U15131 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n11677) );
  NAND2_X1 U15132 ( .A1(n19582), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19478) );
  OR2_X1 U15133 ( .A1(n19594), .A2(n19478), .ZN(n19586) );
  INV_X1 U15134 ( .A(n19586), .ZN(n11674) );
  NOR2_X1 U15135 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n11672) );
  NAND2_X1 U15136 ( .A1(n18988), .A2(n17879), .ZN(n11673) );
  NOR2_X1 U15137 ( .A1(n11674), .A2(n11673), .ZN(n11675) );
  INV_X1 U15138 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19664) );
  INV_X1 U15139 ( .A(n17924), .ZN(n17932) );
  NAND2_X1 U15140 ( .A1(n17628), .A2(n17932), .ZN(n17629) );
  NOR3_X1 U15141 ( .A1(n19666), .A2(n19664), .A3(n17629), .ZN(n11676) );
  AOI21_X1 U15142 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n11676), .A(n17650), 
        .ZN(n17606) );
  AOI221_X1 U15143 ( .B1(n11677), .B2(n17930), .C1(n19670), .C2(n17930), .A(
        n17606), .ZN(n17578) );
  INV_X1 U15144 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19677) );
  INV_X1 U15145 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n21480) );
  OAI22_X1 U15146 ( .A1(n17578), .A2(n19677), .B1(n21480), .B2(n17918), .ZN(
        n11683) );
  AOI211_X4 U15147 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18494), .A(n11679), .B(
        n11678), .ZN(n17916) );
  NOR2_X1 U15148 ( .A1(n17928), .A2(n11680), .ZN(n17570) );
  OAI21_X1 U15149 ( .B1(n17916), .B2(n17570), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n11681) );
  INV_X1 U15150 ( .A(n11681), .ZN(n11682) );
  INV_X1 U15151 ( .A(n11754), .ZN(n11687) );
  NOR2_X2 U15152 ( .A1(n11688), .A2(n11687), .ZN(n16291) );
  NAND2_X1 U15153 ( .A1(n11756), .A2(n11742), .ZN(n16292) );
  OAI21_X1 U15154 ( .B1(n16291), .B2(n16292), .A(n11756), .ZN(n16284) );
  INV_X1 U15155 ( .A(n16281), .ZN(n11689) );
  AOI21_X1 U15156 ( .B1(n16284), .B2(n16282), .A(n11689), .ZN(n11692) );
  NAND2_X1 U15157 ( .A1(n11743), .A2(n11690), .ZN(n11691) );
  XNOR2_X1 U15158 ( .A(n11692), .B(n11691), .ZN(n16279) );
  OR2_X1 U15159 ( .A1(n9653), .A2(n11693), .ZN(n11694) );
  NAND2_X1 U15160 ( .A1(n11173), .A2(n11694), .ZN(n16276) );
  AND2_X1 U15161 ( .A1(n16423), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16272) );
  INV_X1 U15162 ( .A(n16272), .ZN(n11696) );
  OAI211_X1 U15163 ( .C1(n16276), .C2(n19964), .A(n11696), .B(n11695), .ZN(
        n11697) );
  AOI21_X1 U15164 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n11698), .A(
        n11697), .ZN(n11699) );
  INV_X1 U15165 ( .A(n11699), .ZN(n11705) );
  NAND2_X1 U15166 ( .A1(n11700), .A2(n11701), .ZN(n11702) );
  NAND2_X1 U15167 ( .A1(n11703), .A2(n11702), .ZN(n16151) );
  NOR2_X1 U15168 ( .A1(n16151), .A2(n19949), .ZN(n11704) );
  INV_X1 U15169 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16541) );
  OR2_X1 U15170 ( .A1(n16537), .A2(n16541), .ZN(n11735) );
  NAND3_X1 U15171 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11738) );
  NAND2_X1 U15172 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11714) );
  NAND2_X1 U15173 ( .A1(n12555), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U15174 ( .A1(n11720), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11712) );
  INV_X1 U15175 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11717) );
  NAND2_X1 U15176 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11716) );
  AOI22_X1 U15177 ( .A1(n11720), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11715) );
  OAI211_X1 U15178 ( .C1(n11717), .C2(n13776), .A(n11716), .B(n11715), .ZN(
        n16020) );
  AND2_X2 U15179 ( .A1(n15747), .A2(n16020), .ZN(n15731) );
  INV_X1 U15180 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n15738) );
  NAND2_X1 U15181 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11719) );
  AOI22_X1 U15182 ( .A1(n11720), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11718) );
  OAI211_X1 U15183 ( .C1(n15738), .C2(n13776), .A(n11719), .B(n11718), .ZN(
        n15732) );
  NAND2_X1 U15184 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11723) );
  NAND2_X1 U15185 ( .A1(n12555), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U15186 ( .A1(n11720), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11721) );
  NAND2_X1 U15187 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11726) );
  NAND2_X1 U15188 ( .A1(n12555), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U15189 ( .A1(n13774), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11724) );
  NAND2_X1 U15190 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11728) );
  AOI22_X1 U15191 ( .A1(n13774), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11727) );
  OAI211_X1 U15192 ( .C1(n16001), .C2(n13776), .A(n11728), .B(n11727), .ZN(
        n15687) );
  NAND2_X1 U15193 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U15194 ( .A1(n12555), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U15195 ( .A1(n13774), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11729) );
  NAND2_X1 U15196 ( .A1(n11732), .A2(n11733), .ZN(n11734) );
  INV_X1 U15197 ( .A(n11735), .ZN(n16234) );
  INV_X1 U15198 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16515) );
  NOR2_X1 U15199 ( .A1(n10013), .A2(n16515), .ZN(n16510) );
  NAND3_X1 U15200 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11736) );
  OR2_X1 U15201 ( .A1(n16474), .A2(n11736), .ZN(n11737) );
  NAND2_X1 U15202 ( .A1(n11737), .A2(n16475), .ZN(n13721) );
  INV_X1 U15203 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13722) );
  NAND2_X1 U15204 ( .A1(n16665), .A2(n16234), .ZN(n16498) );
  NAND2_X1 U15205 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11739) );
  NAND2_X1 U15206 ( .A1(n16463), .A2(n13722), .ZN(n13720) );
  NAND2_X1 U15207 ( .A1(n16423), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n16206) );
  OAI211_X1 U15208 ( .C1(n13721), .C2(n13722), .A(n13720), .B(n16206), .ZN(
        n11740) );
  AOI21_X1 U15209 ( .B1(n16210), .B2(n19944), .A(n11740), .ZN(n11817) );
  AND4_X1 U15210 ( .A1(n16306), .A2(n11741), .A3(n16323), .A4(n16330), .ZN(
        n11744) );
  AND4_X1 U15211 ( .A1(n16282), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11752) );
  INV_X1 U15212 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n16035) );
  INV_X1 U15213 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11746) );
  INV_X1 U15214 ( .A(n11745), .ZN(n11748) );
  NOR2_X1 U15215 ( .A1(n20006), .A2(n11746), .ZN(n11747) );
  AOI21_X1 U15216 ( .B1(n11748), .B2(n11747), .A(n11778), .ZN(n11749) );
  NAND2_X1 U15217 ( .A1(n11763), .A2(n11749), .ZN(n15750) );
  NOR2_X1 U15218 ( .A1(n15750), .A2(n13768), .ZN(n11753) );
  INV_X1 U15219 ( .A(n11753), .ZN(n11750) );
  NAND2_X1 U15220 ( .A1(n11750), .A2(n16541), .ZN(n16261) );
  NAND2_X1 U15221 ( .A1(n11753), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16262) );
  AND4_X1 U15222 ( .A1(n16307), .A2(n16342), .A3(n16331), .A4(n16345), .ZN(
        n11755) );
  AND4_X1 U15223 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n16322), .ZN(
        n11759) );
  AND4_X1 U15224 ( .A1(n16262), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n11760) );
  NAND2_X1 U15225 ( .A1(n13390), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11761) );
  INV_X1 U15226 ( .A(n11761), .ZN(n11762) );
  NAND2_X1 U15227 ( .A1(n11763), .A2(n11762), .ZN(n11764) );
  NAND2_X1 U15228 ( .A1(n11767), .A2(n11764), .ZN(n17306) );
  OR2_X1 U15229 ( .A1(n17306), .A2(n13768), .ZN(n11765) );
  NAND2_X1 U15230 ( .A1(n11765), .A2(n10013), .ZN(n16253) );
  OR3_X1 U15231 ( .A1(n17306), .A2(n13768), .A3(n10013), .ZN(n16252) );
  INV_X1 U15232 ( .A(n16252), .ZN(n11766) );
  NOR2_X1 U15233 ( .A1(n20006), .A2(n15738), .ZN(n11768) );
  NAND2_X1 U15234 ( .A1(n11767), .A2(n11768), .ZN(n11769) );
  NAND2_X1 U15235 ( .A1(n11773), .A2(n11769), .ZN(n15741) );
  OR2_X1 U15236 ( .A1(n15741), .A2(n13768), .ZN(n11770) );
  XNOR2_X1 U15237 ( .A(n11770), .B(n16515), .ZN(n16244) );
  NAND2_X1 U15238 ( .A1(n11076), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11771) );
  INV_X1 U15239 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16501) );
  NAND2_X1 U15240 ( .A1(n13390), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11776) );
  AND2_X2 U15241 ( .A1(n11775), .A2(n11774), .ZN(n11777) );
  OAI211_X1 U15242 ( .C1(n11775), .C2(n11776), .A(n11779), .B(n11780), .ZN(
        n15725) );
  NOR2_X1 U15243 ( .A1(n15725), .A2(n13768), .ZN(n16239) );
  NAND2_X1 U15244 ( .A1(n11785), .A2(n16227), .ZN(n16223) );
  NOR2_X1 U15245 ( .A1(n20006), .A2(n16001), .ZN(n11781) );
  AND2_X1 U15246 ( .A1(n11782), .A2(n11781), .ZN(n11783) );
  NOR3_X1 U15247 ( .A1(n15694), .A2(n13768), .A3(n16217), .ZN(n16193) );
  INV_X1 U15248 ( .A(n16193), .ZN(n11784) );
  OAI21_X1 U15249 ( .B1(n15694), .B2(n13768), .A(n16217), .ZN(n13380) );
  NAND2_X1 U15250 ( .A1(n11784), .A2(n13380), .ZN(n16215) );
  NOR2_X1 U15251 ( .A1(n11785), .A2(n16227), .ZN(n16212) );
  NAND2_X1 U15252 ( .A1(n13390), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11786) );
  NAND2_X1 U15253 ( .A1(n13766), .A2(n11786), .ZN(n13382) );
  INV_X1 U15254 ( .A(n11786), .ZN(n11787) );
  NAND2_X1 U15255 ( .A1(n11788), .A2(n11787), .ZN(n11789) );
  NAND2_X1 U15256 ( .A1(n13382), .A2(n11789), .ZN(n16194) );
  XNOR2_X1 U15257 ( .A(n16192), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11790) );
  XNOR2_X1 U15258 ( .A(n11791), .B(n11790), .ZN(n16211) );
  AOI22_X1 U15259 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n11794) );
  NAND2_X1 U15260 ( .A1(n12525), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11793) );
  INV_X1 U15261 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U15262 ( .A1(n12524), .A2(P2_EAX_REG_22__SCAN_IN), .ZN(n11797) );
  NAND2_X1 U15263 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11796) );
  OAI211_X1 U15264 ( .C1(n14727), .C2(n11798), .A(n11797), .B(n11796), .ZN(
        n16123) );
  INV_X1 U15265 ( .A(n15728), .ZN(n11802) );
  AOI22_X1 U15266 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11800) );
  NAND2_X1 U15267 ( .A1(n12525), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11799) );
  AND2_X1 U15268 ( .A1(n11800), .A2(n11799), .ZN(n15729) );
  AOI22_X1 U15269 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U15270 ( .A1(n12525), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11803) );
  INV_X1 U15271 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20586) );
  NAND2_X1 U15272 ( .A1(n12524), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n11806) );
  NAND2_X1 U15273 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11805) );
  OAI211_X1 U15274 ( .C1(n14727), .C2(n20586), .A(n11806), .B(n11805), .ZN(
        n15699) );
  INV_X1 U15275 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20588) );
  NAND2_X1 U15276 ( .A1(n12524), .A2(P2_EAX_REG_26__SCAN_IN), .ZN(n11808) );
  NAND2_X1 U15277 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11807) );
  OAI211_X1 U15278 ( .C1(n14727), .C2(n20588), .A(n11808), .B(n11807), .ZN(
        n15686) );
  AOI22_X1 U15279 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11810) );
  NAND2_X1 U15280 ( .A1(n12525), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11809) );
  AND2_X1 U15281 ( .A1(n11810), .A2(n11809), .ZN(n11812) );
  OR2_X2 U15282 ( .A1(n11811), .A2(n11812), .ZN(n15661) );
  NAND2_X1 U15283 ( .A1(n15685), .A2(n11812), .ZN(n11813) );
  NAND2_X1 U15284 ( .A1(n15661), .A2(n11813), .ZN(n16094) );
  INV_X1 U15285 ( .A(n16094), .ZN(n11814) );
  NAND2_X1 U15286 ( .A1(n11814), .A2(n19960), .ZN(n11815) );
  NAND4_X1 U15287 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        P2_U3019) );
  AND2_X2 U15288 ( .A1(n11826), .A2(n14485), .ZN(n11919) );
  INV_X1 U15289 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11820) );
  AND2_X2 U15290 ( .A1(n11827), .A2(n14087), .ZN(n11874) );
  AOI22_X1 U15291 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11825) );
  AND2_X2 U15292 ( .A1(n11826), .A2(n11827), .ZN(n11924) );
  NOR2_X4 U15293 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U15294 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12024), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11824) );
  INV_X1 U15295 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11821) );
  AND2_X2 U15296 ( .A1(n14481), .A2(n11828), .ZN(n11925) );
  AOI22_X1 U15298 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12712), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11823) );
  AND2_X2 U15299 ( .A1(n14481), .A2(n14087), .ZN(n11902) );
  AOI22_X1 U15300 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U15301 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U15302 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12098), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U15303 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U15304 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12712), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U15305 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U15306 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U15307 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U15308 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12024), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U15309 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12098), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U15310 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U15311 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12024), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U15312 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12712), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U15313 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U15314 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U15315 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12098), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U15316 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U15317 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11848) );
  NAND2_X1 U15319 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11857) );
  NAND2_X1 U15320 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U15321 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U15322 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11854) );
  NAND2_X1 U15323 ( .A1(n11931), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11861) );
  NAND2_X1 U15324 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11860) );
  NAND2_X1 U15325 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11859) );
  NAND2_X1 U15326 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11858) );
  NAND2_X1 U15327 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11865) );
  NAND2_X1 U15328 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U15329 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11863) );
  NAND2_X1 U15330 ( .A1(n12712), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11862) );
  NAND2_X1 U15331 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11869) );
  NAND2_X1 U15332 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11868) );
  NAND2_X1 U15333 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11867) );
  NAND2_X1 U15334 ( .A1(n12111), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11866) );
  AOI22_X1 U15335 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n11924), .ZN(n11879) );
  AOI22_X1 U15336 ( .A1(n9581), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9584), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U15337 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U15338 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U15339 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U15340 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12712), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11881) );
  INV_X2 U15341 ( .A(n11961), .ZN(n12591) );
  AOI22_X1 U15342 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12712), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U15343 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12024), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U15344 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U15345 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U15346 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U15347 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12098), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U15348 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11931), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U15349 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U15350 ( .A1(n12591), .A2(n11968), .ZN(n11896) );
  NAND2_X1 U15351 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11901) );
  NAND2_X1 U15352 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11900) );
  NAND2_X1 U15353 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11899) );
  NAND2_X1 U15354 ( .A1(n12712), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11898) );
  NAND2_X1 U15355 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11906) );
  NAND2_X1 U15356 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U15357 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11904) );
  NAND2_X1 U15358 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11903) );
  NAND2_X1 U15359 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11910) );
  NAND2_X1 U15360 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11909) );
  NAND2_X1 U15361 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11908) );
  NAND2_X1 U15362 ( .A1(n11931), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11907) );
  NAND2_X1 U15363 ( .A1(n9586), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11914) );
  NAND2_X1 U15364 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11913) );
  NAND2_X1 U15365 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11912) );
  NAND2_X1 U15366 ( .A1(n12111), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11911) );
  NAND2_X1 U15367 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U15368 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11922) );
  NAND2_X1 U15369 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U15370 ( .A1(n12116), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U15371 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11929) );
  NAND2_X1 U15372 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11928) );
  NAND2_X1 U15373 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11927) );
  NAND2_X1 U15374 ( .A1(n12712), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11926) );
  NAND2_X1 U15375 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11935) );
  NAND2_X1 U15376 ( .A1(n9581), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U15377 ( .A1(n12098), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U15378 ( .A1(n11931), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11932) );
  NAND2_X1 U15379 ( .A1(n12117), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U15380 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11938) );
  NAND2_X1 U15381 ( .A1(n9584), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U15382 ( .A1(n12111), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11936) );
  NAND2_X1 U15383 ( .A1(n12302), .A2(n14187), .ZN(n11948) );
  NAND2_X1 U15384 ( .A1(n12591), .A2(n11960), .ZN(n11970) );
  NAND2_X1 U15385 ( .A1(n11970), .A2(n12149), .ZN(n11983) );
  NAND2_X1 U15386 ( .A1(n11944), .A2(n11968), .ZN(n11972) );
  NAND2_X1 U15387 ( .A1(n11968), .A2(n11961), .ZN(n11949) );
  NAND2_X1 U15388 ( .A1(n11972), .A2(n11949), .ZN(n11945) );
  NAND2_X1 U15389 ( .A1(n11983), .A2(n11945), .ZN(n11963) );
  NAND2_X1 U15390 ( .A1(n11956), .A2(n11960), .ZN(n11953) );
  AND2_X1 U15391 ( .A1(n11966), .A2(n20842), .ZN(n14079) );
  NAND2_X1 U15392 ( .A1(n11951), .A2(n14079), .ZN(n12452) );
  INV_X1 U15393 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21364) );
  INV_X1 U15394 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n13864) );
  NAND2_X1 U15395 ( .A1(n21364), .A2(n13864), .ZN(n12300) );
  NAND2_X1 U15396 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_1__SCAN_IN), 
        .ZN(n15644) );
  NAND2_X1 U15397 ( .A1(n12450), .A2(n9687), .ZN(n11952) );
  AND3_X2 U15398 ( .A1(n12312), .A2(n12452), .A3(n11952), .ZN(n11977) );
  NAND2_X1 U15399 ( .A1(n11955), .A2(n14275), .ZN(n13969) );
  OAI211_X1 U15400 ( .C1(n11955), .C2(n20832), .A(n14080), .B(n13969), .ZN(
        n11986) );
  BUF_X1 U15401 ( .A(n11956), .Z(n11957) );
  OAI21_X1 U15402 ( .B1(n14273), .B2(n11957), .A(n11958), .ZN(n11959) );
  NOR2_X1 U15403 ( .A1(n11986), .A2(n11959), .ZN(n11974) );
  NAND2_X1 U15404 ( .A1(n14666), .A2(n13652), .ZN(n11962) );
  INV_X1 U15405 ( .A(n11963), .ZN(n11964) );
  NAND2_X1 U15406 ( .A1(n11965), .A2(n11964), .ZN(n12291) );
  NAND2_X1 U15407 ( .A1(n12291), .A2(n11966), .ZN(n12322) );
  NAND2_X1 U15408 ( .A1(n11967), .A2(n13652), .ZN(n11969) );
  NAND2_X1 U15409 ( .A1(n12290), .A2(n11957), .ZN(n12286) );
  INV_X1 U15410 ( .A(n12286), .ZN(n11971) );
  NAND2_X1 U15411 ( .A1(n11973), .A2(n15626), .ZN(n11981) );
  NAND4_X1 U15412 ( .A1(n11977), .A2(n11974), .A3(n12322), .A4(n11981), .ZN(
        n11975) );
  NAND2_X1 U15413 ( .A1(n21432), .A2(n21234), .ZN(n21191) );
  NAND2_X1 U15414 ( .A1(n21191), .A2(n21296), .ZN(n21131) );
  INV_X1 U15415 ( .A(n21131), .ZN(n21067) );
  INV_X1 U15416 ( .A(n13009), .ZN(n12043) );
  AND2_X1 U15417 ( .A1(n17355), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11991) );
  AOI21_X1 U15418 ( .B1(n21067), .B2(n12043), .A(n11991), .ZN(n11976) );
  INV_X1 U15419 ( .A(n11977), .ZN(n11978) );
  INV_X1 U15420 ( .A(n17355), .ZN(n11980) );
  MUX2_X1 U15421 ( .A(n11980), .B(n13009), .S(n21234), .Z(n12034) );
  INV_X1 U15422 ( .A(n11981), .ZN(n11982) );
  NAND2_X1 U15423 ( .A1(n11982), .A2(n14275), .ZN(n11989) );
  INV_X1 U15424 ( .A(n11966), .ZN(n13948) );
  AND2_X1 U15425 ( .A1(n13948), .A2(n12390), .ZN(n14745) );
  NAND2_X1 U15426 ( .A1(n14745), .A2(n11983), .ZN(n11985) );
  NAND2_X1 U15427 ( .A1(n15629), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20643) );
  INV_X1 U15428 ( .A(n20643), .ZN(n11984) );
  OR2_X1 U15429 ( .A1(n11958), .A2(n13652), .ZN(n12325) );
  AOI21_X1 U15430 ( .B1(n21398), .B2(n12286), .A(n11986), .ZN(n11987) );
  AOI21_X2 U15431 ( .B1(n12033), .B2(n12034), .A(n9630), .ZN(n12017) );
  NAND2_X1 U15432 ( .A1(n12016), .A2(n12017), .ZN(n12019) );
  INV_X1 U15433 ( .A(n11990), .ZN(n11994) );
  INV_X1 U15434 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U15435 ( .A1(n11992), .A2(n12230), .ZN(n11993) );
  NAND2_X1 U15436 ( .A1(n17355), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11998) );
  XNOR2_X1 U15437 ( .A(n21296), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20823) );
  NAND2_X1 U15438 ( .A1(n12043), .A2(n20823), .ZN(n11997) );
  OAI211_X2 U15439 ( .C1(n11996), .C2(n14101), .A(n11998), .B(n11997), .ZN(
        n11999) );
  AOI22_X1 U15440 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12024), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15441 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15442 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15443 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12001) );
  NAND4_X1 U15444 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12011) );
  AOI22_X1 U15445 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U15446 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15447 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U15448 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12006) );
  NAND4_X1 U15449 ( .A1(n12009), .A2(n12008), .A3(n12007), .A4(n12006), .ZN(
        n12010) );
  INV_X1 U15450 ( .A(n12046), .ZN(n12014) );
  AOI22_X1 U15451 ( .A1(n12277), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12014), .B2(n12013), .ZN(n12015) );
  INV_X1 U15452 ( .A(n12017), .ZN(n12018) );
  INV_X1 U15453 ( .A(n12047), .ZN(n12031) );
  AOI22_X1 U15454 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13698), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15455 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15456 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15457 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12020) );
  NAND4_X1 U15458 ( .A1(n12023), .A2(n12022), .A3(n12021), .A4(n12020), .ZN(
        n12030) );
  AOI22_X1 U15459 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15460 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15461 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15462 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12025) );
  NAND4_X1 U15463 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12029) );
  NAND2_X1 U15464 ( .A1(n12031), .A2(n12132), .ZN(n12032) );
  NAND2_X1 U15465 ( .A1(n12033), .A2(n12034), .ZN(n12035) );
  INV_X1 U15466 ( .A(n12132), .ZN(n12037) );
  NAND2_X1 U15467 ( .A1(n12277), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12036) );
  OAI211_X1 U15468 ( .C1(n12037), .C2(n12046), .A(n12036), .B(n12047), .ZN(
        n12038) );
  INV_X1 U15469 ( .A(n12038), .ZN(n12039) );
  NAND2_X1 U15470 ( .A1(n12148), .A2(n12039), .ZN(n12583) );
  OAI21_X1 U15471 ( .B1(n21296), .B2(n21064), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12042) );
  INV_X1 U15472 ( .A(n21296), .ZN(n12041) );
  NAND2_X1 U15473 ( .A1(n21132), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21007) );
  INV_X1 U15474 ( .A(n21007), .ZN(n12040) );
  NAND2_X1 U15475 ( .A1(n12041), .A2(n12040), .ZN(n21035) );
  NAND2_X1 U15476 ( .A1(n12042), .A2(n21035), .ZN(n21066) );
  AOI22_X1 U15477 ( .A1(n21066), .A2(n12043), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17355), .ZN(n12044) );
  XNOR2_X2 U15478 ( .A(n13976), .B(n20953), .ZN(n14480) );
  AOI22_X1 U15479 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15480 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15481 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15482 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12048) );
  NAND4_X1 U15483 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n12058) );
  INV_X1 U15484 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21518) );
  BUF_X2 U15485 ( .A(n12117), .Z(n12052) );
  AOI22_X1 U15486 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12056) );
  AOI22_X1 U15487 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15488 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15489 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12053) );
  NAND4_X1 U15490 ( .A1(n12056), .A2(n12055), .A3(n12054), .A4(n12053), .ZN(
        n12057) );
  AOI22_X1 U15491 ( .A1(n12264), .A2(n12168), .B1(n12277), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15492 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15493 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15494 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15495 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12060) );
  NAND4_X1 U15496 ( .A1(n12063), .A2(n12062), .A3(n12061), .A4(n12060), .ZN(
        n12069) );
  AOI22_X1 U15497 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15498 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15499 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15500 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12064) );
  NAND4_X1 U15501 ( .A1(n12067), .A2(n12066), .A3(n12065), .A4(n12064), .ZN(
        n12068) );
  NAND2_X1 U15502 ( .A1(n12264), .A2(n12177), .ZN(n12071) );
  NAND2_X1 U15503 ( .A1(n12277), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12070) );
  NAND2_X1 U15504 ( .A1(n12071), .A2(n12070), .ZN(n12175) );
  AOI22_X1 U15505 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15506 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15507 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15508 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12072) );
  NAND4_X1 U15509 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n12072), .ZN(
        n12081) );
  AOI22_X1 U15510 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15511 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15512 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15513 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12076) );
  NAND4_X1 U15514 ( .A1(n12079), .A2(n12078), .A3(n12077), .A4(n12076), .ZN(
        n12080) );
  NAND2_X1 U15515 ( .A1(n12264), .A2(n12188), .ZN(n12083) );
  NAND2_X1 U15516 ( .A1(n12277), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12082) );
  NAND2_X1 U15517 ( .A1(n12083), .A2(n12082), .ZN(n12185) );
  AOI22_X1 U15518 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15519 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15520 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15521 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12084) );
  NAND4_X1 U15522 ( .A1(n12087), .A2(n12086), .A3(n12085), .A4(n12084), .ZN(
        n12093) );
  AOI22_X1 U15523 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15524 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15525 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U15526 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12088) );
  NAND4_X1 U15527 ( .A1(n12091), .A2(n12090), .A3(n12089), .A4(n12088), .ZN(
        n12092) );
  NAND2_X1 U15528 ( .A1(n12264), .A2(n12199), .ZN(n12196) );
  AOI22_X1 U15529 ( .A1(n12024), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15530 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15531 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9587), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U15532 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12094) );
  NAND4_X1 U15533 ( .A1(n12097), .A2(n12096), .A3(n12095), .A4(n12094), .ZN(
        n12104) );
  AOI22_X1 U15534 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12945), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15535 ( .A1(n12052), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15536 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15537 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U15538 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12103) );
  NAND2_X1 U15539 ( .A1(n11957), .A2(n12208), .ZN(n12142) );
  INV_X1 U15540 ( .A(n12142), .ZN(n12105) );
  INV_X1 U15541 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15571) );
  NAND2_X1 U15542 ( .A1(n12217), .A2(n15571), .ZN(n15335) );
  NAND2_X1 U15543 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U15544 ( .A1(n12217), .A2(n12107), .ZN(n15333) );
  AND2_X1 U15545 ( .A1(n15335), .A2(n15333), .ZN(n12108) );
  INV_X1 U15546 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17394) );
  NAND2_X1 U15547 ( .A1(n12217), .A2(n17394), .ZN(n12109) );
  INV_X1 U15548 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15544) );
  NAND2_X1 U15549 ( .A1(n12217), .A2(n15544), .ZN(n15309) );
  INV_X1 U15550 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12213) );
  NAND2_X1 U15551 ( .A1(n12217), .A2(n12213), .ZN(n15298) );
  XNOR2_X1 U15552 ( .A(n12217), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15302) );
  AOI22_X1 U15553 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12945), .B1(
        n12879), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15554 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15555 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15556 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9590), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12112) );
  NAND4_X1 U15557 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(
        n12124) );
  AOI22_X1 U15558 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12024), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15559 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n12884), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15560 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13693), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15561 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12005), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12119) );
  NAND4_X1 U15562 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12119), .ZN(
        n12123) );
  NAND2_X1 U15563 ( .A1(n12132), .A2(n12150), .ZN(n12157) );
  NAND2_X1 U15564 ( .A1(n12157), .A2(n12158), .ZN(n12170) );
  NAND2_X1 U15565 ( .A1(n12170), .A2(n12168), .ZN(n12178) );
  INV_X1 U15566 ( .A(n12177), .ZN(n12125) );
  OR2_X1 U15567 ( .A1(n12178), .A2(n12125), .ZN(n12189) );
  INV_X1 U15568 ( .A(n12189), .ZN(n12126) );
  NAND2_X1 U15569 ( .A1(n12126), .A2(n12188), .ZN(n12200) );
  INV_X1 U15570 ( .A(n12200), .ZN(n12127) );
  NAND2_X1 U15571 ( .A1(n12127), .A2(n12199), .ZN(n12209) );
  INV_X1 U15572 ( .A(n12209), .ZN(n12128) );
  NAND3_X1 U15573 ( .A1(n12128), .A2(n21398), .A3(n12208), .ZN(n12129) );
  INV_X1 U15574 ( .A(n15379), .ZN(n12131) );
  XNOR2_X1 U15575 ( .A(n12132), .B(n12150), .ZN(n12134) );
  OAI211_X1 U15576 ( .C1(n12134), .C2(n14273), .A(n12133), .B(n14666), .ZN(
        n12135) );
  INV_X1 U15577 ( .A(n12135), .ZN(n12136) );
  INV_X1 U15578 ( .A(n12208), .ZN(n12138) );
  NAND2_X1 U15579 ( .A1(n12138), .A2(n11957), .ZN(n12139) );
  MUX2_X1 U15580 ( .A(n12142), .B(n12139), .S(n12150), .Z(n12140) );
  INV_X1 U15581 ( .A(n12140), .ZN(n12141) );
  NAND2_X1 U15582 ( .A1(n12141), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U15583 ( .A1(n12277), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12144) );
  AOI21_X1 U15584 ( .B1(n11955), .B2(n12150), .A(n10287), .ZN(n12143) );
  NAND3_X1 U15585 ( .A1(n12144), .A2(n12143), .A3(n12142), .ZN(n12145) );
  XNOR2_X1 U15586 ( .A(n12146), .B(n12145), .ZN(n12147) );
  NAND2_X1 U15587 ( .A1(n11955), .A2(n12149), .ZN(n12159) );
  OAI21_X1 U15588 ( .B1(n14273), .B2(n12150), .A(n12159), .ZN(n12151) );
  INV_X1 U15589 ( .A(n12151), .ZN(n12152) );
  NAND2_X1 U15590 ( .A1(n12153), .A2(n12152), .ZN(n14107) );
  INV_X1 U15591 ( .A(n12154), .ZN(n14108) );
  NAND2_X1 U15592 ( .A1(n14108), .A2(n12155), .ZN(n12156) );
  INV_X1 U15593 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14262) );
  OAI21_X1 U15594 ( .B1(n12158), .B2(n12157), .A(n12170), .ZN(n12161) );
  INV_X1 U15595 ( .A(n12159), .ZN(n12160) );
  AOI21_X1 U15596 ( .B1(n12161), .B2(n21398), .A(n12160), .ZN(n12162) );
  NAND2_X1 U15597 ( .A1(n12163), .A2(n12162), .ZN(n14253) );
  NAND2_X1 U15598 ( .A1(n14252), .A2(n14253), .ZN(n12166) );
  NAND2_X1 U15599 ( .A1(n12164), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12165) );
  INV_X1 U15600 ( .A(n12168), .ZN(n12169) );
  XNOR2_X1 U15601 ( .A(n12170), .B(n12169), .ZN(n12171) );
  NAND2_X1 U15602 ( .A1(n12171), .A2(n21398), .ZN(n12172) );
  INV_X1 U15603 ( .A(n14463), .ZN(n12174) );
  INV_X1 U15604 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14471) );
  XNOR2_X1 U15605 ( .A(n12176), .B(n12175), .ZN(n12614) );
  NAND2_X1 U15606 ( .A1(n12614), .A2(n12243), .ZN(n12181) );
  XNOR2_X1 U15607 ( .A(n12178), .B(n12177), .ZN(n12179) );
  NAND2_X1 U15608 ( .A1(n12179), .A2(n21398), .ZN(n12180) );
  NAND2_X1 U15609 ( .A1(n12181), .A2(n12180), .ZN(n12183) );
  INV_X1 U15610 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U15611 ( .A1(n12183), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12184) );
  OR2_X1 U15612 ( .A1(n12186), .A2(n12185), .ZN(n12187) );
  XNOR2_X1 U15613 ( .A(n12189), .B(n12188), .ZN(n12190) );
  NAND2_X1 U15614 ( .A1(n12190), .A2(n21398), .ZN(n12191) );
  NAND2_X1 U15615 ( .A1(n12192), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12193) );
  NAND2_X1 U15616 ( .A1(n12277), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12195) );
  AND2_X1 U15617 ( .A1(n12196), .A2(n12195), .ZN(n12197) );
  NAND2_X1 U15618 ( .A1(n12194), .A2(n12197), .ZN(n12627) );
  NAND3_X1 U15619 ( .A1(n12198), .A2(n12627), .A3(n12243), .ZN(n12203) );
  XNOR2_X1 U15620 ( .A(n12200), .B(n12199), .ZN(n12201) );
  NAND2_X1 U15621 ( .A1(n12201), .A2(n21398), .ZN(n12202) );
  NAND2_X1 U15622 ( .A1(n12203), .A2(n12202), .ZN(n12204) );
  OR2_X1 U15623 ( .A1(n12204), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17372) );
  NAND2_X1 U15624 ( .A1(n12204), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17371) );
  NAND2_X1 U15625 ( .A1(n12264), .A2(n12208), .ZN(n12206) );
  NAND2_X1 U15626 ( .A1(n12277), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12205) );
  XNOR2_X1 U15627 ( .A(n12207), .B(n10595), .ZN(n12634) );
  XNOR2_X1 U15628 ( .A(n12209), .B(n12208), .ZN(n12210) );
  NAND2_X1 U15629 ( .A1(n12210), .A2(n21398), .ZN(n12211) );
  OR2_X1 U15630 ( .A1(n17364), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12212) );
  NAND2_X1 U15631 ( .A1(n15292), .A2(n12212), .ZN(n12215) );
  OR2_X1 U15632 ( .A1(n12217), .A2(n12213), .ZN(n15297) );
  NAND2_X1 U15633 ( .A1(n17364), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12214) );
  INV_X1 U15634 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15522) );
  OR2_X1 U15635 ( .A1(n12217), .A2(n15571), .ZN(n15334) );
  NOR2_X1 U15636 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12216) );
  OR2_X1 U15637 ( .A1(n12217), .A2(n12216), .ZN(n15331) );
  NAND2_X1 U15638 ( .A1(n15334), .A2(n15331), .ZN(n15319) );
  NOR2_X1 U15639 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12218) );
  NOR2_X1 U15640 ( .A1(n12217), .A2(n12218), .ZN(n12219) );
  INV_X1 U15641 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15501) );
  INV_X1 U15642 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15240) );
  INV_X1 U15643 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15491) );
  NAND3_X1 U15644 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12222) );
  NAND2_X1 U15645 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15471) );
  NOR2_X1 U15646 ( .A1(n12222), .A2(n15471), .ZN(n12224) );
  NOR2_X1 U15647 ( .A1(n12217), .A2(n15469), .ZN(n12223) );
  NAND3_X1 U15648 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15425) );
  AND2_X1 U15649 ( .A1(n15190), .A2(n12217), .ZN(n15210) );
  INV_X1 U15650 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15433) );
  INV_X1 U15651 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15211) );
  NAND2_X1 U15652 ( .A1(n15433), .A2(n15211), .ZN(n12567) );
  AND2_X1 U15653 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15395) );
  INV_X1 U15654 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15416) );
  INV_X1 U15655 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12572) );
  NAND2_X1 U15656 ( .A1(n15416), .A2(n12572), .ZN(n15404) );
  XNOR2_X1 U15657 ( .A(n12217), .B(n10324), .ZN(n15187) );
  AOI21_X1 U15658 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n10324), .A(
        n15187), .ZN(n12229) );
  INV_X1 U15659 ( .A(n13825), .ZN(n12456) );
  NAND2_X1 U15660 ( .A1(n21432), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12232) );
  NAND2_X1 U15661 ( .A1(n12230), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12231) );
  NAND2_X1 U15662 ( .A1(n12232), .A2(n12231), .ZN(n12240) );
  NAND2_X1 U15663 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21234), .ZN(
        n12244) );
  NAND2_X1 U15664 ( .A1(n21064), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12236) );
  NAND2_X1 U15665 ( .A1(n14101), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12233) );
  NAND2_X1 U15666 ( .A1(n12236), .A2(n12233), .ZN(n12255) );
  INV_X1 U15667 ( .A(n12255), .ZN(n12234) );
  NAND2_X1 U15668 ( .A1(n12235), .A2(n12234), .ZN(n12257) );
  NAND2_X1 U15669 ( .A1(n12257), .A2(n12236), .ZN(n12272) );
  MUX2_X1 U15670 ( .A(n21132), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n15642), .Z(n12271) );
  AOI222_X1 U15671 ( .A1(n12269), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n12269), .B2(n13981), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n13981), .ZN(n12297) );
  NAND2_X1 U15672 ( .A1(n20842), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12237) );
  NAND2_X1 U15673 ( .A1(n12238), .A2(n12237), .ZN(n12251) );
  INV_X1 U15674 ( .A(n12251), .ZN(n12239) );
  NAND2_X1 U15675 ( .A1(n12239), .A2(n14275), .ZN(n12276) );
  NAND2_X1 U15676 ( .A1(n12240), .A2(n12244), .ZN(n12241) );
  NAND2_X1 U15677 ( .A1(n12242), .A2(n12241), .ZN(n12295) );
  INV_X1 U15678 ( .A(n12295), .ZN(n12254) );
  NAND2_X1 U15679 ( .A1(n12251), .A2(n12254), .ZN(n12253) );
  NAND2_X1 U15680 ( .A1(n12277), .A2(n12243), .ZN(n12282) );
  OAI21_X1 U15681 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21234), .A(
        n12244), .ZN(n12245) );
  INV_X1 U15682 ( .A(n12245), .ZN(n12248) );
  NAND2_X1 U15683 ( .A1(n12264), .A2(n12248), .ZN(n12246) );
  NAND2_X1 U15684 ( .A1(n12282), .A2(n12246), .ZN(n12250) );
  NAND2_X1 U15685 ( .A1(n20842), .A2(n14119), .ZN(n12247) );
  NAND2_X1 U15686 ( .A1(n12247), .A2(n20828), .ZN(n12263) );
  OAI211_X1 U15687 ( .C1(n12319), .C2(n11955), .A(n12263), .B(n12248), .ZN(
        n12249) );
  OAI211_X1 U15688 ( .C1(n12251), .C2(n12254), .A(n12250), .B(n12249), .ZN(
        n12252) );
  OAI211_X1 U15689 ( .C1(n12276), .C2(n12254), .A(n12253), .B(n12252), .ZN(
        n12262) );
  NAND2_X1 U15690 ( .A1(n12256), .A2(n12255), .ZN(n12258) );
  NAND2_X1 U15691 ( .A1(n12258), .A2(n12257), .ZN(n12294) );
  INV_X1 U15692 ( .A(n12277), .ZN(n12260) );
  NAND2_X1 U15693 ( .A1(n12264), .A2(n12265), .ZN(n12259) );
  OAI211_X1 U15694 ( .C1(n12265), .C2(n12260), .A(n12263), .B(n12259), .ZN(
        n12261) );
  NAND2_X1 U15695 ( .A1(n12262), .A2(n12261), .ZN(n12268) );
  INV_X1 U15696 ( .A(n12263), .ZN(n12266) );
  NAND3_X1 U15697 ( .A1(n12266), .A2(n12265), .A3(n12264), .ZN(n12267) );
  AND2_X1 U15698 ( .A1(n13981), .A2(n12269), .ZN(n12270) );
  NOR2_X1 U15699 ( .A1(n12272), .A2(n12271), .ZN(n12273) );
  OAI22_X1 U15700 ( .A1(n12298), .A2(n12276), .B1(n12279), .B2(n12275), .ZN(
        n12278) );
  NAND3_X1 U15701 ( .A1(n12280), .A2(n12279), .A3(n12298), .ZN(n12281) );
  INV_X1 U15702 ( .A(n12282), .ZN(n12283) );
  NAND2_X1 U15703 ( .A1(n12297), .A2(n12283), .ZN(n12284) );
  NOR2_X1 U15704 ( .A1(n15626), .A2(n20828), .ZN(n12329) );
  INV_X1 U15705 ( .A(n14208), .ZN(n12285) );
  MUX2_X1 U15706 ( .A(n12286), .B(n20828), .S(n12285), .Z(n12287) );
  NAND2_X1 U15707 ( .A1(n12287), .A2(n14119), .ZN(n12324) );
  AOI21_X1 U15708 ( .B1(n15626), .B2(n11955), .A(n12288), .ZN(n12311) );
  OR2_X1 U15709 ( .A1(n14208), .A2(n12012), .ZN(n12289) );
  AND2_X1 U15710 ( .A1(n12324), .A2(n12310), .ZN(n12293) );
  OR2_X1 U15711 ( .A1(n12319), .A2(n14119), .ZN(n12292) );
  NOR2_X1 U15712 ( .A1(n12293), .A2(n13950), .ZN(n13971) );
  AOI21_X1 U15713 ( .B1(n14096), .B2(n12329), .A(n13971), .ZN(n12308) );
  NOR3_X1 U15714 ( .A1(n12296), .A2(n12295), .A3(n12294), .ZN(n12299) );
  AOI21_X1 U15715 ( .B1(n12299), .B2(n12298), .A(n12297), .ZN(n13955) );
  AND3_X1 U15716 ( .A1(n12300), .A2(n15650), .A3(n15644), .ZN(n17346) );
  INV_X1 U15717 ( .A(n17346), .ZN(n13946) );
  AOI21_X1 U15718 ( .B1(n14275), .B2(n13946), .A(n17352), .ZN(n12301) );
  NAND2_X1 U15719 ( .A1(n13955), .A2(n12301), .ZN(n12307) );
  OAI21_X1 U15720 ( .B1(n14275), .B2(n17346), .A(n21404), .ZN(n13800) );
  INV_X1 U15721 ( .A(n13800), .ZN(n12303) );
  NAND2_X1 U15722 ( .A1(n12302), .A2(n12303), .ZN(n12304) );
  NAND3_X1 U15723 ( .A1(n12304), .A2(n14119), .A3(n13853), .ZN(n12305) );
  NAND2_X1 U15724 ( .A1(n14116), .A2(n12305), .ZN(n12306) );
  NAND2_X1 U15725 ( .A1(n12310), .A2(n12309), .ZN(n17335) );
  NAND2_X1 U15726 ( .A1(n12311), .A2(n11966), .ZN(n14088) );
  NAND2_X1 U15727 ( .A1(n17335), .A2(n14088), .ZN(n13951) );
  OAI21_X1 U15728 ( .B1(n11957), .B2(n12452), .A(n12312), .ZN(n12313) );
  NOR2_X1 U15729 ( .A1(n13951), .A2(n12313), .ZN(n12314) );
  NAND2_X1 U15730 ( .A1(n13950), .A2(n14275), .ZN(n17323) );
  INV_X1 U15731 ( .A(n12315), .ZN(n12318) );
  INV_X1 U15732 ( .A(n12390), .ZN(n12446) );
  OAI21_X1 U15733 ( .B1(n11958), .B2(n20828), .A(n12316), .ZN(n12317) );
  AOI21_X1 U15734 ( .B1(n12318), .B2(n12446), .A(n12317), .ZN(n12323) );
  NAND2_X1 U15735 ( .A1(n14200), .A2(n12288), .ZN(n12321) );
  INV_X1 U15736 ( .A(n13969), .ZN(n15060) );
  NAND2_X1 U15737 ( .A1(n15060), .A2(n12319), .ZN(n12320) );
  NAND4_X1 U15738 ( .A1(n12324), .A2(n12323), .A3(n12328), .A4(n12322), .ZN(
        n14084) );
  OAI21_X1 U15739 ( .B1(n14080), .B2(n14119), .A(n12325), .ZN(n12326) );
  NOR2_X1 U15740 ( .A1(n14084), .A2(n12326), .ZN(n12327) );
  INV_X1 U15741 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15390) );
  NOR2_X1 U15742 ( .A1(n15464), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12330) );
  INV_X1 U15743 ( .A(n14196), .ZN(n15614) );
  NAND3_X1 U15744 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15523) );
  NOR2_X1 U15745 ( .A1(n15523), .A2(n15522), .ZN(n15516) );
  AND2_X1 U15746 ( .A1(n15516), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12346) );
  NAND2_X1 U15747 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15596) );
  INV_X1 U15748 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15580) );
  NOR2_X1 U15749 ( .A1(n15596), .A2(n15580), .ZN(n12331) );
  AND3_X1 U15750 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15589) );
  AND2_X1 U15751 ( .A1(n12331), .A2(n15589), .ZN(n15572) );
  NAND2_X1 U15752 ( .A1(n15572), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12334) );
  NAND2_X1 U15753 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17400) );
  NOR2_X1 U15754 ( .A1(n21471), .A2(n17400), .ZN(n15570) );
  OAI21_X1 U15755 ( .B1(n14194), .B2(n14261), .A(n14262), .ZN(n14468) );
  NAND2_X1 U15756 ( .A1(n15570), .A2(n14468), .ZN(n15561) );
  NOR2_X1 U15757 ( .A1(n12334), .A2(n15561), .ZN(n15460) );
  NAND2_X1 U15758 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15460), .ZN(
        n12342) );
  INV_X1 U15759 ( .A(n12342), .ZN(n15513) );
  AND2_X1 U15760 ( .A1(n12346), .A2(n15513), .ZN(n12332) );
  NOR2_X1 U15761 ( .A1(n15562), .A2(n12332), .ZN(n12333) );
  NOR2_X1 U15762 ( .A1(n14465), .A2(n12333), .ZN(n12336) );
  NAND2_X1 U15763 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12346), .ZN(
        n15466) );
  NOR2_X1 U15764 ( .A1(n14262), .A2(n14261), .ZN(n14467) );
  NAND2_X1 U15765 ( .A1(n14467), .A2(n15570), .ZN(n12341) );
  OR2_X1 U15766 ( .A1(n12334), .A2(n12341), .ZN(n15461) );
  OAI21_X1 U15767 ( .B1(n15466), .B2(n15461), .A(n17401), .ZN(n12335) );
  INV_X1 U15768 ( .A(n15471), .ZN(n15470) );
  NAND2_X1 U15769 ( .A1(n15502), .A2(n15470), .ZN(n12337) );
  INV_X1 U15770 ( .A(n17404), .ZN(n15515) );
  NAND2_X1 U15771 ( .A1(n15515), .A2(n15590), .ZN(n15592) );
  NAND2_X1 U15772 ( .A1(n12337), .A2(n15592), .ZN(n15472) );
  NAND2_X1 U15773 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12344) );
  NAND2_X1 U15774 ( .A1(n17404), .A2(n12344), .ZN(n12338) );
  NOR2_X1 U15775 ( .A1(n15562), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12339) );
  NAND2_X1 U15776 ( .A1(n17404), .A2(n15425), .ZN(n12340) );
  INV_X1 U15777 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15424) );
  NOR2_X1 U15778 ( .A1(n15456), .A2(n17404), .ZN(n15413) );
  AOI21_X1 U15779 ( .B1(n15423), .B2(n15395), .A(n15413), .ZN(n15399) );
  INV_X1 U15780 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14095) );
  NOR3_X1 U15781 ( .A1(n15388), .A2(n15413), .A3(n14095), .ZN(n12350) );
  NAND2_X1 U15782 ( .A1(n17416), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n13823) );
  INV_X1 U15783 ( .A(n13823), .ZN(n12349) );
  NAND2_X1 U15784 ( .A1(n15488), .A2(n14194), .ZN(n14191) );
  INV_X1 U15785 ( .A(n15589), .ZN(n15577) );
  OR3_X1 U15786 ( .A1(n15577), .A2(n12341), .A3(n15596), .ZN(n15564) );
  NAND3_X1 U15787 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17387) );
  NOR2_X1 U15788 ( .A1(n15564), .A2(n17387), .ZN(n15510) );
  NAND2_X1 U15789 ( .A1(n15565), .A2(n15510), .ZN(n15444) );
  OR2_X1 U15790 ( .A1(n15562), .A2(n12342), .ZN(n12343) );
  NAND2_X1 U15791 ( .A1(n15444), .A2(n12343), .ZN(n15535) );
  NOR2_X1 U15792 ( .A1(n15471), .A2(n12344), .ZN(n12345) );
  AND2_X1 U15793 ( .A1(n12346), .A2(n12345), .ZN(n12347) );
  NAND2_X1 U15794 ( .A1(n15535), .A2(n12347), .ZN(n15452) );
  NAND3_X1 U15795 ( .A1(n15417), .A2(n15395), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15389) );
  NOR3_X1 U15796 ( .A1(n15389), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15390), .ZN(n12348) );
  AOI22_X1 U15797 ( .A1(n14200), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n13947), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14674) );
  INV_X1 U15798 ( .A(n12361), .ZN(n12353) );
  INV_X1 U15799 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12352) );
  NAND2_X1 U15800 ( .A1(n12353), .A2(n12352), .ZN(n12357) );
  NAND2_X1 U15801 ( .A1(n12362), .A2(n14261), .ZN(n12355) );
  NAND2_X1 U15802 ( .A1(n14187), .A2(n12352), .ZN(n12354) );
  NAND3_X1 U15803 ( .A1(n12355), .A2(n14671), .A3(n12354), .ZN(n12356) );
  INV_X1 U15804 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n21553) );
  NAND2_X1 U15805 ( .A1(n14671), .A2(n21553), .ZN(n12359) );
  NAND2_X1 U15806 ( .A1(n12362), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12358) );
  AND2_X1 U15807 ( .A1(n12359), .A2(n12358), .ZN(n14201) );
  OR2_X1 U15808 ( .A1(n12361), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12367) );
  INV_X1 U15809 ( .A(n12362), .ZN(n12378) );
  NAND2_X1 U15810 ( .A1(n12362), .A2(n14262), .ZN(n12365) );
  INV_X1 U15811 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12363) );
  NAND2_X1 U15812 ( .A1(n14187), .A2(n12363), .ZN(n12364) );
  NAND3_X1 U15813 ( .A1(n12365), .A2(n14671), .A3(n12364), .ZN(n12366) );
  AND2_X1 U15814 ( .A1(n12367), .A2(n12366), .ZN(n14254) );
  MUX2_X1 U15815 ( .A(n12440), .B(n14671), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12370) );
  OAI21_X1 U15816 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14200), .A(
        n12370), .ZN(n14446) );
  MUX2_X1 U15817 ( .A(n12361), .B(n12362), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12372) );
  NAND2_X1 U15818 ( .A1(n12378), .A2(n13947), .ZN(n12386) );
  NAND2_X1 U15819 ( .A1(n13947), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12371) );
  INV_X1 U15820 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20703) );
  NAND2_X1 U15821 ( .A1(n12413), .A2(n20703), .ZN(n12376) );
  NAND2_X1 U15822 ( .A1(n14187), .A2(n20703), .ZN(n12374) );
  NAND2_X1 U15823 ( .A1(n14671), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12373) );
  NAND3_X1 U15824 ( .A1(n12362), .A2(n12374), .A3(n12373), .ZN(n12375) );
  INV_X1 U15825 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17408) );
  OAI21_X1 U15826 ( .B1(n14187), .B2(n17408), .A(n12386), .ZN(n12377) );
  INV_X1 U15827 ( .A(n12377), .ZN(n12380) );
  MUX2_X1 U15828 ( .A(n12361), .B(n12362), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12379) );
  NAND2_X1 U15829 ( .A1(n12380), .A2(n12379), .ZN(n14635) );
  INV_X1 U15830 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n12381) );
  NAND2_X1 U15831 ( .A1(n12413), .A2(n12381), .ZN(n12385) );
  NAND2_X1 U15832 ( .A1(n14187), .A2(n12381), .ZN(n12383) );
  NAND2_X1 U15833 ( .A1(n12390), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12382) );
  NAND3_X1 U15834 ( .A1(n12362), .A2(n12383), .A3(n12382), .ZN(n12384) );
  AND2_X1 U15835 ( .A1(n12385), .A2(n12384), .ZN(n14628) );
  MUX2_X1 U15836 ( .A(n12361), .B(n12362), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12389) );
  OAI21_X1 U15837 ( .B1(n14187), .B2(n12130), .A(n12386), .ZN(n12387) );
  INV_X1 U15838 ( .A(n12387), .ZN(n12388) );
  AND2_X1 U15839 ( .A1(n12389), .A2(n12388), .ZN(n15049) );
  INV_X1 U15840 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20664) );
  NAND2_X1 U15841 ( .A1(n12413), .A2(n20664), .ZN(n12394) );
  NAND2_X1 U15842 ( .A1(n14187), .A2(n20664), .ZN(n12392) );
  NAND2_X1 U15843 ( .A1(n12390), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12391) );
  NAND3_X1 U15844 ( .A1(n12362), .A2(n12392), .A3(n12391), .ZN(n12393) );
  AND2_X1 U15845 ( .A1(n12394), .A2(n12393), .ZN(n14652) );
  AND2_X2 U15846 ( .A1(n14651), .A2(n14652), .ZN(n15037) );
  OR2_X1 U15847 ( .A1(n12361), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n12398) );
  INV_X1 U15848 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15362) );
  NAND2_X1 U15849 ( .A1(n12362), .A2(n15362), .ZN(n12396) );
  INV_X1 U15850 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15106) );
  NAND2_X1 U15851 ( .A1(n14187), .A2(n15106), .ZN(n12395) );
  NAND3_X1 U15852 ( .A1(n12396), .A2(n14671), .A3(n12395), .ZN(n12397) );
  NAND2_X1 U15853 ( .A1(n12398), .A2(n12397), .ZN(n15036) );
  MUX2_X1 U15854 ( .A(n12440), .B(n14671), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12399) );
  OAI21_X1 U15855 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14200), .A(
        n12399), .ZN(n15023) );
  MUX2_X1 U15856 ( .A(n12361), .B(n12362), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12401) );
  NAND2_X1 U15857 ( .A1(n13947), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12400) );
  AND2_X1 U15858 ( .A1(n12401), .A2(n12400), .ZN(n15007) );
  INV_X1 U15859 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15102) );
  NAND2_X1 U15860 ( .A1(n12413), .A2(n15102), .ZN(n12405) );
  NAND2_X1 U15861 ( .A1(n14187), .A2(n15102), .ZN(n12403) );
  NAND2_X1 U15862 ( .A1(n14671), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12402) );
  NAND3_X1 U15863 ( .A1(n12362), .A2(n12403), .A3(n12402), .ZN(n12404) );
  MUX2_X1 U15864 ( .A(n12361), .B(n12362), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12407) );
  NAND2_X1 U15865 ( .A1(n13947), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12406) );
  NAND2_X1 U15866 ( .A1(n12407), .A2(n12406), .ZN(n14970) );
  NAND2_X1 U15867 ( .A1(n14989), .A2(n14970), .ZN(n14954) );
  MUX2_X1 U15868 ( .A(n12440), .B(n14671), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12408) );
  OAI21_X1 U15869 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14200), .A(
        n12408), .ZN(n14955) );
  OR2_X1 U15870 ( .A1(n12361), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n12411) );
  INV_X1 U15871 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15534) );
  NAND2_X1 U15872 ( .A1(n12362), .A2(n15534), .ZN(n12409) );
  OAI211_X1 U15873 ( .C1(n13947), .C2(P1_EBX_REG_16__SCAN_IN), .A(n14671), .B(
        n12409), .ZN(n12410) );
  AND2_X2 U15874 ( .A1(n14939), .A2(n12412), .ZN(n14942) );
  INV_X1 U15875 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15097) );
  NAND2_X1 U15876 ( .A1(n12413), .A2(n15097), .ZN(n12417) );
  NAND2_X1 U15877 ( .A1(n14187), .A2(n15097), .ZN(n12415) );
  NAND2_X1 U15878 ( .A1(n14671), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12414) );
  NAND3_X1 U15879 ( .A1(n12362), .A2(n12415), .A3(n12414), .ZN(n12416) );
  NAND2_X1 U15880 ( .A1(n12362), .A2(n12221), .ZN(n12418) );
  OAI211_X1 U15881 ( .C1(n13947), .C2(P1_EBX_REG_18__SCAN_IN), .A(n14671), .B(
        n12418), .ZN(n12420) );
  OR2_X1 U15882 ( .A1(n12361), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U15883 ( .A1(n12420), .A2(n12419), .ZN(n14897) );
  MUX2_X1 U15884 ( .A(n12440), .B(n14671), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12421) );
  OAI21_X1 U15885 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14200), .A(
        n12421), .ZN(n14894) );
  MUX2_X1 U15886 ( .A(n12361), .B(n12362), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12423) );
  NAND2_X1 U15887 ( .A1(n13947), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12422) );
  INV_X1 U15888 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n12424) );
  NAND2_X1 U15889 ( .A1(n14187), .A2(n12424), .ZN(n12426) );
  NAND2_X1 U15890 ( .A1(n14671), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12425) );
  NAND3_X1 U15891 ( .A1(n12362), .A2(n12426), .A3(n12425), .ZN(n12427) );
  OAI21_X1 U15892 ( .B1(n12440), .B2(P1_EBX_REG_21__SCAN_IN), .A(n12427), .ZN(
        n14856) );
  NAND2_X1 U15893 ( .A1(n12362), .A2(n15469), .ZN(n12428) );
  OAI211_X1 U15894 ( .C1(n13947), .C2(P1_EBX_REG_22__SCAN_IN), .A(n14671), .B(
        n12428), .ZN(n12430) );
  OR2_X1 U15895 ( .A1(n12361), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n12429) );
  NAND2_X1 U15896 ( .A1(n12430), .A2(n12429), .ZN(n14840) );
  MUX2_X1 U15897 ( .A(n12440), .B(n14671), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12432) );
  OR2_X1 U15898 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12431) );
  AND2_X2 U15899 ( .A1(n14832), .A2(n14833), .ZN(n14835) );
  NAND2_X1 U15900 ( .A1(n12362), .A2(n15211), .ZN(n12433) );
  OAI211_X1 U15901 ( .C1(n13947), .C2(P1_EBX_REG_24__SCAN_IN), .A(n14671), .B(
        n12433), .ZN(n12435) );
  OR2_X1 U15902 ( .A1(n12361), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n12434) );
  NAND2_X1 U15903 ( .A1(n12435), .A2(n12434), .ZN(n14815) );
  MUX2_X1 U15904 ( .A(n12440), .B(n14671), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12436) );
  OAI21_X1 U15905 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14200), .A(
        n12436), .ZN(n14806) );
  OR2_X1 U15906 ( .A1(n12361), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n12439) );
  NAND2_X1 U15907 ( .A1(n12362), .A2(n15424), .ZN(n12437) );
  OAI211_X1 U15908 ( .C1(n13947), .C2(P1_EBX_REG_26__SCAN_IN), .A(n14671), .B(
        n12437), .ZN(n12438) );
  MUX2_X1 U15909 ( .A(n12440), .B(n14671), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12442) );
  OR2_X1 U15910 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12441) );
  AND2_X1 U15911 ( .A1(n12442), .A2(n12441), .ZN(n14774) );
  MUX2_X1 U15912 ( .A(n12361), .B(n12362), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12444) );
  NAND2_X1 U15913 ( .A1(n13947), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12443) );
  NAND2_X1 U15914 ( .A1(n12444), .A2(n12443), .ZN(n13659) );
  NAND2_X1 U15915 ( .A1(n13657), .A2(n13659), .ZN(n13658) );
  OR2_X1 U15916 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12445) );
  INV_X1 U15917 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15086) );
  NAND2_X1 U15918 ( .A1(n14187), .A2(n15086), .ZN(n12447) );
  NAND2_X1 U15919 ( .A1(n12445), .A2(n12447), .ZN(n14670) );
  MUX2_X1 U15920 ( .A(n14670), .B(n12447), .S(n12446), .Z(n14751) );
  AOI22_X1 U15921 ( .A1(n14200), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n13947), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12448) );
  INV_X1 U15922 ( .A(n12452), .ZN(n12453) );
  AOI22_X1 U15923 ( .A1(n12451), .A2(n20828), .B1(n12453), .B2(n11957), .ZN(
        n12454) );
  OAI211_X1 U15924 ( .C1(n12456), .C2(n17397), .A(n12351), .B(n9664), .ZN(
        P1_U3000) );
  NAND2_X1 U15925 ( .A1(n12503), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12506) );
  NAND2_X1 U15926 ( .A1(n12512), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12511) );
  INV_X1 U15927 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12514) );
  INV_X1 U15928 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16200) );
  INV_X1 U15929 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12457) );
  NAND2_X1 U15930 ( .A1(n13781), .A2(n16902), .ZN(n12459) );
  NAND2_X1 U15931 ( .A1(n20619), .A2(n16902), .ZN(n12460) );
  MUX2_X1 U15932 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n15963) );
  INV_X1 U15933 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13939) );
  MUX2_X1 U15934 ( .A(n13939), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n15964) );
  NOR2_X1 U15935 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21437) );
  INV_X1 U15936 ( .A(n21437), .ZN(n12462) );
  NAND2_X1 U15937 ( .A1(n12465), .A2(n12462), .ZN(n15953) );
  NAND2_X1 U15938 ( .A1(n15966), .A2(n15953), .ZN(n15933) );
  AND2_X1 U15939 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  NOR2_X1 U15940 ( .A1(n12463), .A2(n12466), .ZN(n16451) );
  OR2_X1 U15941 ( .A1(n15933), .A2(n16451), .ZN(n19814) );
  OR2_X1 U15942 ( .A1(n12463), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12467) );
  AND2_X1 U15943 ( .A1(n12469), .A2(n12467), .ZN(n19816) );
  NOR2_X1 U15944 ( .A1(n19814), .A2(n19816), .ZN(n19818) );
  NAND2_X1 U15945 ( .A1(n12469), .A2(n12468), .ZN(n12470) );
  NAND2_X1 U15946 ( .A1(n12471), .A2(n12470), .ZN(n19794) );
  NAND2_X1 U15947 ( .A1(n19818), .A2(n19794), .ZN(n15921) );
  NAND2_X1 U15948 ( .A1(n12471), .A2(n21556), .ZN(n12472) );
  NAND2_X1 U15949 ( .A1(n12473), .A2(n12472), .ZN(n15922) );
  INV_X1 U15950 ( .A(n15922), .ZN(n16414) );
  OR2_X1 U15951 ( .A1(n15921), .A2(n16414), .ZN(n15910) );
  AND2_X1 U15952 ( .A1(n12473), .A2(n16403), .ZN(n12474) );
  NOR2_X1 U15953 ( .A1(n12475), .A2(n12474), .ZN(n16405) );
  NOR2_X1 U15954 ( .A1(n15910), .A2(n16405), .ZN(n15899) );
  OR2_X1 U15955 ( .A1(n12475), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12476) );
  NAND2_X1 U15956 ( .A1(n12477), .A2(n12476), .ZN(n16394) );
  AND2_X1 U15957 ( .A1(n15899), .A2(n16394), .ZN(n19778) );
  NAND2_X1 U15958 ( .A1(n12477), .A2(n19788), .ZN(n12478) );
  NAND2_X1 U15959 ( .A1(n9648), .A2(n12478), .ZN(n19779) );
  NAND2_X1 U15960 ( .A1(n19778), .A2(n19779), .ZN(n15885) );
  AND2_X1 U15961 ( .A1(n9648), .A2(n10418), .ZN(n12479) );
  NOR2_X1 U15962 ( .A1(n12482), .A2(n12479), .ZN(n16367) );
  OR2_X1 U15963 ( .A1(n15885), .A2(n16367), .ZN(n19763) );
  NAND2_X1 U15964 ( .A1(n12484), .A2(n12480), .ZN(n12481) );
  NAND2_X1 U15965 ( .A1(n9629), .A2(n12481), .ZN(n16348) );
  OR2_X1 U15966 ( .A1(n12482), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12483) );
  NAND2_X1 U15967 ( .A1(n12484), .A2(n12483), .ZN(n19765) );
  NAND2_X1 U15968 ( .A1(n16348), .A2(n19765), .ZN(n12485) );
  NOR2_X1 U15969 ( .A1(n19763), .A2(n12485), .ZN(n15870) );
  AND2_X1 U15970 ( .A1(n9629), .A2(n12486), .ZN(n12487) );
  OR2_X1 U15971 ( .A1(n12487), .A2(n12488), .ZN(n16338) );
  AND2_X1 U15972 ( .A1(n15870), .A2(n16338), .ZN(n15843) );
  NOR2_X1 U15973 ( .A1(n12488), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12489) );
  OR2_X1 U15974 ( .A1(n12490), .A2(n12489), .ZN(n16318) );
  NAND2_X1 U15975 ( .A1(n15843), .A2(n16318), .ZN(n15845) );
  OR2_X1 U15976 ( .A1(n12490), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12491) );
  AND2_X1 U15977 ( .A1(n9645), .A2(n12491), .ZN(n16314) );
  OR2_X1 U15978 ( .A1(n15845), .A2(n16314), .ZN(n15816) );
  NAND2_X1 U15979 ( .A1(n9645), .A2(n12492), .ZN(n12493) );
  AND2_X1 U15980 ( .A1(n9632), .A2(n12493), .ZN(n15817) );
  NOR2_X1 U15981 ( .A1(n15816), .A2(n15817), .ZN(n15806) );
  NAND2_X1 U15982 ( .A1(n9632), .A2(n12494), .ZN(n12495) );
  NAND2_X1 U15983 ( .A1(n12496), .A2(n12495), .ZN(n16294) );
  NAND2_X1 U15984 ( .A1(n15806), .A2(n16294), .ZN(n15775) );
  AND2_X1 U15985 ( .A1(n12496), .A2(n16285), .ZN(n12497) );
  NOR2_X1 U15986 ( .A1(n12498), .A2(n12497), .ZN(n16288) );
  OR2_X1 U15987 ( .A1(n15775), .A2(n16288), .ZN(n15776) );
  OR2_X1 U15988 ( .A1(n12498), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12499) );
  AND2_X1 U15989 ( .A1(n12499), .A2(n11176), .ZN(n16273) );
  NOR2_X1 U15990 ( .A1(n15776), .A2(n16273), .ZN(n15762) );
  AND2_X1 U15991 ( .A1(n15762), .A2(n15761), .ZN(n15763) );
  AND2_X1 U15992 ( .A1(n12500), .A2(n15755), .ZN(n12501) );
  OR2_X1 U15993 ( .A1(n12501), .A2(n12503), .ZN(n16266) );
  OR2_X1 U15994 ( .A1(n12503), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12504) );
  AND2_X1 U15995 ( .A1(n12506), .A2(n12504), .ZN(n17310) );
  NAND2_X1 U15996 ( .A1(n12506), .A2(n12505), .ZN(n12507) );
  NAND2_X1 U15997 ( .A1(n9760), .A2(n12507), .ZN(n16246) );
  AND2_X1 U15998 ( .A1(n9760), .A2(n16238), .ZN(n12509) );
  NOR2_X1 U15999 ( .A1(n12508), .A2(n12509), .ZN(n16236) );
  NOR2_X1 U16000 ( .A1(n12508), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12510) );
  OR2_X1 U16001 ( .A1(n12512), .A2(n12510), .ZN(n16229) );
  OR2_X1 U16002 ( .A1(n12512), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12513) );
  AND2_X1 U16003 ( .A1(n12511), .A2(n12513), .ZN(n16218) );
  AOI21_X1 U16004 ( .B1(n15706), .B2(n15968), .A(n16218), .ZN(n15678) );
  NAND2_X1 U16005 ( .A1(n12511), .A2(n12514), .ZN(n12515) );
  NAND2_X1 U16006 ( .A1(n12516), .A2(n12515), .ZN(n16207) );
  OAI21_X1 U16007 ( .B1(n15678), .B2(n19815), .A(n16207), .ZN(n15670) );
  NAND2_X1 U16008 ( .A1(n12516), .A2(n16200), .ZN(n12517) );
  AOI21_X1 U16009 ( .B1(n15670), .B2(n15968), .A(n10605), .ZN(n12521) );
  INV_X1 U16010 ( .A(n13734), .ZN(n12520) );
  NAND2_X1 U16011 ( .A1(n9737), .A2(n12518), .ZN(n12519) );
  NAND2_X1 U16012 ( .A1(n12520), .A2(n12519), .ZN(n16187) );
  OAI21_X1 U16013 ( .B1(n12521), .B2(n16187), .A(n19820), .ZN(n12522) );
  OAI21_X1 U16014 ( .B1(n12521), .B2(n19815), .A(n16187), .ZN(n13745) );
  INV_X1 U16015 ( .A(n13745), .ZN(n13742) );
  AOI21_X1 U16016 ( .B1(n17314), .B2(n12522), .A(n13742), .ZN(n12523) );
  AOI22_X1 U16017 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n14723), .B1(
        n12524), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U16018 ( .A1(n12525), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12526) );
  INV_X1 U16019 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20594) );
  NAND2_X1 U16020 ( .A1(n12524), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n12529) );
  NAND2_X1 U16021 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12528) );
  OAI211_X1 U16022 ( .C1(n14727), .C2(n20594), .A(n12529), .B(n12528), .ZN(
        n12530) );
  NOR2_X1 U16023 ( .A1(n15663), .A2(n12530), .ZN(n12531) );
  NOR2_X1 U16024 ( .A1(n14164), .A2(n16888), .ZN(n12533) );
  NAND2_X1 U16025 ( .A1(n12533), .A2(n13910), .ZN(n19837) );
  NAND2_X1 U16026 ( .A1(n13987), .A2(n20408), .ZN(n15653) );
  NOR2_X1 U16027 ( .A1(n15653), .A2(n12534), .ZN(n16880) );
  NAND2_X1 U16028 ( .A1(n16880), .A2(n16856), .ZN(n12535) );
  NAND2_X1 U16029 ( .A1(n13390), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13381) );
  INV_X1 U16030 ( .A(n13381), .ZN(n12536) );
  NAND2_X1 U16031 ( .A1(n13390), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13388) );
  XNOR2_X1 U16032 ( .A(n13389), .B(n13388), .ZN(n13386) );
  AND2_X1 U16033 ( .A1(n16887), .A2(n20408), .ZN(n12537) );
  NOR2_X1 U16034 ( .A1(n13889), .A2(n12537), .ZN(n12540) );
  INV_X1 U16035 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14716) );
  NOR2_X1 U16036 ( .A1(n13987), .A2(n14716), .ZN(n12538) );
  NAND2_X1 U16037 ( .A1(n14358), .A2(n20408), .ZN(n12539) );
  NAND2_X1 U16038 ( .A1(n13926), .A2(n12539), .ZN(n14717) );
  NAND2_X1 U16039 ( .A1(n12540), .A2(n14716), .ZN(n12541) );
  AND2_X1 U16040 ( .A1(n20619), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12542) );
  NAND2_X1 U16041 ( .A1(n12543), .A2(n12542), .ZN(n16886) );
  NAND2_X1 U16042 ( .A1(n19838), .A2(n16886), .ZN(n12544) );
  NOR2_X1 U16043 ( .A1(n12544), .A2(n16423), .ZN(n12545) );
  AOI22_X1 U16044 ( .A1(n19830), .A2(P2_EBX_REG_29__SCAN_IN), .B1(n19827), 
        .B2(P2_REIP_REG_29__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U16045 ( .A1(n19841), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12546) );
  OAI211_X1 U16046 ( .C1(n13386), .C2(n19809), .A(n12547), .B(n12546), .ZN(
        n12548) );
  NAND2_X1 U16047 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12552) );
  NAND2_X1 U16048 ( .A1(n12555), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U16049 ( .A1(n13774), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12550) );
  AND3_X1 U16050 ( .A1(n12552), .A2(n12551), .A3(n12550), .ZN(n15665) );
  NAND2_X1 U16051 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12558) );
  NAND2_X1 U16052 ( .A1(n12555), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U16053 ( .A1(n13774), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12556) );
  AND2_X1 U16054 ( .A1(n12560), .A2(n12559), .ZN(n12561) );
  INV_X1 U16055 ( .A(n16184), .ZN(n12563) );
  NAND2_X1 U16056 ( .A1(n11232), .A2(n16887), .ZN(n12562) );
  NAND3_X1 U16057 ( .A1(n12566), .A2(n12565), .A3(n12564), .ZN(P2_U2826) );
  NOR4_X1 U16058 ( .A1(n12567), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12568) );
  NAND2_X1 U16059 ( .A1(n9928), .A2(n12568), .ZN(n12571) );
  NAND3_X1 U16060 ( .A1(n12569), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12570) );
  XNOR2_X1 U16061 ( .A(n12573), .B(n12572), .ZN(n15412) );
  INV_X1 U16062 ( .A(n15642), .ZN(n14486) );
  INV_X1 U16063 ( .A(n13853), .ZN(n12575) );
  NAND2_X1 U16064 ( .A1(n12575), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12610) );
  NOR2_X1 U16065 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12576), .ZN(
        n12577) );
  NOR2_X1 U16066 ( .A1(n12611), .A2(n12577), .ZN(n20732) );
  INV_X1 U16067 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21447) );
  NAND2_X1 U16068 ( .A1(n12586), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14427) );
  OAI22_X1 U16069 ( .A1(n20732), .A2(n13797), .B1(n21447), .B2(n14427), .ZN(
        n12578) );
  AOI21_X1 U16070 ( .B1(n13787), .B2(P1_EAX_REG_3__SCAN_IN), .A(n12578), .ZN(
        n12579) );
  OAI21_X1 U16071 ( .B1(n14486), .B2(n12610), .A(n12579), .ZN(n12580) );
  AOI21_X1 U16072 ( .B1(n12581), .B2(n12756), .A(n12580), .ZN(n14409) );
  NAND2_X1 U16073 ( .A1(n14507), .A2(n12756), .ZN(n12590) );
  AOI22_X1 U16074 ( .A1(n13787), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n12586), .ZN(n12588) );
  INV_X1 U16075 ( .A(n12610), .ZN(n12602) );
  NAND2_X1 U16076 ( .A1(n12602), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12587) );
  AND2_X1 U16077 ( .A1(n12588), .A2(n12587), .ZN(n12589) );
  NAND2_X1 U16078 ( .A1(n20889), .A2(n12591), .ZN(n12592) );
  NAND2_X1 U16079 ( .A1(n12592), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14103) );
  NAND2_X1 U16080 ( .A1(n12586), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12595) );
  NAND2_X1 U16081 ( .A1(n12621), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12594) );
  OAI211_X1 U16082 ( .C1(n12610), .C2(n12593), .A(n12595), .B(n12594), .ZN(
        n12596) );
  AOI21_X1 U16083 ( .B1(n20921), .B2(n12756), .A(n12596), .ZN(n12597) );
  INV_X1 U16084 ( .A(n12597), .ZN(n14105) );
  OR2_X1 U16085 ( .A1(n14105), .A2(n13797), .ZN(n12598) );
  NAND2_X1 U16086 ( .A1(n14104), .A2(n12598), .ZN(n14185) );
  NAND2_X1 U16087 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12599) );
  INV_X1 U16088 ( .A(n14410), .ZN(n12600) );
  INV_X1 U16089 ( .A(n12756), .ZN(n12664) );
  NAND2_X1 U16090 ( .A1(n12602), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12603) );
  NAND2_X1 U16091 ( .A1(n13787), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n14424) );
  XNOR2_X1 U16092 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15065) );
  NAND2_X1 U16093 ( .A1(n15065), .A2(n13683), .ZN(n14423) );
  NAND3_X1 U16094 ( .A1(n14424), .A2(n14427), .A3(n14423), .ZN(n12606) );
  OR2_X2 U16095 ( .A1(n14426), .A2(n12606), .ZN(n14411) );
  NAND2_X1 U16096 ( .A1(n12607), .A2(n14411), .ZN(n14408) );
  NAND2_X1 U16097 ( .A1(n12586), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12609) );
  NAND2_X1 U16098 ( .A1(n13787), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12608) );
  OAI211_X1 U16099 ( .C1(n12610), .C2(n13981), .A(n12609), .B(n12608), .ZN(
        n12612) );
  NAND2_X1 U16100 ( .A1(n12611), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12615) );
  OAI21_X1 U16101 ( .B1(n12611), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n12615), .ZN(n14537) );
  MUX2_X1 U16102 ( .A(n12612), .B(n14537), .S(n13683), .Z(n12613) );
  AOI21_X1 U16103 ( .B1(n12614), .B2(n12756), .A(n12613), .ZN(n14542) );
  AND2_X1 U16104 ( .A1(n12615), .A2(n20701), .ZN(n12616) );
  OR2_X1 U16105 ( .A1(n12616), .A2(n12622), .ZN(n20712) );
  NAND2_X1 U16106 ( .A1(n20712), .A2(n13683), .ZN(n12617) );
  OAI21_X1 U16107 ( .B1(n14427), .B2(n20701), .A(n12617), .ZN(n12618) );
  AOI21_X1 U16108 ( .B1(n13787), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12618), .ZN(
        n12619) );
  NAND2_X1 U16109 ( .A1(n14541), .A2(n14553), .ZN(n14552) );
  INV_X1 U16110 ( .A(n14552), .ZN(n12629) );
  INV_X1 U16111 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12625) );
  NOR2_X1 U16112 ( .A1(n12622), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12623) );
  OR2_X1 U16113 ( .A1(n12630), .A2(n12623), .ZN(n20691) );
  AOI22_X1 U16114 ( .A1(n20691), .A2(n13683), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13786), .ZN(n12624) );
  OAI21_X1 U16115 ( .B1(n12605), .B2(n12625), .A(n12624), .ZN(n12626) );
  AOI21_X1 U16116 ( .B1(n12627), .B2(n12756), .A(n12626), .ZN(n14634) );
  NOR2_X1 U16117 ( .A1(n12630), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12631) );
  OR2_X1 U16118 ( .A1(n12659), .A2(n12631), .ZN(n20680) );
  AOI22_X1 U16119 ( .A1(n20680), .A2(n13683), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13786), .ZN(n12632) );
  OAI21_X1 U16120 ( .B1(n12605), .B2(n20769), .A(n12632), .ZN(n12633) );
  AOI21_X1 U16121 ( .B1(n12634), .B2(n12756), .A(n12633), .ZN(n14625) );
  AOI22_X1 U16122 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12879), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12638) );
  AOI22_X1 U16123 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n12945), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12637) );
  AOI22_X1 U16124 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n9582), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U16125 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12635) );
  NAND4_X1 U16126 ( .A1(n12638), .A2(n12637), .A3(n12636), .A4(n12635), .ZN(
        n12644) );
  AOI22_X1 U16127 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U16128 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U16129 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12884), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U16130 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12639) );
  NAND4_X1 U16131 ( .A1(n12642), .A2(n12641), .A3(n12640), .A4(n12639), .ZN(
        n12643) );
  OAI21_X1 U16132 ( .B1(n12644), .B2(n12643), .A(n12756), .ZN(n12648) );
  NAND2_X1 U16133 ( .A1(n13787), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12647) );
  XNOR2_X1 U16134 ( .A(n12659), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15383) );
  NAND2_X1 U16135 ( .A1(n15383), .A2(n13683), .ZN(n12646) );
  NAND2_X1 U16136 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12645) );
  AOI22_X1 U16137 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U16138 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U16139 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U16140 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12649) );
  NAND4_X1 U16141 ( .A1(n12652), .A2(n12651), .A3(n12650), .A4(n12649), .ZN(
        n12658) );
  AOI22_X1 U16142 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12945), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U16143 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U16144 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U16145 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12653) );
  NAND4_X1 U16146 ( .A1(n12656), .A2(n12655), .A3(n12654), .A4(n12653), .ZN(
        n12657) );
  NOR2_X1 U16147 ( .A1(n12658), .A2(n12657), .ZN(n12663) );
  XOR2_X1 U16148 ( .A(n20665), .B(n12665), .Z(n20669) );
  INV_X1 U16149 ( .A(n20669), .ZN(n12660) );
  AOI22_X1 U16150 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n13786), .B1(
        n13683), .B2(n12660), .ZN(n12662) );
  NAND2_X1 U16151 ( .A1(n13787), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12661) );
  OAI211_X1 U16152 ( .C1(n12664), .C2(n12663), .A(n12662), .B(n12661), .ZN(
        n14650) );
  XNOR2_X1 U16153 ( .A(n12680), .B(n12679), .ZN(n15369) );
  NAND2_X1 U16154 ( .A1(n15369), .A2(n13683), .ZN(n12678) );
  AOI22_X1 U16155 ( .A1(n13787), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13786), .ZN(n12677) );
  AOI22_X1 U16156 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12945), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U16157 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U16158 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U16159 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12666) );
  NAND4_X1 U16160 ( .A1(n12669), .A2(n12668), .A3(n12667), .A4(n12666), .ZN(
        n12675) );
  AOI22_X1 U16161 ( .A1(n13667), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U16162 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U16163 ( .A1(n12052), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U16164 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12670) );
  NAND4_X1 U16165 ( .A1(n12673), .A2(n12672), .A3(n12671), .A4(n12670), .ZN(
        n12674) );
  OAI21_X1 U16166 ( .B1(n12675), .B2(n12674), .A(n12756), .ZN(n12676) );
  INV_X1 U16167 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14959) );
  XNOR2_X1 U16168 ( .A(n12778), .B(n14959), .ZN(n15315) );
  AOI22_X1 U16169 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U16170 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U16171 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U16172 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12681) );
  NAND4_X1 U16173 ( .A1(n12684), .A2(n12683), .A3(n12682), .A4(n12681), .ZN(
        n12691) );
  AOI22_X1 U16174 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12945), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U16175 ( .A1(n12685), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U16176 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U16177 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12686) );
  NAND4_X1 U16178 ( .A1(n12689), .A2(n12688), .A3(n12687), .A4(n12686), .ZN(
        n12690) );
  OAI21_X1 U16179 ( .B1(n12691), .B2(n12690), .A(n12756), .ZN(n12694) );
  NAND2_X1 U16180 ( .A1(n13787), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12693) );
  NAND2_X1 U16181 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12692) );
  NAND3_X1 U16182 ( .A1(n12694), .A2(n12693), .A3(n12692), .ZN(n12695) );
  AOI21_X1 U16183 ( .B1(n15315), .B2(n13683), .A(n12695), .ZN(n14953) );
  INV_X1 U16184 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12696) );
  XNOR2_X1 U16185 ( .A(n12697), .B(n12696), .ZN(n15326) );
  AOI22_X1 U16186 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U16187 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U16188 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U16189 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12698) );
  NAND4_X1 U16190 ( .A1(n12701), .A2(n12700), .A3(n12699), .A4(n12698), .ZN(
        n12707) );
  AOI22_X1 U16191 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U16192 ( .A1(n11919), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U16193 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U16194 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12702) );
  NAND4_X1 U16195 ( .A1(n12705), .A2(n12704), .A3(n12703), .A4(n12702), .ZN(
        n12706) );
  OAI21_X1 U16196 ( .B1(n12707), .B2(n12706), .A(n12756), .ZN(n12710) );
  NAND2_X1 U16197 ( .A1(n13787), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12709) );
  NAND2_X1 U16198 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12708) );
  NAND3_X1 U16199 ( .A1(n12710), .A2(n12709), .A3(n12708), .ZN(n12711) );
  AOI21_X1 U16200 ( .B1(n15326), .B2(n13683), .A(n12711), .ZN(n14952) );
  AOI22_X1 U16201 ( .A1(n13667), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U16202 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U16203 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U16204 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12713) );
  NAND4_X1 U16205 ( .A1(n12716), .A2(n12715), .A3(n12714), .A4(n12713), .ZN(
        n12722) );
  AOI22_X1 U16206 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12945), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U16207 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U16208 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U16209 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12717) );
  NAND4_X1 U16210 ( .A1(n12720), .A2(n12719), .A3(n12718), .A4(n12717), .ZN(
        n12721) );
  OR2_X1 U16211 ( .A1(n12722), .A2(n12721), .ZN(n12723) );
  AND2_X1 U16212 ( .A1(n12756), .A2(n12723), .ZN(n14949) );
  INV_X1 U16213 ( .A(n12724), .ZN(n12725) );
  INV_X1 U16214 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15026) );
  NAND2_X1 U16215 ( .A1(n12725), .A2(n15026), .ZN(n12726) );
  NAND2_X1 U16216 ( .A1(n12747), .A2(n12726), .ZN(n15356) );
  NAND2_X1 U16217 ( .A1(n15356), .A2(n13683), .ZN(n12728) );
  AOI22_X1 U16218 ( .A1(n13787), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13786), .ZN(n12727) );
  NAND2_X1 U16219 ( .A1(n12728), .A2(n12727), .ZN(n14982) );
  OR2_X1 U16220 ( .A1(n12747), .A2(n12746), .ZN(n12730) );
  XNOR2_X1 U16221 ( .A(n12730), .B(n12729), .ZN(n15338) );
  NAND2_X1 U16222 ( .A1(n15338), .A2(n13683), .ZN(n12745) );
  AOI22_X1 U16223 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U16224 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U16225 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U16226 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12731) );
  NAND4_X1 U16227 ( .A1(n12734), .A2(n12733), .A3(n12732), .A4(n12731), .ZN(
        n12740) );
  AOI22_X1 U16228 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U16229 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U16230 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U16231 ( .A1(n12052), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12735) );
  NAND4_X1 U16232 ( .A1(n12738), .A2(n12737), .A3(n12736), .A4(n12735), .ZN(
        n12739) );
  OAI21_X1 U16233 ( .B1(n12740), .B2(n12739), .A(n12756), .ZN(n12743) );
  NAND2_X1 U16234 ( .A1(n13787), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12742) );
  NAND2_X1 U16235 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12741) );
  AND3_X1 U16236 ( .A1(n12743), .A2(n12742), .A3(n12741), .ZN(n12744) );
  NAND2_X1 U16237 ( .A1(n12745), .A2(n12744), .ZN(n14984) );
  XNOR2_X1 U16238 ( .A(n12747), .B(n12746), .ZN(n15346) );
  NAND2_X1 U16239 ( .A1(n15346), .A2(n13683), .ZN(n12762) );
  AOI22_X1 U16240 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U16241 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U16242 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U16243 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12748) );
  NAND4_X1 U16244 ( .A1(n12751), .A2(n12750), .A3(n12749), .A4(n12748), .ZN(
        n12758) );
  AOI22_X1 U16245 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12945), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U16246 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U16247 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U16248 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12752) );
  NAND4_X1 U16249 ( .A1(n12755), .A2(n12754), .A3(n12753), .A4(n12752), .ZN(
        n12757) );
  OAI21_X1 U16250 ( .B1(n12758), .B2(n12757), .A(n12756), .ZN(n12761) );
  NAND2_X1 U16251 ( .A1(n13787), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12760) );
  NAND2_X1 U16252 ( .A1(n13786), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12759) );
  NAND2_X1 U16253 ( .A1(n12762), .A2(n10601), .ZN(n15005) );
  OAI211_X1 U16254 ( .C1(n14949), .C2(n14982), .A(n14984), .B(n15005), .ZN(
        n12763) );
  INV_X1 U16255 ( .A(n15626), .ZN(n12765) );
  AOI22_X1 U16256 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U16257 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U16258 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U16259 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12005), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12766) );
  NAND4_X1 U16260 ( .A1(n12769), .A2(n12768), .A3(n12767), .A4(n12766), .ZN(
        n12775) );
  AOI22_X1 U16261 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n12945), .B1(
        n13698), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U16262 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n12884), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12772) );
  AOI22_X1 U16263 ( .A1(n12052), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U16264 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n9587), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12770) );
  NAND4_X1 U16265 ( .A1(n12773), .A2(n12772), .A3(n12771), .A4(n12770), .ZN(
        n12774) );
  NOR2_X1 U16266 ( .A1(n12775), .A2(n12774), .ZN(n12777) );
  AOI22_X1 U16267 ( .A1(n13787), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12586), .ZN(n12776) );
  OAI21_X1 U16268 ( .B1(n13709), .B2(n12777), .A(n12776), .ZN(n12783) );
  NAND2_X1 U16269 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  NAND2_X1 U16270 ( .A1(n12812), .A2(n12782), .ZN(n15304) );
  MUX2_X1 U16271 ( .A(n12783), .B(n15304), .S(n13683), .Z(n14929) );
  INV_X1 U16272 ( .A(n14911), .ZN(n12799) );
  INV_X1 U16273 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12784) );
  XNOR2_X1 U16274 ( .A(n12812), .B(n12784), .ZN(n15288) );
  AOI22_X1 U16275 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U16276 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U16277 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U16278 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12785) );
  NAND4_X1 U16279 ( .A1(n12788), .A2(n12787), .A3(n12786), .A4(n12785), .ZN(
        n12794) );
  AOI22_X1 U16280 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U16281 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U16282 ( .A1(n12052), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U16283 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12789) );
  NAND4_X1 U16284 ( .A1(n12792), .A2(n12791), .A3(n12790), .A4(n12789), .ZN(
        n12793) );
  NOR2_X1 U16285 ( .A1(n12794), .A2(n12793), .ZN(n12796) );
  AOI22_X1 U16286 ( .A1(n13787), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n13786), .ZN(n12795) );
  OAI21_X1 U16287 ( .B1(n13709), .B2(n12796), .A(n12795), .ZN(n12797) );
  AOI21_X1 U16288 ( .B1(n15288), .B2(n13683), .A(n12797), .ZN(n14914) );
  AOI22_X1 U16289 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U16290 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U16291 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U16292 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12800) );
  NAND4_X1 U16293 ( .A1(n12803), .A2(n12802), .A3(n12801), .A4(n12800), .ZN(
        n12809) );
  AOI22_X1 U16294 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U16295 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U16296 ( .A1(n12052), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U16297 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12804) );
  NAND4_X1 U16298 ( .A1(n12807), .A2(n12806), .A3(n12805), .A4(n12804), .ZN(
        n12808) );
  NOR2_X1 U16299 ( .A1(n12809), .A2(n12808), .ZN(n12811) );
  AOI22_X1 U16300 ( .A1(n13787), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12586), .ZN(n12810) );
  OAI21_X1 U16301 ( .B1(n13709), .B2(n12811), .A(n12810), .ZN(n12815) );
  NAND2_X1 U16302 ( .A1(n12813), .A2(n14903), .ZN(n12814) );
  NAND2_X1 U16303 ( .A1(n12829), .A2(n12814), .ZN(n15277) );
  MUX2_X1 U16304 ( .A(n12815), .B(n15277), .S(n13683), .Z(n14901) );
  XNOR2_X1 U16305 ( .A(n12829), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15271) );
  AOI22_X1 U16306 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12945), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U16307 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U16308 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U16309 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12816) );
  NAND4_X1 U16310 ( .A1(n12819), .A2(n12818), .A3(n12817), .A4(n12816), .ZN(
        n12825) );
  AOI22_X1 U16311 ( .A1(n13667), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U16312 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U16313 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U16314 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12820) );
  NAND4_X1 U16315 ( .A1(n12823), .A2(n12822), .A3(n12821), .A4(n12820), .ZN(
        n12824) );
  OR2_X1 U16316 ( .A1(n12825), .A2(n12824), .ZN(n12827) );
  INV_X1 U16317 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15152) );
  INV_X1 U16318 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15273) );
  OAI22_X1 U16319 ( .A1(n12605), .A2(n15152), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15273), .ZN(n12826) );
  AOI21_X1 U16320 ( .B1(n13679), .B2(n12827), .A(n12826), .ZN(n12828) );
  MUX2_X1 U16321 ( .A(n15271), .B(n12828), .S(n13797), .Z(n14880) );
  NAND2_X1 U16322 ( .A1(n12831), .A2(n12830), .ZN(n12832) );
  NAND2_X1 U16323 ( .A1(n12860), .A2(n12832), .ZN(n15263) );
  AOI22_X1 U16324 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U16325 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U16326 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U16327 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9585), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12833) );
  NAND4_X1 U16328 ( .A1(n12836), .A2(n12835), .A3(n12834), .A4(n12833), .ZN(
        n12842) );
  AOI22_X1 U16329 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U16330 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U16331 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U16332 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12837) );
  NAND4_X1 U16333 ( .A1(n12840), .A2(n12839), .A3(n12838), .A4(n12837), .ZN(
        n12841) );
  NOR2_X1 U16334 ( .A1(n12842), .A2(n12841), .ZN(n12844) );
  AOI22_X1 U16335 ( .A1(n13787), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12586), .ZN(n12843) );
  OAI21_X1 U16336 ( .B1(n13709), .B2(n12844), .A(n12843), .ZN(n12845) );
  MUX2_X1 U16337 ( .A(n15263), .B(n12845), .S(n13797), .Z(n14863) );
  INV_X1 U16338 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12846) );
  XNOR2_X1 U16339 ( .A(n12860), .B(n12846), .ZN(n15250) );
  AOI22_X1 U16340 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U16341 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U16342 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12848) );
  AOI22_X1 U16343 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12847) );
  NAND4_X1 U16344 ( .A1(n12850), .A2(n12849), .A3(n12848), .A4(n12847), .ZN(
        n12856) );
  AOI22_X1 U16345 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U16346 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U16347 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U16348 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9590), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12851) );
  NAND4_X1 U16349 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n12855) );
  NOR2_X1 U16350 ( .A1(n12856), .A2(n12855), .ZN(n12858) );
  AOI22_X1 U16351 ( .A1(n13787), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12586), .ZN(n12857) );
  OAI21_X1 U16352 ( .B1(n13709), .B2(n12858), .A(n12857), .ZN(n12859) );
  MUX2_X1 U16353 ( .A(n15250), .B(n12859), .S(n13797), .Z(n14854) );
  NAND2_X1 U16354 ( .A1(n12862), .A2(n12861), .ZN(n12863) );
  NAND2_X1 U16355 ( .A1(n12905), .A2(n12863), .ZN(n15245) );
  AOI22_X1 U16356 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U16357 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U16358 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12865) );
  AOI22_X1 U16359 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12864) );
  NAND4_X1 U16360 ( .A1(n12867), .A2(n12866), .A3(n12865), .A4(n12864), .ZN(
        n12873) );
  AOI22_X1 U16361 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U16362 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13698), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U16363 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12869) );
  AOI22_X1 U16364 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12868) );
  NAND4_X1 U16365 ( .A1(n12871), .A2(n12870), .A3(n12869), .A4(n12868), .ZN(
        n12872) );
  NOR2_X1 U16366 ( .A1(n12873), .A2(n12872), .ZN(n12875) );
  AOI22_X1 U16367 ( .A1(n13787), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12586), .ZN(n12874) );
  OAI21_X1 U16368 ( .B1(n13709), .B2(n12875), .A(n12874), .ZN(n12876) );
  MUX2_X1 U16369 ( .A(n15245), .B(n12876), .S(n13797), .Z(n12877) );
  AOI22_X1 U16370 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12883) );
  AOI22_X1 U16371 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12882) );
  AOI22_X1 U16372 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12881) );
  AOI22_X1 U16373 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12880) );
  NAND4_X1 U16374 ( .A1(n12883), .A2(n12882), .A3(n12881), .A4(n12880), .ZN(
        n12890) );
  AOI22_X1 U16375 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U16376 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U16377 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U16378 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12885) );
  NAND4_X1 U16379 ( .A1(n12888), .A2(n12887), .A3(n12886), .A4(n12885), .ZN(
        n12889) );
  NOR2_X1 U16380 ( .A1(n12890), .A2(n12889), .ZN(n12909) );
  AOI22_X1 U16381 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U16382 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U16383 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12892) );
  AOI22_X1 U16384 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12891) );
  NAND4_X1 U16385 ( .A1(n12894), .A2(n12893), .A3(n12892), .A4(n12891), .ZN(
        n12900) );
  AOI22_X1 U16386 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n12945), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U16387 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12897) );
  AOI22_X1 U16388 ( .A1(n12052), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U16389 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n9587), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12895) );
  NAND4_X1 U16390 ( .A1(n12898), .A2(n12897), .A3(n12896), .A4(n12895), .ZN(
        n12899) );
  NOR2_X1 U16391 ( .A1(n12900), .A2(n12899), .ZN(n12910) );
  XOR2_X1 U16392 ( .A(n12909), .B(n12910), .Z(n12903) );
  INV_X1 U16393 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12901) );
  INV_X1 U16394 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15235) );
  OAI22_X1 U16395 ( .A1(n12605), .A2(n12901), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15235), .ZN(n12902) );
  AOI21_X1 U16396 ( .B1(n13679), .B2(n12903), .A(n12902), .ZN(n12904) );
  XNOR2_X1 U16397 ( .A(n12905), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15233) );
  MUX2_X1 U16398 ( .A(n12904), .B(n15233), .S(n13683), .Z(n14824) );
  INV_X1 U16399 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12906) );
  NAND2_X1 U16400 ( .A1(n12907), .A2(n12906), .ZN(n12908) );
  NAND2_X1 U16401 ( .A1(n12959), .A2(n12908), .ZN(n15223) );
  NOR2_X1 U16402 ( .A1(n12910), .A2(n12909), .ZN(n12926) );
  INV_X1 U16403 ( .A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n21450) );
  AOI22_X1 U16404 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U16405 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U16406 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12913) );
  AOI22_X1 U16407 ( .A1(n12931), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12912) );
  NAND4_X1 U16408 ( .A1(n12915), .A2(n12914), .A3(n12913), .A4(n12912), .ZN(
        n12921) );
  AOI22_X1 U16409 ( .A1(n12884), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U16410 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16411 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16412 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12916) );
  NAND4_X1 U16413 ( .A1(n12919), .A2(n12918), .A3(n12917), .A4(n12916), .ZN(
        n12920) );
  OR2_X1 U16414 ( .A1(n12921), .A2(n12920), .ZN(n12925) );
  XNOR2_X1 U16415 ( .A(n12926), .B(n12925), .ZN(n12923) );
  AOI22_X1 U16416 ( .A1(n13787), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12586), .ZN(n12922) );
  OAI21_X1 U16417 ( .B1(n12923), .B2(n13709), .A(n12922), .ZN(n12924) );
  MUX2_X1 U16418 ( .A(n15223), .B(n12924), .S(n13797), .Z(n14813) );
  XNOR2_X1 U16419 ( .A(n12959), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15219) );
  NAND2_X1 U16420 ( .A1(n12926), .A2(n12925), .ZN(n12943) );
  AOI22_X1 U16421 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U16422 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U16423 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U16424 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12927) );
  NAND4_X1 U16425 ( .A1(n12930), .A2(n12929), .A3(n12928), .A4(n12927), .ZN(
        n12937) );
  AOI22_X1 U16426 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U16427 ( .A1(n12911), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U16428 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12933) );
  AOI22_X1 U16429 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12932) );
  NAND4_X1 U16430 ( .A1(n12935), .A2(n12934), .A3(n12933), .A4(n12932), .ZN(
        n12936) );
  NOR2_X1 U16431 ( .A1(n12937), .A2(n12936), .ZN(n12944) );
  XOR2_X1 U16432 ( .A(n12943), .B(n12944), .Z(n12939) );
  INV_X1 U16433 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15130) );
  OAI22_X1 U16434 ( .A1(n12605), .A2(n15130), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15217), .ZN(n12938) );
  AOI21_X1 U16435 ( .B1(n12939), .B2(n13679), .A(n12938), .ZN(n12940) );
  MUX2_X1 U16436 ( .A(n15219), .B(n12940), .S(n13797), .Z(n14800) );
  NOR2_X1 U16437 ( .A1(n12944), .A2(n12943), .ZN(n12965) );
  AOI22_X1 U16438 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U16439 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U16440 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12911), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U16441 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12116), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12946) );
  NAND4_X1 U16442 ( .A1(n12949), .A2(n12948), .A3(n12947), .A4(n12946), .ZN(
        n12955) );
  AOI22_X1 U16443 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U16444 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12952) );
  AOI22_X1 U16445 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U16446 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9590), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12950) );
  NAND4_X1 U16447 ( .A1(n12953), .A2(n12952), .A3(n12951), .A4(n12950), .ZN(
        n12954) );
  INV_X1 U16448 ( .A(n12964), .ZN(n12956) );
  XNOR2_X1 U16449 ( .A(n12965), .B(n12956), .ZN(n12958) );
  INV_X1 U16450 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15125) );
  INV_X1 U16451 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15205) );
  OAI22_X1 U16452 ( .A1(n12605), .A2(n15125), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15205), .ZN(n12957) );
  AOI21_X1 U16453 ( .B1(n12958), .B2(n13679), .A(n12957), .ZN(n12963) );
  INV_X1 U16454 ( .A(n12960), .ZN(n12961) );
  NAND2_X1 U16455 ( .A1(n12961), .A2(n15205), .ZN(n12962) );
  AND2_X1 U16456 ( .A1(n12997), .A2(n12962), .ZN(n15207) );
  MUX2_X1 U16457 ( .A(n12963), .B(n15207), .S(n13683), .Z(n14789) );
  XNOR2_X1 U16458 ( .A(n12997), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15194) );
  NAND2_X1 U16459 ( .A1(n15194), .A2(n13683), .ZN(n12982) );
  NAND2_X1 U16460 ( .A1(n12965), .A2(n12964), .ZN(n12983) );
  AOI22_X1 U16461 ( .A1(n13667), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U16462 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U16463 ( .A1(n12052), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16464 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12966) );
  NAND4_X1 U16465 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        n12975) );
  AOI22_X1 U16466 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12945), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16467 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16468 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16469 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12970) );
  NAND4_X1 U16470 ( .A1(n12973), .A2(n12972), .A3(n12971), .A4(n12970), .ZN(
        n12974) );
  NOR2_X1 U16471 ( .A1(n12975), .A2(n12974), .ZN(n12984) );
  XOR2_X1 U16472 ( .A(n12983), .B(n12984), .Z(n12976) );
  NAND2_X1 U16473 ( .A1(n12976), .A2(n13679), .ZN(n12980) );
  INV_X1 U16474 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12977) );
  AOI21_X1 U16475 ( .B1(n12977), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12978) );
  AOI21_X1 U16476 ( .B1(n13787), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12978), .ZN(
        n12979) );
  NAND2_X1 U16477 ( .A1(n12980), .A2(n12979), .ZN(n12981) );
  NAND2_X1 U16478 ( .A1(n12982), .A2(n12981), .ZN(n14777) );
  NOR2_X1 U16479 ( .A1(n12984), .A2(n12983), .ZN(n13666) );
  AOI22_X1 U16480 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12024), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16481 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16482 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U16483 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12985) );
  NAND4_X1 U16484 ( .A1(n12988), .A2(n12987), .A3(n12986), .A4(n12985), .ZN(
        n12994) );
  AOI22_X1 U16485 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16486 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16487 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16488 ( .A1(n12118), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12989) );
  NAND4_X1 U16489 ( .A1(n12992), .A2(n12991), .A3(n12990), .A4(n12989), .ZN(
        n12993) );
  OR2_X1 U16490 ( .A1(n12994), .A2(n12993), .ZN(n13665) );
  XNOR2_X1 U16491 ( .A(n13666), .B(n13665), .ZN(n12996) );
  AOI22_X1 U16492 ( .A1(n13787), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n12586), .ZN(n12995) );
  OAI21_X1 U16493 ( .B1(n12996), .B2(n13709), .A(n12995), .ZN(n13001) );
  INV_X1 U16494 ( .A(n12997), .ZN(n12998) );
  INV_X1 U16495 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16496 ( .A1(n9702), .A2(n12999), .ZN(n13000) );
  NAND2_X1 U16497 ( .A1(n13686), .A2(n13000), .ZN(n14770) );
  MUX2_X1 U16498 ( .A(n13001), .B(n14770), .S(n13683), .Z(n13003) );
  INV_X1 U16499 ( .A(n13002), .ZN(n13005) );
  INV_X1 U16500 ( .A(n13003), .ZN(n13004) );
  NAND3_X1 U16501 ( .A1(n10287), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17434) );
  INV_X1 U16502 ( .A(n17434), .ZN(n13008) );
  NAND2_X1 U16503 ( .A1(n21302), .A2(n13009), .ZN(n21403) );
  NAND2_X1 U16504 ( .A1(n21403), .A2(n10287), .ZN(n13010) );
  NAND2_X1 U16505 ( .A1(n10287), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17347) );
  NAND2_X1 U16506 ( .A1(n21397), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13011) );
  NAND2_X1 U16507 ( .A1(n17347), .A2(n13011), .ZN(n14110) );
  INV_X1 U16508 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n13880) );
  NOR2_X1 U16509 ( .A1(n20716), .A2(n13880), .ZN(n15405) );
  AOI21_X1 U16510 ( .B1(n17370), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15405), .ZN(n13012) );
  OAI21_X1 U16511 ( .B1(n14770), .B2(n17377), .A(n13012), .ZN(n13013) );
  OAI21_X1 U16512 ( .B1(n15412), .B2(n20646), .A(n13014), .ZN(P1_U2971) );
  NAND2_X1 U16513 ( .A1(n20015), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13015) );
  NAND2_X1 U16514 ( .A1(n20078), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19977) );
  NAND2_X1 U16515 ( .A1(n19977), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13017) );
  NAND2_X1 U16516 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20618), .ZN(
        n20145) );
  INV_X1 U16517 ( .A(n20145), .ZN(n13016) );
  NAND2_X1 U16518 ( .A1(n20078), .A2(n13016), .ZN(n20228) );
  AOI21_X1 U16519 ( .B1(n13017), .B2(n20228), .A(n20614), .ZN(n20334) );
  AOI21_X1 U16520 ( .B1(n13034), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n20334), .ZN(n13018) );
  NAND2_X1 U16521 ( .A1(n13020), .A2(n13021), .ZN(n13023) );
  INV_X1 U16522 ( .A(n13021), .ZN(n13022) );
  NAND2_X1 U16523 ( .A1(n13039), .A2(n13022), .ZN(n16177) );
  NAND2_X1 U16524 ( .A1(n13024), .A2(n10020), .ZN(n13028) );
  INV_X1 U16525 ( .A(n20078), .ZN(n13031) );
  NAND2_X1 U16526 ( .A1(n13031), .A2(n16860), .ZN(n13025) );
  NAND2_X1 U16527 ( .A1(n19977), .A2(n13025), .ZN(n20110) );
  NOR2_X1 U16528 ( .A1(n20110), .A2(n20614), .ZN(n13026) );
  AOI21_X1 U16529 ( .B1(n13034), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13026), .ZN(n13027) );
  NAND2_X1 U16530 ( .A1(n20627), .A2(n20335), .ZN(n20113) );
  NAND2_X1 U16531 ( .A1(n20113), .A2(n13031), .ZN(n20111) );
  NOR2_X1 U16532 ( .A1(n20111), .A2(n20614), .ZN(n16777) );
  AOI21_X1 U16533 ( .B1(n13034), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n16777), .ZN(n13032) );
  AOI22_X1 U16534 ( .A1(n13034), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20266), .B2(n20627), .ZN(n13035) );
  INV_X1 U16535 ( .A(n13036), .ZN(n13037) );
  NAND2_X1 U16536 ( .A1(n14236), .A2(n14235), .ZN(n14237) );
  NAND2_X1 U16537 ( .A1(n20015), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13038) );
  NAND2_X1 U16538 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14415) );
  INV_X1 U16539 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14593) );
  NOR2_X1 U16540 ( .A1(n14415), .A2(n14593), .ZN(n13040) );
  NAND4_X1 U16541 ( .A1(n16062), .A2(n19854), .A3(n16058), .A4(n13040), .ZN(
        n13042) );
  NAND2_X1 U16542 ( .A1(n14600), .A2(n14595), .ZN(n13041) );
  NOR2_X1 U16543 ( .A1(n13042), .A2(n13041), .ZN(n14605) );
  AOI22_X1 U16544 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U16545 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U16546 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13044) );
  AOI22_X1 U16547 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13043) );
  NAND4_X1 U16548 ( .A1(n13046), .A2(n13045), .A3(n13044), .A4(n13043), .ZN(
        n13052) );
  AOI22_X1 U16549 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16550 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U16551 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U16552 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13047) );
  NAND4_X1 U16553 ( .A1(n13050), .A2(n13049), .A3(n13048), .A4(n13047), .ZN(
        n13051) );
  OR2_X1 U16554 ( .A1(n13052), .A2(n13051), .ZN(n19846) );
  NAND3_X1 U16555 ( .A1(n14616), .A2(n19846), .A3(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U16556 ( .A1(n19847), .A2(n14620), .ZN(n13053) );
  NOR2_X1 U16557 ( .A1(n13054), .A2(n13053), .ZN(n13055) );
  AND3_X1 U16558 ( .A1(n14369), .A2(n14605), .A3(n13055), .ZN(n13056) );
  AOI22_X1 U16559 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U16560 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U16561 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U16562 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13057) );
  NAND4_X1 U16563 ( .A1(n13060), .A2(n13059), .A3(n13058), .A4(n13057), .ZN(
        n13066) );
  AOI22_X1 U16564 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16565 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U16566 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U16567 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13061) );
  NAND4_X1 U16568 ( .A1(n13064), .A2(n13063), .A3(n13062), .A4(n13061), .ZN(
        n13065) );
  OR2_X1 U16569 ( .A1(n13066), .A2(n13065), .ZN(n16030) );
  AOI22_X1 U16570 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10947), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U16571 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U16572 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U16573 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13067) );
  NAND4_X1 U16574 ( .A1(n13070), .A2(n13069), .A3(n13068), .A4(n13067), .ZN(
        n13076) );
  AOI22_X1 U16575 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13074) );
  AOI22_X1 U16576 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U16577 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U16578 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10882), .B1(
        n10931), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13071) );
  NAND4_X1 U16579 ( .A1(n13074), .A2(n13073), .A3(n13072), .A4(n13071), .ZN(
        n13075) );
  OR2_X1 U16580 ( .A1(n13076), .A2(n13075), .ZN(n16029) );
  AOI22_X1 U16581 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U16582 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13079) );
  AOI22_X1 U16583 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13078) );
  AOI22_X1 U16584 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13077) );
  NAND4_X1 U16585 ( .A1(n13080), .A2(n13079), .A3(n13078), .A4(n13077), .ZN(
        n13086) );
  AOI22_X1 U16586 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U16587 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U16588 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13082) );
  AOI22_X1 U16589 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13081) );
  NAND4_X1 U16590 ( .A1(n13084), .A2(n13083), .A3(n13082), .A4(n13081), .ZN(
        n13085) );
  OR2_X1 U16591 ( .A1(n13086), .A2(n13085), .ZN(n16042) );
  AOI22_X1 U16592 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16593 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U16594 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U16595 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13087) );
  NAND4_X1 U16596 ( .A1(n13090), .A2(n13089), .A3(n13088), .A4(n13087), .ZN(
        n13096) );
  AOI22_X1 U16597 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16598 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16599 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16600 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13091) );
  NAND4_X1 U16601 ( .A1(n13094), .A2(n13093), .A3(n13092), .A4(n13091), .ZN(
        n13095) );
  OR2_X1 U16602 ( .A1(n13096), .A2(n13095), .ZN(n16033) );
  AOI22_X1 U16603 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16604 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13099) );
  AOI22_X1 U16605 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U16606 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13097) );
  NAND4_X1 U16607 ( .A1(n13100), .A2(n13099), .A3(n13098), .A4(n13097), .ZN(
        n13106) );
  AOI22_X1 U16608 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U16609 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U16610 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13102) );
  AOI22_X1 U16611 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13101) );
  NAND4_X1 U16612 ( .A1(n13104), .A2(n13103), .A3(n13102), .A4(n13101), .ZN(
        n13105) );
  INV_X1 U16613 ( .A(n16024), .ZN(n13118) );
  AOI22_X1 U16614 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10948), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13110) );
  AOI22_X1 U16615 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U16616 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13108) );
  AOI22_X1 U16617 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13107) );
  NAND4_X1 U16618 ( .A1(n13110), .A2(n13109), .A3(n13108), .A4(n13107), .ZN(
        n13116) );
  AOI22_X1 U16619 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16620 ( .A1(n10873), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13113) );
  AOI22_X1 U16621 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13112) );
  AOI22_X1 U16622 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10931), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13111) );
  NAND4_X1 U16623 ( .A1(n13114), .A2(n13113), .A3(n13112), .A4(n13111), .ZN(
        n13115) );
  NOR2_X1 U16624 ( .A1(n13116), .A2(n13115), .ZN(n16022) );
  INV_X1 U16625 ( .A(n16022), .ZN(n13117) );
  AOI22_X1 U16626 ( .A1(n10947), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10873), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16627 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10852), .B1(
        n10832), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13123) );
  AOI22_X1 U16628 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13120), .B1(
        n13119), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16629 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10833), .B1(
        n10834), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13121) );
  NAND4_X1 U16630 ( .A1(n13124), .A2(n13123), .A3(n13122), .A4(n13121), .ZN(
        n13131) );
  AOI22_X1 U16631 ( .A1(n10846), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10881), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U16632 ( .A1(n10948), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16633 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10908), .B1(
        n10839), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13127) );
  AOI22_X1 U16634 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10931), .B1(
        n10847), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13126) );
  NAND4_X1 U16635 ( .A1(n13129), .A2(n13128), .A3(n13127), .A4(n13126), .ZN(
        n13130) );
  NOR2_X1 U16636 ( .A1(n13131), .A2(n13130), .ZN(n13159) );
  AOI22_X1 U16637 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13144) );
  AOI22_X1 U16638 ( .A1(n13326), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13143) );
  INV_X1 U16639 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13136) );
  AND2_X1 U16640 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13134) );
  OR2_X1 U16641 ( .A1(n13134), .A2(n13133), .ZN(n13295) );
  INV_X1 U16642 ( .A(n13295), .ZN(n13332) );
  INV_X1 U16643 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13135) );
  OAI211_X1 U16644 ( .C1(n13322), .C2(n13136), .A(n13332), .B(n9768), .ZN(
        n13137) );
  INV_X1 U16645 ( .A(n13137), .ZN(n13142) );
  INV_X1 U16646 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16838) );
  INV_X1 U16647 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16824) );
  OAI22_X1 U16648 ( .A1(n16755), .A2(n16838), .B1(n13331), .B2(n16824), .ZN(
        n13140) );
  INV_X1 U16649 ( .A(n13140), .ZN(n13141) );
  NAND4_X1 U16650 ( .A1(n13144), .A2(n13143), .A3(n13142), .A4(n13141), .ZN(
        n13156) );
  INV_X1 U16651 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13147) );
  INV_X1 U16652 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13146) );
  OAI22_X1 U16653 ( .A1(n13322), .A2(n13147), .B1(n13306), .B2(n13146), .ZN(
        n13148) );
  INV_X1 U16654 ( .A(n13148), .ZN(n13154) );
  AOI22_X1 U16655 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13153) );
  AOI22_X1 U16656 ( .A1(n13335), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13338), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13152) );
  INV_X1 U16657 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16796) );
  INV_X1 U16658 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13149) );
  OAI211_X1 U16659 ( .C1(n16796), .C2(n13331), .A(n9769), .B(n13295), .ZN(
        n13150) );
  INV_X1 U16660 ( .A(n13150), .ZN(n13151) );
  NAND4_X1 U16661 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n13151), .ZN(
        n13155) );
  NAND2_X1 U16662 ( .A1(n13156), .A2(n13155), .ZN(n13184) );
  NOR2_X1 U16663 ( .A1(n13987), .A2(n13184), .ZN(n13157) );
  XOR2_X1 U16664 ( .A(n13159), .B(n13157), .Z(n13185) );
  INV_X1 U16665 ( .A(n13184), .ZN(n13160) );
  NAND2_X1 U16666 ( .A1(n13987), .A2(n13160), .ZN(n16015) );
  INV_X1 U16667 ( .A(n13185), .ZN(n13158) );
  INV_X1 U16668 ( .A(n13159), .ZN(n13161) );
  NAND2_X1 U16669 ( .A1(n13161), .A2(n13160), .ZN(n13188) );
  AOI22_X1 U16670 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13279), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13170) );
  AOI22_X1 U16671 ( .A1(n13338), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13169) );
  INV_X1 U16672 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13162) );
  OAI22_X1 U16673 ( .A1(n13322), .A2(n21485), .B1(n13331), .B2(n13162), .ZN(
        n13163) );
  INV_X1 U16674 ( .A(n13163), .ZN(n13168) );
  INV_X1 U16675 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13165) );
  OAI211_X1 U16676 ( .C1(n13306), .C2(n13165), .A(n13295), .B(n9741), .ZN(
        n13166) );
  INV_X1 U16677 ( .A(n13166), .ZN(n13167) );
  NAND4_X1 U16678 ( .A1(n13170), .A2(n13169), .A3(n13168), .A4(n13167), .ZN(
        n13181) );
  AOI22_X1 U16679 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13179) );
  INV_X1 U16680 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13171) );
  OAI211_X1 U16681 ( .C1(n13306), .C2(n10811), .A(n13332), .B(n9742), .ZN(
        n13172) );
  INV_X1 U16682 ( .A(n13172), .ZN(n13178) );
  AOI22_X1 U16683 ( .A1(n13338), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13177) );
  INV_X1 U16684 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13174) );
  INV_X1 U16685 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13173) );
  OAI22_X1 U16686 ( .A1(n13322), .A2(n13174), .B1(n13331), .B2(n13173), .ZN(
        n13175) );
  INV_X1 U16687 ( .A(n13175), .ZN(n13176) );
  NAND4_X1 U16688 ( .A1(n13179), .A2(n13178), .A3(n13177), .A4(n13176), .ZN(
        n13180) );
  NAND2_X1 U16689 ( .A1(n13181), .A2(n13180), .ZN(n13187) );
  XOR2_X1 U16690 ( .A(n13188), .B(n13187), .Z(n13182) );
  NAND2_X1 U16691 ( .A1(n13182), .A2(n14369), .ZN(n16009) );
  INV_X1 U16692 ( .A(n13187), .ZN(n13183) );
  NAND2_X1 U16693 ( .A1(n13987), .A2(n13183), .ZN(n16011) );
  NOR3_X1 U16694 ( .A1(n13185), .A2(n13184), .A3(n16011), .ZN(n13186) );
  INV_X1 U16695 ( .A(n13236), .ZN(n13211) );
  NOR2_X1 U16696 ( .A1(n13188), .A2(n13187), .ZN(n13210) );
  AOI22_X1 U16697 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13198) );
  INV_X1 U16698 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13190) );
  OAI211_X1 U16699 ( .C1(n13322), .C2(n13190), .A(n13332), .B(n9743), .ZN(
        n13191) );
  INV_X1 U16700 ( .A(n13191), .ZN(n13197) );
  AOI22_X1 U16701 ( .A1(n13338), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13196) );
  INV_X1 U16702 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13193) );
  INV_X1 U16703 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13192) );
  OAI22_X1 U16704 ( .A1(n13306), .A2(n13193), .B1(n13331), .B2(n13192), .ZN(
        n13194) );
  INV_X1 U16705 ( .A(n13194), .ZN(n13195) );
  NAND4_X1 U16706 ( .A1(n13198), .A2(n13197), .A3(n13196), .A4(n13195), .ZN(
        n13209) );
  AOI22_X1 U16707 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U16708 ( .A1(n13335), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13338), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13206) );
  OAI211_X1 U16709 ( .C1(n13306), .C2(n13199), .A(n13295), .B(n9744), .ZN(
        n13200) );
  INV_X1 U16710 ( .A(n13200), .ZN(n13205) );
  INV_X1 U16711 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13201) );
  OAI22_X1 U16712 ( .A1(n13322), .A2(n13202), .B1(n13331), .B2(n13201), .ZN(
        n13203) );
  INV_X1 U16713 ( .A(n13203), .ZN(n13204) );
  NAND4_X1 U16714 ( .A1(n13207), .A2(n13206), .A3(n13205), .A4(n13204), .ZN(
        n13208) );
  NAND2_X1 U16715 ( .A1(n13210), .A2(n13233), .ZN(n13237) );
  OAI211_X1 U16716 ( .C1(n13210), .C2(n13233), .A(n14369), .B(n13237), .ZN(
        n13235) );
  XNOR2_X2 U16717 ( .A(n13211), .B(n13235), .ZN(n16005) );
  AOI22_X1 U16718 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13220) );
  AOI22_X1 U16719 ( .A1(n13338), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13219) );
  INV_X1 U16720 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13213) );
  INV_X1 U16721 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13212) );
  OAI22_X1 U16722 ( .A1(n13322), .A2(n13213), .B1(n13331), .B2(n13212), .ZN(
        n13214) );
  INV_X1 U16723 ( .A(n13214), .ZN(n13218) );
  INV_X1 U16724 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13215) );
  OAI211_X1 U16725 ( .C1(n13306), .C2(n13215), .A(n13295), .B(n9745), .ZN(
        n13216) );
  INV_X1 U16726 ( .A(n13216), .ZN(n13217) );
  NAND4_X1 U16727 ( .A1(n13220), .A2(n13219), .A3(n13218), .A4(n13217), .ZN(
        n13232) );
  AOI22_X1 U16728 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13230) );
  OAI211_X1 U16729 ( .C1(n13306), .C2(n13222), .A(n13332), .B(n9776), .ZN(
        n13223) );
  INV_X1 U16730 ( .A(n13223), .ZN(n13229) );
  AOI22_X1 U16731 ( .A1(n13338), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13228) );
  INV_X1 U16732 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13225) );
  INV_X1 U16733 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13224) );
  OAI22_X1 U16734 ( .A1(n13322), .A2(n13225), .B1(n13331), .B2(n13224), .ZN(
        n13226) );
  INV_X1 U16735 ( .A(n13226), .ZN(n13227) );
  NAND4_X1 U16736 ( .A1(n13230), .A2(n13229), .A3(n13228), .A4(n13227), .ZN(
        n13231) );
  AND2_X1 U16737 ( .A1(n13232), .A2(n13231), .ZN(n13239) );
  INV_X1 U16738 ( .A(n13233), .ZN(n13234) );
  NOR2_X1 U16739 ( .A1(n11232), .A2(n13234), .ZN(n16004) );
  NAND3_X1 U16740 ( .A1(n16005), .A2(n13239), .A3(n16004), .ZN(n13240) );
  OR2_X1 U16741 ( .A1(n13236), .A2(n13235), .ZN(n15995) );
  INV_X1 U16742 ( .A(n13237), .ZN(n13238) );
  INV_X1 U16743 ( .A(n13239), .ZN(n15996) );
  OR2_X1 U16744 ( .A1(n13237), .A2(n15996), .ZN(n13264) );
  OAI211_X1 U16745 ( .C1(n13239), .C2(n13238), .A(n13264), .B(n14369), .ZN(
        n15998) );
  AOI22_X1 U16746 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U16747 ( .A1(n13338), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13249) );
  INV_X1 U16748 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13242) );
  INV_X1 U16749 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13241) );
  OAI22_X1 U16750 ( .A1(n13322), .A2(n13242), .B1(n13331), .B2(n13241), .ZN(
        n13243) );
  INV_X1 U16751 ( .A(n13243), .ZN(n13248) );
  INV_X1 U16752 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13245) );
  OAI211_X1 U16753 ( .C1(n13306), .C2(n13245), .A(n13295), .B(n9777), .ZN(
        n13246) );
  INV_X1 U16754 ( .A(n13246), .ZN(n13247) );
  NAND4_X1 U16755 ( .A1(n13250), .A2(n13249), .A3(n13248), .A4(n13247), .ZN(
        n13262) );
  AOI22_X1 U16756 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13260) );
  INV_X1 U16757 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13252) );
  OAI211_X1 U16758 ( .C1(n13306), .C2(n13252), .A(n13332), .B(n9778), .ZN(
        n13253) );
  INV_X1 U16759 ( .A(n13253), .ZN(n13259) );
  AOI22_X1 U16760 ( .A1(n13338), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13258) );
  INV_X1 U16761 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13255) );
  INV_X1 U16762 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13254) );
  OAI22_X1 U16763 ( .A1(n13322), .A2(n13255), .B1(n13331), .B2(n13254), .ZN(
        n13256) );
  INV_X1 U16764 ( .A(n13256), .ZN(n13257) );
  NAND4_X1 U16765 ( .A1(n13260), .A2(n13259), .A3(n13258), .A4(n13257), .ZN(
        n13261) );
  NAND2_X1 U16766 ( .A1(n13262), .A2(n13261), .ZN(n13267) );
  NOR2_X1 U16767 ( .A1(n13264), .A2(n13267), .ZN(n13293) );
  AOI211_X1 U16768 ( .C1(n13267), .C2(n13264), .A(n13263), .B(n13293), .ZN(
        n13265) );
  INV_X1 U16769 ( .A(n13267), .ZN(n13268) );
  NAND2_X1 U16770 ( .A1(n13987), .A2(n13268), .ZN(n15990) );
  INV_X1 U16771 ( .A(n13269), .ZN(n13292) );
  AOI22_X1 U16772 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U16773 ( .A1(n13338), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13277) );
  INV_X1 U16774 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13271) );
  INV_X1 U16775 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13270) );
  OAI22_X1 U16776 ( .A1(n13322), .A2(n13271), .B1(n13331), .B2(n13270), .ZN(
        n13272) );
  INV_X1 U16777 ( .A(n13272), .ZN(n13276) );
  INV_X1 U16778 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13273) );
  OAI211_X1 U16779 ( .C1(n13306), .C2(n13273), .A(n13295), .B(n9779), .ZN(
        n13274) );
  INV_X1 U16780 ( .A(n13274), .ZN(n13275) );
  NAND4_X1 U16781 ( .A1(n13278), .A2(n13277), .A3(n13276), .A4(n13275), .ZN(
        n13291) );
  AOI22_X1 U16782 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13289) );
  OAI211_X1 U16783 ( .C1(n13306), .C2(n13281), .A(n13332), .B(n9780), .ZN(
        n13282) );
  INV_X1 U16784 ( .A(n13282), .ZN(n13288) );
  AOI22_X1 U16785 ( .A1(n13338), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13287) );
  INV_X1 U16786 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13284) );
  INV_X1 U16787 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13283) );
  OAI22_X1 U16788 ( .A1(n13322), .A2(n13284), .B1(n13331), .B2(n13283), .ZN(
        n13285) );
  INV_X1 U16789 ( .A(n13285), .ZN(n13286) );
  NAND4_X1 U16790 ( .A1(n13289), .A2(n13288), .A3(n13287), .A4(n13286), .ZN(
        n13290) );
  INV_X1 U16791 ( .A(n13293), .ZN(n15985) );
  NAND2_X1 U16792 ( .A1(n11232), .A2(n15986), .ZN(n13294) );
  NOR2_X1 U16793 ( .A1(n15985), .A2(n13294), .ZN(n13318) );
  INV_X1 U16794 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13296) );
  OAI211_X1 U16795 ( .C1(n13322), .C2(n13296), .A(n13295), .B(n9781), .ZN(
        n13300) );
  INV_X1 U16796 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13298) );
  INV_X1 U16797 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13297) );
  OAI22_X1 U16798 ( .A1(n16755), .A2(n13298), .B1(n13331), .B2(n13297), .ZN(
        n13299) );
  NOR2_X1 U16799 ( .A1(n13300), .A2(n13299), .ZN(n13303) );
  AOI22_X1 U16800 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U16801 ( .A1(n13326), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13301) );
  NAND3_X1 U16802 ( .A1(n13303), .A2(n13302), .A3(n13301), .ZN(n13316) );
  OAI211_X1 U16803 ( .C1(n13306), .C2(n13305), .A(n13332), .B(n9782), .ZN(
        n13307) );
  INV_X1 U16804 ( .A(n13307), .ZN(n13314) );
  AOI22_X1 U16805 ( .A1(n13335), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13338), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U16806 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13312) );
  INV_X1 U16807 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13309) );
  INV_X1 U16808 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13308) );
  OAI22_X1 U16809 ( .A1(n13322), .A2(n13309), .B1(n13331), .B2(n13308), .ZN(
        n13310) );
  INV_X1 U16810 ( .A(n13310), .ZN(n13311) );
  NAND4_X1 U16811 ( .A1(n13314), .A2(n13313), .A3(n13312), .A4(n13311), .ZN(
        n13315) );
  AND2_X1 U16812 ( .A1(n13316), .A2(n13315), .ZN(n13317) );
  NAND2_X1 U16813 ( .A1(n13318), .A2(n13317), .ZN(n13319) );
  OAI21_X1 U16814 ( .B1(n13318), .B2(n13317), .A(n13319), .ZN(n15981) );
  INV_X1 U16815 ( .A(n13319), .ZN(n13320) );
  NOR2_X1 U16816 ( .A1(n15980), .A2(n13320), .ZN(n13347) );
  INV_X1 U16817 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13321) );
  OAI22_X1 U16818 ( .A1(n13322), .A2(n21492), .B1(n16755), .B2(n13321), .ZN(
        n13325) );
  INV_X1 U16819 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13323) );
  AOI211_X1 U16820 ( .C1(n13326), .C2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n13325), .B(n13324), .ZN(n13330) );
  AOI22_X1 U16821 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U16822 ( .A1(n13335), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13327), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13328) );
  NAND3_X1 U16823 ( .A1(n13330), .A2(n13329), .A3(n13328), .ZN(n13345) );
  INV_X1 U16824 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n20076) );
  NOR2_X1 U16825 ( .A1(n13331), .A2(n20076), .ZN(n13333) );
  AOI211_X1 U16826 ( .C1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .C2(n13334), .A(
        n13333), .B(n13332), .ZN(n13343) );
  AOI22_X1 U16827 ( .A1(n13279), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13335), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U16828 ( .A1(n13337), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13336), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U16829 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13338), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13340) );
  NAND4_X1 U16830 ( .A1(n13343), .A2(n13342), .A3(n13341), .A4(n13340), .ZN(
        n13344) );
  NAND2_X1 U16831 ( .A1(n13345), .A2(n13344), .ZN(n13346) );
  XNOR2_X1 U16832 ( .A(n13347), .B(n13346), .ZN(n15979) );
  INV_X1 U16833 ( .A(n15979), .ZN(n13354) );
  INV_X1 U16834 ( .A(n13348), .ZN(n13349) );
  NAND2_X1 U16835 ( .A1(n13354), .A2(n19903), .ZN(n13379) );
  INV_X1 U16836 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n13357) );
  NAND2_X1 U16837 ( .A1(n12524), .A2(P2_EAX_REG_30__SCAN_IN), .ZN(n13356) );
  NAND2_X1 U16838 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13355) );
  OAI211_X1 U16839 ( .C1(n14727), .C2(n13357), .A(n13356), .B(n13355), .ZN(
        n13358) );
  NAND2_X1 U16840 ( .A1(n20022), .A2(n20015), .ZN(n13362) );
  NOR4_X1 U16841 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13366) );
  NOR4_X1 U16842 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13365) );
  NOR4_X1 U16843 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13364) );
  NOR4_X1 U16844 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13363) );
  AND4_X1 U16845 ( .A1(n13366), .A2(n13365), .A3(n13364), .A4(n13363), .ZN(
        n13371) );
  NOR4_X1 U16846 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13369) );
  NOR4_X1 U16847 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13368) );
  NOR4_X1 U16848 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n13367) );
  AND4_X1 U16849 ( .A1(n13369), .A2(n13368), .A3(n13367), .A4(n20544), .ZN(
        n13370) );
  NAND2_X1 U16850 ( .A1(n13371), .A2(n13370), .ZN(n13372) );
  NAND2_X1 U16851 ( .A1(n19869), .A2(BUF1_REG_30__SCAN_IN), .ZN(n13377) );
  NAND2_X1 U16852 ( .A1(n13390), .A2(n20022), .ZN(n13373) );
  INV_X1 U16853 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n13375) );
  NAND2_X1 U16854 ( .A1(n16790), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13374) );
  OAI21_X1 U16855 ( .B1(n16790), .B2(n13375), .A(n13374), .ZN(n14588) );
  AOI22_X1 U16856 ( .A1(n19868), .A2(n14588), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19898), .ZN(n13376) );
  NAND2_X1 U16857 ( .A1(n13377), .A2(n13376), .ZN(n13378) );
  NOR2_X2 U16858 ( .A1(n14269), .A2(n16790), .ZN(n19870) );
  NAND3_X1 U16859 ( .A1(n13379), .A2(n10607), .A3(n10594), .ZN(P2_U2889) );
  AND2_X1 U16860 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13399) );
  XNOR2_X1 U16861 ( .A(n13382), .B(n13381), .ZN(n16196) );
  OAI211_X1 U16862 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n16196), .B(n11076), .ZN(
        n13383) );
  OAI21_X1 U16863 ( .B1(n13386), .B2(n13768), .A(n13730), .ZN(n13718) );
  INV_X1 U16864 ( .A(n13386), .ZN(n13387) );
  NAND3_X1 U16865 ( .A1(n13387), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11076), .ZN(n13760) );
  NAND2_X1 U16866 ( .A1(n13763), .A2(n13760), .ZN(n13395) );
  NAND2_X1 U16867 ( .A1(n13389), .A2(n13388), .ZN(n13764) );
  NAND2_X1 U16868 ( .A1(n13390), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13391) );
  XNOR2_X1 U16869 ( .A(n13764), .B(n13391), .ZN(n13392) );
  AOI21_X1 U16870 ( .B1(n13392), .B2(n11076), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13762) );
  INV_X1 U16871 ( .A(n13762), .ZN(n13393) );
  INV_X1 U16872 ( .A(n13392), .ZN(n13750) );
  NAND2_X1 U16873 ( .A1(n13393), .A2(n13761), .ZN(n13394) );
  NAND2_X1 U16874 ( .A1(n13733), .A2(n17444), .ZN(n13404) );
  INV_X1 U16875 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n13398) );
  NAND2_X1 U16876 ( .A1(n13778), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13397) );
  AOI22_X1 U16877 ( .A1(n13774), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n13396) );
  OAI211_X1 U16878 ( .C1(n13398), .C2(n13776), .A(n13397), .B(n13396), .ZN(
        n13772) );
  XNOR2_X1 U16879 ( .A(n13773), .B(n13772), .ZN(n15976) );
  NAND2_X1 U16880 ( .A1(n16423), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13736) );
  AND2_X1 U16881 ( .A1(n13399), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14734) );
  AND2_X1 U16882 ( .A1(n16463), .A2(n14734), .ZN(n13400) );
  OAI211_X1 U16883 ( .C1(n19970), .C2(n14734), .A(n13721), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14732) );
  OAI21_X1 U16884 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13400), .A(
        n14732), .ZN(n13401) );
  OAI211_X1 U16885 ( .C1(n15976), .C2(n19964), .A(n13736), .B(n13401), .ZN(
        n13402) );
  INV_X1 U16886 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13408) );
  NAND2_X1 U16887 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13407) );
  NAND2_X1 U16888 ( .A1(n11604), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13406) );
  OAI211_X1 U16889 ( .C1(n18251), .C2(n13408), .A(n13407), .B(n13406), .ZN(
        n13409) );
  INV_X1 U16890 ( .A(n13409), .ZN(n13413) );
  AOI22_X1 U16891 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U16892 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U16893 ( .A1(n11549), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13410) );
  NAND4_X1 U16894 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n13410), .ZN(
        n13419) );
  AOI22_X1 U16895 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11524), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U16896 ( .A1(n13511), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U16897 ( .A1(n13513), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13512), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U16898 ( .A1(n11607), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13514), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13414) );
  NAND4_X1 U16899 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13418) );
  INV_X1 U16900 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13422) );
  NAND2_X1 U16901 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13421) );
  NAND2_X1 U16902 ( .A1(n11604), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13420) );
  OAI211_X1 U16903 ( .C1(n18251), .C2(n13422), .A(n13421), .B(n13420), .ZN(
        n13423) );
  INV_X1 U16904 ( .A(n13423), .ZN(n13427) );
  AOI22_X1 U16905 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U16906 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13425) );
  NAND2_X1 U16907 ( .A1(n11549), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13424) );
  AOI22_X1 U16908 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11524), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U16909 ( .A1(n13511), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U16910 ( .A1(n13513), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13512), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13429) );
  AOI22_X1 U16911 ( .A1(n11607), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13514), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13428) );
  NAND2_X1 U16912 ( .A1(n13607), .A2(n13609), .ZN(n13525) );
  INV_X1 U16913 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17182) );
  NAND2_X1 U16914 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n13433) );
  NAND2_X1 U16915 ( .A1(n18236), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n13432) );
  AOI22_X1 U16916 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13514), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U16917 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13437) );
  INV_X1 U16918 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13435) );
  OR2_X1 U16919 ( .A1(n18251), .A2(n13435), .ZN(n13436) );
  NAND4_X1 U16920 ( .A1(n9705), .A2(n13438), .A3(n13437), .A4(n13436), .ZN(
        n13444) );
  AOI22_X1 U16921 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13442) );
  AOI22_X1 U16922 ( .A1(n13511), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13441) );
  AOI22_X1 U16923 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13512), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U16924 ( .A1(n11524), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13439) );
  NAND4_X1 U16925 ( .A1(n13442), .A2(n13441), .A3(n13440), .A4(n13439), .ZN(
        n13443) );
  NOR2_X2 U16926 ( .A1(n13525), .A2(n18426), .ZN(n13536) );
  INV_X1 U16927 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13447) );
  NAND2_X1 U16928 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13446) );
  NAND2_X1 U16929 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13445) );
  OAI211_X1 U16930 ( .C1(n18251), .C2(n13447), .A(n13446), .B(n13445), .ZN(
        n13448) );
  INV_X1 U16931 ( .A(n13448), .ZN(n13452) );
  AOI22_X1 U16932 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13451) );
  AOI22_X1 U16933 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13450) );
  NAND2_X1 U16934 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13449) );
  NAND4_X1 U16935 ( .A1(n13452), .A2(n13451), .A3(n13450), .A4(n13449), .ZN(
        n13458) );
  AOI22_X1 U16936 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U16937 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U16938 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U16939 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13453) );
  NAND4_X1 U16940 ( .A1(n13456), .A2(n13455), .A3(n13454), .A4(n13453), .ZN(
        n13457) );
  AOI22_X1 U16941 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18192), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13462) );
  AOI22_X1 U16942 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13461) );
  AOI22_X1 U16943 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13460) );
  AOI22_X1 U16944 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13459) );
  AOI22_X1 U16945 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13467) );
  INV_X1 U16946 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13463) );
  NAND2_X1 U16947 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n13465) );
  NAND2_X1 U16948 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13464) );
  NAND4_X1 U16949 ( .A1(n13467), .A2(n13466), .A3(n13465), .A4(n13464), .ZN(
        n13472) );
  INV_X1 U16950 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13470) );
  NAND2_X1 U16951 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13469) );
  NAND2_X1 U16952 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n13468) );
  OAI211_X1 U16953 ( .C1(n18251), .C2(n13470), .A(n13469), .B(n13468), .ZN(
        n13471) );
  NOR2_X1 U16954 ( .A1(n13472), .A2(n13471), .ZN(n13473) );
  NOR2_X1 U16955 ( .A1(n18421), .A2(n18418), .ZN(n13475) );
  AOI22_X1 U16956 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13479) );
  AOI22_X1 U16957 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13478) );
  AOI22_X1 U16958 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13477) );
  AOI22_X1 U16959 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13476) );
  AOI22_X1 U16960 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13483) );
  NAND2_X1 U16961 ( .A1(n18243), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13481) );
  NAND2_X1 U16962 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13480) );
  NAND4_X1 U16963 ( .A1(n13483), .A2(n13482), .A3(n13481), .A4(n13480), .ZN(
        n13488) );
  INV_X1 U16964 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13486) );
  NAND2_X1 U16965 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13485) );
  NAND2_X1 U16966 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13484) );
  OAI211_X1 U16967 ( .C1(n18251), .C2(n13486), .A(n13485), .B(n13484), .ZN(
        n13487) );
  NOR2_X1 U16968 ( .A1(n13488), .A2(n13487), .ZN(n13489) );
  INV_X1 U16969 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18141) );
  NAND2_X1 U16970 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13491) );
  AOI22_X1 U16971 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13495) );
  AOI22_X1 U16972 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13494) );
  INV_X1 U16973 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13492) );
  OR2_X1 U16974 ( .A1(n18216), .A2(n13492), .ZN(n13493) );
  NAND4_X1 U16975 ( .A1(n9709), .A2(n13495), .A3(n13494), .A4(n13493), .ZN(
        n13501) );
  AOI22_X1 U16976 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13499) );
  AOI22_X1 U16977 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13498) );
  AOI22_X1 U16978 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U16979 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13496) );
  NAND4_X1 U16980 ( .A1(n13499), .A2(n13498), .A3(n13497), .A4(n13496), .ZN(
        n13500) );
  INV_X1 U16981 ( .A(n13599), .ZN(n18414) );
  XNOR2_X1 U16982 ( .A(n13609), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14214) );
  INV_X1 U16983 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13505) );
  NAND2_X1 U16984 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13504) );
  NAND2_X1 U16985 ( .A1(n11604), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13503) );
  OAI211_X1 U16986 ( .C1(n18251), .C2(n13505), .A(n13504), .B(n13503), .ZN(
        n13506) );
  INV_X1 U16987 ( .A(n13506), .ZN(n13510) );
  AOI22_X1 U16988 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13509) );
  AOI22_X1 U16989 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13508) );
  NAND2_X1 U16990 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13507) );
  NAND4_X1 U16991 ( .A1(n13510), .A2(n13509), .A3(n13508), .A4(n13507), .ZN(
        n13520) );
  AOI22_X1 U16992 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11524), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U16993 ( .A1(n13511), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U16994 ( .A1(n13513), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13512), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U16995 ( .A1(n11607), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13514), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13515) );
  NAND4_X1 U16996 ( .A1(n13518), .A2(n13517), .A3(n13516), .A4(n13515), .ZN(
        n13519) );
  AND2_X1 U16997 ( .A1(n14215), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14226) );
  NAND2_X1 U16998 ( .A1(n14214), .A2(n14226), .ZN(n14216) );
  INV_X1 U16999 ( .A(n13609), .ZN(n14206) );
  NAND2_X1 U17000 ( .A1(n14206), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13521) );
  NAND2_X1 U17001 ( .A1(n14216), .A2(n13521), .ZN(n18803) );
  XNOR2_X1 U17002 ( .A(n13522), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18804) );
  NAND2_X1 U17003 ( .A1(n18803), .A2(n18804), .ZN(n18802) );
  INV_X1 U17004 ( .A(n13522), .ZN(n13523) );
  NAND2_X1 U17005 ( .A1(n13523), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13524) );
  AND2_X1 U17006 ( .A1(n13525), .A2(n18426), .ZN(n13526) );
  NAND2_X1 U17007 ( .A1(n18788), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13531) );
  INV_X1 U17008 ( .A(n13527), .ZN(n13528) );
  NAND2_X1 U17009 ( .A1(n13529), .A2(n13528), .ZN(n13530) );
  NAND2_X1 U17010 ( .A1(n13531), .A2(n13530), .ZN(n18772) );
  XNOR2_X1 U17011 ( .A(n13536), .B(n13603), .ZN(n13532) );
  XNOR2_X1 U17012 ( .A(n13532), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18771) );
  NAND2_X1 U17013 ( .A1(n18772), .A2(n18771), .ZN(n18770) );
  INV_X1 U17014 ( .A(n13532), .ZN(n13533) );
  NAND2_X1 U17015 ( .A1(n13533), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13534) );
  NAND2_X2 U17016 ( .A1(n18770), .A2(n13534), .ZN(n13540) );
  INV_X1 U17017 ( .A(n18418), .ZN(n13535) );
  AOI21_X1 U17018 ( .B1(n13536), .B2(n13603), .A(n13535), .ZN(n13537) );
  OR2_X1 U17019 ( .A1(n13545), .A2(n13537), .ZN(n13538) );
  INV_X1 U17020 ( .A(n13538), .ZN(n13539) );
  XNOR2_X1 U17021 ( .A(n13545), .B(n13599), .ZN(n13542) );
  XNOR2_X1 U17022 ( .A(n13542), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18748) );
  INV_X1 U17023 ( .A(n13542), .ZN(n13543) );
  NAND2_X1 U17024 ( .A1(n13543), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13544) );
  AOI21_X1 U17025 ( .B1(n13545), .B2(n13599), .A(n17098), .ZN(n13546) );
  NAND2_X1 U17026 ( .A1(n13548), .A2(n10074), .ZN(n13549) );
  NOR2_X1 U17027 ( .A1(n19000), .A2(n18724), .ZN(n18976) );
  NAND2_X1 U17028 ( .A1(n18977), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16994) );
  NAND2_X1 U17029 ( .A1(n18939), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18927) );
  INV_X1 U17030 ( .A(n18927), .ZN(n18712) );
  NAND2_X1 U17031 ( .A1(n18712), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18917) );
  NAND2_X1 U17032 ( .A1(n19000), .A2(n18724), .ZN(n16991) );
  INV_X1 U17033 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17029) );
  INV_X1 U17034 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18969) );
  NAND4_X1 U17035 ( .A1(n17029), .A2(n18940), .A3(n18912), .A4(n18969), .ZN(
        n13552) );
  NAND2_X1 U17036 ( .A1(n13553), .A2(n10083), .ZN(n18669) );
  NAND2_X1 U17037 ( .A1(n18669), .A2(n17131), .ZN(n18617) );
  INV_X1 U17038 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18629) );
  NOR2_X1 U17039 ( .A1(n18895), .A2(n18629), .ZN(n18884) );
  NAND2_X1 U17040 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18884), .ZN(
        n18875) );
  NAND2_X1 U17041 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13554) );
  NOR2_X1 U17042 ( .A1(n18875), .A2(n13554), .ZN(n13555) );
  AND2_X1 U17043 ( .A1(n18614), .A2(n13555), .ZN(n18577) );
  NAND2_X1 U17044 ( .A1(n18669), .A2(n17121), .ZN(n13559) );
  NOR2_X1 U17045 ( .A1(n18694), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18649) );
  NAND2_X1 U17046 ( .A1(n18649), .A2(n18895), .ZN(n13556) );
  NOR2_X1 U17047 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13556), .ZN(
        n18618) );
  NOR3_X1 U17048 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13557) );
  NAND2_X1 U17049 ( .A1(n18618), .A2(n13557), .ZN(n13558) );
  NAND2_X1 U17050 ( .A1(n13559), .A2(n13558), .ZN(n13560) );
  INV_X1 U17051 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17124) );
  NAND2_X1 U17052 ( .A1(n13561), .A2(n18694), .ZN(n18560) );
  INV_X1 U17053 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13563) );
  INV_X1 U17054 ( .A(n13564), .ZN(n13565) );
  OR2_X1 U17055 ( .A1(n18694), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16955) );
  INV_X1 U17056 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17073) );
  NAND2_X1 U17057 ( .A1(n17073), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13636) );
  INV_X1 U17058 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17148) );
  NAND2_X1 U17059 ( .A1(n17148), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13642) );
  XNOR2_X1 U17060 ( .A(n18694), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13567) );
  INV_X1 U17061 ( .A(n13568), .ZN(n13573) );
  INV_X1 U17062 ( .A(n13569), .ZN(n13571) );
  NAND2_X1 U17063 ( .A1(n14453), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13570) );
  NAND2_X1 U17064 ( .A1(n13571), .A2(n13570), .ZN(n13586) );
  NAND3_X1 U17065 ( .A1(n13575), .A2(n13587), .A3(n13574), .ZN(n14141) );
  NAND2_X1 U17066 ( .A1(n19117), .A2(n13576), .ZN(n13584) );
  NOR2_X1 U17067 ( .A1(n13626), .A2(n9674), .ZN(n13596) );
  NAND2_X1 U17068 ( .A1(n13596), .A2(n13577), .ZN(n13580) );
  INV_X1 U17069 ( .A(n13578), .ZN(n13579) );
  AOI21_X1 U17070 ( .B1(n13580), .B2(n17546), .A(n13579), .ZN(n14391) );
  INV_X1 U17071 ( .A(n19708), .ZN(n14386) );
  AOI21_X1 U17072 ( .B1(n19709), .B2(n13582), .A(n14386), .ZN(n13581) );
  NAND2_X1 U17073 ( .A1(n19117), .A2(n18494), .ZN(n13589) );
  AOI21_X1 U17074 ( .B1(n13581), .B2(n13589), .A(n19705), .ZN(n17545) );
  OAI211_X1 U17075 ( .C1(n19131), .C2(n13582), .A(n14140), .B(n17545), .ZN(
        n13583) );
  OAI211_X1 U17076 ( .C1(n14141), .C2(n13584), .A(n14391), .B(n13583), .ZN(
        n13585) );
  INV_X1 U17077 ( .A(n13585), .ZN(n13592) );
  NOR2_X1 U17078 ( .A1(n13587), .A2(n13586), .ZN(n13588) );
  OR2_X1 U17079 ( .A1(n13589), .A2(n19135), .ZN(n13594) );
  INV_X1 U17080 ( .A(n13594), .ZN(n13590) );
  NAND2_X1 U17081 ( .A1(n16907), .A2(n13590), .ZN(n13591) );
  NAND2_X1 U17082 ( .A1(n13592), .A2(n13591), .ZN(n13593) );
  NOR2_X1 U17083 ( .A1(n13594), .A2(n14143), .ZN(n13595) );
  NAND2_X1 U17084 ( .A1(n16909), .A2(n18997), .ZN(n13650) );
  INV_X1 U17085 ( .A(n13607), .ZN(n14243) );
  NAND2_X1 U17086 ( .A1(n13608), .A2(n14243), .ZN(n13605) );
  NAND2_X1 U17087 ( .A1(n13604), .A2(n13603), .ZN(n13601) );
  NOR2_X1 U17088 ( .A1(n18418), .A2(n13601), .ZN(n13600) );
  NAND2_X1 U17089 ( .A1(n13600), .A2(n13599), .ZN(n13598) );
  NOR2_X1 U17090 ( .A1(n18411), .A2(n13598), .ZN(n13622) );
  XOR2_X1 U17091 ( .A(n13598), .B(n18411), .Z(n18738) );
  XOR2_X1 U17092 ( .A(n13600), .B(n13599), .Z(n13615) );
  XOR2_X1 U17093 ( .A(n13601), .B(n18418), .Z(n13602) );
  NAND2_X1 U17094 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13602), .ZN(
        n13614) );
  XOR2_X1 U17095 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n13602), .Z(
        n18759) );
  INV_X1 U17096 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19042) );
  XOR2_X1 U17097 ( .A(n13604), .B(n13603), .Z(n18777) );
  XNOR2_X1 U17098 ( .A(n13605), .B(n18426), .ZN(n13606) );
  NAND2_X1 U17099 ( .A1(n13606), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13613) );
  XOR2_X1 U17100 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13606), .Z(
        n18786) );
  INV_X1 U17101 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19089) );
  OR2_X1 U17102 ( .A1(n13611), .A2(n19089), .ZN(n13612) );
  AOI21_X1 U17103 ( .B1(n14206), .B2(n21541), .A(n13610), .ZN(n18801) );
  NAND2_X1 U17104 ( .A1(n18801), .A2(n18800), .ZN(n18799) );
  NAND2_X1 U17105 ( .A1(n13612), .A2(n18799), .ZN(n18785) );
  NAND2_X1 U17106 ( .A1(n18786), .A2(n18785), .ZN(n18784) );
  NAND2_X1 U17107 ( .A1(n13615), .A2(n13616), .ZN(n13617) );
  NOR2_X1 U17108 ( .A1(n18738), .A2(n18737), .ZN(n18736) );
  INV_X1 U17109 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13618) );
  NAND2_X1 U17110 ( .A1(n13622), .A2(n13619), .ZN(n13623) );
  NAND2_X1 U17111 ( .A1(n13622), .A2(n13621), .ZN(n13620) );
  NOR2_X1 U17112 ( .A1(n18845), .A2(n18854), .ZN(n18557) );
  AND2_X1 U17113 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16947) );
  AND2_X1 U17114 ( .A1(n16947), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17069) );
  NAND2_X1 U17115 ( .A1(n16959), .A2(n17069), .ZN(n17071) );
  OAI21_X1 U17116 ( .B1(n17071), .B2(n13642), .A(n13636), .ZN(n13624) );
  AOI21_X1 U17117 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17071), .A(
        n13624), .ZN(n16923) );
  NOR2_X2 U17118 ( .A1(n13625), .A2(n17153), .ZN(n18877) );
  NAND2_X1 U17119 ( .A1(n19135), .A2(n14143), .ZN(n14400) );
  NAND2_X1 U17120 ( .A1(n18494), .A2(n18432), .ZN(n17179) );
  NAND2_X1 U17121 ( .A1(n14145), .A2(n17179), .ZN(n19721) );
  NOR2_X2 U17122 ( .A1(n18914), .A2(n18916), .ZN(n18978) );
  NOR2_X1 U17123 ( .A1(n19709), .A2(n13627), .ZN(n13629) );
  INV_X1 U17124 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19041) );
  NAND3_X1 U17125 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19036) );
  NOR2_X1 U17126 ( .A1(n19041), .A2(n19036), .ZN(n19022) );
  AND2_X1 U17127 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n19022), .ZN(
        n19006) );
  NAND2_X1 U17128 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19006), .ZN(
        n13630) );
  NAND2_X1 U17129 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19003) );
  OR2_X1 U17130 ( .A1(n13630), .A2(n19003), .ZN(n18913) );
  NOR2_X1 U17131 ( .A1(n18668), .A2(n18913), .ZN(n18866) );
  NAND2_X1 U17132 ( .A1(n18877), .A2(n18991), .ZN(n19075) );
  AOI21_X1 U17133 ( .B1(n17096), .B2(n18866), .A(n17135), .ZN(n17115) );
  INV_X1 U17134 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18856) );
  NOR2_X1 U17135 ( .A1(n18856), .A2(n18854), .ZN(n17116) );
  AND2_X1 U17136 ( .A1(n17120), .A2(n17116), .ZN(n13631) );
  INV_X1 U17137 ( .A(n13631), .ZN(n17097) );
  OAI21_X1 U17138 ( .B1(n10220), .B2(n21541), .A(n19089), .ZN(n19002) );
  INV_X1 U17139 ( .A(n13630), .ZN(n17137) );
  NAND2_X1 U17140 ( .A1(n19002), .A2(n17137), .ZN(n18915) );
  NOR2_X1 U17141 ( .A1(n18668), .A2(n18915), .ZN(n13641) );
  NOR2_X1 U17142 ( .A1(n19546), .A2(n13641), .ZN(n18834) );
  INV_X1 U17143 ( .A(n18834), .ZN(n18870) );
  OAI21_X1 U17144 ( .B1(n17096), .B2(n19546), .A(n18870), .ZN(n18848) );
  AOI21_X1 U17145 ( .B1(n18916), .B2(n17097), .A(n18848), .ZN(n17119) );
  NOR2_X1 U17146 ( .A1(n18991), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19076) );
  INV_X1 U17147 ( .A(n19076), .ZN(n17130) );
  OAI211_X1 U17148 ( .C1(n17135), .C2(n13631), .A(n17119), .B(n17130), .ZN(
        n13632) );
  AOI211_X1 U17149 ( .C1(n18973), .C2(n18830), .A(n17115), .B(n13632), .ZN(
        n17083) );
  INV_X1 U17150 ( .A(n17069), .ZN(n16929) );
  AOI21_X1 U17151 ( .B1(n19005), .B2(n16929), .A(n19082), .ZN(n13634) );
  INV_X2 U17152 ( .A(n18992), .ZN(n18905) );
  AOI21_X1 U17153 ( .B1(n17083), .B2(n13634), .A(n18905), .ZN(n17078) );
  AND2_X1 U17154 ( .A1(n19005), .A2(n19062), .ZN(n19030) );
  INV_X1 U17155 ( .A(n19030), .ZN(n19055) );
  AND2_X1 U17156 ( .A1(n18905), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n16911) );
  INV_X1 U17157 ( .A(n16911), .ZN(n13635) );
  OAI21_X1 U17158 ( .B1(n19055), .B2(n13636), .A(n13635), .ZN(n13646) );
  INV_X1 U17159 ( .A(n17121), .ZN(n18571) );
  INV_X1 U17160 ( .A(n17120), .ZN(n13638) );
  NOR2_X1 U17161 ( .A1(n18550), .A2(n13638), .ZN(n16958) );
  INV_X1 U17162 ( .A(n16958), .ZN(n17117) );
  NOR2_X1 U17163 ( .A1(n17117), .A2(n16929), .ZN(n16926) );
  NAND2_X1 U17164 ( .A1(n16926), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13639) );
  XNOR2_X1 U17165 ( .A(n13639), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16920) );
  AOI21_X1 U17166 ( .B1(n18973), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18914), .ZN(n19074) );
  INV_X1 U17167 ( .A(n19074), .ZN(n13640) );
  AOI22_X1 U17168 ( .A1(n18916), .A2(n13641), .B1(n13640), .B2(n18866), .ZN(
        n17095) );
  NAND2_X1 U17169 ( .A1(n17096), .A2(n17116), .ZN(n18835) );
  NOR2_X1 U17170 ( .A1(n17095), .A2(n18835), .ZN(n18838) );
  NAND2_X1 U17171 ( .A1(n18838), .A2(n17120), .ZN(n17067) );
  NOR3_X1 U17172 ( .A1(n17067), .A2(n13642), .A3(n16929), .ZN(n13643) );
  AOI21_X1 U17173 ( .B1(n16920), .B2(n18971), .A(n13643), .ZN(n13644) );
  NOR2_X1 U17174 ( .A1(n13644), .A2(n19082), .ZN(n13645) );
  AOI211_X1 U17175 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17078), .A(
        n13646), .B(n13645), .ZN(n13647) );
  INV_X1 U17176 ( .A(n13648), .ZN(n13649) );
  NAND2_X1 U17177 ( .A1(n13650), .A2(n13649), .ZN(P3_U2831) );
  INV_X1 U17178 ( .A(n11958), .ZN(n14085) );
  INV_X1 U17179 ( .A(n13651), .ZN(n13654) );
  NOR2_X1 U17180 ( .A1(n14207), .A2(n20640), .ZN(n13653) );
  NAND4_X1 U17181 ( .A1(n14085), .A2(n13654), .A3(n13653), .A4(n13652), .ZN(
        n13835) );
  OR2_X1 U17182 ( .A1(n13835), .A2(n13947), .ZN(n13655) );
  OAI21_X1 U17183 ( .B1(n13657), .B2(n13659), .A(n13658), .ZN(n14764) );
  NAND2_X1 U17184 ( .A1(n13660), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n13661) );
  NAND2_X1 U17185 ( .A1(n13666), .A2(n13665), .ZN(n13688) );
  AOI22_X1 U17186 ( .A1(n12879), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13667), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13671) );
  AOI22_X1 U17187 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13670) );
  AOI22_X1 U17188 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13669) );
  AOI22_X1 U17189 ( .A1(n9585), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13668) );
  NAND4_X1 U17190 ( .A1(n13671), .A2(n13670), .A3(n13669), .A4(n13668), .ZN(
        n13678) );
  AOI22_X1 U17191 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13676) );
  AOI22_X1 U17192 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12931), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13675) );
  AOI22_X1 U17193 ( .A1(n9587), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12005), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U17194 ( .A1(n13672), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13673) );
  NAND4_X1 U17195 ( .A1(n13676), .A2(n13675), .A3(n13674), .A4(n13673), .ZN(
        n13677) );
  NOR2_X1 U17196 ( .A1(n13678), .A2(n13677), .ZN(n13689) );
  XOR2_X1 U17197 ( .A(n13688), .B(n13689), .Z(n13680) );
  NAND2_X1 U17198 ( .A1(n13680), .A2(n13679), .ZN(n13682) );
  AOI22_X1 U17199 ( .A1(n13787), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n12586), .ZN(n13681) );
  NAND2_X1 U17200 ( .A1(n13682), .A2(n13681), .ZN(n13684) );
  INV_X1 U17201 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14755) );
  XNOR2_X1 U17202 ( .A(n13686), .B(n14755), .ZN(n15185) );
  MUX2_X1 U17203 ( .A(n13684), .B(n15185), .S(n13683), .Z(n14748) );
  INV_X1 U17204 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13687) );
  XNOR2_X1 U17205 ( .A(n13791), .B(n13687), .ZN(n14686) );
  NOR2_X1 U17206 ( .A1(n13689), .A2(n13688), .ZN(n13707) );
  AOI22_X1 U17207 ( .A1(n11924), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12024), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U17208 ( .A1(n11925), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U17209 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13692), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13695) );
  AOI22_X1 U17210 ( .A1(n12005), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9590), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13694) );
  NAND4_X1 U17211 ( .A1(n13697), .A2(n13696), .A3(n13695), .A4(n13694), .ZN(
        n13705) );
  AOI22_X1 U17212 ( .A1(n13698), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U17213 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12685), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U17214 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12052), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U17215 ( .A1(n9582), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12118), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13700) );
  NAND4_X1 U17216 ( .A1(n13703), .A2(n13702), .A3(n13701), .A4(n13700), .ZN(
        n13704) );
  NOR2_X1 U17217 ( .A1(n13705), .A2(n13704), .ZN(n13706) );
  XOR2_X1 U17218 ( .A(n13707), .B(n13706), .Z(n13710) );
  AOI22_X1 U17219 ( .A1(n13787), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n12586), .ZN(n13708) );
  OAI21_X1 U17220 ( .B1(n13710), .B2(n13709), .A(n13708), .ZN(n13711) );
  INV_X1 U17221 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n13882) );
  NOR2_X1 U17222 ( .A1(n20716), .A2(n13882), .ZN(n15391) );
  NOR2_X1 U17223 ( .A1(n14686), .A2(n17377), .ZN(n13715) );
  AOI211_X1 U17224 ( .C1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n17370), .A(
        n15391), .B(n13715), .ZN(n13716) );
  OAI211_X1 U17225 ( .C1(n14689), .C2(n20811), .A(n13717), .B(n13716), .ZN(
        P1_U2969) );
  NOR2_X1 U17226 ( .A1(n16080), .A2(n19949), .ZN(n13729) );
  OAI21_X1 U17227 ( .B1(n13722), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13724) );
  INV_X1 U17228 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16462) );
  NAND2_X1 U17229 ( .A1(n13730), .A2(n16462), .ZN(n13723) );
  NAND3_X1 U17230 ( .A1(n16463), .A2(n13724), .A3(n13723), .ZN(n13725) );
  NAND2_X1 U17231 ( .A1(n16423), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16186) );
  NAND2_X1 U17232 ( .A1(n13725), .A2(n16186), .ZN(n13726) );
  AOI21_X1 U17233 ( .B1(n16465), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13726), .ZN(n13727) );
  OAI21_X1 U17234 ( .B1(n16184), .B2(n19964), .A(n13727), .ZN(n13728) );
  NAND3_X1 U17235 ( .A1(n9706), .A2(n13732), .A3(n13731), .ZN(P2_U3017) );
  NOR2_X1 U17236 ( .A1(n15976), .A2(n16455), .ZN(n13738) );
  XNOR2_X1 U17237 ( .A(n13734), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13743) );
  NAND2_X1 U17238 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13735) );
  OAI211_X1 U17239 ( .C1(n13743), .C2(n16441), .A(n13736), .B(n13735), .ZN(
        n13737) );
  NAND3_X1 U17240 ( .A1(n13741), .A2(n13740), .A3(n13739), .ZN(P2_U2984) );
  INV_X1 U17241 ( .A(n13743), .ZN(n13744) );
  AOI21_X1 U17242 ( .B1(n13745), .B2(n15968), .A(n13744), .ZN(n14722) );
  AOI21_X1 U17243 ( .B1(n17314), .B2(n13746), .A(n14722), .ZN(n13747) );
  INV_X1 U17244 ( .A(n13747), .ZN(n13757) );
  AOI22_X1 U17245 ( .A1(n19830), .A2(P2_EBX_REG_30__SCAN_IN), .B1(n19827), 
        .B2(P2_REIP_REG_30__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U17246 ( .A1(n19841), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13748) );
  OAI211_X1 U17247 ( .C1(n13750), .C2(n19809), .A(n13749), .B(n13748), .ZN(
        n13751) );
  INV_X1 U17248 ( .A(n13751), .ZN(n13752) );
  NAND3_X1 U17249 ( .A1(n13757), .A2(n13756), .A3(n13755), .ZN(P2_U2825) );
  INV_X1 U17250 ( .A(n13764), .ZN(n13765) );
  MUX2_X1 U17251 ( .A(n13767), .B(n13766), .S(n20006), .Z(n14720) );
  XNOR2_X1 U17252 ( .A(n13769), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13770) );
  NAND2_X1 U17253 ( .A1(n14740), .A2(n16435), .ZN(n13785) );
  AOI22_X1 U17254 ( .A1(n13774), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13775) );
  OAI21_X1 U17255 ( .B1(n13776), .B2(n14716), .A(n13775), .ZN(n13777) );
  AOI21_X1 U17256 ( .B1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13778), .A(
        n13777), .ZN(n13779) );
  NOR2_X1 U17257 ( .A1(n14738), .A2(n16455), .ZN(n13783) );
  NAND2_X1 U17258 ( .A1(n16423), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14736) );
  NAND2_X1 U17259 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13780) );
  OAI211_X1 U17260 ( .C1(n13781), .C2(n16441), .A(n14736), .B(n13780), .ZN(
        n13782) );
  OAI211_X1 U17261 ( .C1(n14743), .C2(n16446), .A(n13785), .B(n13784), .ZN(
        P2_U2983) );
  AOI22_X1 U17262 ( .A1(n13787), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13786), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13788) );
  INV_X1 U17263 ( .A(n13788), .ZN(n13789) );
  XNOR2_X2 U17264 ( .A(n13790), .B(n13789), .ZN(n13839) );
  NAND2_X1 U17265 ( .A1(n13792), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13793) );
  NAND2_X1 U17266 ( .A1(n13955), .A2(n13950), .ZN(n13943) );
  NAND2_X1 U17267 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n10287), .ZN(n13796) );
  NOR2_X1 U17268 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n17359) );
  NOR2_X1 U17269 ( .A1(n21197), .A2(n21399), .ZN(n17351) );
  INV_X1 U17270 ( .A(n17351), .ZN(n13795) );
  OAI22_X1 U17271 ( .A1(n13797), .A2(n13796), .B1(n10287), .B2(n13795), .ZN(
        n13798) );
  NAND2_X1 U17272 ( .A1(n13839), .A2(n9887), .ZN(n13821) );
  NAND2_X1 U17273 ( .A1(n14187), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13809) );
  AND2_X1 U17274 ( .A1(n21404), .A2(n21397), .ZN(n17345) );
  NOR2_X1 U17275 ( .A1(n13809), .A2(n17345), .ZN(n13799) );
  AND2_X1 U17276 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n13808) );
  OR2_X1 U17277 ( .A1(n13800), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13811) );
  NOR2_X1 U17278 ( .A1(n13811), .A2(n11955), .ZN(n13801) );
  NAND2_X1 U17279 ( .A1(n20726), .A2(n15059), .ZN(n20676) );
  NAND3_X1 U17280 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_26__SCAN_IN), .ZN(n13804) );
  NAND2_X1 U17281 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14827) );
  INV_X1 U17282 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20727) );
  INV_X1 U17283 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21386) );
  INV_X1 U17284 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n14257) );
  NOR4_X1 U17285 ( .A1(n20727), .A2(n20739), .A3(n21386), .A4(n14257), .ZN(
        n15046) );
  INV_X1 U17286 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13904) );
  INV_X1 U17287 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20688) );
  INV_X1 U17288 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20699) );
  INV_X1 U17289 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20692) );
  NOR4_X1 U17290 ( .A1(n13904), .A2(n20688), .A3(n20699), .A4(n20692), .ZN(
        n14881) );
  AND2_X1 U17291 ( .A1(n15046), .A2(n14881), .ZN(n14825) );
  AND2_X1 U17292 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n14995) );
  AND2_X1 U17293 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14994) );
  NAND3_X1 U17294 ( .A1(n14995), .A2(n14994), .A3(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14973) );
  AND2_X1 U17295 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14933) );
  NAND3_X1 U17296 ( .A1(n14933), .A2(P1_REIP_REG_14__SCAN_IN), .A3(
        P1_REIP_REG_17__SCAN_IN), .ZN(n13802) );
  NOR2_X1 U17297 ( .A1(n14973), .A2(n13802), .ZN(n14884) );
  AND4_X1 U17298 ( .A1(n14884), .A2(P1_REIP_REG_20__SCAN_IN), .A3(
        P1_REIP_REG_19__SCAN_IN), .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n14826) );
  NAND2_X1 U17299 ( .A1(n14825), .A2(n14826), .ZN(n14844) );
  NOR2_X1 U17300 ( .A1(n14827), .A2(n14844), .ZN(n13803) );
  NAND2_X1 U17301 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n13803), .ZN(n14816) );
  NOR2_X1 U17302 ( .A1(n13804), .A2(n14816), .ZN(n13805) );
  AND2_X1 U17303 ( .A1(n15059), .A2(n13805), .ZN(n14778) );
  AND2_X1 U17304 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n13806) );
  NAND2_X1 U17305 ( .A1(n14778), .A2(n13806), .ZN(n13807) );
  NAND2_X1 U17306 ( .A1(n20676), .A2(n13807), .ZN(n14754) );
  OAI21_X1 U17307 ( .B1(n13808), .B2(n20726), .A(n14754), .ZN(n14682) );
  AND3_X1 U17308 ( .A1(n13811), .A2(n13810), .A3(n13809), .ZN(n13812) );
  NAND2_X1 U17309 ( .A1(n21402), .A2(n13812), .ZN(n20702) );
  INV_X1 U17310 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15085) );
  OAI22_X1 U17311 ( .A1(n13813), .A2(n20718), .B1(n20702), .B2(n15085), .ZN(
        n13817) );
  INV_X1 U17312 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n15222) );
  NOR2_X1 U17313 ( .A1(n14816), .A2(n15222), .ZN(n13814) );
  NAND2_X1 U17314 ( .A1(n15071), .A2(n13814), .ZN(n14805) );
  INV_X1 U17315 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15216) );
  NOR2_X1 U17316 ( .A1(n14805), .A2(n15216), .ZN(n14790) );
  AND2_X1 U17317 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n13815) );
  NAND2_X1 U17318 ( .A1(n14790), .A2(n13815), .ZN(n14765) );
  OR2_X1 U17319 ( .A1(n14765), .A2(n13880), .ZN(n14756) );
  INV_X1 U17320 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n15184) );
  NOR4_X1 U17321 ( .A1(n14756), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n13882), 
        .A4(n15184), .ZN(n13816) );
  AOI211_X1 U17322 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14682), .A(n13817), 
        .B(n13816), .ZN(n13818) );
  NAND2_X1 U17323 ( .A1(n13821), .A2(n13820), .ZN(P1_U2809) );
  NAND2_X1 U17324 ( .A1(n13839), .A2(n17381), .ZN(n13827) );
  NAND2_X1 U17325 ( .A1(n17370), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13822) );
  OAI211_X1 U17326 ( .C1(n14681), .C2(n17377), .A(n13823), .B(n13822), .ZN(
        n13824) );
  NAND2_X1 U17327 ( .A1(n13827), .A2(n13826), .ZN(P1_U2968) );
  AND2_X1 U17328 ( .A1(n14275), .A2(n21404), .ZN(n14276) );
  NAND2_X1 U17329 ( .A1(n12451), .A2(n14276), .ZN(n13828) );
  NAND2_X1 U17330 ( .A1(n13828), .A2(n14088), .ZN(n13829) );
  NAND2_X1 U17331 ( .A1(n14116), .A2(n13829), .ZN(n13834) );
  NOR2_X1 U17332 ( .A1(n13831), .A2(n17352), .ZN(n13832) );
  NAND2_X1 U17333 ( .A1(n13955), .A2(n13832), .ZN(n13833) );
  AND2_X1 U17334 ( .A1(n15151), .A2(n20851), .ZN(n13838) );
  NAND2_X1 U17335 ( .A1(n13839), .A2(n13838), .ZN(n13858) );
  NOR4_X1 U17336 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13843) );
  NOR4_X1 U17337 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n13842) );
  NOR4_X1 U17338 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13841) );
  NOR4_X1 U17339 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13840) );
  AND4_X1 U17340 ( .A1(n13843), .A2(n13842), .A3(n13841), .A4(n13840), .ZN(
        n13848) );
  NOR4_X1 U17341 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13846) );
  NOR4_X1 U17342 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n13845) );
  NOR4_X1 U17343 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n13844) );
  AND4_X1 U17344 ( .A1(n13846), .A2(n13845), .A3(n13844), .A4(n13869), .ZN(
        n13847) );
  NAND2_X1 U17345 ( .A1(n13848), .A2(n13847), .ZN(n13849) );
  NOR3_X1 U17346 ( .A1(n15179), .A2(n20812), .A3(n13853), .ZN(n13850) );
  AOI22_X1 U17347 ( .A1(n15165), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15179), .ZN(n13851) );
  INV_X1 U17348 ( .A(n13851), .ZN(n13856) );
  INV_X1 U17349 ( .A(n20812), .ZN(n13852) );
  NOR2_X1 U17350 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  INV_X1 U17351 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17456) );
  NOR2_X1 U17352 ( .A1(n15153), .A2(n17456), .ZN(n13855) );
  NOR2_X1 U17353 ( .A1(n13856), .A2(n13855), .ZN(n13857) );
  NAND2_X1 U17354 ( .A1(n13858), .A2(n13857), .ZN(P1_U2873) );
  NOR2_X1 U17355 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13860) );
  NOR4_X1 U17356 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13859) );
  NAND4_X1 U17357 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13860), .A4(n13859), .ZN(n13863) );
  NOR2_X4 U17358 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13863), .ZN(n17532)
         );
  INV_X2 U17359 ( .A(n17532), .ZN(U215) );
  NOR3_X1 U17360 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21395), .ZN(n13862) );
  NOR4_X1 U17361 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13861) );
  AOI22_X1 U17362 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n13865) );
  NOR2_X1 U17363 ( .A1(n13864), .A2(n21363), .ZN(n21366) );
  NAND2_X1 U17364 ( .A1(n17352), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n15647) );
  OAI211_X1 U17365 ( .C1(n13865), .C2(n21366), .A(n13946), .B(n15647), .ZN(
        P1_U3195) );
  MUX2_X1 U17366 ( .A(n16887), .B(P2_STATEBS16_REG_SCAN_IN), .S(n16902), .Z(
        n13866) );
  AOI21_X1 U17367 ( .B1(n13866), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n13868) );
  INV_X1 U17368 ( .A(n14169), .ZN(n13867) );
  NOR2_X1 U17369 ( .A1(n13868), .A2(n16904), .ZN(P2_U3178) );
  OAI222_X1 U17370 ( .A1(n13891), .A2(n21386), .B1(n14257), .B2(n21376), .C1(
        n21396), .C2(n13869), .ZN(P1_U3197) );
  INV_X1 U17371 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n13871) );
  INV_X1 U17372 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15324) );
  INV_X1 U17373 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13870) );
  OAI222_X1 U17374 ( .A1(n13891), .A2(n13871), .B1(n15324), .B2(n21376), .C1(
        n13870), .C2(n21396), .ZN(P1_U3209) );
  INV_X1 U17375 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15345) );
  INV_X1 U17376 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21514) );
  OAI222_X1 U17377 ( .A1(n13891), .A2(n15345), .B1(n21396), .B2(n21514), .C1(
        n21376), .C2(n13871), .ZN(P1_U3208) );
  INV_X1 U17378 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21499) );
  INV_X1 U17379 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15313) );
  OAI222_X1 U17380 ( .A1(n13891), .A2(n15324), .B1(n21499), .B2(n21396), .C1(
        n15313), .C2(n21376), .ZN(P1_U3210) );
  INV_X1 U17381 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n13873) );
  OAI21_X1 U17382 ( .B1(n21364), .B2(P1_STATE_REG_2__SCAN_IN), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n13872) );
  AND2_X1 U17383 ( .A1(n13872), .A2(n21407), .ZN(n21385) );
  OAI21_X1 U17384 ( .B1(n21396), .B2(n13873), .A(n21361), .ZN(P1_U2802) );
  INV_X1 U17385 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14871) );
  AOI22_X1 U17386 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n13905), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n13907), .ZN(n13874) );
  OAI21_X1 U17387 ( .B1(n14871), .B2(n13891), .A(n13874), .ZN(P1_U3215) );
  AOI22_X1 U17388 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n13905), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n13907), .ZN(n13875) );
  OAI21_X1 U17389 ( .B1(n15313), .B2(n13891), .A(n13875), .ZN(P1_U3211) );
  AOI22_X1 U17390 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n13905), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n13907), .ZN(n13876) );
  OAI21_X1 U17391 ( .B1(n20699), .B2(n13891), .A(n13876), .ZN(P1_U3202) );
  INV_X1 U17392 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21377) );
  AOI22_X1 U17393 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n13905), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n13907), .ZN(n13877) );
  OAI21_X1 U17394 ( .B1(n21377), .B2(n13891), .A(n13877), .ZN(P1_U3223) );
  AOI22_X1 U17395 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n13878), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n13907), .ZN(n13879) );
  OAI21_X1 U17396 ( .B1(n13880), .B2(n13891), .A(n13879), .ZN(P1_U3224) );
  AOI22_X1 U17397 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(n13878), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n13907), .ZN(n13881) );
  OAI21_X1 U17398 ( .B1(n13882), .B2(n13891), .A(n13881), .ZN(P1_U3226) );
  INV_X1 U17399 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21373) );
  AOI22_X1 U17400 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n13878), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n13907), .ZN(n13883) );
  OAI21_X1 U17401 ( .B1(n21373), .B2(n13891), .A(n13883), .ZN(P1_U3219) );
  INV_X1 U17402 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15355) );
  AOI22_X1 U17403 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n13878), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21407), .ZN(n13884) );
  OAI21_X1 U17404 ( .B1(n15355), .B2(n13891), .A(n13884), .ZN(P1_U3207) );
  INV_X1 U17405 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U17406 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n13878), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21407), .ZN(n13885) );
  OAI21_X1 U17407 ( .B1(n13886), .B2(n13891), .A(n13885), .ZN(P1_U3216) );
  INV_X1 U17408 ( .A(n13891), .ZN(n21374) );
  AOI222_X1 U17409 ( .A1(n21374), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13905), .C1(P1_ADDRESS_REG_1__SCAN_IN), 
        .C2(n21407), .ZN(n13887) );
  INV_X1 U17410 ( .A(n13887), .ZN(P1_U3198) );
  INV_X1 U17411 ( .A(n19837), .ZN(n19813) );
  INV_X1 U17412 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13890) );
  NOR2_X1 U17413 ( .A1(n20614), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13912) );
  INV_X1 U17414 ( .A(n13912), .ZN(n13888) );
  OAI211_X1 U17415 ( .C1(n19813), .C2(n13890), .A(n13889), .B(n13888), .ZN(
        P2_U2814) );
  AOI22_X1 U17416 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(n21407), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(n13878), .ZN(n13892) );
  OAI21_X1 U17417 ( .B1(n15216), .B2(n13891), .A(n13892), .ZN(P1_U3221) );
  INV_X1 U17418 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21371) );
  AOI22_X1 U17419 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n13905), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n21407), .ZN(n13893) );
  OAI21_X1 U17420 ( .B1(n21371), .B2(n13891), .A(n13893), .ZN(P1_U3214) );
  AOI22_X1 U17421 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n13878), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n13907), .ZN(n13894) );
  OAI21_X1 U17422 ( .B1(n15222), .B2(n13891), .A(n13894), .ZN(P1_U3220) );
  INV_X1 U17423 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U17424 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21407), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n13905), .ZN(n13895) );
  OAI21_X1 U17425 ( .B1(n13896), .B2(n13891), .A(n13895), .ZN(P1_U3212) );
  INV_X1 U17426 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20739) );
  AOI22_X1 U17427 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n13878), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n21407), .ZN(n13897) );
  OAI21_X1 U17428 ( .B1(n20739), .B2(n13891), .A(n13897), .ZN(P1_U3199) );
  AOI22_X1 U17429 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13905), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n13907), .ZN(n13898) );
  OAI21_X1 U17430 ( .B1(n20688), .B2(n13891), .A(n13898), .ZN(P1_U3203) );
  INV_X1 U17431 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17432 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n13905), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21407), .ZN(n13899) );
  OAI21_X1 U17433 ( .B1(n13900), .B2(n13891), .A(n13899), .ZN(P1_U3206) );
  AOI22_X1 U17434 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n13878), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n13907), .ZN(n13901) );
  OAI21_X1 U17435 ( .B1(n20692), .B2(n13891), .A(n13901), .ZN(P1_U3201) );
  AOI22_X1 U17436 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n13905), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n13907), .ZN(n13902) );
  OAI21_X1 U17437 ( .B1(n20727), .B2(n13891), .A(n13902), .ZN(P1_U3200) );
  AOI22_X1 U17438 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n21407), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n13905), .ZN(n13903) );
  OAI21_X1 U17439 ( .B1(n13904), .B2(n13891), .A(n13903), .ZN(P1_U3204) );
  INV_X1 U17440 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15249) );
  AOI22_X1 U17441 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n21407), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n13905), .ZN(n13906) );
  OAI21_X1 U17442 ( .B1(n15249), .B2(n13891), .A(n13906), .ZN(P1_U3217) );
  AOI22_X1 U17443 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n13878), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n13907), .ZN(n13908) );
  OAI21_X1 U17444 ( .B1(n15184), .B2(n13891), .A(n13908), .ZN(P1_U3225) );
  AOI21_X1 U17445 ( .B1(n15652), .B2(n16887), .A(n14358), .ZN(n13909) );
  NAND3_X1 U17446 ( .A1(n16848), .A2(n13910), .A3(n13909), .ZN(n16851) );
  AND2_X1 U17447 ( .A1(n16851), .A2(n16899), .ZN(n20636) );
  OAI21_X1 U17448 ( .B1(n20636), .B2(n16853), .A(n13911), .ZN(P2_U2819) );
  INV_X1 U17449 ( .A(n15652), .ZN(n13914) );
  OAI21_X1 U17450 ( .B1(n13912), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19728), 
        .ZN(n13913) );
  OAI21_X1 U17451 ( .B1(n13914), .B2(n19728), .A(n13913), .ZN(P2_U3612) );
  AND2_X1 U17452 ( .A1(n21265), .A2(n21357), .ZN(n14744) );
  AOI21_X1 U17453 ( .B1(n13915), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14744), 
        .ZN(n13916) );
  NAND2_X1 U17454 ( .A1(n14278), .A2(n13916), .ZN(P1_U2801) );
  NAND2_X1 U17455 ( .A1(n13917), .A2(n17446), .ZN(n13918) );
  NAND2_X1 U17456 ( .A1(n13919), .A2(n13918), .ZN(n17448) );
  OAI21_X1 U17457 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19828), .A(
        n13935), .ZN(n17442) );
  NAND2_X1 U17458 ( .A1(n16423), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U17459 ( .B1(n16459), .B2(n17442), .A(n17447), .ZN(n13920) );
  OAI21_X1 U17460 ( .B1(n16450), .B2(n13921), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13922) );
  OAI211_X1 U17461 ( .C1(n17448), .C2(n16446), .A(n13923), .B(n13922), .ZN(
        P2_U3014) );
  INV_X1 U17462 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13929) );
  INV_X1 U17463 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n13925) );
  INV_X1 U17464 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13924) );
  MUX2_X1 U17465 ( .A(n13925), .B(n13924), .S(n16790), .Z(n14643) );
  INV_X1 U17466 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13927) );
  OAI222_X1 U17467 ( .A1(n13993), .A2(n13929), .B1(n13928), .B2(n14643), .C1(
        n13927), .C2(n14077), .ZN(P2_U2982) );
  OR2_X1 U17468 ( .A1(n13930), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13932) );
  NAND2_X1 U17469 ( .A1(n13932), .A2(n13931), .ZN(n19962) );
  XNOR2_X1 U17470 ( .A(n15969), .B(n13933), .ZN(n13934) );
  XNOR2_X1 U17471 ( .A(n13935), .B(n13934), .ZN(n19975) );
  INV_X1 U17472 ( .A(n19975), .ZN(n13936) );
  NAND2_X1 U17473 ( .A1(n16435), .A2(n13936), .ZN(n13937) );
  NAND2_X1 U17474 ( .A1(n16423), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19972) );
  OAI211_X1 U17475 ( .C1(n19962), .C2(n16446), .A(n13937), .B(n19972), .ZN(
        n13938) );
  INV_X1 U17476 ( .A(n13938), .ZN(n13941) );
  MUX2_X1 U17477 ( .A(n16424), .B(n16441), .S(n13939), .Z(n13940) );
  OAI211_X1 U17478 ( .C1(n19965), .C2(n16455), .A(n13941), .B(n13940), .ZN(
        P2_U3013) );
  OR2_X1 U17479 ( .A1(n14116), .A2(n11966), .ZN(n13945) );
  INV_X1 U17480 ( .A(n12451), .ZN(n13942) );
  NAND2_X1 U17481 ( .A1(n13943), .A2(n13942), .ZN(n13944) );
  NAND2_X1 U17482 ( .A1(n13945), .A2(n13944), .ZN(n20641) );
  NAND3_X1 U17483 ( .A1(n13948), .A2(n13947), .A3(n13946), .ZN(n13949) );
  AND2_X1 U17484 ( .A1(n13949), .A2(n21404), .ZN(n21401) );
  NOR2_X1 U17485 ( .A1(n20641), .A2(n21401), .ZN(n17339) );
  NOR2_X1 U17486 ( .A1(n17339), .A2(n20640), .ZN(n20648) );
  INV_X1 U17487 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13957) );
  INV_X1 U17488 ( .A(n13950), .ZN(n13954) );
  NOR2_X1 U17489 ( .A1(n13951), .A2(n12451), .ZN(n13952) );
  MUX2_X1 U17490 ( .A(n13952), .B(n14089), .S(n14116), .Z(n13953) );
  OAI21_X1 U17491 ( .B1(n13955), .B2(n13954), .A(n13953), .ZN(n17336) );
  NAND2_X1 U17492 ( .A1(n20648), .A2(n17336), .ZN(n13956) );
  OAI21_X1 U17493 ( .B1(n20648), .B2(n13957), .A(n13956), .ZN(P1_U3484) );
  XOR2_X1 U17494 ( .A(n13959), .B(n13958), .Z(n19945) );
  XNOR2_X1 U17495 ( .A(n13961), .B(n13960), .ZN(n19942) );
  NOR2_X1 U17496 ( .A1(n16459), .A2(n19942), .ZN(n13964) );
  NAND2_X1 U17497 ( .A1(n16423), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19947) );
  NAND2_X1 U17498 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13962) );
  OAI211_X1 U17499 ( .C1(n16441), .C2(n15953), .A(n19947), .B(n13962), .ZN(
        n13963) );
  AOI211_X1 U17500 ( .C1(n19945), .C2(n16457), .A(n13964), .B(n13963), .ZN(
        n13965) );
  OAI21_X1 U17501 ( .B1(n16768), .B2(n16455), .A(n13965), .ZN(P2_U3012) );
  INV_X1 U17502 ( .A(n14089), .ZN(n13968) );
  INV_X1 U17503 ( .A(n12302), .ZN(n14082) );
  NAND2_X1 U17504 ( .A1(n17346), .A2(n21404), .ZN(n13966) );
  AOI21_X1 U17505 ( .B1(n17323), .B2(n14082), .A(n13966), .ZN(n13967) );
  MUX2_X1 U17506 ( .A(n13968), .B(n13967), .S(n14116), .Z(n13974) );
  OR2_X1 U17507 ( .A1(n13971), .A2(n13970), .ZN(n13972) );
  INV_X1 U17508 ( .A(n14504), .ZN(n17436) );
  NAND2_X1 U17509 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17436), .ZN(n17440) );
  INV_X1 U17510 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20647) );
  NOR2_X1 U17511 ( .A1(n17440), .A2(n20647), .ZN(n13975) );
  AOI21_X1 U17512 ( .B1(n17324), .B2(n14115), .A(n13975), .ZN(n13978) );
  INV_X1 U17513 ( .A(n20953), .ZN(n21188) );
  NOR2_X1 U17514 ( .A1(n13976), .A2(n21188), .ZN(n13977) );
  XOR2_X1 U17515 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n13977), .Z(
        n20715) );
  INV_X1 U17516 ( .A(n13831), .ZN(n14499) );
  INV_X1 U17517 ( .A(n13978), .ZN(n13979) );
  NAND4_X1 U17518 ( .A1(n20715), .A2(n15629), .A3(n14499), .A4(n13979), .ZN(
        n13980) );
  OAI21_X1 U17519 ( .B1(n13981), .B2(n15640), .A(n13980), .ZN(P1_U3468) );
  INV_X1 U17520 ( .A(n16844), .ZN(n13983) );
  INV_X1 U17521 ( .A(n16845), .ZN(n13982) );
  NAND2_X1 U17522 ( .A1(n13983), .A2(n13982), .ZN(n14361) );
  NAND2_X1 U17523 ( .A1(n14361), .A2(n11470), .ZN(n13984) );
  NOR2_X1 U17524 ( .A1(n16902), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13985) );
  OAI211_X1 U17525 ( .C1(n13987), .C2(n13149), .A(n13986), .B(n13985), .ZN(
        n13988) );
  INV_X1 U17526 ( .A(n13988), .ZN(n13989) );
  NAND2_X1 U17527 ( .A1(n16813), .A2(n19863), .ZN(n13991) );
  OAI211_X1 U17528 ( .C1(n13992), .C2(n19866), .A(n13991), .B(n13990), .ZN(
        P2_U2887) );
  INV_X1 U17529 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13996) );
  NAND2_X1 U17530 ( .A1(n14073), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13995) );
  NAND2_X1 U17531 ( .A1(n16790), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13994) );
  OAI21_X1 U17532 ( .B1(n16790), .B2(n19105), .A(n13994), .ZN(n19867) );
  NAND2_X1 U17533 ( .A1(n14048), .A2(n19867), .ZN(n14016) );
  OAI211_X1 U17534 ( .C1(n14077), .C2(n13996), .A(n13995), .B(n14016), .ZN(
        P2_U2952) );
  INV_X1 U17535 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14517) );
  NAND2_X1 U17536 ( .A1(n14073), .A2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13999) );
  NAND2_X1 U17537 ( .A1(n16788), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13998) );
  NAND2_X1 U17538 ( .A1(n16790), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13997) );
  AND2_X1 U17539 ( .A1(n13998), .A2(n13997), .ZN(n19908) );
  NAND2_X1 U17540 ( .A1(n14048), .A2(n19989), .ZN(n14037) );
  OAI211_X1 U17541 ( .C1(n14077), .C2(n14517), .A(n13999), .B(n14037), .ZN(
        P2_U2953) );
  INV_X1 U17542 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19926) );
  NAND2_X1 U17543 ( .A1(n14073), .A2(P2_LWORD_REG_6__SCAN_IN), .ZN(n14002) );
  INV_X1 U17544 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n14001) );
  NAND2_X1 U17545 ( .A1(n16790), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14000) );
  OAI21_X1 U17546 ( .B1(n16790), .B2(n14001), .A(n14000), .ZN(n20016) );
  NAND2_X1 U17547 ( .A1(n14048), .A2(n20016), .ZN(n14050) );
  OAI211_X1 U17548 ( .C1(n14077), .C2(n19926), .A(n14002), .B(n14050), .ZN(
        P2_U2973) );
  INV_X1 U17549 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n14004) );
  NAND2_X1 U17550 ( .A1(n14073), .A2(P2_LWORD_REG_5__SCAN_IN), .ZN(n14003) );
  MUX2_X1 U17551 ( .A(BUF2_REG_5__SCAN_IN), .B(BUF1_REG_5__SCAN_IN), .S(n16790), .Z(n20007) );
  NAND2_X1 U17552 ( .A1(n14048), .A2(n20007), .ZN(n14053) );
  OAI211_X1 U17553 ( .C1(n14077), .C2(n14004), .A(n14003), .B(n14053), .ZN(
        P2_U2972) );
  INV_X1 U17554 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n14008) );
  NAND2_X1 U17555 ( .A1(n14073), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n14007) );
  NAND2_X1 U17556 ( .A1(n16788), .A2(BUF2_REG_4__SCAN_IN), .ZN(n14006) );
  NAND2_X1 U17557 ( .A1(n16790), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14005) );
  AND2_X1 U17558 ( .A1(n14006), .A2(n14005), .ZN(n19882) );
  INV_X1 U17559 ( .A(n19882), .ZN(n20003) );
  NAND2_X1 U17560 ( .A1(n14048), .A2(n20003), .ZN(n14055) );
  OAI211_X1 U17561 ( .C1(n14077), .C2(n14008), .A(n14007), .B(n14055), .ZN(
        P2_U2971) );
  INV_X1 U17562 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n14012) );
  NAND2_X1 U17563 ( .A1(n14073), .A2(P2_LWORD_REG_3__SCAN_IN), .ZN(n14011) );
  NAND2_X1 U17564 ( .A1(n16788), .A2(BUF2_REG_3__SCAN_IN), .ZN(n14010) );
  NAND2_X1 U17565 ( .A1(n16790), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14009) );
  AND2_X1 U17566 ( .A1(n14010), .A2(n14009), .ZN(n19889) );
  INV_X1 U17567 ( .A(n19889), .ZN(n19998) );
  NAND2_X1 U17568 ( .A1(n14048), .A2(n19998), .ZN(n14041) );
  OAI211_X1 U17569 ( .C1(n14077), .C2(n14012), .A(n14011), .B(n14041), .ZN(
        P2_U2970) );
  INV_X1 U17570 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14477) );
  NAND2_X1 U17571 ( .A1(n14073), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14015) );
  INV_X1 U17572 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n14014) );
  NAND2_X1 U17573 ( .A1(n16790), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14013) );
  OAI21_X1 U17574 ( .B1(n16790), .B2(n14014), .A(n14013), .ZN(n16074) );
  NAND2_X1 U17575 ( .A1(n14048), .A2(n16074), .ZN(n14020) );
  OAI211_X1 U17576 ( .C1(n14077), .C2(n14477), .A(n14015), .B(n14020), .ZN(
        P2_U2965) );
  INV_X1 U17577 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n14018) );
  NAND2_X1 U17578 ( .A1(n14073), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n14017) );
  OAI211_X1 U17579 ( .C1(n14077), .C2(n14018), .A(n14017), .B(n14016), .ZN(
        P2_U2967) );
  INV_X1 U17580 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14515) );
  NAND2_X1 U17581 ( .A1(n14073), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14019) );
  NAND2_X1 U17582 ( .A1(n14048), .A2(n14588), .ZN(n14062) );
  OAI211_X1 U17583 ( .C1(n14515), .C2(n14077), .A(n14019), .B(n14062), .ZN(
        P2_U2966) );
  INV_X1 U17584 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n14022) );
  NAND2_X1 U17585 ( .A1(n14073), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n14021) );
  OAI211_X1 U17586 ( .C1(n14077), .C2(n14022), .A(n14021), .B(n14020), .ZN(
        P2_U2980) );
  INV_X1 U17587 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n14026) );
  NAND2_X1 U17588 ( .A1(n14073), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n14025) );
  INV_X1 U17589 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n14024) );
  NAND2_X1 U17590 ( .A1(n16790), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14023) );
  OAI21_X1 U17591 ( .B1(n16790), .B2(n14024), .A(n14023), .ZN(n16081) );
  NAND2_X1 U17592 ( .A1(n14048), .A2(n16081), .ZN(n14066) );
  OAI211_X1 U17593 ( .C1(n14077), .C2(n14026), .A(n14025), .B(n14066), .ZN(
        P2_U2979) );
  INV_X1 U17594 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14184) );
  NAND2_X1 U17595 ( .A1(n14073), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14029) );
  INV_X1 U17596 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U17597 ( .A1(n16790), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14027) );
  OAI21_X1 U17598 ( .B1(n16790), .B2(n14028), .A(n14027), .ZN(n16102) );
  NAND2_X1 U17599 ( .A1(n14048), .A2(n16102), .ZN(n14074) );
  OAI211_X1 U17600 ( .C1(n14077), .C2(n14184), .A(n14029), .B(n14074), .ZN(
        P2_U2961) );
  INV_X1 U17601 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14177) );
  NAND2_X1 U17602 ( .A1(n14073), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n14032) );
  INV_X1 U17603 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n14031) );
  NAND2_X1 U17604 ( .A1(n16790), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14030) );
  OAI21_X1 U17605 ( .B1(n16790), .B2(n14031), .A(n14030), .ZN(n16109) );
  NAND2_X1 U17606 ( .A1(n14048), .A2(n16109), .ZN(n14068) );
  OAI211_X1 U17607 ( .C1(n14077), .C2(n14177), .A(n14032), .B(n14068), .ZN(
        P2_U2960) );
  INV_X1 U17608 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n14036) );
  NAND2_X1 U17609 ( .A1(n14073), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n14035) );
  INV_X1 U17610 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n14034) );
  NAND2_X1 U17611 ( .A1(n16790), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14033) );
  OAI21_X1 U17612 ( .B1(n16790), .B2(n14034), .A(n14033), .ZN(n16088) );
  NAND2_X1 U17613 ( .A1(n14048), .A2(n16088), .ZN(n14060) );
  OAI211_X1 U17614 ( .C1(n14077), .C2(n14036), .A(n14035), .B(n14060), .ZN(
        P2_U2978) );
  INV_X1 U17615 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19936) );
  NAND2_X1 U17616 ( .A1(n14073), .A2(P2_LWORD_REG_1__SCAN_IN), .ZN(n14038) );
  OAI211_X1 U17617 ( .C1(n14077), .C2(n19936), .A(n14038), .B(n14037), .ZN(
        P2_U2968) );
  INV_X1 U17618 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14181) );
  NAND2_X1 U17619 ( .A1(n14073), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14040) );
  INV_X1 U17620 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18525) );
  NAND2_X1 U17621 ( .A1(n16790), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14039) );
  OAI21_X1 U17622 ( .B1(n16790), .B2(n18525), .A(n14039), .ZN(n16095) );
  NAND2_X1 U17623 ( .A1(n14048), .A2(n16095), .ZN(n14064) );
  OAI211_X1 U17624 ( .C1(n14181), .C2(n14077), .A(n14040), .B(n14064), .ZN(
        P2_U2962) );
  INV_X1 U17625 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14179) );
  NAND2_X1 U17626 ( .A1(n14073), .A2(P2_UWORD_REG_3__SCAN_IN), .ZN(n14042) );
  OAI211_X1 U17627 ( .C1(n14077), .C2(n14179), .A(n14042), .B(n14041), .ZN(
        P2_U2955) );
  INV_X1 U17628 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14175) );
  NAND2_X1 U17629 ( .A1(n14073), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n14045) );
  NAND2_X1 U17630 ( .A1(n16788), .A2(BUF2_REG_2__SCAN_IN), .ZN(n14044) );
  NAND2_X1 U17631 ( .A1(n16790), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14043) );
  AND2_X1 U17632 ( .A1(n14044), .A2(n14043), .ZN(n19897) );
  NAND2_X1 U17633 ( .A1(n14048), .A2(n19993), .ZN(n14058) );
  OAI211_X1 U17634 ( .C1(n14077), .C2(n14175), .A(n14045), .B(n14058), .ZN(
        P2_U2954) );
  INV_X1 U17635 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14173) );
  NAND2_X1 U17636 ( .A1(n14073), .A2(P2_UWORD_REG_7__SCAN_IN), .ZN(n14049) );
  INV_X1 U17637 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n14047) );
  NAND2_X1 U17638 ( .A1(n16790), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14046) );
  OAI21_X1 U17639 ( .B1(n16790), .B2(n14047), .A(n14046), .ZN(n20026) );
  NAND2_X1 U17640 ( .A1(n14048), .A2(n20026), .ZN(n14071) );
  OAI211_X1 U17641 ( .C1(n14077), .C2(n14173), .A(n14049), .B(n14071), .ZN(
        P2_U2959) );
  INV_X1 U17642 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14052) );
  NAND2_X1 U17643 ( .A1(n14073), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n14051) );
  OAI211_X1 U17644 ( .C1(n14077), .C2(n14052), .A(n14051), .B(n14050), .ZN(
        P2_U2958) );
  INV_X1 U17645 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14171) );
  NAND2_X1 U17646 ( .A1(n14073), .A2(P2_UWORD_REG_5__SCAN_IN), .ZN(n14054) );
  OAI211_X1 U17647 ( .C1(n14077), .C2(n14171), .A(n14054), .B(n14053), .ZN(
        P2_U2957) );
  INV_X1 U17648 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14057) );
  NAND2_X1 U17649 ( .A1(n14073), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n14056) );
  OAI211_X1 U17650 ( .C1(n14077), .C2(n14057), .A(n14056), .B(n14055), .ZN(
        P2_U2956) );
  INV_X1 U17651 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19934) );
  NAND2_X1 U17652 ( .A1(n14073), .A2(P2_LWORD_REG_2__SCAN_IN), .ZN(n14059) );
  OAI211_X1 U17653 ( .C1(n14077), .C2(n19934), .A(n14059), .B(n14058), .ZN(
        P2_U2969) );
  INV_X1 U17654 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14513) );
  NAND2_X1 U17655 ( .A1(n14073), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14061) );
  OAI211_X1 U17656 ( .C1(n14077), .C2(n14513), .A(n14061), .B(n14060), .ZN(
        P2_U2963) );
  INV_X1 U17657 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19915) );
  NAND2_X1 U17658 ( .A1(n14073), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n14063) );
  OAI211_X1 U17659 ( .C1(n19915), .C2(n14077), .A(n14063), .B(n14062), .ZN(
        P2_U2981) );
  INV_X1 U17660 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19920) );
  NAND2_X1 U17661 ( .A1(n14073), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14065) );
  OAI211_X1 U17662 ( .C1(n19920), .C2(n14077), .A(n14065), .B(n14064), .ZN(
        P2_U2977) );
  INV_X1 U17663 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14519) );
  NAND2_X1 U17664 ( .A1(n14073), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14067) );
  OAI211_X1 U17665 ( .C1(n14077), .C2(n14519), .A(n14067), .B(n14066), .ZN(
        P2_U2964) );
  INV_X1 U17666 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n14070) );
  NAND2_X1 U17667 ( .A1(n14073), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n14069) );
  OAI211_X1 U17668 ( .C1(n14077), .C2(n14070), .A(n14069), .B(n14068), .ZN(
        P2_U2975) );
  INV_X1 U17669 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19924) );
  NAND2_X1 U17670 ( .A1(n14073), .A2(P2_LWORD_REG_7__SCAN_IN), .ZN(n14072) );
  OAI211_X1 U17671 ( .C1(n14077), .C2(n19924), .A(n14072), .B(n14071), .ZN(
        P2_U2974) );
  INV_X1 U17672 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n14076) );
  NAND2_X1 U17673 ( .A1(n14073), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n14075) );
  OAI211_X1 U17674 ( .C1(n14077), .C2(n14076), .A(n14075), .B(n14074), .ZN(
        P2_U2976) );
  INV_X1 U17675 ( .A(n14079), .ZN(n14081) );
  NAND3_X1 U17676 ( .A1(n14082), .A2(n14081), .A3(n14080), .ZN(n14083) );
  NOR2_X1 U17677 ( .A1(n14084), .A2(n14083), .ZN(n14086) );
  NAND2_X1 U17678 ( .A1(n14086), .A2(n13831), .ZN(n15628) );
  INV_X1 U17679 ( .A(n15628), .ZN(n14709) );
  OR2_X1 U17680 ( .A1(n14078), .A2(n14709), .ZN(n14094) );
  NAND2_X1 U17681 ( .A1(n14086), .A2(n14085), .ZN(n14482) );
  XNOR2_X1 U17682 ( .A(n14087), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14097) );
  INV_X1 U17683 ( .A(n17323), .ZN(n14708) );
  XNOR2_X1 U17684 ( .A(n14101), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14090) );
  NAND2_X1 U17685 ( .A1(n14089), .A2(n14088), .ZN(n14490) );
  AOI22_X1 U17686 ( .A1(n14708), .A2(n14090), .B1(n14490), .B2(n14097), .ZN(
        n14091) );
  OAI21_X1 U17687 ( .B1(n14482), .B2(n14097), .A(n14091), .ZN(n14092) );
  INV_X1 U17688 ( .A(n14092), .ZN(n14093) );
  NAND2_X1 U17689 ( .A1(n14094), .A2(n14093), .ZN(n14479) );
  OAI22_X1 U17690 ( .A1(n14095), .A2(n14261), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15631) );
  INV_X1 U17691 ( .A(n15631), .ZN(n14099) );
  NOR2_X1 U17692 ( .A1(n21357), .A2(n14194), .ZN(n15632) );
  INV_X1 U17693 ( .A(n14097), .ZN(n14098) );
  AOI222_X1 U17694 ( .A1(n14479), .A2(n15629), .B1(n14099), .B2(n15632), .C1(
        n17358), .C2(n14098), .ZN(n14100) );
  MUX2_X1 U17695 ( .A(n14101), .B(n14100), .S(n15640), .Z(n14102) );
  INV_X1 U17696 ( .A(n14102), .ZN(P1_U3472) );
  INV_X1 U17697 ( .A(n14103), .ZN(n14106) );
  OAI21_X1 U17698 ( .B1(n14106), .B2(n14105), .A(n14104), .ZN(n15083) );
  INV_X1 U17699 ( .A(n14107), .ZN(n14109) );
  AOI21_X1 U17700 ( .B1(n14109), .B2(n14194), .A(n14108), .ZN(n15613) );
  INV_X1 U17701 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21392) );
  NOR2_X1 U17702 ( .A1(n20716), .A2(n21392), .ZN(n15612) );
  INV_X1 U17703 ( .A(n14110), .ZN(n14112) );
  INV_X1 U17704 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14111) );
  AOI21_X1 U17705 ( .B1(n17385), .B2(n14112), .A(n14111), .ZN(n14113) );
  AOI211_X1 U17706 ( .C1(n15613), .C2(n17382), .A(n15612), .B(n14113), .ZN(
        n14114) );
  OAI21_X1 U17707 ( .B1(n20811), .B2(n15083), .A(n14114), .ZN(P1_U2999) );
  NAND3_X1 U17708 ( .A1(n14116), .A2(n14115), .A3(n14708), .ZN(n14117) );
  OAI21_X1 U17709 ( .B1(n14278), .B2(n14275), .A(n14117), .ZN(n14118) );
  NAND2_X1 U17710 ( .A1(n10287), .A2(n17436), .ZN(n20774) );
  INV_X2 U17711 ( .A(n20774), .ZN(n20784) );
  AOI22_X1 U17712 ( .A1(n20784), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14120) );
  OAI21_X1 U17713 ( .B1(n12901), .B2(n14135), .A(n14120), .ZN(P1_U2913) );
  INV_X1 U17714 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14311) );
  AOI22_X1 U17715 ( .A1(n20784), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14121) );
  OAI21_X1 U17716 ( .B1(n14311), .B2(n14135), .A(n14121), .ZN(P1_U2918) );
  INV_X1 U17717 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21454) );
  AOI22_X1 U17718 ( .A1(n20784), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14122) );
  OAI21_X1 U17719 ( .B1(n21454), .B2(n14135), .A(n14122), .ZN(P1_U2915) );
  INV_X1 U17720 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14337) );
  AOI22_X1 U17721 ( .A1(n20784), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14123) );
  OAI21_X1 U17722 ( .B1(n14337), .B2(n14135), .A(n14123), .ZN(P1_U2908) );
  AOI22_X1 U17723 ( .A1(n20784), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14124) );
  OAI21_X1 U17724 ( .B1(n15130), .B2(n14135), .A(n14124), .ZN(P1_U2911) );
  INV_X1 U17725 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U17726 ( .A1(n20784), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14125) );
  OAI21_X1 U17727 ( .B1(n14341), .B2(n14135), .A(n14125), .ZN(P1_U2912) );
  AOI22_X1 U17728 ( .A1(n20784), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14126) );
  OAI21_X1 U17729 ( .B1(n15152), .B2(n14135), .A(n14126), .ZN(P1_U2917) );
  AOI22_X1 U17730 ( .A1(n20784), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14127) );
  OAI21_X1 U17731 ( .B1(n15125), .B2(n14135), .A(n14127), .ZN(P1_U2910) );
  INV_X1 U17732 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14282) );
  AOI22_X1 U17733 ( .A1(n20784), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14128) );
  OAI21_X1 U17734 ( .B1(n14282), .B2(n14135), .A(n14128), .ZN(P1_U2914) );
  INV_X1 U17735 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U17736 ( .A1(n20784), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14129) );
  OAI21_X1 U17737 ( .B1(n14323), .B2(n14135), .A(n14129), .ZN(P1_U2906) );
  INV_X1 U17738 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14327) );
  AOI22_X1 U17739 ( .A1(n20784), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14130) );
  OAI21_X1 U17740 ( .B1(n14327), .B2(n14135), .A(n14130), .ZN(P1_U2907) );
  INV_X1 U17741 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14295) );
  AOI22_X1 U17742 ( .A1(n20784), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14131) );
  OAI21_X1 U17743 ( .B1(n14295), .B2(n14135), .A(n14131), .ZN(P1_U2920) );
  INV_X1 U17744 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14299) );
  AOI22_X1 U17745 ( .A1(n20784), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14132) );
  OAI21_X1 U17746 ( .B1(n14299), .B2(n14135), .A(n14132), .ZN(P1_U2909) );
  INV_X1 U17747 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14292) );
  AOI22_X1 U17748 ( .A1(n20784), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14133) );
  OAI21_X1 U17749 ( .B1(n14292), .B2(n14135), .A(n14133), .ZN(P1_U2919) );
  INV_X1 U17750 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U17751 ( .A1(n20784), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14134) );
  OAI21_X1 U17752 ( .B1(n14333), .B2(n14135), .A(n14134), .ZN(P1_U2916) );
  NOR2_X1 U17753 ( .A1(n19965), .A2(n16065), .ZN(n14138) );
  AOI21_X1 U17754 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n16065), .A(n14138), .ZN(
        n14139) );
  OAI21_X1 U17755 ( .B1(n16798), .B2(n19855), .A(n14139), .ZN(P2_U2886) );
  NAND2_X1 U17756 ( .A1(n14140), .A2(n19710), .ZN(n14392) );
  NOR3_X1 U17757 ( .A1(n14143), .A2(n18277), .A3(n14142), .ZN(n14144) );
  NOR2_X1 U17758 ( .A1(n17180), .A2(n14145), .ZN(n14146) );
  NOR2_X1 U17759 ( .A1(n14147), .A2(n18293), .ZN(n18398) );
  INV_X1 U17760 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18491) );
  NOR2_X1 U17761 ( .A1(n18277), .A2(n18293), .ZN(n18379) );
  INV_X1 U17762 ( .A(n18379), .ZN(n18294) );
  OAI22_X1 U17763 ( .A1(n14241), .A2(n18491), .B1(P3_EAX_REG_0__SCAN_IN), .B2(
        n18294), .ZN(n14148) );
  AOI21_X1 U17764 ( .B1(n14215), .B2(n18382), .A(n14148), .ZN(n14149) );
  OAI21_X1 U17765 ( .B1(n19105), .B2(n18430), .A(n14149), .ZN(P3_U2735) );
  INV_X1 U17766 ( .A(n14437), .ZN(n20621) );
  OR2_X1 U17767 ( .A1(n20614), .A2(n20408), .ZN(n16786) );
  OAI21_X1 U17768 ( .B1(n16798), .B2(n20621), .A(n16786), .ZN(n14155) );
  NAND2_X1 U17769 ( .A1(n16797), .A2(n14150), .ZN(n14438) );
  OR2_X1 U17770 ( .A1(n14152), .A2(n14151), .ZN(n14153) );
  NAND2_X1 U17771 ( .A1(n14154), .A2(n14153), .ZN(n19959) );
  AOI22_X1 U17772 ( .A1(n14155), .A2(n14438), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19959), .ZN(n14163) );
  NAND2_X1 U17773 ( .A1(n16902), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14156) );
  NAND2_X1 U17774 ( .A1(n20629), .A2(n16853), .ZN(n14160) );
  NAND2_X1 U17775 ( .A1(n14160), .A2(n16904), .ZN(n14161) );
  NAND2_X1 U17776 ( .A1(n20119), .A2(n14161), .ZN(n20626) );
  INV_X1 U17777 ( .A(n20626), .ZN(n20625) );
  NAND2_X1 U17778 ( .A1(n20625), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14162) );
  OAI21_X1 U17779 ( .B1(n14163), .B2(n20625), .A(n14162), .ZN(P2_U3604) );
  NAND2_X1 U17780 ( .A1(n14359), .A2(n16899), .ZN(n14166) );
  NAND2_X1 U17781 ( .A1(n14166), .A2(n14077), .ZN(n14167) );
  NOR2_X4 U17782 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14169), .ZN(n19927) );
  NOR2_X4 U17783 ( .A1(n19928), .A2(n19927), .ZN(n14475) );
  AOI22_X1 U17784 ( .A1(n19927), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14170) );
  OAI21_X1 U17785 ( .B1(n14171), .B2(n19910), .A(n14170), .ZN(P2_U2930) );
  AOI22_X1 U17786 ( .A1(n19927), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14172) );
  OAI21_X1 U17787 ( .B1(n14173), .B2(n19910), .A(n14172), .ZN(P2_U2928) );
  AOI22_X1 U17788 ( .A1(n19927), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14174) );
  OAI21_X1 U17789 ( .B1(n14175), .B2(n19910), .A(n14174), .ZN(P2_U2933) );
  AOI22_X1 U17790 ( .A1(n19927), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14176) );
  OAI21_X1 U17791 ( .B1(n14177), .B2(n19910), .A(n14176), .ZN(P2_U2927) );
  AOI22_X1 U17792 ( .A1(n19927), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14178) );
  OAI21_X1 U17793 ( .B1(n14179), .B2(n19910), .A(n14178), .ZN(P2_U2932) );
  AOI22_X1 U17794 ( .A1(n19927), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14180) );
  OAI21_X1 U17795 ( .B1(n14181), .B2(n19910), .A(n14180), .ZN(P2_U2925) );
  AOI22_X1 U17796 ( .A1(n19927), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14182) );
  OAI21_X1 U17797 ( .B1(n14057), .B2(n19910), .A(n14182), .ZN(P2_U2931) );
  AOI22_X1 U17798 ( .A1(n19927), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14183) );
  OAI21_X1 U17799 ( .B1(n14184), .B2(n19910), .A(n14183), .ZN(P2_U2926) );
  OAI21_X1 U17800 ( .B1(n14186), .B2(n14185), .A(n14430), .ZN(n15075) );
  OAI22_X1 U17801 ( .A1(n15114), .A2(n14193), .B1(n12352), .B2(n15113), .ZN(
        n14188) );
  INV_X1 U17802 ( .A(n14188), .ZN(n14189) );
  OAI21_X1 U17803 ( .B1(n15075), .B2(n15101), .A(n14189), .ZN(P1_U2871) );
  XNOR2_X1 U17804 ( .A(n14190), .B(n14261), .ZN(n14250) );
  NAND3_X1 U17805 ( .A1(n17404), .A2(n14261), .A3(n14191), .ZN(n14192) );
  NAND2_X1 U17806 ( .A1(n17416), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14248) );
  OAI211_X1 U17807 ( .C1(n17390), .C2(n14193), .A(n14192), .B(n14248), .ZN(
        n14198) );
  INV_X1 U17808 ( .A(n15464), .ZN(n14195) );
  OAI21_X1 U17809 ( .B1(n14469), .B2(n14195), .A(n14194), .ZN(n15617) );
  AOI21_X1 U17810 ( .B1(n14196), .B2(n15617), .A(n14261), .ZN(n14197) );
  AOI211_X1 U17811 ( .C1(n17429), .C2(n14250), .A(n14198), .B(n14197), .ZN(
        n14199) );
  INV_X1 U17812 ( .A(n14199), .ZN(P1_U3030) );
  NOR2_X1 U17813 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14202) );
  OR2_X1 U17814 ( .A1(n14202), .A2(n14201), .ZN(n15610) );
  OAI222_X1 U17815 ( .A1(n15610), .A2(n15114), .B1(n15113), .B2(n21553), .C1(
        n15083), .C2(n15111), .ZN(P1_U2872) );
  OAI21_X1 U17816 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n18277), .A(n14241), .ZN(
        n14203) );
  AOI22_X1 U17817 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18398), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n14203), .ZN(n14205) );
  INV_X1 U17818 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18515) );
  NAND3_X1 U17819 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18379), .A3(n18515), .ZN(
        n14204) );
  OAI211_X1 U17820 ( .C1(n14206), .C2(n18427), .A(n14205), .B(n14204), .ZN(
        P3_U2734) );
  NAND2_X1 U17821 ( .A1(n14208), .A2(n14207), .ZN(n14209) );
  INV_X1 U17822 ( .A(DATAI_1_), .ZN(n14211) );
  NAND2_X1 U17823 ( .A1(n20812), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14210) );
  OAI21_X1 U17824 ( .B1(n20812), .B2(n14211), .A(n14210), .ZN(n15160) );
  INV_X1 U17825 ( .A(n15160), .ZN(n20829) );
  INV_X1 U17826 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20782) );
  OAI222_X1 U17827 ( .A1(n15075), .A2(n15182), .B1(n14639), .B2(n20829), .C1(
        n15151), .C2(n20782), .ZN(P1_U2903) );
  INV_X1 U17828 ( .A(DATAI_0_), .ZN(n14213) );
  NAND2_X1 U17829 ( .A1(n20812), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14212) );
  OAI21_X1 U17830 ( .B1(n20812), .B2(n14213), .A(n14212), .ZN(n20821) );
  INV_X1 U17831 ( .A(n20821), .ZN(n14293) );
  INV_X1 U17832 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20787) );
  OAI222_X1 U17833 ( .A1(n15083), .A2(n15182), .B1(n14639), .B2(n14293), .C1(
        n15151), .C2(n20787), .ZN(P1_U2904) );
  NOR2_X1 U17834 ( .A1(n14215), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14227) );
  XNOR2_X1 U17835 ( .A(n14214), .B(n14227), .ZN(n18812) );
  INV_X1 U17836 ( .A(n19086), .ZN(n17075) );
  OAI21_X1 U17837 ( .B1(n14214), .B2(n14226), .A(n14216), .ZN(n18816) );
  NAND2_X1 U17838 ( .A1(n18905), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18814) );
  OAI21_X1 U17839 ( .B1(n17075), .B2(n18816), .A(n18814), .ZN(n14217) );
  INV_X1 U17840 ( .A(n14217), .ZN(n14222) );
  OAI21_X1 U17841 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18914), .A(
        n19030), .ZN(n14220) );
  NAND2_X1 U17842 ( .A1(n19546), .A2(n18991), .ZN(n18874) );
  INV_X1 U17843 ( .A(n18874), .ZN(n18894) );
  NAND2_X1 U17844 ( .A1(n19062), .A2(n10220), .ZN(n14218) );
  NOR2_X1 U17845 ( .A1(n18894), .A2(n14218), .ZN(n14231) );
  NOR2_X1 U17846 ( .A1(n14231), .A2(n19066), .ZN(n14219) );
  MUX2_X1 U17847 ( .A(n14220), .B(n14219), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n14221) );
  OAI211_X1 U17848 ( .C1(n19095), .C2(n18812), .A(n14222), .B(n14221), .ZN(
        P3_U2861) );
  INV_X1 U17849 ( .A(n16799), .ZN(n16769) );
  MUX2_X1 U17850 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n19943), .S(n19866), .Z(
        n14224) );
  AOI21_X1 U17851 ( .B1(n16769), .B2(n19863), .A(n14224), .ZN(n14225) );
  INV_X1 U17852 ( .A(n14225), .ZN(P2_U2885) );
  INV_X1 U17853 ( .A(n14226), .ZN(n14229) );
  INV_X1 U17854 ( .A(n14227), .ZN(n14228) );
  NAND2_X1 U17855 ( .A1(n14229), .A2(n14228), .ZN(n17062) );
  INV_X1 U17856 ( .A(n17062), .ZN(n17061) );
  INV_X1 U17857 ( .A(n18914), .ZN(n14230) );
  OAI21_X1 U17858 ( .B1(n18905), .B2(n14230), .A(n19090), .ZN(n14233) );
  INV_X1 U17859 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19696) );
  OAI22_X1 U17860 ( .A1(n17075), .A2(n17062), .B1(n19696), .B2(n18992), .ZN(
        n14232) );
  AOI211_X1 U17861 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n14233), .A(
        n14232), .B(n14231), .ZN(n14234) );
  OAI21_X1 U17862 ( .B1(n17061), .B2(n19095), .A(n14234), .ZN(P3_U2862) );
  NOR2_X1 U17863 ( .A1(n16733), .A2(n16065), .ZN(n14239) );
  AOI21_X1 U17864 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16065), .A(n14239), .ZN(
        n14240) );
  OAI21_X1 U17865 ( .B1(n16775), .B2(n19855), .A(n14240), .ZN(P2_U2884) );
  NOR3_X1 U17866 ( .A1(n18515), .A2(n18491), .A3(n18294), .ZN(n14242) );
  AOI21_X1 U17867 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18425), .A(n14242), .ZN(
        n14246) );
  AND2_X1 U17868 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n14242), .ZN(n18424) );
  INV_X1 U17869 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19116) );
  OAI22_X1 U17870 ( .A1(n18427), .A2(n14243), .B1(n18430), .B2(n19116), .ZN(
        n14244) );
  INV_X1 U17871 ( .A(n14244), .ZN(n14245) );
  OAI21_X1 U17872 ( .B1(n14246), .B2(n18424), .A(n14245), .ZN(P3_U2733) );
  MUX2_X1 U17873 ( .A(n17377), .B(n17385), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14247) );
  OAI211_X1 U17874 ( .C1(n15075), .C2(n20811), .A(n14248), .B(n14247), .ZN(
        n14249) );
  AOI21_X1 U17875 ( .B1(n17382), .B2(n14250), .A(n14249), .ZN(n14251) );
  INV_X1 U17876 ( .A(n14251), .ZN(P1_U2998) );
  XOR2_X1 U17877 ( .A(n14253), .B(n14252), .Z(n14435) );
  NAND2_X1 U17878 ( .A1(n14255), .A2(n14254), .ZN(n14256) );
  NAND2_X1 U17879 ( .A1(n14447), .A2(n14256), .ZN(n14431) );
  OAI22_X1 U17880 ( .A1(n17390), .A2(n14431), .B1(n14257), .B2(n20716), .ZN(
        n14260) );
  NAND2_X1 U17881 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14258) );
  AOI221_X1 U17882 ( .B1(n14262), .B2(n14468), .C1(n14258), .C2(n14468), .A(
        n15562), .ZN(n14259) );
  AOI211_X1 U17883 ( .C1(n14435), .C2(n17429), .A(n14260), .B(n14259), .ZN(
        n14266) );
  AOI21_X1 U17884 ( .B1(n14261), .B2(n17401), .A(n14465), .ZN(n14264) );
  NAND2_X1 U17885 ( .A1(n15565), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14263) );
  MUX2_X1 U17886 ( .A(n14264), .B(n14263), .S(n14262), .Z(n14265) );
  NAND2_X1 U17887 ( .A1(n14266), .A2(n14265), .ZN(P1_U3029) );
  XOR2_X1 U17888 ( .A(n14267), .B(n14268), .Z(n19826) );
  XNOR2_X1 U17889 ( .A(n16813), .B(n19826), .ZN(n14272) );
  AOI22_X1 U17890 ( .A1(n19899), .A2(n19826), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19898), .ZN(n14271) );
  INV_X1 U17891 ( .A(n19907), .ZN(n16180) );
  NAND2_X1 U17892 ( .A1(n16180), .A2(n19867), .ZN(n14270) );
  OAI211_X1 U17893 ( .C1(n14272), .C2(n16164), .A(n14271), .B(n14270), .ZN(
        P2_U2919) );
  INV_X1 U17894 ( .A(n14276), .ZN(n14277) );
  INV_X1 U17895 ( .A(DATAI_6_), .ZN(n14280) );
  NAND2_X1 U17896 ( .A1(n20812), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14279) );
  OAI21_X1 U17897 ( .B1(n20812), .B2(n14280), .A(n14279), .ZN(n20846) );
  INV_X1 U17898 ( .A(n20846), .ZN(n14638) );
  NOR2_X1 U17899 ( .A1(n14383), .A2(n14638), .ZN(n14289) );
  AOI21_X1 U17900 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n20797), .A(n14289), 
        .ZN(n14281) );
  OAI21_X1 U17901 ( .B1(n14282), .B2(n14533), .A(n14281), .ZN(P1_U2943) );
  INV_X1 U17902 ( .A(DATAI_3_), .ZN(n14284) );
  NAND2_X1 U17903 ( .A1(n20812), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14283) );
  OAI21_X1 U17904 ( .B1(n20812), .B2(n14284), .A(n14283), .ZN(n20836) );
  INV_X1 U17905 ( .A(n20836), .ZN(n14414) );
  NOR2_X1 U17906 ( .A1(n14383), .A2(n14414), .ZN(n14307) );
  AOI21_X1 U17907 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n20797), .A(n14307), 
        .ZN(n14285) );
  OAI21_X1 U17908 ( .B1(n15152), .B2(n14533), .A(n14285), .ZN(P1_U2940) );
  INV_X1 U17909 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20769) );
  INV_X1 U17910 ( .A(DATAI_7_), .ZN(n14287) );
  NAND2_X1 U17911 ( .A1(n20812), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14286) );
  OAI21_X1 U17912 ( .B1(n20812), .B2(n14287), .A(n14286), .ZN(n20854) );
  INV_X1 U17913 ( .A(n20854), .ZN(n14637) );
  NOR2_X1 U17914 ( .A1(n14383), .A2(n14637), .ZN(n14312) );
  AOI21_X1 U17915 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n20797), .A(n14312), 
        .ZN(n14288) );
  OAI21_X1 U17916 ( .B1(n20769), .B2(n14533), .A(n14288), .ZN(P1_U2959) );
  AOI21_X1 U17917 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n20804), .A(n14289), 
        .ZN(n14290) );
  OAI21_X1 U17918 ( .B1(n12625), .B2(n14533), .A(n14290), .ZN(P1_U2958) );
  NOR2_X1 U17919 ( .A1(n14383), .A2(n20829), .ZN(n14302) );
  AOI21_X1 U17920 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n20804), .A(n14302), 
        .ZN(n14291) );
  OAI21_X1 U17921 ( .B1(n14292), .B2(n14533), .A(n14291), .ZN(P1_U2938) );
  NOR2_X1 U17922 ( .A1(n14383), .A2(n14293), .ZN(n14300) );
  AOI21_X1 U17923 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n20804), .A(n14300), 
        .ZN(n14294) );
  OAI21_X1 U17924 ( .B1(n14295), .B2(n14533), .A(n14294), .ZN(P1_U2937) );
  INV_X1 U17925 ( .A(DATAI_11_), .ZN(n14297) );
  NAND2_X1 U17926 ( .A1(n20812), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14296) );
  OAI21_X1 U17927 ( .B1(n20812), .B2(n14297), .A(n14296), .ZN(n20794) );
  AOI22_X1 U17928 ( .A1(n20807), .A2(n20794), .B1(P1_UWORD_REG_11__SCAN_IN), 
        .B2(n20804), .ZN(n14298) );
  OAI21_X1 U17929 ( .B1(n14299), .B2(n14533), .A(n14298), .ZN(P1_U2948) );
  AOI21_X1 U17930 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n20804), .A(n14300), 
        .ZN(n14301) );
  OAI21_X1 U17931 ( .B1(n20787), .B2(n14533), .A(n14301), .ZN(P1_U2952) );
  AOI21_X1 U17932 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n20804), .A(n14302), 
        .ZN(n14303) );
  OAI21_X1 U17933 ( .B1(n20782), .B2(n14533), .A(n14303), .ZN(P1_U2953) );
  INV_X1 U17934 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20780) );
  INV_X1 U17935 ( .A(DATAI_2_), .ZN(n14305) );
  NAND2_X1 U17936 ( .A1(n20812), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14304) );
  OAI21_X1 U17937 ( .B1(n20812), .B2(n14305), .A(n14304), .ZN(n20833) );
  INV_X1 U17938 ( .A(n20833), .ZN(n14456) );
  NOR2_X1 U17939 ( .A1(n14383), .A2(n14456), .ZN(n14309) );
  AOI21_X1 U17940 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n20804), .A(n14309), 
        .ZN(n14306) );
  OAI21_X1 U17941 ( .B1(n20780), .B2(n14533), .A(n14306), .ZN(P1_U2954) );
  INV_X1 U17942 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20778) );
  AOI21_X1 U17943 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n20804), .A(n14307), 
        .ZN(n14308) );
  OAI21_X1 U17944 ( .B1(n20778), .B2(n14533), .A(n14308), .ZN(P1_U2955) );
  AOI21_X1 U17945 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n20804), .A(n14309), 
        .ZN(n14310) );
  OAI21_X1 U17946 ( .B1(n14311), .B2(n14533), .A(n14310), .ZN(P1_U2939) );
  AOI21_X1 U17947 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n20797), .A(n14312), 
        .ZN(n14313) );
  OAI21_X1 U17948 ( .B1(n12901), .B2(n14533), .A(n14313), .ZN(P1_U2944) );
  INV_X1 U17949 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20776) );
  INV_X1 U17950 ( .A(DATAI_4_), .ZN(n14315) );
  NAND2_X1 U17951 ( .A1(n20812), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14314) );
  OAI21_X1 U17952 ( .B1(n20812), .B2(n14315), .A(n14314), .ZN(n20839) );
  INV_X1 U17953 ( .A(n20839), .ZN(n14547) );
  NOR2_X1 U17954 ( .A1(n14383), .A2(n14547), .ZN(n14331) );
  AOI21_X1 U17955 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n20804), .A(n14331), 
        .ZN(n14316) );
  OAI21_X1 U17956 ( .B1(n20776), .B2(n14533), .A(n14316), .ZN(P1_U2956) );
  INV_X1 U17957 ( .A(DATAI_9_), .ZN(n14318) );
  NAND2_X1 U17958 ( .A1(n20812), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14317) );
  OAI21_X1 U17959 ( .B1(n20812), .B2(n14318), .A(n14317), .ZN(n20788) );
  AOI22_X1 U17960 ( .A1(n20807), .A2(n20788), .B1(P1_UWORD_REG_9__SCAN_IN), 
        .B2(n20804), .ZN(n14319) );
  OAI21_X1 U17961 ( .B1(n15130), .B2(n14533), .A(n14319), .ZN(P1_U2946) );
  INV_X1 U17962 ( .A(DATAI_14_), .ZN(n14321) );
  NAND2_X1 U17963 ( .A1(n20812), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14320) );
  OAI21_X1 U17964 ( .B1(n20812), .B2(n14321), .A(n14320), .ZN(n20806) );
  AOI22_X1 U17965 ( .A1(n20807), .A2(n20806), .B1(P1_UWORD_REG_14__SCAN_IN), 
        .B2(n20804), .ZN(n14322) );
  OAI21_X1 U17966 ( .B1(n14323), .B2(n14533), .A(n14322), .ZN(P1_U2951) );
  INV_X1 U17967 ( .A(DATAI_13_), .ZN(n14325) );
  NAND2_X1 U17968 ( .A1(n20812), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14324) );
  OAI21_X1 U17969 ( .B1(n20812), .B2(n14325), .A(n14324), .ZN(n20801) );
  AOI22_X1 U17970 ( .A1(n20807), .A2(n20801), .B1(P1_UWORD_REG_13__SCAN_IN), 
        .B2(n20804), .ZN(n14326) );
  OAI21_X1 U17971 ( .B1(n14327), .B2(n14533), .A(n14326), .ZN(P1_U2950) );
  INV_X1 U17972 ( .A(DATAI_10_), .ZN(n14329) );
  NAND2_X1 U17973 ( .A1(n20812), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14328) );
  OAI21_X1 U17974 ( .B1(n20812), .B2(n14329), .A(n14328), .ZN(n20791) );
  AOI22_X1 U17975 ( .A1(n20807), .A2(n20791), .B1(P1_UWORD_REG_10__SCAN_IN), 
        .B2(n20797), .ZN(n14330) );
  OAI21_X1 U17976 ( .B1(n15125), .B2(n14533), .A(n14330), .ZN(P1_U2947) );
  AOI21_X1 U17977 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n20804), .A(n14331), 
        .ZN(n14332) );
  OAI21_X1 U17978 ( .B1(n14333), .B2(n14533), .A(n14332), .ZN(P1_U2941) );
  INV_X1 U17979 ( .A(DATAI_12_), .ZN(n14335) );
  NAND2_X1 U17980 ( .A1(n20812), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14334) );
  OAI21_X1 U17981 ( .B1(n20812), .B2(n14335), .A(n14334), .ZN(n20798) );
  AOI22_X1 U17982 ( .A1(n20807), .A2(n20798), .B1(P1_UWORD_REG_12__SCAN_IN), 
        .B2(n20804), .ZN(n14336) );
  OAI21_X1 U17983 ( .B1(n14337), .B2(n14533), .A(n14336), .ZN(P1_U2949) );
  INV_X1 U17984 ( .A(DATAI_8_), .ZN(n14339) );
  NAND2_X1 U17985 ( .A1(n20812), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14338) );
  OAI21_X1 U17986 ( .B1(n20812), .B2(n14339), .A(n14338), .ZN(n15136) );
  NAND2_X1 U17987 ( .A1(n20807), .A2(n15136), .ZN(n14534) );
  NAND2_X1 U17988 ( .A1(n20797), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14340) );
  OAI211_X1 U17989 ( .C1(n14533), .C2(n14341), .A(n14534), .B(n14340), .ZN(
        P1_U2945) );
  INV_X1 U17990 ( .A(DATAI_5_), .ZN(n14343) );
  NAND2_X1 U17991 ( .A1(n20812), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14342) );
  OAI21_X1 U17992 ( .B1(n20812), .B2(n14343), .A(n14342), .ZN(n20843) );
  NAND2_X1 U17993 ( .A1(n20807), .A2(n20843), .ZN(n14346) );
  NAND2_X1 U17994 ( .A1(n20797), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14344) );
  OAI211_X1 U17995 ( .C1(n14533), .C2(n21454), .A(n14346), .B(n14344), .ZN(
        P1_U2942) );
  INV_X1 U17996 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20773) );
  NAND2_X1 U17997 ( .A1(n20797), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n14345) );
  OAI211_X1 U17998 ( .C1(n14533), .C2(n20773), .A(n14346), .B(n14345), .ZN(
        P1_U2957) );
  INV_X1 U17999 ( .A(n14702), .ZN(n16767) );
  OR2_X1 U18000 ( .A1(n16733), .A2(n16767), .ZN(n14357) );
  NAND2_X1 U18001 ( .A1(n11484), .A2(n11470), .ZN(n16762) );
  INV_X1 U18002 ( .A(n16757), .ZN(n14347) );
  NAND2_X1 U18003 ( .A1(n16759), .A2(n14347), .ZN(n14349) );
  NAND2_X1 U18004 ( .A1(n14348), .A2(n10958), .ZN(n16756) );
  NAND2_X1 U18005 ( .A1(n14349), .A2(n16756), .ZN(n14350) );
  AOI21_X1 U18006 ( .B1(n16762), .B2(n16755), .A(n14350), .ZN(n14355) );
  INV_X1 U18007 ( .A(n14351), .ZN(n16846) );
  NAND2_X1 U18008 ( .A1(n16846), .A2(n16845), .ZN(n16764) );
  NAND2_X1 U18009 ( .A1(n16759), .A2(n16757), .ZN(n14352) );
  NAND2_X1 U18010 ( .A1(n14352), .A2(n16755), .ZN(n14353) );
  AOI21_X1 U18011 ( .B1(n16764), .B2(n16756), .A(n14353), .ZN(n14354) );
  MUX2_X1 U18012 ( .A(n14355), .B(n14354), .S(n10635), .Z(n14356) );
  NAND2_X1 U18013 ( .A1(n14357), .A2(n14356), .ZN(n16841) );
  AOI22_X1 U18014 ( .A1(n20610), .A2(n16883), .B1(n19730), .B2(n16841), .ZN(
        n14367) );
  NAND2_X1 U18015 ( .A1(n14359), .A2(n14358), .ZN(n14364) );
  AND3_X1 U18016 ( .A1(n14362), .A2(n14361), .A3(n14360), .ZN(n14363) );
  NAND2_X1 U18017 ( .A1(n16863), .A2(n16899), .ZN(n14366) );
  AOI22_X1 U18018 ( .A1(n16904), .A2(P2_FLUSH_REG_SCAN_IN), .B1(n16902), .B2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14365) );
  MUX2_X1 U18019 ( .A(n14367), .B(n10543), .S(n16773), .Z(n14368) );
  INV_X1 U18020 ( .A(n14368), .ZN(P2_U3596) );
  AND2_X1 U18021 ( .A1(n14369), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n16175) );
  XOR2_X1 U18022 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n16179), .Z(n14379)
         );
  NAND2_X1 U18023 ( .A1(n14373), .A2(n14374), .ZN(n14375) );
  INV_X1 U18024 ( .A(n19800), .ZN(n14377) );
  MUX2_X1 U18025 ( .A(n14377), .B(n14376), .S(n16065), .Z(n14378) );
  OAI21_X1 U18026 ( .B1(n14379), .B2(n19855), .A(n14378), .ZN(P2_U2882) );
  INV_X1 U18027 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14384) );
  INV_X1 U18028 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20753) );
  INV_X1 U18029 ( .A(DATAI_15_), .ZN(n14381) );
  NAND2_X1 U18030 ( .A1(n20812), .A2(BUF1_REG_15__SCAN_IN), .ZN(n14380) );
  OAI21_X1 U18031 ( .B1(n20812), .B2(n14381), .A(n14380), .ZN(n15170) );
  INV_X1 U18032 ( .A(n15170), .ZN(n14382) );
  OAI222_X1 U18033 ( .A1(n14533), .A2(n14384), .B1(n14536), .B2(n20753), .C1(
        n14383), .C2(n14382), .ZN(P1_U2967) );
  NAND2_X1 U18034 ( .A1(n19709), .A2(n14385), .ZN(n19581) );
  INV_X1 U18035 ( .A(n19581), .ZN(n14387) );
  AOI21_X1 U18036 ( .B1(n14389), .B2(n19547), .A(n14388), .ZN(n14390) );
  INV_X1 U18037 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19097) );
  NOR3_X1 U18038 ( .A1(n19592), .A2(n19591), .A3(n19582), .ZN(n19599) );
  INV_X1 U18039 ( .A(n19599), .ZN(n19688) );
  NOR2_X1 U18040 ( .A1(n19097), .A2(n19688), .ZN(n14393) );
  INV_X1 U18041 ( .A(n14394), .ZN(n17154) );
  NAND2_X1 U18042 ( .A1(n17154), .A2(n9940), .ZN(n17164) );
  NAND2_X1 U18043 ( .A1(n17164), .A2(n18916), .ZN(n14397) );
  NOR2_X1 U18044 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18914), .ZN(
        n17147) );
  INV_X1 U18045 ( .A(n17147), .ZN(n14395) );
  NAND2_X1 U18046 ( .A1(n14401), .A2(n14395), .ZN(n14396) );
  AOI21_X1 U18047 ( .B1(n14397), .B2(n14396), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19554) );
  INV_X1 U18048 ( .A(n19554), .ZN(n14403) );
  NAND2_X1 U18049 ( .A1(n14401), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17163) );
  OAI21_X1 U18050 ( .B1(n14400), .B2(n14399), .A(n14398), .ZN(n17156) );
  OAI21_X1 U18051 ( .B1(n14401), .B2(n18877), .A(n17164), .ZN(n14402) );
  AOI21_X1 U18052 ( .B1(n17163), .B2(n17156), .A(n14402), .ZN(n19552) );
  OAI22_X1 U18053 ( .A1(n17178), .A2(n14403), .B1(n19552), .B2(n14407), .ZN(
        n14404) );
  NAND2_X1 U18054 ( .A1(n14404), .A2(n17540), .ZN(n14406) );
  AOI21_X1 U18055 ( .B1(n14407), .B2(n17163), .A(n17208), .ZN(n17885) );
  NAND3_X1 U18056 ( .A1(n17174), .A2(n19578), .A3(n17885), .ZN(n14405) );
  OAI211_X1 U18057 ( .C1(n17174), .C2(n14407), .A(n14406), .B(n14405), .ZN(
        P3_U3285) );
  NAND2_X1 U18058 ( .A1(n14411), .A2(n14410), .ZN(n14412) );
  NAND2_X1 U18059 ( .A1(n14409), .A2(n14412), .ZN(n14413) );
  NAND2_X1 U18060 ( .A1(n14408), .A2(n14413), .ZN(n20743) );
  OAI222_X1 U18061 ( .A1(n20743), .A2(n15182), .B1(n14639), .B2(n14414), .C1(
        n15151), .C2(n20778), .ZN(P1_U2901) );
  NOR2_X1 U18062 ( .A1(n16179), .A2(n20010), .ZN(n14416) );
  OAI211_X1 U18063 ( .C1(n14416), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19863), .B(n14594), .ZN(n14422) );
  NAND2_X1 U18064 ( .A1(n14371), .A2(n14418), .ZN(n14419) );
  NAND2_X1 U18065 ( .A1(n14417), .A2(n14419), .ZN(n16703) );
  MUX2_X1 U18066 ( .A(n16703), .B(n14420), .S(n16065), .Z(n14421) );
  NAND2_X1 U18067 ( .A1(n14422), .A2(n14421), .ZN(P2_U2881) );
  NAND2_X1 U18068 ( .A1(n14424), .A2(n14423), .ZN(n14425) );
  NOR2_X1 U18069 ( .A1(n14426), .A2(n14425), .ZN(n14428) );
  MUX2_X1 U18070 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(n14428), .S(n14427), .Z(n14429) );
  XNOR2_X1 U18071 ( .A(n14430), .B(n14429), .ZN(n15069) );
  INV_X1 U18072 ( .A(n14431), .ZN(n15061) );
  AOI22_X1 U18073 ( .A1(n15104), .A2(n15061), .B1(n13660), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14432) );
  OAI21_X1 U18074 ( .B1(n15069), .B2(n15111), .A(n14432), .ZN(P1_U2870) );
  AOI22_X1 U18075 ( .A1(n17370), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n17416), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14433) );
  OAI21_X1 U18076 ( .B1(n15065), .B2(n17377), .A(n14433), .ZN(n14434) );
  AOI21_X1 U18077 ( .B1(n14435), .B2(n17382), .A(n14434), .ZN(n14436) );
  OAI21_X1 U18078 ( .B1(n15069), .B2(n20811), .A(n14436), .ZN(P1_U2997) );
  OR2_X1 U18079 ( .A1(n20079), .A2(n16786), .ZN(n20609) );
  INV_X1 U18080 ( .A(n20609), .ZN(n14444) );
  NAND2_X1 U18081 ( .A1(n14438), .A2(n14437), .ZN(n20608) );
  OR2_X1 U18082 ( .A1(n14440), .A2(n14439), .ZN(n14441) );
  NAND2_X1 U18083 ( .A1(n14442), .A2(n14441), .ZN(n19890) );
  INV_X1 U18084 ( .A(n19890), .ZN(n19950) );
  OAI22_X1 U18085 ( .A1(n16799), .A2(n20608), .B1(n19950), .B2(n16814), .ZN(
        n14443) );
  OAI21_X1 U18086 ( .B1(n14444), .B2(n14443), .A(n20626), .ZN(n14445) );
  OAI21_X1 U18087 ( .B1(n20626), .B2(n16860), .A(n14445), .ZN(P2_U3603) );
  NAND2_X1 U18088 ( .A1(n14447), .A2(n14446), .ZN(n14448) );
  NAND2_X1 U18089 ( .A1(n14527), .A2(n14448), .ZN(n20733) );
  INV_X1 U18090 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14449) );
  OAI222_X1 U18091 ( .A1(n20733), .A2(n15114), .B1(n14449), .B2(n15113), .C1(
        n20743), .C2(n15111), .ZN(P1_U2869) );
  NOR2_X1 U18092 ( .A1(n14450), .A2(n18973), .ZN(n17146) );
  MUX2_X1 U18093 ( .A(n18877), .B(n17146), .S(n14453), .Z(n19559) );
  INV_X1 U18094 ( .A(n17540), .ZN(n19719) );
  NAND2_X1 U18095 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n10220), .ZN(n14451) );
  OAI211_X1 U18096 ( .C1(n19559), .C2(n19719), .A(n17174), .B(n14451), .ZN(
        n14452) );
  OAI21_X1 U18097 ( .B1(n17174), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n14452), .ZN(n14455) );
  NAND3_X1 U18098 ( .A1(n17174), .A2(n19578), .A3(n14453), .ZN(n14454) );
  NAND2_X1 U18099 ( .A1(n14455), .A2(n14454), .ZN(P3_U3290) );
  OAI222_X1 U18100 ( .A1(n15182), .A2(n15069), .B1(n14639), .B2(n14456), .C1(
        n15151), .C2(n20780), .ZN(P1_U2902) );
  XOR2_X1 U18101 ( .A(n14594), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n14462)
         );
  AND2_X1 U18102 ( .A1(n14417), .A2(n14457), .ZN(n14459) );
  OR2_X1 U18103 ( .A1(n14459), .A2(n14458), .ZN(n16407) );
  MUX2_X1 U18104 ( .A(n16407), .B(n14460), .S(n16065), .Z(n14461) );
  OAI21_X1 U18105 ( .B1(n14462), .B2(n19855), .A(n14461), .ZN(P2_U2880) );
  XNOR2_X1 U18106 ( .A(n9761), .B(n14471), .ZN(n14464) );
  XNOR2_X1 U18107 ( .A(n14464), .B(n14463), .ZN(n14521) );
  INV_X1 U18108 ( .A(n14467), .ZN(n17402) );
  AOI21_X1 U18109 ( .B1(n17401), .B2(n17402), .A(n14465), .ZN(n14466) );
  OAI21_X1 U18110 ( .B1(n15562), .B2(n14468), .A(n14466), .ZN(n14531) );
  NAND2_X1 U18111 ( .A1(n15565), .A2(n14467), .ZN(n17403) );
  NAND2_X1 U18112 ( .A1(n14469), .A2(n14468), .ZN(n14470) );
  NAND2_X1 U18113 ( .A1(n17403), .A2(n14470), .ZN(n17422) );
  AOI22_X1 U18114 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14531), .B1(
        n17422), .B2(n14471), .ZN(n14472) );
  OR2_X1 U18115 ( .A1(n20716), .A2(n20739), .ZN(n14522) );
  OAI211_X1 U18116 ( .C1(n17390), .C2(n20733), .A(n14472), .B(n14522), .ZN(
        n14473) );
  AOI21_X1 U18117 ( .B1(n14521), .B2(n17429), .A(n14473), .ZN(n14474) );
  INV_X1 U18118 ( .A(n14474), .ZN(P1_U3028) );
  AOI22_X1 U18119 ( .A1(n19927), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14476) );
  OAI21_X1 U18120 ( .B1(n14477), .B2(n19910), .A(n14476), .ZN(P2_U2922) );
  NOR2_X1 U18121 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21357), .ZN(n14496) );
  MUX2_X1 U18122 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14479), .S(
        n17324), .Z(n17320) );
  AOI22_X1 U18123 ( .A1(n14496), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21357), .B2(n17320), .ZN(n14498) );
  INV_X1 U18124 ( .A(n14087), .ZN(n15624) );
  AOI211_X1 U18125 ( .C1(n15642), .C2(n15624), .A(n14481), .B(n11874), .ZN(
        n15637) );
  NOR2_X1 U18126 ( .A1(n14482), .A2(n15637), .ZN(n14494) );
  NAND2_X1 U18127 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14484) );
  INV_X1 U18128 ( .A(n14484), .ZN(n14483) );
  MUX2_X1 U18129 ( .A(n14484), .B(n14483), .S(n15642), .Z(n14492) );
  INV_X1 U18130 ( .A(n14485), .ZN(n14489) );
  MUX2_X1 U18131 ( .A(n14487), .B(n14486), .S(n14087), .Z(n14488) );
  NAND3_X1 U18132 ( .A1(n14490), .A2(n14489), .A3(n14488), .ZN(n14491) );
  OAI21_X1 U18133 ( .B1(n17323), .B2(n14492), .A(n14491), .ZN(n14493) );
  AOI211_X1 U18134 ( .C1(n21063), .C2(n15628), .A(n14494), .B(n14493), .ZN(
        n15639) );
  NOR2_X1 U18135 ( .A1(n17324), .A2(n15642), .ZN(n14495) );
  AOI21_X1 U18136 ( .B1(n15639), .B2(n17324), .A(n14495), .ZN(n17334) );
  AOI22_X1 U18137 ( .A1(n14496), .A2(n15642), .B1(n17334), .B2(n21357), .ZN(
        n14497) );
  NOR2_X1 U18138 ( .A1(n14498), .A2(n14497), .ZN(n17344) );
  INV_X1 U18139 ( .A(n11829), .ZN(n15625) );
  NAND2_X1 U18140 ( .A1(n17344), .A2(n15625), .ZN(n15620) );
  NAND3_X1 U18141 ( .A1(n20715), .A2(n14499), .A3(n14500), .ZN(n14503) );
  INV_X1 U18142 ( .A(n14500), .ZN(n14501) );
  NAND3_X1 U18143 ( .A1(n14501), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n20647), .ZN(n14502) );
  NAND2_X1 U18144 ( .A1(n14503), .A2(n14502), .ZN(n17343) );
  INV_X1 U18145 ( .A(n17343), .ZN(n15619) );
  NAND3_X1 U18146 ( .A1(n15620), .A2(n15619), .A3(n20647), .ZN(n14506) );
  INV_X1 U18147 ( .A(n17440), .ZN(n14505) );
  INV_X1 U18148 ( .A(n20810), .ZN(n14698) );
  NAND2_X1 U18149 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21197), .ZN(n15621) );
  NAND2_X1 U18150 ( .A1(n14698), .A2(n15621), .ZN(n14693) );
  NOR2_X1 U18151 ( .A1(n14508), .A2(n21397), .ZN(n20862) );
  AOI21_X1 U18152 ( .B1(n14508), .B2(n21397), .A(n20862), .ZN(n14509) );
  NOR3_X1 U18153 ( .A1(n20810), .A2(n14509), .A3(n21302), .ZN(n14510) );
  AOI21_X1 U18154 ( .B1(n20810), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n14510), .ZN(n14511) );
  OAI21_X1 U18155 ( .B1(n21065), .B2(n14693), .A(n14511), .ZN(P1_U3477) );
  AOI22_X1 U18156 ( .A1(n19927), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14512) );
  OAI21_X1 U18157 ( .B1(n14513), .B2(n19910), .A(n14512), .ZN(P2_U2924) );
  AOI22_X1 U18158 ( .A1(n19927), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14514) );
  OAI21_X1 U18159 ( .B1(n14515), .B2(n19910), .A(n14514), .ZN(P2_U2921) );
  AOI22_X1 U18160 ( .A1(n19927), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14516) );
  OAI21_X1 U18161 ( .B1(n14517), .B2(n19910), .A(n14516), .ZN(P2_U2934) );
  AOI22_X1 U18162 ( .A1(n19927), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14518) );
  OAI21_X1 U18163 ( .B1(n14519), .B2(n19910), .A(n14518), .ZN(P2_U2923) );
  AOI22_X1 U18164 ( .A1(n19927), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n14520) );
  OAI21_X1 U18165 ( .B1(n13996), .B2(n19910), .A(n14520), .ZN(P2_U2935) );
  NAND2_X1 U18166 ( .A1(n14521), .A2(n17382), .ZN(n14525) );
  OAI21_X1 U18167 ( .B1(n17385), .B2(n21447), .A(n14522), .ZN(n14523) );
  AOI21_X1 U18168 ( .B1(n17379), .B2(n20732), .A(n14523), .ZN(n14524) );
  OAI211_X1 U18169 ( .C1(n20811), .C2(n20743), .A(n14525), .B(n14524), .ZN(
        P1_U2996) );
  INV_X1 U18170 ( .A(n14527), .ZN(n14528) );
  OAI21_X1 U18171 ( .B1(n14528), .B2(n9788), .A(n9774), .ZN(n20713) );
  OAI211_X1 U18172 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n17422), .B(n17400), .ZN(n14529) );
  OR2_X1 U18173 ( .A1(n20716), .A2(n20727), .ZN(n14538) );
  OAI211_X1 U18174 ( .C1(n17390), .C2(n20713), .A(n14529), .B(n14538), .ZN(
        n14530) );
  AOI21_X1 U18175 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14531), .A(
        n14530), .ZN(n14532) );
  OAI21_X1 U18176 ( .B1(n17397), .B2(n14546), .A(n14532), .ZN(P1_U3027) );
  INV_X1 U18177 ( .A(P1_LWORD_REG_8__SCAN_IN), .ZN(n21527) );
  NAND2_X1 U18178 ( .A1(n20805), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n14535) );
  OAI211_X1 U18179 ( .C1(n14536), .C2(n21527), .A(n14535), .B(n14534), .ZN(
        P1_U2960) );
  INV_X1 U18180 ( .A(n14537), .ZN(n20720) );
  INV_X1 U18181 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14539) );
  OAI21_X1 U18182 ( .B1(n17385), .B2(n14539), .A(n14538), .ZN(n14540) );
  AOI21_X1 U18183 ( .B1(n17379), .B2(n20720), .A(n14540), .ZN(n14545) );
  AND2_X1 U18184 ( .A1(n14408), .A2(n14542), .ZN(n14543) );
  NOR2_X1 U18185 ( .A1(n14541), .A2(n14543), .ZN(n20724) );
  NAND2_X1 U18186 ( .A1(n20724), .A2(n17381), .ZN(n14544) );
  OAI211_X1 U18187 ( .C1(n14546), .C2(n20646), .A(n14545), .B(n14544), .ZN(
        P1_U2995) );
  INV_X1 U18188 ( .A(n20724), .ZN(n14559) );
  OAI222_X1 U18189 ( .A1(n14559), .A2(n15182), .B1(n14639), .B2(n14547), .C1(
        n15151), .C2(n20776), .ZN(P1_U2900) );
  OAI21_X1 U18190 ( .B1(n14548), .B2(n14550), .A(n14549), .ZN(n16653) );
  AOI22_X1 U18191 ( .A1(n16180), .A2(n16095), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19898), .ZN(n14551) );
  OAI21_X1 U18192 ( .B1(n16653), .B2(n16183), .A(n14551), .ZN(P2_U2909) );
  OR2_X1 U18193 ( .A1(n14541), .A2(n14553), .ZN(n14554) );
  AND2_X1 U18194 ( .A1(n14552), .A2(n14554), .ZN(n20709) );
  INV_X1 U18195 ( .A(n20709), .ZN(n14558) );
  INV_X1 U18196 ( .A(n14555), .ZN(n14629) );
  AOI21_X1 U18197 ( .B1(n9785), .B2(n9774), .A(n14629), .ZN(n20707) );
  AOI22_X1 U18198 ( .A1(n20707), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n14556) );
  OAI21_X1 U18199 ( .B1(n14558), .B2(n15101), .A(n14556), .ZN(P1_U2867) );
  AOI22_X1 U18200 ( .A1(n15180), .A2(n20843), .B1(P1_EAX_REG_5__SCAN_IN), .B2(
        n15179), .ZN(n14557) );
  OAI21_X1 U18201 ( .B1(n14558), .B2(n15182), .A(n14557), .ZN(P1_U2899) );
  INV_X1 U18202 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14560) );
  OAI222_X1 U18203 ( .A1(n20713), .A2(n15114), .B1(n14560), .B2(n15113), .C1(
        n14559), .C2(n15111), .ZN(P1_U2868) );
  NAND2_X1 U18204 ( .A1(n14561), .A2(n14562), .ZN(n14563) );
  NAND2_X1 U18205 ( .A1(n9617), .A2(n14563), .ZN(n16681) );
  INV_X1 U18206 ( .A(n16109), .ZN(n14564) );
  OAI222_X1 U18207 ( .A1(n16681), .A2(n16183), .B1(n14644), .B2(n14070), .C1(
        n19907), .C2(n14564), .ZN(P2_U2911) );
  AOI21_X1 U18208 ( .B1(n14565), .B2(n9617), .A(n14548), .ZN(n19785) );
  INV_X1 U18209 ( .A(n19785), .ZN(n14567) );
  INV_X1 U18210 ( .A(n16102), .ZN(n14566) );
  OAI222_X1 U18211 ( .A1(n14567), .A2(n16183), .B1(n14644), .B2(n14076), .C1(
        n19907), .C2(n14566), .ZN(P2_U2910) );
  NAND2_X1 U18212 ( .A1(n14549), .A2(n14569), .ZN(n14570) );
  NAND2_X1 U18213 ( .A1(n14568), .A2(n14570), .ZN(n19755) );
  INV_X1 U18214 ( .A(n16088), .ZN(n14571) );
  OAI222_X1 U18215 ( .A1(n19755), .A2(n16183), .B1(n14571), .B2(n19907), .C1(
        n14036), .C2(n14644), .ZN(P2_U2908) );
  AOI21_X1 U18216 ( .B1(n14572), .B2(n14568), .A(n9599), .ZN(n16628) );
  INV_X1 U18217 ( .A(n16628), .ZN(n14574) );
  INV_X1 U18218 ( .A(n16081), .ZN(n14573) );
  OAI222_X1 U18219 ( .A1(n14574), .A2(n16183), .B1(n14644), .B2(n14026), .C1(
        n19907), .C2(n14573), .ZN(P2_U2907) );
  OAI21_X1 U18220 ( .B1(n14576), .B2(n14575), .A(n14561), .ZN(n16689) );
  INV_X1 U18221 ( .A(n20026), .ZN(n14577) );
  OAI222_X1 U18222 ( .A1(n16689), .A2(n16183), .B1(n19924), .B2(n14644), .C1(
        n19907), .C2(n14577), .ZN(P2_U2912) );
  CLKBUF_X1 U18223 ( .A(n14578), .Z(n14587) );
  NOR2_X1 U18224 ( .A1(n9599), .A2(n14579), .ZN(n14580) );
  OR2_X1 U18225 ( .A1(n14587), .A2(n14580), .ZN(n16614) );
  INV_X1 U18226 ( .A(n16074), .ZN(n14581) );
  OAI222_X1 U18227 ( .A1(n16614), .A2(n16183), .B1(n14581), .B2(n19907), .C1(
        n14022), .C2(n14644), .ZN(P2_U2906) );
  XOR2_X1 U18228 ( .A(n14582), .B(n14583), .Z(n16708) );
  INV_X1 U18229 ( .A(n16708), .ZN(n15932) );
  INV_X1 U18230 ( .A(n20016), .ZN(n14584) );
  OAI222_X1 U18231 ( .A1(n15932), .A2(n16183), .B1(n19926), .B2(n14644), .C1(
        n19907), .C2(n14584), .ZN(P2_U2913) );
  OAI21_X1 U18232 ( .B1(n14587), .B2(n14586), .A(n14585), .ZN(n16599) );
  AOI22_X1 U18233 ( .A1(n16180), .A2(n14588), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19898), .ZN(n14589) );
  OAI21_X1 U18234 ( .B1(n16599), .B2(n16183), .A(n14589), .ZN(P2_U2905) );
  OR2_X1 U18235 ( .A1(n14458), .A2(n14590), .ZN(n14592) );
  INV_X1 U18236 ( .A(n16678), .ZN(n14599) );
  NOR2_X1 U18237 ( .A1(n14594), .A2(n14593), .ZN(n14596) );
  NAND2_X1 U18238 ( .A1(n14596), .A2(n14595), .ZN(n16054) );
  OAI211_X1 U18239 ( .C1(n14596), .C2(n14595), .A(n16054), .B(n19863), .ZN(
        n14598) );
  NAND2_X1 U18240 ( .A1(n16065), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14597) );
  OAI211_X1 U18241 ( .C1(n14599), .C2(n16065), .A(n14598), .B(n14597), .ZN(
        P2_U2879) );
  INV_X1 U18242 ( .A(n14600), .ZN(n16053) );
  XNOR2_X1 U18243 ( .A(n16054), .B(n16053), .ZN(n14604) );
  INV_X1 U18244 ( .A(n14601), .ZN(n15890) );
  AOI21_X1 U18245 ( .B1(n14602), .B2(n14591), .A(n14601), .ZN(n16667) );
  INV_X1 U18246 ( .A(n16667), .ZN(n19777) );
  MUX2_X1 U18247 ( .A(n19772), .B(n19777), .S(n19866), .Z(n14603) );
  OAI21_X1 U18248 ( .B1(n14604), .B2(n19855), .A(n14603), .ZN(P2_U2878) );
  INV_X1 U18249 ( .A(n14605), .ZN(n14606) );
  NOR2_X1 U18250 ( .A1(n16179), .A2(n14606), .ZN(n16056) );
  XNOR2_X1 U18251 ( .A(n16056), .B(n14616), .ZN(n14612) );
  NAND2_X1 U18252 ( .A1(n14607), .A2(n14608), .ZN(n14609) );
  AND2_X1 U18253 ( .A1(n9746), .A2(n14609), .ZN(n16611) );
  NOR2_X1 U18254 ( .A1(n19866), .A2(n15862), .ZN(n14610) );
  AOI21_X1 U18255 ( .B1(n16611), .B2(n19866), .A(n14610), .ZN(n14611) );
  OAI21_X1 U18256 ( .B1(n14612), .B2(n19855), .A(n14611), .ZN(P2_U2874) );
  AND2_X1 U18257 ( .A1(n9746), .A2(n14613), .ZN(n14615) );
  OR2_X1 U18258 ( .A1(n14615), .A2(n14614), .ZN(n16601) );
  NAND2_X1 U18259 ( .A1(n16056), .A2(n14616), .ZN(n14618) );
  INV_X1 U18260 ( .A(n14618), .ZN(n14621) );
  INV_X1 U18261 ( .A(n14620), .ZN(n14617) );
  NOR2_X1 U18262 ( .A1(n14618), .A2(n14617), .ZN(n19848) );
  INV_X1 U18263 ( .A(n19848), .ZN(n14619) );
  OAI211_X1 U18264 ( .C1(n14621), .C2(n14620), .A(n14619), .B(n19863), .ZN(
        n14623) );
  NAND2_X1 U18265 ( .A1(n16065), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14622) );
  OAI211_X1 U18266 ( .C1(n16601), .C2(n16065), .A(n14623), .B(n14622), .ZN(
        P2_U2873) );
  AND2_X1 U18267 ( .A1(n14625), .A2(n14624), .ZN(n14627) );
  OR2_X1 U18268 ( .A1(n14627), .A2(n14626), .ZN(n17367) );
  AOI21_X1 U18269 ( .B1(n14629), .B2(n14635), .A(n14628), .ZN(n14631) );
  INV_X1 U18270 ( .A(n15050), .ZN(n14630) );
  NOR2_X1 U18271 ( .A1(n14631), .A2(n14630), .ZN(n20678) );
  AOI22_X1 U18272 ( .A1(n20678), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n14632) );
  OAI21_X1 U18273 ( .B1(n17367), .B2(n15101), .A(n14632), .ZN(P1_U2865) );
  INV_X1 U18274 ( .A(n14624), .ZN(n14633) );
  AOI21_X1 U18275 ( .B1(n14634), .B2(n14552), .A(n14633), .ZN(n20697) );
  INV_X1 U18276 ( .A(n20697), .ZN(n14640) );
  XNOR2_X1 U18277 ( .A(n14555), .B(n14635), .ZN(n20689) );
  AOI22_X1 U18278 ( .A1(n20689), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n14636) );
  OAI21_X1 U18279 ( .B1(n14640), .B2(n15111), .A(n14636), .ZN(P1_U2866) );
  OAI222_X1 U18280 ( .A1(n17367), .A2(n15182), .B1(n14639), .B2(n14637), .C1(
        n20769), .C2(n15151), .ZN(P1_U2897) );
  OAI222_X1 U18281 ( .A1(n14640), .A2(n15182), .B1(n14639), .B2(n14638), .C1(
        n15151), .C2(n12625), .ZN(P1_U2898) );
  NAND2_X1 U18282 ( .A1(n14585), .A2(n14641), .ZN(n14642) );
  AND2_X1 U18283 ( .A1(n15830), .A2(n14642), .ZN(n16588) );
  INV_X1 U18284 ( .A(n16588), .ZN(n14645) );
  OAI222_X1 U18285 ( .A1(n14645), .A2(n16183), .B1(n14644), .B2(n13927), .C1(
        n14643), .C2(n19907), .ZN(P2_U2904) );
  INV_X1 U18286 ( .A(n14626), .ZN(n14647) );
  AOI21_X1 U18287 ( .B1(n9775), .B2(n14647), .A(n14646), .ZN(n15385) );
  INV_X1 U18288 ( .A(n15385), .ZN(n15110) );
  AOI22_X1 U18289 ( .A1(n15180), .A2(n15136), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15179), .ZN(n14648) );
  OAI21_X1 U18290 ( .B1(n15110), .B2(n15182), .A(n14648), .ZN(P1_U2896) );
  OAI21_X1 U18291 ( .B1(n14646), .B2(n14650), .A(n14649), .ZN(n20668) );
  NOR2_X1 U18292 ( .A1(n14651), .A2(n14652), .ZN(n14653) );
  OR2_X1 U18293 ( .A1(n15037), .A2(n14653), .ZN(n15604) );
  INV_X1 U18294 ( .A(n15604), .ZN(n20667) );
  AOI22_X1 U18295 ( .A1(n20667), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n14654) );
  OAI21_X1 U18296 ( .B1(n20668), .B2(n15111), .A(n14654), .ZN(P1_U2863) );
  AOI22_X1 U18297 ( .A1(n15180), .A2(n20788), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15179), .ZN(n14655) );
  OAI21_X1 U18298 ( .B1(n20668), .B2(n15182), .A(n14655), .ZN(P1_U2895) );
  NOR2_X1 U18299 ( .A1(n14656), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14658) );
  OR2_X1 U18300 ( .A1(n19538), .A2(n14658), .ZN(n19550) );
  NOR2_X1 U18301 ( .A1(n19719), .A2(n19550), .ZN(n14657) );
  MUX2_X1 U18302 ( .A(n14657), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n17178), .Z(P3_U3284) );
  NAND2_X1 U18303 ( .A1(n14659), .A2(n14658), .ZN(n19098) );
  NOR2_X1 U18304 ( .A1(n19098), .A2(P3_FLUSH_REG_SCAN_IN), .ZN(n14662) );
  NOR2_X1 U18305 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19712) );
  INV_X1 U18306 ( .A(n19712), .ZN(n14660) );
  AOI21_X1 U18307 ( .B1(n14660), .B2(n19096), .A(n19578), .ZN(n14661) );
  INV_X1 U18308 ( .A(n14661), .ZN(n19106) );
  OAI21_X1 U18309 ( .B1(n14662), .B2(n19688), .A(n19252), .ZN(n19103) );
  INV_X1 U18310 ( .A(n19103), .ZN(n14663) );
  NAND2_X1 U18311 ( .A1(n19690), .A2(n19096), .ZN(n19702) );
  NOR2_X1 U18312 ( .A1(n18790), .A2(n19702), .ZN(n17293) );
  AOI21_X1 U18313 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n17293), .ZN(n17294) );
  NOR2_X1 U18314 ( .A1(n14663), .A2(n17294), .ZN(n14665) );
  NAND3_X1 U18315 ( .A1(n19582), .A2(n19690), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19390) );
  INV_X1 U18316 ( .A(n19390), .ZN(n19450) );
  NOR2_X1 U18317 ( .A1(n19690), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19144) );
  OR2_X1 U18318 ( .A1(n19144), .A2(n14663), .ZN(n17292) );
  OR2_X1 U18319 ( .A1(n19450), .A2(n17292), .ZN(n14664) );
  MUX2_X1 U18320 ( .A(n14665), .B(n14664), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AOI22_X1 U18321 ( .A1(n15164), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15179), .ZN(n14669) );
  NOR3_X1 U18322 ( .A1(n15179), .A2(n20851), .A3(n14666), .ZN(n14667) );
  AOI22_X1 U18323 ( .A1(n15166), .A2(n20806), .B1(n15165), .B2(DATAI_30_), 
        .ZN(n14668) );
  OAI211_X1 U18324 ( .C1(n14689), .C2(n15182), .A(n14669), .B(n14668), .ZN(
        P1_U2874) );
  INV_X1 U18325 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14678) );
  INV_X1 U18326 ( .A(n14753), .ZN(n14672) );
  OAI22_X1 U18327 ( .A1(n14672), .A2(n14671), .B1(n13658), .B2(n14670), .ZN(
        n14673) );
  INV_X1 U18328 ( .A(n14674), .ZN(n14675) );
  OAI222_X1 U18329 ( .A1(n15111), .A2(n14689), .B1(n15113), .B2(n14678), .C1(
        n14677), .C2(n15114), .ZN(P1_U2842) );
  INV_X1 U18330 ( .A(n14679), .ZN(n14680) );
  AOI22_X1 U18331 ( .A1(n20736), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20738), .ZN(n14685) );
  NOR2_X1 U18332 ( .A1(n14756), .A2(n15184), .ZN(n14683) );
  OAI21_X1 U18333 ( .B1(n14683), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14682), 
        .ZN(n14684) );
  OAI211_X1 U18334 ( .C1(n20750), .C2(n14686), .A(n14685), .B(n14684), .ZN(
        n14687) );
  AOI21_X1 U18335 ( .B1(n15392), .B2(n20735), .A(n14687), .ZN(n14688) );
  OAI21_X1 U18336 ( .B1(n14689), .B2(n15058), .A(n14688), .ZN(P1_U2810) );
  NAND2_X1 U18337 ( .A1(n14508), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21160) );
  NOR3_X1 U18338 ( .A1(n20810), .A2(n21302), .A3(n14690), .ZN(n14691) );
  AOI21_X1 U18339 ( .B1(n20810), .B2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n14691), .ZN(n14692) );
  OAI21_X1 U18340 ( .B1(n14078), .B2(n14693), .A(n14692), .ZN(P1_U3476) );
  INV_X1 U18341 ( .A(n14693), .ZN(n14694) );
  NAND2_X1 U18342 ( .A1(n14694), .A2(n21063), .ZN(n14697) );
  INV_X1 U18343 ( .A(n21160), .ZN(n20917) );
  AOI21_X1 U18344 ( .B1(n21264), .B2(n20917), .A(n21302), .ZN(n21303) );
  NAND3_X1 U18345 ( .A1(n14698), .A2(n21303), .A3(n14695), .ZN(n14696) );
  OAI211_X1 U18346 ( .C1(n21132), .C2(n14698), .A(n14697), .B(n14696), .ZN(
        P1_U3475) );
  NAND2_X1 U18347 ( .A1(n15968), .A2(n15963), .ZN(n19839) );
  NAND2_X1 U18348 ( .A1(n19815), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16749) );
  AND3_X1 U18349 ( .A1(n19839), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n16749), 
        .ZN(n14706) );
  INV_X1 U18350 ( .A(n11445), .ZN(n14700) );
  NAND2_X1 U18351 ( .A1(n14700), .A2(n14699), .ZN(n16744) );
  MUX2_X1 U18352 ( .A(n16744), .B(n16759), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14701) );
  INV_X1 U18353 ( .A(n16883), .ZN(n14703) );
  OAI22_X1 U18354 ( .A1(n16868), .A2(n17296), .B1(n14704), .B2(n14703), .ZN(
        n14705) );
  OAI21_X1 U18355 ( .B1(n14706), .B2(n14705), .A(n17302), .ZN(n14707) );
  OAI21_X1 U18356 ( .B1(n17302), .B2(n10093), .A(n14707), .ZN(P2_U3601) );
  INV_X1 U18357 ( .A(n15640), .ZN(n14713) );
  AOI21_X1 U18358 ( .B1(n14708), .B2(n15629), .A(n14713), .ZN(n14714) );
  INV_X1 U18359 ( .A(n20921), .ZN(n14710) );
  OAI22_X1 U18360 ( .A1(n14710), .A2(n14709), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15626), .ZN(n17321) );
  INV_X1 U18361 ( .A(n17358), .ZN(n15636) );
  OAI22_X1 U18362 ( .A1(n15636), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21357), .ZN(n14711) );
  AOI21_X1 U18363 ( .B1(n15629), .B2(n17321), .A(n14711), .ZN(n14712) );
  OAI22_X1 U18364 ( .A1(n14714), .A2(n12593), .B1(n14713), .B2(n14712), .ZN(
        P1_U3474) );
  NAND2_X1 U18365 ( .A1(n16065), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14715) );
  OAI21_X1 U18366 ( .B1(n14738), .B2(n16065), .A(n14715), .ZN(P2_U2856) );
  INV_X1 U18367 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n14726) );
  OAI22_X1 U18368 ( .A1(n14717), .A2(n14716), .B1(n19804), .B2(n14726), .ZN(
        n14718) );
  AOI21_X1 U18369 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19841), .A(
        n14718), .ZN(n14719) );
  OAI21_X1 U18370 ( .B1(n14720), .B2(n19809), .A(n14719), .ZN(n14721) );
  AOI21_X1 U18371 ( .B1(n14722), .B2(n15952), .A(n14721), .ZN(n14731) );
  NAND2_X1 U18372 ( .A1(n14723), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14725) );
  NAND2_X1 U18373 ( .A1(n12524), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n14724) );
  OAI211_X1 U18374 ( .C1(n14727), .C2(n14726), .A(n14725), .B(n14724), .ZN(
        n14728) );
  NAND2_X1 U18375 ( .A1(n16069), .A2(n19812), .ZN(n14730) );
  OAI211_X1 U18376 ( .C1(n14738), .C2(n19776), .A(n14731), .B(n14730), .ZN(
        P2_U2824) );
  NAND3_X1 U18377 ( .A1(n14732), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16475), .ZN(n14737) );
  NAND4_X1 U18378 ( .A1(n16463), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14734), .A4(n14733), .ZN(n14735) );
  OAI21_X1 U18379 ( .B1(n14738), .B2(n19964), .A(n10608), .ZN(n14739) );
  NAND2_X1 U18380 ( .A1(n14740), .A2(n17444), .ZN(n14741) );
  OAI211_X1 U18381 ( .C1(n19963), .C2(n14743), .A(n14742), .B(n14741), .ZN(
        P2_U3015) );
  OR2_X1 U18382 ( .A1(n14744), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14747) );
  INV_X1 U18383 ( .A(n14745), .ZN(n14746) );
  MUX2_X1 U18384 ( .A(n14747), .B(n14746), .S(n21402), .Z(P1_U3487) );
  INV_X1 U18385 ( .A(n13712), .ZN(n14750) );
  NAND2_X1 U18386 ( .A1(n13658), .A2(n14751), .ZN(n14752) );
  NAND2_X1 U18387 ( .A1(n14753), .A2(n14752), .ZN(n15402) );
  INV_X1 U18388 ( .A(n15402), .ZN(n14761) );
  INV_X1 U18389 ( .A(n14754), .ZN(n14766) );
  OAI22_X1 U18390 ( .A1(n14755), .A2(n20718), .B1(n20702), .B2(n15086), .ZN(
        n14758) );
  NOR2_X1 U18391 ( .A1(n14756), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14757) );
  AOI211_X1 U18392 ( .C1(n14766), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14758), 
        .B(n14757), .ZN(n14759) );
  OAI21_X1 U18393 ( .B1(n20750), .B2(n15185), .A(n14759), .ZN(n14760) );
  AOI21_X1 U18394 ( .B1(n14761), .B2(n20735), .A(n14760), .ZN(n14762) );
  OAI21_X1 U18395 ( .B1(n15189), .B2(n15058), .A(n14762), .ZN(P1_U2811) );
  INV_X1 U18396 ( .A(n14764), .ZN(n15410) );
  AOI22_X1 U18397 ( .A1(n20736), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20738), .ZN(n14769) );
  INV_X1 U18398 ( .A(n14765), .ZN(n14767) );
  OAI21_X1 U18399 ( .B1(n14767), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14766), 
        .ZN(n14768) );
  OAI211_X1 U18400 ( .C1(n20750), .C2(n14770), .A(n14769), .B(n14768), .ZN(
        n14771) );
  AOI21_X1 U18401 ( .B1(n15410), .B2(n20735), .A(n14771), .ZN(n14772) );
  OAI21_X1 U18402 ( .B1(n15121), .B2(n15058), .A(n14772), .ZN(P1_U2812) );
  INV_X1 U18403 ( .A(n13657), .ZN(n14773) );
  OAI21_X1 U18404 ( .B1(n14774), .B2(n9647), .A(n14773), .ZN(n15418) );
  AOI21_X1 U18405 ( .B1(n14777), .B2(n14776), .A(n13002), .ZN(n15198) );
  NAND2_X1 U18406 ( .A1(n15198), .A2(n9887), .ZN(n14784) );
  INV_X1 U18407 ( .A(n14778), .ZN(n14779) );
  NAND2_X1 U18408 ( .A1(n20676), .A2(n14779), .ZN(n14791) );
  NAND3_X1 U18409 ( .A1(n14790), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n21377), 
        .ZN(n14781) );
  AOI22_X1 U18410 ( .A1(n20736), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20738), .ZN(n14780) );
  OAI211_X1 U18411 ( .C1(n14791), .C2(n21377), .A(n14781), .B(n14780), .ZN(
        n14782) );
  AOI21_X1 U18412 ( .B1(n20721), .B2(n15194), .A(n14782), .ZN(n14783) );
  OAI211_X1 U18413 ( .C1(n15079), .C2(n15418), .A(n14784), .B(n14783), .ZN(
        P1_U2813) );
  AND2_X1 U18414 ( .A1(n14808), .A2(n14785), .ZN(n14786) );
  OR2_X1 U18415 ( .A1(n14786), .A2(n9647), .ZN(n15426) );
  INV_X1 U18416 ( .A(n14776), .ZN(n14788) );
  NAND2_X1 U18417 ( .A1(n15203), .A2(n9887), .ZN(n14796) );
  INV_X1 U18418 ( .A(n14790), .ZN(n14792) );
  INV_X1 U18419 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15204) );
  AOI21_X1 U18420 ( .B1(n14792), .B2(n15204), .A(n14791), .ZN(n14794) );
  INV_X1 U18421 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15088) );
  OAI22_X1 U18422 ( .A1(n15205), .A2(n20718), .B1(n20702), .B2(n15088), .ZN(
        n14793) );
  AOI211_X1 U18423 ( .C1(n20721), .C2(n15207), .A(n14794), .B(n14793), .ZN(
        n14795) );
  OAI211_X1 U18424 ( .C1(n15426), .C2(n15079), .A(n14796), .B(n14795), .ZN(
        P1_U2814) );
  INV_X1 U18425 ( .A(n14787), .ZN(n14799) );
  AOI21_X1 U18426 ( .B1(n14800), .B2(n14798), .A(n14799), .ZN(n15215) );
  INV_X1 U18427 ( .A(n15215), .ZN(n15135) );
  INV_X1 U18428 ( .A(n15059), .ZN(n14801) );
  AOI21_X1 U18429 ( .B1(n15071), .B2(n14816), .A(n14801), .ZN(n14830) );
  OAI21_X1 U18430 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n20726), .A(n14830), 
        .ZN(n14802) );
  NAND2_X1 U18431 ( .A1(n14802), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14804) );
  AOI22_X1 U18432 ( .A1(n20736), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20738), .ZN(n14803) );
  OAI211_X1 U18433 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14805), .A(n14804), 
        .B(n14803), .ZN(n14810) );
  NAND2_X1 U18434 ( .A1(n14814), .A2(n14806), .ZN(n14807) );
  NAND2_X1 U18435 ( .A1(n14808), .A2(n14807), .ZN(n15435) );
  NOR2_X1 U18436 ( .A1(n15435), .A2(n15079), .ZN(n14809) );
  AOI211_X1 U18437 ( .C1(n20721), .C2(n15219), .A(n14810), .B(n14809), .ZN(
        n14811) );
  OAI21_X1 U18438 ( .B1(n15135), .B2(n15058), .A(n14811), .ZN(P1_U2815) );
  OAI21_X1 U18439 ( .B1(n14812), .B2(n14813), .A(n14798), .ZN(n15230) );
  OAI21_X1 U18440 ( .B1(n14835), .B2(n14815), .A(n14814), .ZN(n15450) );
  INV_X1 U18441 ( .A(n15450), .ZN(n14821) );
  NOR2_X1 U18442 ( .A1(n20750), .A2(n15223), .ZN(n14820) );
  AOI22_X1 U18443 ( .A1(n20736), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20738), .ZN(n14818) );
  OR3_X1 U18444 ( .A1(n20726), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14816), .ZN(
        n14817) );
  OAI211_X1 U18445 ( .C1(n14830), .C2(n15222), .A(n14818), .B(n14817), .ZN(
        n14819) );
  AOI211_X1 U18446 ( .C1(n14821), .C2(n20735), .A(n14820), .B(n14819), .ZN(
        n14822) );
  OAI21_X1 U18447 ( .B1(n15230), .B2(n15058), .A(n14822), .ZN(P1_U2816) );
  AOI21_X1 U18448 ( .B1(n14824), .B2(n14823), .A(n14812), .ZN(n15237) );
  INV_X1 U18449 ( .A(n15237), .ZN(n15141) );
  AND2_X1 U18450 ( .A1(n20672), .A2(n14826), .ZN(n14858) );
  INV_X1 U18451 ( .A(n14827), .ZN(n14828) );
  AOI21_X1 U18452 ( .B1(n14858), .B2(n14828), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14831) );
  AOI22_X1 U18453 ( .A1(n20736), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20738), .ZN(n14829) );
  OAI21_X1 U18454 ( .B1(n14831), .B2(n14830), .A(n14829), .ZN(n14837) );
  NOR2_X1 U18455 ( .A1(n14832), .A2(n14833), .ZN(n14834) );
  OR2_X1 U18456 ( .A1(n14835), .A2(n14834), .ZN(n15453) );
  NOR2_X1 U18457 ( .A1(n15453), .A2(n15079), .ZN(n14836) );
  AOI211_X1 U18458 ( .C1(n20721), .C2(n15233), .A(n14837), .B(n14836), .ZN(
        n14838) );
  OAI21_X1 U18459 ( .B1(n15141), .B2(n15058), .A(n14838), .ZN(P1_U2817) );
  INV_X1 U18460 ( .A(n14832), .ZN(n14839) );
  OAI21_X1 U18461 ( .B1(n14855), .B2(n14840), .A(n14839), .ZN(n15459) );
  INV_X1 U18462 ( .A(n14823), .ZN(n14842) );
  AOI21_X1 U18463 ( .B1(n10572), .B2(n14841), .A(n14842), .ZN(n15247) );
  NAND2_X1 U18464 ( .A1(n15247), .A2(n9887), .ZN(n14852) );
  INV_X1 U18465 ( .A(n15245), .ZN(n14850) );
  INV_X1 U18466 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14843) );
  NAND3_X1 U18467 ( .A1(n14858), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14843), 
        .ZN(n14848) );
  AOI22_X1 U18468 ( .A1(n20736), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20738), .ZN(n14847) );
  INV_X1 U18469 ( .A(n14844), .ZN(n14845) );
  AND2_X1 U18470 ( .A1(n15059), .A2(n14845), .ZN(n14872) );
  NAND2_X1 U18471 ( .A1(n14872), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14857) );
  NAND3_X1 U18472 ( .A1(n20676), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n14857), 
        .ZN(n14846) );
  NAND3_X1 U18473 ( .A1(n14848), .A2(n14847), .A3(n14846), .ZN(n14849) );
  AOI21_X1 U18474 ( .B1(n20721), .B2(n14850), .A(n14849), .ZN(n14851) );
  OAI211_X1 U18475 ( .C1(n15459), .C2(n15079), .A(n14852), .B(n14851), .ZN(
        P1_U2818) );
  OAI21_X1 U18476 ( .B1(n14853), .B2(n14854), .A(n14841), .ZN(n15257) );
  AOI21_X1 U18477 ( .B1(n14856), .B2(n14867), .A(n14855), .ZN(n15480) );
  AOI22_X1 U18478 ( .A1(n20736), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20738), .ZN(n14860) );
  OAI211_X1 U18479 ( .C1(n14858), .C2(P1_REIP_REG_21__SCAN_IN), .A(n20676), 
        .B(n14857), .ZN(n14859) );
  OAI211_X1 U18480 ( .C1(n20750), .C2(n15250), .A(n14860), .B(n14859), .ZN(
        n14861) );
  AOI21_X1 U18481 ( .B1(n15480), .B2(n20735), .A(n14861), .ZN(n14862) );
  OAI21_X1 U18482 ( .B1(n15257), .B2(n15058), .A(n14862), .ZN(P1_U2819) );
  INV_X1 U18483 ( .A(n14863), .ZN(n14866) );
  INV_X1 U18484 ( .A(n14864), .ZN(n14865) );
  AOI21_X1 U18485 ( .B1(n14866), .B2(n14865), .A(n14853), .ZN(n15265) );
  INV_X1 U18486 ( .A(n15265), .ZN(n15150) );
  INV_X1 U18487 ( .A(n14867), .ZN(n14868) );
  AOI21_X1 U18488 ( .B1(n14869), .B2(n14892), .A(n14868), .ZN(n15496) );
  AOI22_X1 U18489 ( .A1(n20736), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20738), .ZN(n14876) );
  NOR2_X1 U18490 ( .A1(n14973), .A2(n15324), .ZN(n14930) );
  AND2_X1 U18491 ( .A1(n20672), .A2(n14930), .ZN(n14958) );
  AND2_X1 U18492 ( .A1(n14933), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n14870) );
  NAND2_X1 U18493 ( .A1(n14958), .A2(n14870), .ZN(n14906) );
  NOR3_X1 U18494 ( .A1(n14906), .A2(n14871), .A3(n21371), .ZN(n14874) );
  INV_X1 U18495 ( .A(n14872), .ZN(n14873) );
  OAI211_X1 U18496 ( .C1(n14874), .C2(P1_REIP_REG_20__SCAN_IN), .A(n20676), 
        .B(n14873), .ZN(n14875) );
  OAI211_X1 U18497 ( .C1(n20750), .C2(n15263), .A(n14876), .B(n14875), .ZN(
        n14877) );
  AOI21_X1 U18498 ( .B1(n15496), .B2(n20735), .A(n14877), .ZN(n14878) );
  OAI21_X1 U18499 ( .B1(n15150), .B2(n15058), .A(n14878), .ZN(P1_U2820) );
  AOI21_X1 U18500 ( .B1(n14880), .B2(n14879), .A(n14864), .ZN(n15275) );
  INV_X1 U18501 ( .A(n15275), .ZN(n15157) );
  XNOR2_X1 U18502 ( .A(P1_REIP_REG_19__SCAN_IN), .B(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14890) );
  NAND2_X1 U18503 ( .A1(n15059), .A2(n15046), .ZN(n20677) );
  NAND2_X1 U18504 ( .A1(n20676), .A2(n20677), .ZN(n20708) );
  INV_X1 U18505 ( .A(n14881), .ZN(n14882) );
  NAND2_X1 U18506 ( .A1(n20676), .A2(n14882), .ZN(n14883) );
  INV_X1 U18507 ( .A(n14884), .ZN(n14885) );
  NAND2_X1 U18508 ( .A1(n15071), .A2(n14885), .ZN(n14886) );
  NAND2_X1 U18509 ( .A1(n15053), .A2(n14886), .ZN(n14922) );
  NAND2_X1 U18510 ( .A1(n14922), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14889) );
  OAI21_X1 U18511 ( .B1(n20718), .B2(n15273), .A(n20716), .ZN(n14887) );
  AOI21_X1 U18512 ( .B1(n20736), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14887), .ZN(
        n14888) );
  OAI211_X1 U18513 ( .C1(n14906), .C2(n14890), .A(n14889), .B(n14888), .ZN(
        n14891) );
  AOI21_X1 U18514 ( .B1(n20721), .B2(n15271), .A(n14891), .ZN(n14896) );
  INV_X1 U18515 ( .A(n14892), .ZN(n14893) );
  AOI21_X1 U18516 ( .B1(n14894), .B2(n14899), .A(n14893), .ZN(n15505) );
  NAND2_X1 U18517 ( .A1(n15505), .A2(n20735), .ZN(n14895) );
  OAI211_X1 U18518 ( .C1(n15157), .C2(n15058), .A(n14896), .B(n14895), .ZN(
        P1_U2821) );
  OR2_X1 U18519 ( .A1(n14917), .A2(n14897), .ZN(n14898) );
  NAND2_X1 U18520 ( .A1(n14899), .A2(n14898), .ZN(n15521) );
  INV_X1 U18521 ( .A(n14900), .ZN(n14913) );
  OAI21_X1 U18522 ( .B1(n14913), .B2(n14901), .A(n14879), .ZN(n15282) );
  INV_X1 U18523 ( .A(n15282), .ZN(n14902) );
  NAND2_X1 U18524 ( .A1(n14902), .A2(n9887), .ZN(n14910) );
  OAI21_X1 U18525 ( .B1(n20718), .B2(n14903), .A(n20716), .ZN(n14904) );
  AOI21_X1 U18526 ( .B1(n20736), .B2(P1_EBX_REG_18__SCAN_IN), .A(n14904), .ZN(
        n14905) );
  OAI21_X1 U18527 ( .B1(n14906), .B2(P1_REIP_REG_18__SCAN_IN), .A(n14905), 
        .ZN(n14908) );
  NOR2_X1 U18528 ( .A1(n20750), .A2(n15277), .ZN(n14907) );
  AOI211_X1 U18529 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n14922), .A(n14908), 
        .B(n14907), .ZN(n14909) );
  OAI211_X1 U18530 ( .C1(n15521), .C2(n15079), .A(n14910), .B(n14909), .ZN(
        P1_U2822) );
  AOI21_X1 U18531 ( .B1(n14914), .B2(n14912), .A(n14913), .ZN(n15290) );
  NOR2_X1 U18532 ( .A1(n14942), .A2(n14915), .ZN(n14916) );
  OR2_X1 U18533 ( .A1(n14917), .A2(n14916), .ZN(n15525) );
  NOR2_X1 U18534 ( .A1(n15525), .A2(n15079), .ZN(n14925) );
  NAND2_X1 U18535 ( .A1(n14958), .A2(n14933), .ZN(n14918) );
  INV_X1 U18536 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15286) );
  NAND2_X1 U18537 ( .A1(n14918), .A2(n15286), .ZN(n14921) );
  NAND2_X1 U18538 ( .A1(n20738), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14919) );
  OAI211_X1 U18539 ( .C1(n20702), .C2(n15097), .A(n20716), .B(n14919), .ZN(
        n14920) );
  AOI21_X1 U18540 ( .B1(n14922), .B2(n14921), .A(n14920), .ZN(n14923) );
  OAI21_X1 U18541 ( .B1(n20750), .B2(n15288), .A(n14923), .ZN(n14924) );
  AOI211_X1 U18542 ( .C1(n15290), .C2(n9887), .A(n14925), .B(n14924), .ZN(
        n14926) );
  INV_X1 U18543 ( .A(n14926), .ZN(P1_U2823) );
  OAI21_X1 U18544 ( .B1(n14928), .B2(n14929), .A(n14912), .ZN(n15169) );
  INV_X1 U18545 ( .A(n15169), .ZN(n15306) );
  INV_X1 U18546 ( .A(n14930), .ZN(n14931) );
  NAND2_X1 U18547 ( .A1(n15071), .A2(n14931), .ZN(n14932) );
  NAND2_X1 U18548 ( .A1(n15053), .A2(n14932), .ZN(n14975) );
  INV_X1 U18549 ( .A(n14933), .ZN(n14934) );
  OAI211_X1 U18550 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14958), .B(n14934), .ZN(n14937) );
  NAND2_X1 U18551 ( .A1(n20736), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n14936) );
  NAND2_X1 U18552 ( .A1(n20738), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14935) );
  NAND4_X1 U18553 ( .A1(n14937), .A2(n20716), .A3(n14936), .A4(n14935), .ZN(
        n14938) );
  AOI21_X1 U18554 ( .B1(n14975), .B2(P1_REIP_REG_16__SCAN_IN), .A(n14938), 
        .ZN(n14944) );
  INV_X1 U18555 ( .A(n14939), .ZN(n14957) );
  AND2_X1 U18556 ( .A1(n14957), .A2(n14940), .ZN(n14941) );
  NOR2_X1 U18557 ( .A1(n14942), .A2(n14941), .ZN(n15540) );
  NAND2_X1 U18558 ( .A1(n15540), .A2(n20735), .ZN(n14943) );
  OAI211_X1 U18559 ( .C1(n20750), .C2(n15304), .A(n14944), .B(n14943), .ZN(
        n14945) );
  AOI21_X1 U18560 ( .B1(n15306), .B2(n9887), .A(n14945), .ZN(n14946) );
  INV_X1 U18561 ( .A(n14946), .ZN(P1_U2824) );
  INV_X1 U18562 ( .A(n14982), .ZN(n14948) );
  OR2_X1 U18563 ( .A1(n14947), .A2(n15019), .ZN(n14951) );
  NAND2_X1 U18564 ( .A1(n14984), .A2(n15005), .ZN(n14950) );
  INV_X1 U18565 ( .A(n14952), .ZN(n14967) );
  NAND2_X1 U18566 ( .A1(n14985), .A2(n14967), .ZN(n14968) );
  AOI21_X1 U18567 ( .B1(n14968), .B2(n14953), .A(n14928), .ZN(n15317) );
  INV_X1 U18568 ( .A(n15317), .ZN(n15172) );
  NAND2_X1 U18569 ( .A1(n14954), .A2(n14955), .ZN(n14956) );
  AND2_X1 U18570 ( .A1(n14957), .A2(n14956), .ZN(n15548) );
  INV_X1 U18571 ( .A(n14958), .ZN(n14963) );
  NAND2_X1 U18572 ( .A1(n14975), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14962) );
  OAI21_X1 U18573 ( .B1(n20718), .B2(n14959), .A(n20716), .ZN(n14960) );
  AOI21_X1 U18574 ( .B1(n20736), .B2(P1_EBX_REG_15__SCAN_IN), .A(n14960), .ZN(
        n14961) );
  OAI211_X1 U18575 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n14963), .A(n14962), 
        .B(n14961), .ZN(n14965) );
  NOR2_X1 U18576 ( .A1(n20750), .A2(n15315), .ZN(n14964) );
  AOI211_X1 U18577 ( .C1(n15548), .C2(n20735), .A(n14965), .B(n14964), .ZN(
        n14966) );
  OAI21_X1 U18578 ( .B1(n15172), .B2(n15058), .A(n14966), .ZN(P1_U2825) );
  OR2_X1 U18579 ( .A1(n14985), .A2(n14967), .ZN(n14969) );
  INV_X1 U18580 ( .A(n15326), .ZN(n14980) );
  OR2_X1 U18581 ( .A1(n14989), .A2(n14970), .ZN(n14971) );
  NAND2_X1 U18582 ( .A1(n14954), .A2(n14971), .ZN(n17391) );
  INV_X1 U18583 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15100) );
  NOR2_X1 U18584 ( .A1(n20702), .A2(n15100), .ZN(n14972) );
  AOI211_X1 U18585 ( .C1(n20738), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17416), .B(n14972), .ZN(n14978) );
  INV_X1 U18586 ( .A(n20672), .ZN(n14974) );
  NOR2_X1 U18587 ( .A1(n14974), .A2(n14973), .ZN(n14976) );
  OAI21_X1 U18588 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14976), .A(n14975), 
        .ZN(n14977) );
  OAI211_X1 U18589 ( .C1(n17391), .C2(n15079), .A(n14978), .B(n14977), .ZN(
        n14979) );
  AOI21_X1 U18590 ( .B1(n20721), .B2(n14980), .A(n14979), .ZN(n14981) );
  OAI21_X1 U18591 ( .B1(n15174), .B2(n15058), .A(n14981), .ZN(P1_U2826) );
  INV_X1 U18592 ( .A(n14947), .ZN(n15034) );
  OAI21_X1 U18593 ( .B1(n15034), .B2(n14982), .A(n14983), .ZN(n15020) );
  OAI21_X1 U18594 ( .B1(n15020), .B2(n15019), .A(n14983), .ZN(n15006) );
  NAND2_X1 U18595 ( .A1(n15006), .A2(n15005), .ZN(n15004) );
  INV_X1 U18596 ( .A(n14984), .ZN(n14986) );
  AOI21_X1 U18597 ( .B1(n15004), .B2(n14986), .A(n14985), .ZN(n15340) );
  INV_X1 U18598 ( .A(n15340), .ZN(n15176) );
  INV_X1 U18599 ( .A(n15338), .ZN(n15002) );
  NOR2_X1 U18600 ( .A1(n15009), .A2(n14987), .ZN(n14988) );
  OR2_X1 U18601 ( .A1(n14989), .A2(n14988), .ZN(n15551) );
  INV_X1 U18602 ( .A(n14994), .ZN(n14990) );
  NAND2_X1 U18603 ( .A1(n15071), .A2(n14990), .ZN(n14991) );
  AND2_X1 U18604 ( .A1(n15053), .A2(n14991), .ZN(n15041) );
  INV_X1 U18605 ( .A(n14995), .ZN(n14992) );
  NAND2_X1 U18606 ( .A1(n20676), .A2(n14992), .ZN(n14993) );
  NAND2_X1 U18607 ( .A1(n15041), .A2(n14993), .ZN(n15013) );
  NAND2_X1 U18608 ( .A1(n15013), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15000) );
  AND2_X1 U18609 ( .A1(n20672), .A2(n14994), .ZN(n15021) );
  AND2_X1 U18610 ( .A1(n14995), .A2(n13871), .ZN(n14998) );
  NAND2_X1 U18611 ( .A1(n20738), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14996) );
  OAI211_X1 U18612 ( .C1(n20702), .C2(n15102), .A(n20716), .B(n14996), .ZN(
        n14997) );
  AOI21_X1 U18613 ( .B1(n15021), .B2(n14998), .A(n14997), .ZN(n14999) );
  OAI211_X1 U18614 ( .C1(n15551), .C2(n15079), .A(n15000), .B(n14999), .ZN(
        n15001) );
  AOI21_X1 U18615 ( .B1(n20721), .B2(n15002), .A(n15001), .ZN(n15003) );
  OAI21_X1 U18616 ( .B1(n15176), .B2(n15058), .A(n15003), .ZN(P1_U2827) );
  OAI21_X1 U18617 ( .B1(n15006), .B2(n15005), .A(n15004), .ZN(n15350) );
  AND2_X1 U18618 ( .A1(n10469), .A2(n15007), .ZN(n15008) );
  NOR2_X1 U18619 ( .A1(n15009), .A2(n15008), .ZN(n15569) );
  INV_X1 U18620 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15011) );
  NAND2_X1 U18621 ( .A1(n20738), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15010) );
  OAI211_X1 U18622 ( .C1(n20702), .C2(n15011), .A(n20716), .B(n15010), .ZN(
        n15012) );
  AOI21_X1 U18623 ( .B1(n15569), .B2(n20735), .A(n15012), .ZN(n15016) );
  AND2_X1 U18624 ( .A1(n15021), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15014) );
  OAI21_X1 U18625 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n15014), .A(n15013), 
        .ZN(n15015) );
  OAI211_X1 U18626 ( .C1(n20750), .C2(n15346), .A(n15016), .B(n15015), .ZN(
        n15017) );
  INV_X1 U18627 ( .A(n15017), .ZN(n15018) );
  OAI21_X1 U18628 ( .B1(n15350), .B2(n15058), .A(n15018), .ZN(P1_U2828) );
  XNOR2_X1 U18629 ( .A(n15020), .B(n15019), .ZN(n15360) );
  INV_X1 U18630 ( .A(n15041), .ZN(n15032) );
  INV_X1 U18631 ( .A(n15021), .ZN(n15029) );
  NAND2_X1 U18632 ( .A1(n15022), .A2(n15023), .ZN(n15024) );
  AND2_X1 U18633 ( .A1(n10469), .A2(n15024), .ZN(n15584) );
  NAND2_X1 U18634 ( .A1(n20736), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n15025) );
  OAI211_X1 U18635 ( .C1(n20718), .C2(n15026), .A(n15025), .B(n20716), .ZN(
        n15027) );
  AOI21_X1 U18636 ( .B1(n15584), .B2(n20735), .A(n15027), .ZN(n15028) );
  OAI21_X1 U18637 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15029), .A(n15028), 
        .ZN(n15031) );
  NOR2_X1 U18638 ( .A1(n20750), .A2(n15356), .ZN(n15030) );
  AOI211_X1 U18639 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15032), .A(n15031), 
        .B(n15030), .ZN(n15033) );
  OAI21_X1 U18640 ( .B1(n15360), .B2(n15058), .A(n15033), .ZN(P1_U2829) );
  AOI21_X1 U18641 ( .B1(n15035), .B2(n14649), .A(n15034), .ZN(n15371) );
  INV_X1 U18642 ( .A(n15371), .ZN(n15183) );
  INV_X1 U18643 ( .A(n15369), .ZN(n15044) );
  OR2_X1 U18644 ( .A1(n15037), .A2(n15036), .ZN(n15038) );
  NAND2_X1 U18645 ( .A1(n15022), .A2(n15038), .ZN(n15594) );
  NOR2_X1 U18646 ( .A1(n20702), .A2(n15106), .ZN(n15039) );
  AOI211_X1 U18647 ( .C1(n20738), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17416), .B(n15039), .ZN(n15040) );
  OAI21_X1 U18648 ( .B1(n15079), .B2(n15594), .A(n15040), .ZN(n15043) );
  NAND2_X1 U18649 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15053), .ZN(n20671) );
  AOI21_X1 U18650 ( .B1(n13900), .B2(n20671), .A(n15041), .ZN(n15042) );
  AOI211_X1 U18651 ( .C1(n20721), .C2(n15044), .A(n15043), .B(n15042), .ZN(
        n15045) );
  OAI21_X1 U18652 ( .B1(n15183), .B2(n15058), .A(n15045), .ZN(P1_U2830) );
  NAND3_X1 U18653 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n15047) );
  NAND2_X1 U18654 ( .A1(n15071), .A2(n15046), .ZN(n20704) );
  NOR3_X1 U18655 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n15047), .A3(n20704), .ZN(
        n15048) );
  AOI211_X1 U18656 ( .C1(n20738), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17416), .B(n15048), .ZN(n15057) );
  INV_X1 U18657 ( .A(n15383), .ZN(n15055) );
  AND2_X1 U18658 ( .A1(n15050), .A2(n15049), .ZN(n15051) );
  NOR2_X1 U18659 ( .A1(n14651), .A2(n15051), .ZN(n17407) );
  AOI22_X1 U18660 ( .A1(n17407), .A2(n20735), .B1(n20736), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n15052) );
  OAI21_X1 U18661 ( .B1(n15053), .B2(n13904), .A(n15052), .ZN(n15054) );
  AOI21_X1 U18662 ( .B1(n20721), .B2(n15055), .A(n15054), .ZN(n15056) );
  OAI211_X1 U18663 ( .C1(n15110), .C2(n15058), .A(n15057), .B(n15056), .ZN(
        P1_U2832) );
  NAND2_X1 U18664 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20725) );
  NAND2_X1 U18665 ( .A1(n15071), .A2(n20725), .ZN(n15064) );
  NAND2_X1 U18666 ( .A1(n15064), .A2(n15059), .ZN(n20737) );
  NAND2_X1 U18667 ( .A1(n15059), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n15070) );
  INV_X1 U18668 ( .A(n14078), .ZN(n20817) );
  AND2_X1 U18669 ( .A1(n21402), .A2(n15060), .ZN(n20747) );
  AOI22_X1 U18670 ( .A1(n20817), .A2(n20747), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20738), .ZN(n15063) );
  AOI22_X1 U18671 ( .A1(n20736), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n20735), .B2(
        n15061), .ZN(n15062) );
  OAI211_X1 U18672 ( .C1(n15064), .C2(n15070), .A(n15063), .B(n15062), .ZN(
        n15067) );
  NOR2_X1 U18673 ( .A1(n20750), .A2(n15065), .ZN(n15066) );
  AOI211_X1 U18674 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n20737), .A(n15067), .B(
        n15066), .ZN(n15068) );
  OAI21_X1 U18675 ( .B1(n15069), .B2(n20744), .A(n15068), .ZN(P1_U2838) );
  OAI21_X1 U18676 ( .B1(n15071), .B2(P1_REIP_REG_1__SCAN_IN), .A(n15070), .ZN(
        n15072) );
  AOI22_X1 U18677 ( .A1(n20736), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n20747), .B2(
        n21273), .ZN(n15074) );
  MUX2_X1 U18678 ( .A(n20750), .B(n20718), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15073) );
  OAI211_X1 U18679 ( .C1(n20744), .C2(n15075), .A(n15074), .B(n15073), .ZN(
        n15076) );
  OR2_X1 U18680 ( .A1(n15077), .A2(n15076), .ZN(P1_U2839) );
  OAI21_X1 U18681 ( .B1(n20721), .B2(n20738), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15082) );
  AOI22_X1 U18682 ( .A1(n20736), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n20747), .B2(
        n20921), .ZN(n15078) );
  OAI21_X1 U18683 ( .B1(n15079), .B2(n15610), .A(n15078), .ZN(n15080) );
  AOI21_X1 U18684 ( .B1(n20676), .B2(P1_REIP_REG_0__SCAN_IN), .A(n15080), .ZN(
        n15081) );
  OAI211_X1 U18685 ( .C1(n20744), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        P1_U2840) );
  OAI22_X1 U18686 ( .A1(n15084), .A2(n15114), .B1(n15085), .B2(n15113), .ZN(
        P1_U2841) );
  OAI222_X1 U18687 ( .A1(n15086), .A2(n15113), .B1(n15114), .B2(n15402), .C1(
        n15189), .C2(n15111), .ZN(P1_U2843) );
  INV_X1 U18688 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15087) );
  INV_X1 U18689 ( .A(n15198), .ZN(n15124) );
  OAI222_X1 U18690 ( .A1(n15087), .A2(n15113), .B1(n15114), .B2(n15418), .C1(
        n15124), .C2(n15101), .ZN(P1_U2845) );
  INV_X1 U18691 ( .A(n15203), .ZN(n15129) );
  OAI222_X1 U18692 ( .A1(n15088), .A2(n15113), .B1(n15114), .B2(n15426), .C1(
        n15129), .C2(n15101), .ZN(P1_U2846) );
  INV_X1 U18693 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15089) );
  OAI222_X1 U18694 ( .A1(n15089), .A2(n15113), .B1(n15114), .B2(n15435), .C1(
        n15135), .C2(n15101), .ZN(P1_U2847) );
  INV_X1 U18695 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15090) );
  OAI222_X1 U18696 ( .A1(n15090), .A2(n15113), .B1(n15114), .B2(n15450), .C1(
        n15230), .C2(n15101), .ZN(P1_U2848) );
  INV_X1 U18697 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15091) );
  OAI222_X1 U18698 ( .A1(n15453), .A2(n15114), .B1(n15091), .B2(n15113), .C1(
        n15141), .C2(n15101), .ZN(P1_U2849) );
  INV_X1 U18699 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15092) );
  INV_X1 U18700 ( .A(n15247), .ZN(n15144) );
  OAI222_X1 U18701 ( .A1(n15459), .A2(n15114), .B1(n15092), .B2(n15113), .C1(
        n15144), .C2(n15101), .ZN(P1_U2850) );
  AOI22_X1 U18702 ( .A1(n15480), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n15093) );
  OAI21_X1 U18703 ( .B1(n15257), .B2(n15111), .A(n15093), .ZN(P1_U2851) );
  AOI22_X1 U18704 ( .A1(n15496), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n15094) );
  OAI21_X1 U18705 ( .B1(n15150), .B2(n15101), .A(n15094), .ZN(P1_U2852) );
  AOI22_X1 U18706 ( .A1(n15505), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n15095) );
  OAI21_X1 U18707 ( .B1(n15157), .B2(n15101), .A(n15095), .ZN(P1_U2853) );
  INV_X1 U18708 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15096) );
  OAI222_X1 U18709 ( .A1(n15521), .A2(n15114), .B1(n15096), .B2(n15113), .C1(
        n15282), .C2(n15101), .ZN(P1_U2854) );
  INV_X1 U18710 ( .A(n15290), .ZN(n15163) );
  OAI222_X1 U18711 ( .A1(n15525), .A2(n15114), .B1(n15097), .B2(n15113), .C1(
        n15163), .C2(n15101), .ZN(P1_U2855) );
  AOI22_X1 U18712 ( .A1(n15540), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n15098) );
  OAI21_X1 U18713 ( .B1(n15169), .B2(n15111), .A(n15098), .ZN(P1_U2856) );
  AOI22_X1 U18714 ( .A1(n15548), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n15099) );
  OAI21_X1 U18715 ( .B1(n15172), .B2(n15101), .A(n15099), .ZN(P1_U2857) );
  OAI222_X1 U18716 ( .A1(n17391), .A2(n15114), .B1(n15100), .B2(n15113), .C1(
        n15111), .C2(n15174), .ZN(P1_U2858) );
  OAI222_X1 U18717 ( .A1(n15551), .A2(n15114), .B1(n15102), .B2(n15113), .C1(
        n15176), .C2(n15101), .ZN(P1_U2859) );
  AOI22_X1 U18718 ( .A1(n15569), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n15103) );
  OAI21_X1 U18719 ( .B1(n15350), .B2(n15111), .A(n15103), .ZN(P1_U2860) );
  AOI22_X1 U18720 ( .A1(n15584), .A2(n15104), .B1(n13660), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15105) );
  OAI21_X1 U18721 ( .B1(n15360), .B2(n15111), .A(n15105), .ZN(P1_U2861) );
  OAI22_X1 U18722 ( .A1(n15594), .A2(n15114), .B1(n15106), .B2(n15113), .ZN(
        n15107) );
  AOI21_X1 U18723 ( .B1(n15371), .B2(n15108), .A(n15107), .ZN(n15109) );
  INV_X1 U18724 ( .A(n15109), .ZN(P1_U2862) );
  INV_X1 U18725 ( .A(n17407), .ZN(n15115) );
  INV_X1 U18726 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15112) );
  OAI222_X1 U18727 ( .A1(n15115), .A2(n15114), .B1(n15113), .B2(n15112), .C1(
        n15111), .C2(n15110), .ZN(P1_U2864) );
  AOI22_X1 U18728 ( .A1(n15164), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n15179), .ZN(n15117) );
  AOI22_X1 U18729 ( .A1(n15166), .A2(n20801), .B1(n15165), .B2(DATAI_29_), 
        .ZN(n15116) );
  OAI211_X1 U18730 ( .C1(n15189), .C2(n15182), .A(n15117), .B(n15116), .ZN(
        P1_U2875) );
  INV_X1 U18731 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n17460) );
  OAI22_X1 U18732 ( .A1(n15153), .A2(n17460), .B1(n14337), .B2(n15151), .ZN(
        n15118) );
  INV_X1 U18733 ( .A(n15118), .ZN(n15120) );
  AOI22_X1 U18734 ( .A1(n15166), .A2(n20798), .B1(n15165), .B2(DATAI_28_), 
        .ZN(n15119) );
  OAI211_X1 U18735 ( .C1(n15121), .C2(n15182), .A(n15120), .B(n15119), .ZN(
        P1_U2876) );
  AOI22_X1 U18736 ( .A1(n15164), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n15179), .ZN(n15123) );
  AOI22_X1 U18737 ( .A1(n15166), .A2(n20794), .B1(n15165), .B2(DATAI_27_), 
        .ZN(n15122) );
  OAI211_X1 U18738 ( .C1(n15124), .C2(n15182), .A(n15123), .B(n15122), .ZN(
        P1_U2877) );
  INV_X1 U18739 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16097) );
  OAI22_X1 U18740 ( .A1(n15153), .A2(n16097), .B1(n15125), .B2(n15151), .ZN(
        n15126) );
  INV_X1 U18741 ( .A(n15126), .ZN(n15128) );
  AOI22_X1 U18742 ( .A1(n15166), .A2(n20791), .B1(n15165), .B2(DATAI_26_), 
        .ZN(n15127) );
  OAI211_X1 U18743 ( .C1(n15129), .C2(n15182), .A(n15128), .B(n15127), .ZN(
        P1_U2878) );
  INV_X1 U18744 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n15131) );
  OAI22_X1 U18745 ( .A1(n15153), .A2(n15131), .B1(n15130), .B2(n15151), .ZN(
        n15132) );
  INV_X1 U18746 ( .A(n15132), .ZN(n15134) );
  AOI22_X1 U18747 ( .A1(n15166), .A2(n20788), .B1(n15165), .B2(DATAI_25_), 
        .ZN(n15133) );
  OAI211_X1 U18748 ( .C1(n15135), .C2(n15182), .A(n15134), .B(n15133), .ZN(
        P1_U2879) );
  AOI22_X1 U18749 ( .A1(n15164), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n15179), .ZN(n15138) );
  AOI22_X1 U18750 ( .A1(n15166), .A2(n15136), .B1(n15165), .B2(DATAI_24_), 
        .ZN(n15137) );
  OAI211_X1 U18751 ( .C1(n15230), .C2(n15182), .A(n15138), .B(n15137), .ZN(
        P1_U2880) );
  AOI22_X1 U18752 ( .A1(n15164), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n15179), .ZN(n15140) );
  AOI22_X1 U18753 ( .A1(n15166), .A2(n20854), .B1(n15165), .B2(DATAI_23_), 
        .ZN(n15139) );
  OAI211_X1 U18754 ( .C1(n15141), .C2(n15182), .A(n15140), .B(n15139), .ZN(
        P1_U2881) );
  AOI22_X1 U18755 ( .A1(n15164), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15179), .ZN(n15143) );
  AOI22_X1 U18756 ( .A1(n15166), .A2(n20846), .B1(n15165), .B2(DATAI_22_), 
        .ZN(n15142) );
  OAI211_X1 U18757 ( .C1(n15144), .C2(n15182), .A(n15143), .B(n15142), .ZN(
        P1_U2882) );
  AOI22_X1 U18758 ( .A1(n15164), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15179), .ZN(n15146) );
  AOI22_X1 U18759 ( .A1(n15166), .A2(n20843), .B1(n15165), .B2(DATAI_21_), 
        .ZN(n15145) );
  OAI211_X1 U18760 ( .C1(n15257), .C2(n15182), .A(n15146), .B(n15145), .ZN(
        P1_U2883) );
  INV_X1 U18761 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n17473) );
  OAI22_X1 U18762 ( .A1(n15153), .A2(n17473), .B1(n14333), .B2(n15151), .ZN(
        n15147) );
  INV_X1 U18763 ( .A(n15147), .ZN(n15149) );
  AOI22_X1 U18764 ( .A1(n15166), .A2(n20839), .B1(n15165), .B2(DATAI_20_), 
        .ZN(n15148) );
  OAI211_X1 U18765 ( .C1(n15150), .C2(n15182), .A(n15149), .B(n15148), .ZN(
        P1_U2884) );
  INV_X1 U18766 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16147) );
  OAI22_X1 U18767 ( .A1(n15153), .A2(n16147), .B1(n15152), .B2(n15151), .ZN(
        n15154) );
  INV_X1 U18768 ( .A(n15154), .ZN(n15156) );
  AOI22_X1 U18769 ( .A1(n15166), .A2(n20836), .B1(n15165), .B2(DATAI_19_), 
        .ZN(n15155) );
  OAI211_X1 U18770 ( .C1(n15157), .C2(n15182), .A(n15156), .B(n15155), .ZN(
        P1_U2885) );
  AOI22_X1 U18771 ( .A1(n15164), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15179), .ZN(n15159) );
  AOI22_X1 U18772 ( .A1(n15166), .A2(n20833), .B1(n15165), .B2(DATAI_18_), 
        .ZN(n15158) );
  OAI211_X1 U18773 ( .C1(n15282), .C2(n15182), .A(n15159), .B(n15158), .ZN(
        P1_U2886) );
  AOI22_X1 U18774 ( .A1(n15164), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n15179), .ZN(n15162) );
  AOI22_X1 U18775 ( .A1(n15166), .A2(n15160), .B1(n15165), .B2(DATAI_17_), 
        .ZN(n15161) );
  OAI211_X1 U18776 ( .C1(n15163), .C2(n15182), .A(n15162), .B(n15161), .ZN(
        P1_U2887) );
  AOI22_X1 U18777 ( .A1(n15164), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n15179), .ZN(n15168) );
  AOI22_X1 U18778 ( .A1(n15166), .A2(n20821), .B1(n15165), .B2(DATAI_16_), 
        .ZN(n15167) );
  OAI211_X1 U18779 ( .C1(n15169), .C2(n15182), .A(n15168), .B(n15167), .ZN(
        P1_U2888) );
  AOI22_X1 U18780 ( .A1(n15180), .A2(n15170), .B1(P1_EAX_REG_15__SCAN_IN), 
        .B2(n15179), .ZN(n15171) );
  OAI21_X1 U18781 ( .B1(n15172), .B2(n15182), .A(n15171), .ZN(P1_U2889) );
  AOI22_X1 U18782 ( .A1(n15180), .A2(n20806), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15179), .ZN(n15173) );
  OAI21_X1 U18783 ( .B1(n15174), .B2(n15182), .A(n15173), .ZN(P1_U2890) );
  AOI22_X1 U18784 ( .A1(n15180), .A2(n20801), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15179), .ZN(n15175) );
  OAI21_X1 U18785 ( .B1(n15176), .B2(n15182), .A(n15175), .ZN(P1_U2891) );
  AOI22_X1 U18786 ( .A1(n15180), .A2(n20798), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15179), .ZN(n15177) );
  OAI21_X1 U18787 ( .B1(n15350), .B2(n15182), .A(n15177), .ZN(P1_U2892) );
  AOI22_X1 U18788 ( .A1(n15180), .A2(n20794), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15179), .ZN(n15178) );
  OAI21_X1 U18789 ( .B1(n15360), .B2(n15182), .A(n15178), .ZN(P1_U2893) );
  AOI22_X1 U18790 ( .A1(n15180), .A2(n20791), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15179), .ZN(n15181) );
  OAI21_X1 U18791 ( .B1(n15183), .B2(n15182), .A(n15181), .ZN(P1_U2894) );
  NOR2_X1 U18792 ( .A1(n20716), .A2(n15184), .ZN(n15398) );
  NOR2_X1 U18793 ( .A1(n15185), .A2(n17377), .ZN(n15186) );
  AOI211_X1 U18794 ( .C1(n17370), .C2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15398), .B(n15186), .ZN(n15188) );
  MUX2_X1 U18795 ( .A(n15192), .B(n15191), .S(n15351), .Z(n15193) );
  XNOR2_X1 U18796 ( .A(n15193), .B(n15416), .ZN(n15422) );
  INV_X1 U18797 ( .A(n15194), .ZN(n15196) );
  NOR2_X1 U18798 ( .A1(n20716), .A2(n21377), .ZN(n15415) );
  AOI21_X1 U18799 ( .B1(n17370), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15415), .ZN(n15195) );
  OAI21_X1 U18800 ( .B1(n15196), .B2(n17377), .A(n15195), .ZN(n15197) );
  AOI21_X1 U18801 ( .B1(n15198), .B2(n17381), .A(n15197), .ZN(n15199) );
  OAI21_X1 U18802 ( .B1(n20646), .B2(n15422), .A(n15199), .ZN(P1_U2972) );
  OAI21_X1 U18803 ( .B1(n12227), .B2(n15425), .A(n12217), .ZN(n15200) );
  NAND2_X1 U18804 ( .A1(n15201), .A2(n15200), .ZN(n15202) );
  XNOR2_X1 U18805 ( .A(n15202), .B(n15424), .ZN(n15432) );
  NAND2_X1 U18806 ( .A1(n15203), .A2(n17381), .ZN(n15209) );
  NOR2_X1 U18807 ( .A1(n20716), .A2(n15204), .ZN(n15428) );
  NOR2_X1 U18808 ( .A1(n17385), .A2(n15205), .ZN(n15206) );
  AOI211_X1 U18809 ( .C1(n15207), .C2(n17379), .A(n15428), .B(n15206), .ZN(
        n15208) );
  OAI211_X1 U18810 ( .C1(n15432), .C2(n20646), .A(n15209), .B(n15208), .ZN(
        P1_U2973) );
  MUX2_X1 U18811 ( .A(n15212), .B(n15211), .S(n12217), .Z(n15213) );
  AOI21_X1 U18812 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15225), .A(
        n15213), .ZN(n15214) );
  XNOR2_X1 U18813 ( .A(n15214), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15441) );
  NAND2_X1 U18814 ( .A1(n15215), .A2(n17381), .ZN(n15221) );
  NOR2_X1 U18815 ( .A1(n20716), .A2(n15216), .ZN(n15437) );
  NOR2_X1 U18816 ( .A1(n17385), .A2(n15217), .ZN(n15218) );
  AOI211_X1 U18817 ( .C1(n15219), .C2(n17379), .A(n15437), .B(n15218), .ZN(
        n15220) );
  OAI211_X1 U18818 ( .C1(n15441), .C2(n20646), .A(n15221), .B(n15220), .ZN(
        P1_U2974) );
  NOR2_X1 U18819 ( .A1(n20716), .A2(n15222), .ZN(n15446) );
  NOR2_X1 U18820 ( .A1(n15223), .A2(n17377), .ZN(n15224) );
  AOI211_X1 U18821 ( .C1(n17370), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15446), .B(n15224), .ZN(n15229) );
  NAND2_X1 U18822 ( .A1(n12227), .A2(n15225), .ZN(n15226) );
  MUX2_X1 U18823 ( .A(n15226), .B(n15225), .S(n12217), .Z(n15227) );
  XNOR2_X1 U18824 ( .A(n15227), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15442) );
  NAND2_X1 U18825 ( .A1(n15442), .A2(n17382), .ZN(n15228) );
  OAI211_X1 U18826 ( .C1(n15230), .C2(n20811), .A(n15229), .B(n15228), .ZN(
        P1_U2975) );
  XNOR2_X1 U18827 ( .A(n12217), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15232) );
  XNOR2_X1 U18828 ( .A(n15231), .B(n15232), .ZN(n15458) );
  NAND2_X1 U18829 ( .A1(n15233), .A2(n17379), .ZN(n15234) );
  NAND2_X1 U18830 ( .A1(n17416), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15451) );
  OAI211_X1 U18831 ( .C1(n17385), .C2(n15235), .A(n15234), .B(n15451), .ZN(
        n15236) );
  AOI21_X1 U18832 ( .B1(n15237), .B2(n17381), .A(n15236), .ZN(n15238) );
  OAI21_X1 U18833 ( .B1(n15458), .B2(n20646), .A(n15238), .ZN(P1_U2976) );
  XNOR2_X1 U18834 ( .A(n12217), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15279) );
  NAND2_X1 U18835 ( .A1(n15239), .A2(n15279), .ZN(n15508) );
  NOR3_X1 U18836 ( .A1(n15508), .A2(n15471), .A3(n15240), .ZN(n15242) );
  OAI21_X1 U18837 ( .B1(n15242), .B2(n15351), .A(n15241), .ZN(n15243) );
  XNOR2_X1 U18838 ( .A(n15243), .B(n15469), .ZN(n15479) );
  NAND2_X1 U18839 ( .A1(n17416), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15473) );
  NAND2_X1 U18840 ( .A1(n17370), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15244) );
  OAI211_X1 U18841 ( .C1(n15245), .C2(n17377), .A(n15473), .B(n15244), .ZN(
        n15246) );
  AOI21_X1 U18842 ( .B1(n15247), .B2(n17381), .A(n15246), .ZN(n15248) );
  OAI21_X1 U18843 ( .B1(n20646), .B2(n15479), .A(n15248), .ZN(P1_U2977) );
  NOR2_X1 U18844 ( .A1(n20716), .A2(n15249), .ZN(n15483) );
  NOR2_X1 U18845 ( .A1(n15250), .A2(n17377), .ZN(n15251) );
  AOI211_X1 U18846 ( .C1(n17370), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15483), .B(n15251), .ZN(n15256) );
  INV_X1 U18847 ( .A(n15508), .ZN(n15252) );
  AOI21_X1 U18848 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15351), .A(
        n15252), .ZN(n15269) );
  NAND2_X1 U18849 ( .A1(n15351), .A2(n15501), .ZN(n15268) );
  NOR2_X1 U18850 ( .A1(n15268), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15253) );
  NAND2_X1 U18851 ( .A1(n12217), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15267) );
  NOR2_X1 U18852 ( .A1(n15508), .A2(n15267), .ZN(n15259) );
  AOI22_X1 U18853 ( .A1(n15269), .A2(n15253), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15259), .ZN(n15254) );
  XNOR2_X1 U18854 ( .A(n15254), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15481) );
  NAND2_X1 U18855 ( .A1(n15481), .A2(n17382), .ZN(n15255) );
  OAI211_X1 U18856 ( .C1(n15257), .C2(n20811), .A(n15256), .B(n15255), .ZN(
        P1_U2978) );
  INV_X1 U18857 ( .A(n15259), .ZN(n15260) );
  OAI21_X1 U18858 ( .B1(n15268), .B2(n15258), .A(n15260), .ZN(n15261) );
  XNOR2_X1 U18859 ( .A(n15261), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15498) );
  NAND2_X1 U18860 ( .A1(n17416), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15492) );
  NAND2_X1 U18861 ( .A1(n17370), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15262) );
  OAI211_X1 U18862 ( .C1(n17377), .C2(n15263), .A(n15492), .B(n15262), .ZN(
        n15264) );
  AOI21_X1 U18863 ( .B1(n15265), .B2(n17381), .A(n15264), .ZN(n15266) );
  OAI21_X1 U18864 ( .B1(n15498), .B2(n20646), .A(n15266), .ZN(P1_U2979) );
  NAND2_X1 U18865 ( .A1(n15268), .A2(n15267), .ZN(n15270) );
  XOR2_X1 U18866 ( .A(n15270), .B(n15269), .Z(n15507) );
  NAND2_X1 U18867 ( .A1(n17379), .A2(n15271), .ZN(n15272) );
  NAND2_X1 U18868 ( .A1(n17416), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15500) );
  OAI211_X1 U18869 ( .C1(n17385), .C2(n15273), .A(n15272), .B(n15500), .ZN(
        n15274) );
  AOI21_X1 U18870 ( .B1(n15275), .B2(n17381), .A(n15274), .ZN(n15276) );
  OAI21_X1 U18871 ( .B1(n20646), .B2(n15507), .A(n15276), .ZN(P1_U2980) );
  NOR2_X1 U18872 ( .A1(n20716), .A2(n21371), .ZN(n15518) );
  NOR2_X1 U18873 ( .A1(n17377), .A2(n15277), .ZN(n15278) );
  AOI211_X1 U18874 ( .C1(n17370), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15518), .B(n15278), .ZN(n15281) );
  OR2_X1 U18875 ( .A1(n15239), .A2(n15279), .ZN(n15509) );
  NAND3_X1 U18876 ( .A1(n15509), .A2(n17382), .A3(n15508), .ZN(n15280) );
  OAI211_X1 U18877 ( .C1(n15282), .C2(n20811), .A(n15281), .B(n15280), .ZN(
        P1_U2981) );
  NOR2_X1 U18878 ( .A1(n9675), .A2(n15300), .ZN(n15284) );
  NAND3_X1 U18879 ( .A1(n15284), .A2(n15351), .A3(n15534), .ZN(n15283) );
  OAI21_X1 U18880 ( .B1(n15284), .B2(n15351), .A(n15283), .ZN(n15285) );
  XNOR2_X1 U18881 ( .A(n15285), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15531) );
  NOR2_X1 U18882 ( .A1(n20716), .A2(n15286), .ZN(n15527) );
  AOI21_X1 U18883 ( .B1(n17370), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15527), .ZN(n15287) );
  OAI21_X1 U18884 ( .B1(n15288), .B2(n17377), .A(n15287), .ZN(n15289) );
  AOI21_X1 U18885 ( .B1(n15290), .B2(n17381), .A(n15289), .ZN(n15291) );
  OAI21_X1 U18886 ( .B1(n15531), .B2(n20646), .A(n15291), .ZN(P1_U2982) );
  INV_X1 U18887 ( .A(n17366), .ZN(n15295) );
  INV_X1 U18888 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15294) );
  OAI21_X1 U18889 ( .B1(n17366), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17364), .ZN(n15293) );
  OAI21_X1 U18890 ( .B1(n15295), .B2(n15294), .A(n15293), .ZN(n15381) );
  OAI21_X1 U18891 ( .B1(n15381), .B2(n9609), .A(n15296), .ZN(n15374) );
  NAND2_X1 U18892 ( .A1(n15374), .A2(n15297), .ZN(n15361) );
  AND2_X2 U18893 ( .A1(n15361), .A2(n15298), .ZN(n15363) );
  INV_X1 U18894 ( .A(n15363), .ZN(n15352) );
  NOR2_X1 U18895 ( .A1(n15352), .A2(n15299), .ZN(n15308) );
  OAI21_X1 U18896 ( .B1(n15308), .B2(n15300), .A(n15309), .ZN(n15301) );
  XOR2_X1 U18897 ( .A(n15302), .B(n15301), .Z(n15542) );
  NAND2_X1 U18898 ( .A1(n17416), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15536) );
  NAND2_X1 U18899 ( .A1(n17370), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15303) );
  OAI211_X1 U18900 ( .C1(n17377), .C2(n15304), .A(n15536), .B(n15303), .ZN(
        n15305) );
  AOI21_X1 U18901 ( .B1(n15306), .B2(n17381), .A(n15305), .ZN(n15307) );
  OAI21_X1 U18902 ( .B1(n15542), .B2(n20646), .A(n15307), .ZN(P1_U2983) );
  NOR2_X1 U18903 ( .A1(n15308), .A2(n9974), .ZN(n15312) );
  NAND2_X1 U18904 ( .A1(n15310), .A2(n15309), .ZN(n15311) );
  XNOR2_X1 U18905 ( .A(n15312), .B(n15311), .ZN(n15550) );
  NOR2_X1 U18906 ( .A1(n20716), .A2(n15313), .ZN(n15547) );
  AOI21_X1 U18907 ( .B1(n17370), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15547), .ZN(n15314) );
  OAI21_X1 U18908 ( .B1(n15315), .B2(n17377), .A(n15314), .ZN(n15316) );
  AOI21_X1 U18909 ( .B1(n15317), .B2(n17381), .A(n15316), .ZN(n15318) );
  OAI21_X1 U18910 ( .B1(n15550), .B2(n20646), .A(n15318), .ZN(P1_U2984) );
  OR2_X1 U18911 ( .A1(n15363), .A2(n15319), .ZN(n15321) );
  AOI22_X1 U18912 ( .A1(n15321), .A2(n15320), .B1(n15351), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15323) );
  XNOR2_X1 U18913 ( .A(n12217), .B(n17394), .ZN(n15322) );
  XNOR2_X1 U18914 ( .A(n15323), .B(n15322), .ZN(n17398) );
  NOR2_X1 U18915 ( .A1(n20716), .A2(n15324), .ZN(n17388) );
  AOI21_X1 U18916 ( .B1(n17370), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17388), .ZN(n15325) );
  OAI21_X1 U18917 ( .B1(n15326), .B2(n17377), .A(n15325), .ZN(n15327) );
  AOI21_X1 U18918 ( .B1(n15328), .B2(n17381), .A(n15327), .ZN(n15329) );
  OAI21_X1 U18919 ( .B1(n17398), .B2(n20646), .A(n15329), .ZN(P1_U2985) );
  INV_X1 U18920 ( .A(n15331), .ZN(n15332) );
  AOI21_X1 U18921 ( .B1(n15363), .B2(n15333), .A(n15332), .ZN(n15344) );
  AND2_X1 U18922 ( .A1(n15334), .A2(n15335), .ZN(n15343) );
  NAND2_X1 U18923 ( .A1(n15344), .A2(n15343), .ZN(n15342) );
  NAND2_X1 U18924 ( .A1(n15342), .A2(n15335), .ZN(n15336) );
  XOR2_X1 U18925 ( .A(n15330), .B(n15336), .Z(n15559) );
  AND2_X1 U18926 ( .A1(n17416), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15553) );
  AOI21_X1 U18927 ( .B1(n17370), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15553), .ZN(n15337) );
  OAI21_X1 U18928 ( .B1(n15338), .B2(n17377), .A(n15337), .ZN(n15339) );
  AOI21_X1 U18929 ( .B1(n15340), .B2(n17381), .A(n15339), .ZN(n15341) );
  OAI21_X1 U18930 ( .B1(n15559), .B2(n20646), .A(n15341), .ZN(P1_U2986) );
  OAI21_X1 U18931 ( .B1(n15344), .B2(n15343), .A(n15342), .ZN(n15560) );
  NAND2_X1 U18932 ( .A1(n15560), .A2(n17382), .ZN(n15349) );
  NOR2_X1 U18933 ( .A1(n20716), .A2(n15345), .ZN(n15568) );
  NOR2_X1 U18934 ( .A1(n17377), .A2(n15346), .ZN(n15347) );
  AOI211_X1 U18935 ( .C1(n17370), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15568), .B(n15347), .ZN(n15348) );
  OAI211_X1 U18936 ( .C1(n20811), .C2(n15350), .A(n15349), .B(n15348), .ZN(
        P1_U2987) );
  NOR3_X1 U18937 ( .A1(n15352), .A2(n15351), .A3(n15362), .ZN(n15353) );
  NOR3_X1 U18938 ( .A1(n15361), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n12217), .ZN(n15366) );
  NOR2_X1 U18939 ( .A1(n15353), .A2(n15366), .ZN(n15354) );
  XNOR2_X1 U18940 ( .A(n15354), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15579) );
  NAND2_X1 U18941 ( .A1(n15579), .A2(n17382), .ZN(n15359) );
  NOR2_X1 U18942 ( .A1(n20716), .A2(n15355), .ZN(n15583) );
  NOR2_X1 U18943 ( .A1(n17377), .A2(n15356), .ZN(n15357) );
  AOI211_X1 U18944 ( .C1(n17370), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15583), .B(n15357), .ZN(n15358) );
  OAI211_X1 U18945 ( .C1(n20811), .C2(n15360), .A(n15359), .B(n15358), .ZN(
        P1_U2988) );
  AND2_X1 U18946 ( .A1(n15361), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15365) );
  XNOR2_X1 U18947 ( .A(n15363), .B(n15362), .ZN(n15364) );
  MUX2_X1 U18948 ( .A(n15365), .B(n15364), .S(n12217), .Z(n15367) );
  NOR2_X1 U18949 ( .A1(n15367), .A2(n15366), .ZN(n15599) );
  NAND2_X1 U18950 ( .A1(n17416), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15593) );
  NAND2_X1 U18951 ( .A1(n17370), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15368) );
  OAI211_X1 U18952 ( .C1(n17377), .C2(n15369), .A(n15593), .B(n15368), .ZN(
        n15370) );
  AOI21_X1 U18953 ( .B1(n15371), .B2(n17381), .A(n15370), .ZN(n15372) );
  OAI21_X1 U18954 ( .B1(n15599), .B2(n20646), .A(n15372), .ZN(P1_U2989) );
  XNOR2_X1 U18955 ( .A(n12217), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15373) );
  XNOR2_X1 U18956 ( .A(n15374), .B(n15373), .ZN(n15601) );
  NAND2_X1 U18957 ( .A1(n15601), .A2(n17382), .ZN(n15378) );
  INV_X1 U18958 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15375) );
  NOR2_X1 U18959 ( .A1(n20716), .A2(n15375), .ZN(n15602) );
  NOR2_X1 U18960 ( .A1(n17385), .A2(n20665), .ZN(n15376) );
  AOI211_X1 U18961 ( .C1(n17379), .C2(n20669), .A(n15602), .B(n15376), .ZN(
        n15377) );
  OAI211_X1 U18962 ( .C1(n20811), .C2(n20668), .A(n15378), .B(n15377), .ZN(
        P1_U2990) );
  XOR2_X1 U18963 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n15379), .Z(
        n15380) );
  XNOR2_X1 U18964 ( .A(n15381), .B(n15380), .ZN(n17405) );
  AOI22_X1 U18965 ( .A1(n17370), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n17416), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15382) );
  OAI21_X1 U18966 ( .B1(n15383), .B2(n17377), .A(n15382), .ZN(n15384) );
  AOI21_X1 U18967 ( .B1(n15385), .B2(n17381), .A(n15384), .ZN(n15386) );
  OAI21_X1 U18968 ( .B1(n17405), .B2(n20646), .A(n15386), .ZN(P1_U2991) );
  INV_X1 U18969 ( .A(n15387), .ZN(n15393) );
  NAND2_X1 U18970 ( .A1(n15394), .A2(n17429), .ZN(n15401) );
  NOR3_X1 U18971 ( .A1(n15396), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10320), .ZN(n15397) );
  AOI211_X1 U18972 ( .C1(n15399), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15398), .B(n15397), .ZN(n15400) );
  OAI211_X1 U18973 ( .C1(n17390), .C2(n15402), .A(n15401), .B(n15400), .ZN(
        P1_U3002) );
  INV_X1 U18974 ( .A(n15413), .ZN(n15403) );
  NAND2_X1 U18975 ( .A1(n15403), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15408) );
  NAND3_X1 U18976 ( .A1(n15417), .A2(n10320), .A3(n15404), .ZN(n15407) );
  INV_X1 U18977 ( .A(n15405), .ZN(n15406) );
  OAI211_X1 U18978 ( .C1(n15423), .C2(n15408), .A(n15407), .B(n15406), .ZN(
        n15409) );
  AOI21_X1 U18979 ( .B1(n15410), .B2(n17424), .A(n15409), .ZN(n15411) );
  OAI21_X1 U18980 ( .B1(n15412), .B2(n17397), .A(n15411), .ZN(P1_U3003) );
  NOR3_X1 U18981 ( .A1(n15423), .A2(n15413), .A3(n15416), .ZN(n15414) );
  AOI211_X1 U18982 ( .C1(n15417), .C2(n15416), .A(n15415), .B(n15414), .ZN(
        n15421) );
  INV_X1 U18983 ( .A(n15418), .ZN(n15419) );
  NAND2_X1 U18984 ( .A1(n15419), .A2(n17424), .ZN(n15420) );
  OAI211_X1 U18985 ( .C1(n15422), .C2(n17397), .A(n15421), .B(n15420), .ZN(
        P1_U3004) );
  INV_X1 U18986 ( .A(n15423), .ZN(n15430) );
  OAI21_X1 U18987 ( .B1(n15452), .B2(n15425), .A(n15424), .ZN(n15429) );
  NOR2_X1 U18988 ( .A1(n15426), .A2(n17390), .ZN(n15427) );
  AOI211_X1 U18989 ( .C1(n15430), .C2(n15429), .A(n15428), .B(n15427), .ZN(
        n15431) );
  OAI21_X1 U18990 ( .B1(n15432), .B2(n17397), .A(n15431), .ZN(P1_U3005) );
  NAND2_X1 U18991 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15434) );
  OAI21_X1 U18992 ( .B1(n15452), .B2(n15434), .A(n15433), .ZN(n15438) );
  NOR2_X1 U18993 ( .A1(n15435), .A2(n17390), .ZN(n15436) );
  AOI211_X1 U18994 ( .C1(n15439), .C2(n15438), .A(n15437), .B(n15436), .ZN(
        n15440) );
  OAI21_X1 U18995 ( .B1(n15441), .B2(n17397), .A(n15440), .ZN(P1_U3006) );
  NAND2_X1 U18996 ( .A1(n15442), .A2(n17429), .ZN(n15449) );
  OAI21_X1 U18997 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15444), .A(
        n15443), .ZN(n15447) );
  NOR3_X1 U18998 ( .A1(n15452), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n12226), .ZN(n15445) );
  AOI211_X1 U18999 ( .C1(n15447), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15446), .B(n15445), .ZN(n15448) );
  OAI211_X1 U19000 ( .C1(n17390), .C2(n15450), .A(n15449), .B(n15448), .ZN(
        P1_U3007) );
  OAI21_X1 U19001 ( .B1(n15452), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15451), .ZN(n15455) );
  NOR2_X1 U19002 ( .A1(n15453), .A2(n17390), .ZN(n15454) );
  AOI211_X1 U19003 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15456), .A(
        n15455), .B(n15454), .ZN(n15457) );
  OAI21_X1 U19004 ( .B1(n15458), .B2(n17397), .A(n15457), .ZN(P1_U3008) );
  INV_X1 U19005 ( .A(n15459), .ZN(n15477) );
  NOR2_X1 U19006 ( .A1(n15488), .A2(n15461), .ZN(n15555) );
  INV_X1 U19007 ( .A(n15466), .ZN(n15468) );
  INV_X1 U19008 ( .A(n15460), .ZN(n15465) );
  INV_X1 U19009 ( .A(n15461), .ZN(n15462) );
  NAND2_X1 U19010 ( .A1(n15462), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15463) );
  OAI22_X1 U19011 ( .A1(n15562), .A2(n15465), .B1(n15464), .B2(n15463), .ZN(
        n15556) );
  INV_X1 U19012 ( .A(n15556), .ZN(n15467) );
  NOR2_X1 U19013 ( .A1(n15467), .A2(n15466), .ZN(n15489) );
  AOI21_X1 U19014 ( .B1(n15555), .B2(n15468), .A(n15489), .ZN(n15499) );
  NAND3_X1 U19015 ( .A1(n15470), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15469), .ZN(n15475) );
  NOR3_X1 U19016 ( .A1(n15499), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15471), .ZN(n15482) );
  INV_X1 U19017 ( .A(n15472), .ZN(n15484) );
  OAI21_X1 U19018 ( .B1(n15482), .B2(n15484), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15474) );
  OAI211_X1 U19019 ( .C1(n15499), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        n15476) );
  AOI21_X1 U19020 ( .B1(n15477), .B2(n17424), .A(n15476), .ZN(n15478) );
  OAI21_X1 U19021 ( .B1(n15479), .B2(n17397), .A(n15478), .ZN(P1_U3009) );
  INV_X1 U19022 ( .A(n15480), .ZN(n15487) );
  NAND2_X1 U19023 ( .A1(n15481), .A2(n17429), .ZN(n15486) );
  AOI211_X1 U19024 ( .C1(n15484), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15483), .B(n15482), .ZN(n15485) );
  OAI211_X1 U19025 ( .C1(n17390), .C2(n15487), .A(n15486), .B(n15485), .ZN(
        P1_U3010) );
  INV_X1 U19026 ( .A(n15488), .ZN(n15615) );
  OAI21_X1 U19027 ( .B1(n15489), .B2(n15615), .A(n15501), .ZN(n15490) );
  AOI21_X1 U19028 ( .B1(n15490), .B2(n15502), .A(n15491), .ZN(n15495) );
  NAND2_X1 U19029 ( .A1(n15491), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15493) );
  OAI21_X1 U19030 ( .B1(n15499), .B2(n15493), .A(n15492), .ZN(n15494) );
  AOI211_X1 U19031 ( .C1(n15496), .C2(n17424), .A(n15495), .B(n15494), .ZN(
        n15497) );
  OAI21_X1 U19032 ( .B1(n15498), .B2(n17397), .A(n15497), .ZN(P1_U3011) );
  NOR2_X1 U19033 ( .A1(n15499), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15504) );
  OAI21_X1 U19034 ( .B1(n15502), .B2(n15501), .A(n15500), .ZN(n15503) );
  AOI211_X1 U19035 ( .C1(n15505), .C2(n17424), .A(n15504), .B(n15503), .ZN(
        n15506) );
  OAI21_X1 U19036 ( .B1(n15507), .B2(n17397), .A(n15506), .ZN(P1_U3012) );
  NAND3_X1 U19037 ( .A1(n15509), .A2(n17429), .A3(n15508), .ZN(n15520) );
  INV_X1 U19038 ( .A(n15510), .ZN(n15511) );
  NAND2_X1 U19039 ( .A1(n17401), .A2(n15511), .ZN(n15512) );
  OAI211_X1 U19040 ( .C1(n15562), .C2(n15513), .A(n15590), .B(n15512), .ZN(
        n17393) );
  INV_X1 U19041 ( .A(n17393), .ZN(n15514) );
  OAI21_X1 U19042 ( .B1(n15515), .B2(n15516), .A(n15514), .ZN(n15529) );
  AND3_X1 U19043 ( .A1(n15535), .A2(n15516), .A3(n12221), .ZN(n15517) );
  AOI211_X1 U19044 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15529), .A(
        n15518), .B(n15517), .ZN(n15519) );
  OAI211_X1 U19045 ( .C1(n17390), .C2(n15521), .A(n15520), .B(n15519), .ZN(
        P1_U3013) );
  INV_X1 U19046 ( .A(n15535), .ZN(n15524) );
  OAI21_X1 U19047 ( .B1(n15524), .B2(n15523), .A(n15522), .ZN(n15528) );
  NOR2_X1 U19048 ( .A1(n15525), .A2(n17390), .ZN(n15526) );
  AOI211_X1 U19049 ( .C1(n15529), .C2(n15528), .A(n15527), .B(n15526), .ZN(
        n15530) );
  OAI21_X1 U19050 ( .B1(n15531), .B2(n17397), .A(n15530), .ZN(P1_U3014) );
  AND2_X1 U19051 ( .A1(n17404), .A2(n17394), .ZN(n15532) );
  NOR2_X1 U19052 ( .A1(n17393), .A2(n15532), .ZN(n15545) );
  AND2_X1 U19053 ( .A1(n15544), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15533) );
  NAND2_X1 U19054 ( .A1(n15535), .A2(n15533), .ZN(n15543) );
  AOI21_X1 U19055 ( .B1(n15545), .B2(n15543), .A(n15534), .ZN(n15539) );
  NAND4_X1 U19056 ( .A1(n15535), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(n15534), .ZN(n15537) );
  NAND2_X1 U19057 ( .A1(n15537), .A2(n15536), .ZN(n15538) );
  AOI211_X1 U19058 ( .C1(n15540), .C2(n17424), .A(n15539), .B(n15538), .ZN(
        n15541) );
  OAI21_X1 U19059 ( .B1(n15542), .B2(n17397), .A(n15541), .ZN(P1_U3015) );
  OAI21_X1 U19060 ( .B1(n15545), .B2(n15544), .A(n15543), .ZN(n15546) );
  AOI211_X1 U19061 ( .C1(n15548), .C2(n17424), .A(n15547), .B(n15546), .ZN(
        n15549) );
  OAI21_X1 U19062 ( .B1(n15550), .B2(n17397), .A(n15549), .ZN(P1_U3016) );
  INV_X1 U19063 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15554) );
  NOR2_X1 U19064 ( .A1(n15551), .A2(n17390), .ZN(n15552) );
  AOI211_X1 U19065 ( .C1(n15555), .C2(n15554), .A(n15553), .B(n15552), .ZN(
        n15558) );
  OAI21_X1 U19066 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15556), .A(
        n17393), .ZN(n15557) );
  OAI211_X1 U19067 ( .C1(n15559), .C2(n17397), .A(n15558), .B(n15557), .ZN(
        P1_U3018) );
  INV_X1 U19068 ( .A(n15560), .ZN(n15576) );
  NOR2_X1 U19069 ( .A1(n15562), .A2(n15572), .ZN(n15563) );
  INV_X1 U19070 ( .A(n15561), .ZN(n15587) );
  OAI21_X1 U19071 ( .B1(n15562), .B2(n15587), .A(n15590), .ZN(n17399) );
  AOI211_X1 U19072 ( .C1(n17401), .C2(n15564), .A(n15563), .B(n17399), .ZN(
        n15581) );
  NAND2_X1 U19073 ( .A1(n15565), .A2(n15580), .ZN(n15566) );
  AOI21_X1 U19074 ( .B1(n15581), .B2(n15566), .A(n15571), .ZN(n15567) );
  AOI211_X1 U19075 ( .C1(n17424), .C2(n15569), .A(n15568), .B(n15567), .ZN(
        n15575) );
  NAND2_X1 U19076 ( .A1(n17422), .A2(n15570), .ZN(n17421) );
  INV_X1 U19077 ( .A(n17421), .ZN(n15573) );
  NAND3_X1 U19078 ( .A1(n15573), .A2(n15572), .A3(n15571), .ZN(n15574) );
  OAI211_X1 U19079 ( .C1(n15576), .C2(n17397), .A(n15575), .B(n15574), .ZN(
        P1_U3019) );
  NOR2_X1 U19080 ( .A1(n17421), .A2(n15577), .ZN(n15600) );
  INV_X1 U19081 ( .A(n15596), .ZN(n15578) );
  NAND2_X1 U19082 ( .A1(n15600), .A2(n15578), .ZN(n17386) );
  NAND2_X1 U19083 ( .A1(n15579), .A2(n17429), .ZN(n15586) );
  NOR2_X1 U19084 ( .A1(n15581), .A2(n15580), .ZN(n15582) );
  AOI211_X1 U19085 ( .C1(n17424), .C2(n15584), .A(n15583), .B(n15582), .ZN(
        n15585) );
  OAI211_X1 U19086 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n17386), .A(
        n15586), .B(n15585), .ZN(P1_U3020) );
  NAND2_X1 U19087 ( .A1(n17401), .A2(n17402), .ZN(n15588) );
  NAND4_X1 U19088 ( .A1(n15590), .A2(n15589), .A3(n15588), .A4(n15587), .ZN(
        n15591) );
  AND2_X1 U19089 ( .A1(n15592), .A2(n15591), .ZN(n15606) );
  OAI21_X1 U19090 ( .B1(n15594), .B2(n17390), .A(n15593), .ZN(n15595) );
  AOI21_X1 U19091 ( .B1(n15606), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15595), .ZN(n15598) );
  OAI211_X1 U19092 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15600), .B(n15596), .ZN(
        n15597) );
  OAI211_X1 U19093 ( .C1(n15599), .C2(n17397), .A(n15598), .B(n15597), .ZN(
        P1_U3021) );
  INV_X1 U19094 ( .A(n15600), .ZN(n15609) );
  NAND2_X1 U19095 ( .A1(n15601), .A2(n17429), .ZN(n15608) );
  INV_X1 U19096 ( .A(n15602), .ZN(n15603) );
  OAI21_X1 U19097 ( .B1(n15604), .B2(n17390), .A(n15603), .ZN(n15605) );
  AOI21_X1 U19098 ( .B1(n15606), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15605), .ZN(n15607) );
  OAI211_X1 U19099 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15609), .A(
        n15608), .B(n15607), .ZN(P1_U3022) );
  NOR2_X1 U19100 ( .A1(n17390), .A2(n15610), .ZN(n15611) );
  AOI211_X1 U19101 ( .C1(n15613), .C2(n17429), .A(n15612), .B(n15611), .ZN(
        n15618) );
  OAI21_X1 U19102 ( .B1(n15615), .B2(n15614), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15616) );
  NAND3_X1 U19103 ( .A1(n15618), .A2(n15617), .A3(n15616), .ZN(P1_U3031) );
  NAND3_X1 U19104 ( .A1(n15620), .A2(n15619), .A3(n17436), .ZN(n17353) );
  NAND2_X1 U19105 ( .A1(n20921), .A2(n15621), .ZN(n15622) );
  OAI211_X1 U19106 ( .C1(n21302), .C2(n20889), .A(n17353), .B(n15622), .ZN(
        n15623) );
  MUX2_X1 U19107 ( .A(n15623), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(
        n20810), .Z(P1_U3478) );
  NAND2_X1 U19108 ( .A1(n15625), .A2(n15624), .ZN(n15630) );
  OAI22_X1 U19109 ( .A1(n17323), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n15630), .B2(n15626), .ZN(n15627) );
  AOI21_X1 U19110 ( .B1(n21273), .B2(n15628), .A(n15627), .ZN(n17325) );
  INV_X1 U19111 ( .A(n15629), .ZN(n15638) );
  INV_X1 U19112 ( .A(n15630), .ZN(n15633) );
  AOI22_X1 U19113 ( .A1(n17358), .A2(n15633), .B1(n15632), .B2(n15631), .ZN(
        n15634) );
  OAI21_X1 U19114 ( .B1(n17325), .B2(n15638), .A(n15634), .ZN(n15635) );
  MUX2_X1 U19115 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15635), .S(
        n15640), .Z(P1_U3473) );
  OAI22_X1 U19116 ( .A1(n15639), .A2(n15638), .B1(n15637), .B2(n15636), .ZN(
        n15641) );
  MUX2_X1 U19117 ( .A(n15642), .B(n15641), .S(n15640), .Z(P1_U3469) );
  OAI21_X1 U19118 ( .B1(n21404), .B2(NA), .A(P1_STATE_REG_1__SCAN_IN), .ZN(
        n15643) );
  INV_X1 U19119 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21515) );
  AOI21_X1 U19120 ( .B1(n15643), .B2(n21515), .A(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n15651) );
  INV_X1 U19121 ( .A(n15644), .ZN(n15645) );
  INV_X1 U19122 ( .A(NA), .ZN(n21362) );
  NOR2_X1 U19123 ( .A1(n15645), .A2(n21362), .ZN(n15649) );
  NOR2_X1 U19124 ( .A1(n15650), .A2(n21515), .ZN(n15646) );
  NOR2_X1 U19125 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n15646), .ZN(n15648) );
  AND2_X1 U19126 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n15647), .ZN(n21368) );
  OAI33_X1 U19127 ( .A1(n21363), .A2(n15651), .A3(n15650), .B1(n15649), .B2(
        n15648), .B3(n21368), .ZN(P1_U3196) );
  AOI211_X1 U19128 ( .C1(n15653), .C2(n20526), .A(n16902), .B(n15652), .ZN(
        n15655) );
  AOI21_X1 U19129 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n16887), .A(n16884), 
        .ZN(n15654) );
  OR2_X1 U19130 ( .A1(n15655), .A2(n15654), .ZN(n15659) );
  NOR2_X1 U19131 ( .A1(n15656), .A2(n20619), .ZN(n16881) );
  NAND2_X1 U19132 ( .A1(n16887), .A2(n19927), .ZN(n15657) );
  OAI211_X1 U19133 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n16881), .A(n19728), 
        .B(n15657), .ZN(n15658) );
  MUX2_X1 U19134 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n15659), .S(n15658), 
        .Z(P2_U3610) );
  AND2_X1 U19135 ( .A1(n15661), .A2(n15660), .ZN(n15662) );
  NOR2_X1 U19136 ( .A1(n15663), .A2(n15662), .ZN(n16461) );
  INV_X1 U19137 ( .A(n16461), .ZN(n15675) );
  INV_X1 U19138 ( .A(n19841), .ZN(n19803) );
  AOI22_X1 U19139 ( .A1(n19830), .A2(P2_EBX_REG_28__SCAN_IN), .B1(n19827), 
        .B2(P2_REIP_REG_28__SCAN_IN), .ZN(n15664) );
  OAI21_X1 U19140 ( .B1(n19803), .B2(n16200), .A(n15664), .ZN(n15669) );
  NAND2_X1 U19141 ( .A1(n15666), .A2(n15665), .ZN(n15667) );
  NOR2_X1 U19142 ( .A1(n16466), .A2(n19776), .ZN(n15668) );
  AOI211_X1 U19143 ( .C1(n19829), .C2(n16196), .A(n15669), .B(n15668), .ZN(
        n15674) );
  AOI21_X1 U19144 ( .B1(n15670), .B2(n10605), .A(n19838), .ZN(n15672) );
  INV_X1 U19145 ( .A(n12521), .ZN(n15671) );
  OAI21_X1 U19146 ( .B1(n19842), .B2(n15672), .A(n15671), .ZN(n15673) );
  OAI211_X1 U19147 ( .C1(n19833), .C2(n15675), .A(n15674), .B(n15673), .ZN(
        P2_U2827) );
  AOI22_X1 U19148 ( .A1(n19830), .A2(P2_EBX_REG_27__SCAN_IN), .B1(n19827), 
        .B2(P2_REIP_REG_27__SCAN_IN), .ZN(n15677) );
  NAND2_X1 U19149 ( .A1(n19841), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15676) );
  OAI211_X1 U19150 ( .C1(n16194), .C2(n19809), .A(n15677), .B(n15676), .ZN(
        n15682) );
  OAI21_X1 U19151 ( .B1(n15688), .B2(n16207), .A(n19820), .ZN(n15680) );
  INV_X1 U19152 ( .A(n15670), .ZN(n15679) );
  AOI21_X1 U19153 ( .B1(n17314), .B2(n15680), .A(n15679), .ZN(n15681) );
  AOI211_X1 U19154 ( .C1(n19836), .C2(n16210), .A(n15682), .B(n15681), .ZN(
        n15683) );
  OAI21_X1 U19155 ( .B1(n16094), .B2(n19833), .A(n15683), .ZN(P2_U2828) );
  OAI21_X1 U19156 ( .B1(n15684), .B2(n15686), .A(n15685), .ZN(n16473) );
  OAI21_X1 U19157 ( .B1(n9646), .B2(n15687), .A(n11732), .ZN(n16481) );
  INV_X1 U19158 ( .A(n16481), .ZN(n15696) );
  AOI21_X1 U19159 ( .B1(n15706), .B2(n16218), .A(n19838), .ZN(n15690) );
  INV_X1 U19160 ( .A(n15688), .ZN(n15689) );
  OAI21_X1 U19161 ( .B1(n19842), .B2(n15690), .A(n15689), .ZN(n15693) );
  OAI22_X1 U19162 ( .A1(n19773), .A2(n16001), .B1(n20588), .B2(n19804), .ZN(
        n15691) );
  AOI21_X1 U19163 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19841), .A(
        n15691), .ZN(n15692) );
  OAI211_X1 U19164 ( .C1(n19809), .C2(n15694), .A(n15693), .B(n15692), .ZN(
        n15695) );
  AOI21_X1 U19165 ( .B1(n15696), .B2(n19836), .A(n15695), .ZN(n15697) );
  OAI21_X1 U19166 ( .B1(n16473), .B2(n19833), .A(n15697), .ZN(P2_U2829) );
  INV_X1 U19167 ( .A(n15684), .ZN(n15698) );
  OAI21_X1 U19168 ( .B1(n9644), .B2(n15699), .A(n15698), .ZN(n16486) );
  AND2_X1 U19169 ( .A1(n15717), .A2(n15700), .ZN(n15701) );
  OR2_X1 U19170 ( .A1(n15701), .A2(n9646), .ZN(n16492) );
  INV_X1 U19171 ( .A(n16492), .ZN(n15711) );
  OAI22_X1 U19172 ( .A1(n19773), .A2(n16006), .B1(n20586), .B2(n19804), .ZN(
        n15702) );
  AOI21_X1 U19173 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19841), .A(
        n15702), .ZN(n15703) );
  OAI21_X1 U19174 ( .B1(n15704), .B2(n19809), .A(n15703), .ZN(n15710) );
  OAI21_X1 U19175 ( .B1(n15705), .B2(n16229), .A(n19820), .ZN(n15708) );
  INV_X1 U19176 ( .A(n15706), .ZN(n15707) );
  AOI21_X1 U19177 ( .B1(n17314), .B2(n15708), .A(n15707), .ZN(n15709) );
  AOI211_X1 U19178 ( .C1(n15711), .C2(n19836), .A(n15710), .B(n15709), .ZN(
        n15712) );
  OAI21_X1 U19179 ( .B1(n16486), .B2(n19833), .A(n15712), .ZN(P2_U2830) );
  AND2_X1 U19180 ( .A1(n15713), .A2(n15714), .ZN(n15715) );
  OR2_X1 U19181 ( .A1(n15715), .A2(n9644), .ZN(n16497) );
  INV_X1 U19182 ( .A(n15717), .ZN(n15718) );
  AOI21_X1 U19183 ( .B1(n15719), .B2(n15716), .A(n15718), .ZN(n16505) );
  AOI21_X1 U19184 ( .B1(n15735), .B2(n16236), .A(n19838), .ZN(n15721) );
  INV_X1 U19185 ( .A(n15705), .ZN(n15720) );
  OAI21_X1 U19186 ( .B1(n19842), .B2(n15721), .A(n15720), .ZN(n15724) );
  INV_X1 U19187 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20584) );
  OAI22_X1 U19188 ( .A1(n19773), .A2(n11774), .B1(n20584), .B2(n19804), .ZN(
        n15722) );
  AOI21_X1 U19189 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19841), .A(
        n15722), .ZN(n15723) );
  OAI211_X1 U19190 ( .C1(n19809), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        n15726) );
  AOI21_X1 U19191 ( .B1(n16505), .B2(n19836), .A(n15726), .ZN(n15727) );
  OAI21_X1 U19192 ( .B1(n16497), .B2(n19833), .A(n15727), .ZN(P2_U2831) );
  NAND2_X1 U19193 ( .A1(n16125), .A2(n15729), .ZN(n15730) );
  AND2_X1 U19194 ( .A1(n15713), .A2(n15730), .ZN(n16518) );
  OR2_X1 U19195 ( .A1(n15731), .A2(n15732), .ZN(n15733) );
  AND2_X1 U19196 ( .A1(n15716), .A2(n15733), .ZN(n16517) );
  OAI21_X1 U19197 ( .B1(n15734), .B2(n16246), .A(n19820), .ZN(n15737) );
  INV_X1 U19198 ( .A(n15735), .ZN(n15736) );
  AOI21_X1 U19199 ( .B1(n17314), .B2(n15737), .A(n15736), .ZN(n15743) );
  INV_X1 U19200 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20582) );
  OAI22_X1 U19201 ( .A1(n19773), .A2(n15738), .B1(n20582), .B2(n19804), .ZN(
        n15739) );
  AOI21_X1 U19202 ( .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19841), .A(
        n15739), .ZN(n15740) );
  OAI21_X1 U19203 ( .B1(n15741), .B2(n19809), .A(n15740), .ZN(n15742) );
  AOI211_X1 U19204 ( .C1(n16517), .C2(n19836), .A(n15743), .B(n15742), .ZN(
        n15744) );
  OAI21_X1 U19205 ( .B1(n19833), .B2(n16122), .A(n15744), .ZN(P2_U2832) );
  AOI21_X1 U19206 ( .B1(n15746), .B2(n11795), .A(n15745), .ZN(n16546) );
  INV_X1 U19207 ( .A(n16546), .ZN(n16138) );
  AOI21_X1 U19208 ( .B1(n15749), .B2(n15748), .A(n15747), .ZN(n16270) );
  NOR2_X1 U19209 ( .A1(n15750), .A2(n19809), .ZN(n15757) );
  OAI21_X1 U19210 ( .B1(n15763), .B2(n16266), .A(n19820), .ZN(n15751) );
  NAND2_X1 U19211 ( .A1(n17314), .A2(n15751), .ZN(n15752) );
  NAND2_X1 U19212 ( .A1(n17309), .A2(n15752), .ZN(n15754) );
  AOI22_X1 U19213 ( .A1(n19830), .A2(P2_EBX_REG_21__SCAN_IN), .B1(n19827), 
        .B2(P2_REIP_REG_21__SCAN_IN), .ZN(n15753) );
  OAI211_X1 U19214 ( .C1(n19803), .C2(n15755), .A(n15754), .B(n15753), .ZN(
        n15756) );
  AOI211_X1 U19215 ( .C1(n16270), .C2(n19836), .A(n15757), .B(n15756), .ZN(
        n15758) );
  OAI21_X1 U19216 ( .B1(n16138), .B2(n19833), .A(n15758), .ZN(P2_U2834) );
  AOI22_X1 U19217 ( .A1(n19830), .A2(P2_EBX_REG_20__SCAN_IN), .B1(n19827), 
        .B2(P2_REIP_REG_20__SCAN_IN), .ZN(n15760) );
  NAND2_X1 U19218 ( .A1(n19841), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15759) );
  OAI211_X1 U19219 ( .C1(n17314), .C2(n15761), .A(n15760), .B(n15759), .ZN(
        n15767) );
  INV_X1 U19220 ( .A(n15761), .ZN(n15765) );
  INV_X1 U19221 ( .A(n15762), .ZN(n15764) );
  INV_X1 U19222 ( .A(n15952), .ZN(n15844) );
  AOI211_X1 U19223 ( .C1(n15765), .C2(n15764), .A(n15763), .B(n15844), .ZN(
        n15766) );
  AOI211_X1 U19224 ( .C1(n19829), .C2(n15768), .A(n15767), .B(n15766), .ZN(
        n15770) );
  NAND2_X1 U19225 ( .A1(n16139), .A2(n19812), .ZN(n15769) );
  OAI211_X1 U19226 ( .C1(n19776), .C2(n16034), .A(n15770), .B(n15769), .ZN(
        P2_U2835) );
  INV_X1 U19227 ( .A(n16276), .ZN(n15781) );
  INV_X1 U19228 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20575) );
  OAI21_X1 U19229 ( .B1(n19804), .B2(n20575), .A(n10176), .ZN(n15771) );
  AOI21_X1 U19230 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19830), .A(n15771), .ZN(
        n15773) );
  NAND2_X1 U19231 ( .A1(n19841), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15772) );
  OAI211_X1 U19232 ( .C1(n15774), .C2(n19809), .A(n15773), .B(n15772), .ZN(
        n15780) );
  INV_X1 U19233 ( .A(n16288), .ZN(n15786) );
  AND2_X1 U19234 ( .A1(n15968), .A2(n15775), .ZN(n15787) );
  NAND2_X1 U19235 ( .A1(n15787), .A2(n19820), .ZN(n15804) );
  OAI21_X1 U19236 ( .B1(n15844), .B2(n15786), .A(n15804), .ZN(n15778) );
  OAI21_X1 U19237 ( .B1(n15776), .B2(n19838), .A(n17314), .ZN(n15777) );
  MUX2_X1 U19238 ( .A(n15778), .B(n15777), .S(n16273), .Z(n15779) );
  AOI211_X1 U19239 ( .C1(n19836), .C2(n15781), .A(n15780), .B(n15779), .ZN(
        n15782) );
  OAI21_X1 U19240 ( .B1(n16151), .B2(n19833), .A(n15782), .ZN(P2_U2836) );
  OR2_X1 U19241 ( .A1(n15783), .A2(n15784), .ZN(n15785) );
  NAND2_X1 U19242 ( .A1(n11700), .A2(n15785), .ZN(n16552) );
  XNOR2_X1 U19243 ( .A(n15787), .B(n15786), .ZN(n15797) );
  AND2_X1 U19244 ( .A1(n15788), .A2(n15789), .ZN(n15790) );
  OR2_X1 U19245 ( .A1(n15790), .A2(n9653), .ZN(n16558) );
  OAI21_X1 U19246 ( .B1(n19804), .B2(n20573), .A(n10176), .ZN(n15791) );
  AOI21_X1 U19247 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n19830), .A(n15791), .ZN(
        n15792) );
  OAI21_X1 U19248 ( .B1(n16285), .B2(n19803), .A(n15792), .ZN(n15793) );
  AOI21_X1 U19249 ( .B1(n15794), .B2(n19829), .A(n15793), .ZN(n15795) );
  OAI21_X1 U19250 ( .B1(n16558), .B2(n19776), .A(n15795), .ZN(n15796) );
  AOI21_X1 U19251 ( .B1(n19820), .B2(n15797), .A(n15796), .ZN(n15798) );
  OAI21_X1 U19252 ( .B1(n16552), .B2(n19833), .A(n15798), .ZN(P2_U2837) );
  NOR2_X1 U19253 ( .A1(n9635), .A2(n15799), .ZN(n15800) );
  OR2_X1 U19254 ( .A1(n15783), .A2(n15800), .ZN(n16573) );
  NAND2_X1 U19255 ( .A1(n15821), .A2(n15802), .ZN(n15803) );
  INV_X1 U19256 ( .A(n15804), .ZN(n15805) );
  OAI21_X1 U19257 ( .B1(n15806), .B2(n16294), .A(n15805), .ZN(n15813) );
  AOI21_X1 U19258 ( .B1(n19827), .B2(P2_REIP_REG_17__SCAN_IN), .A(n16423), 
        .ZN(n15807) );
  OAI21_X1 U19259 ( .B1(n19773), .B2(n15808), .A(n15807), .ZN(n15811) );
  NOR2_X1 U19260 ( .A1(n15809), .A2(n19809), .ZN(n15810) );
  AOI211_X1 U19261 ( .C1(n19841), .C2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15811), .B(n15810), .ZN(n15812) );
  OAI211_X1 U19262 ( .C1(n17314), .C2(n16294), .A(n15813), .B(n15812), .ZN(
        n15814) );
  AOI21_X1 U19263 ( .B1(n16571), .B2(n19836), .A(n15814), .ZN(n15815) );
  OAI21_X1 U19264 ( .B1(n16573), .B2(n19833), .A(n15815), .ZN(P2_U2838) );
  NAND2_X1 U19265 ( .A1(n15968), .A2(n15816), .ZN(n15818) );
  INV_X1 U19266 ( .A(n15817), .ZN(n16302) );
  XNOR2_X1 U19267 ( .A(n15818), .B(n16302), .ZN(n15834) );
  AOI21_X1 U19268 ( .B1(n15822), .B2(n15820), .A(n15801), .ZN(n19851) );
  AOI21_X1 U19269 ( .B1(n19827), .B2(P2_REIP_REG_16__SCAN_IN), .A(n16423), 
        .ZN(n15823) );
  OAI21_X1 U19270 ( .B1(n19773), .B2(n15824), .A(n15823), .ZN(n15825) );
  AOI21_X1 U19271 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19841), .A(
        n15825), .ZN(n15826) );
  OAI21_X1 U19272 ( .B1(n15827), .B2(n19809), .A(n15826), .ZN(n15828) );
  AOI21_X1 U19273 ( .B1(n19851), .B2(n19836), .A(n15828), .ZN(n15833) );
  AND2_X1 U19274 ( .A1(n15830), .A2(n15829), .ZN(n15831) );
  NOR2_X1 U19275 ( .A1(n9635), .A2(n15831), .ZN(n19871) );
  NAND2_X1 U19276 ( .A1(n19871), .A2(n19812), .ZN(n15832) );
  OAI211_X1 U19277 ( .C1(n19838), .C2(n15834), .A(n15833), .B(n15832), .ZN(
        P2_U2839) );
  OR2_X1 U19278 ( .A1(n14614), .A2(n15835), .ZN(n15836) );
  NAND2_X1 U19279 ( .A1(n15820), .A2(n15836), .ZN(n16591) );
  AOI21_X1 U19280 ( .B1(n19827), .B2(P2_REIP_REG_15__SCAN_IN), .A(n16423), 
        .ZN(n15837) );
  OAI21_X1 U19281 ( .B1(n19773), .B2(n15838), .A(n15837), .ZN(n15841) );
  NOR2_X1 U19282 ( .A1(n15839), .A2(n19809), .ZN(n15840) );
  AOI211_X1 U19283 ( .C1(n19841), .C2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15841), .B(n15840), .ZN(n15842) );
  OAI21_X1 U19284 ( .B1(n16591), .B2(n19776), .A(n15842), .ZN(n15849) );
  NOR2_X1 U19285 ( .A1(n19815), .A2(n15843), .ZN(n15851) );
  NAND2_X1 U19286 ( .A1(n15851), .A2(n19820), .ZN(n15868) );
  OAI21_X1 U19287 ( .B1(n15844), .B2(n16318), .A(n15868), .ZN(n15847) );
  OAI21_X1 U19288 ( .B1(n15845), .B2(n19838), .A(n17314), .ZN(n15846) );
  MUX2_X1 U19289 ( .A(n15847), .B(n15846), .S(n16314), .Z(n15848) );
  AOI211_X1 U19290 ( .C1(n16588), .C2(n19812), .A(n15849), .B(n15848), .ZN(
        n15850) );
  INV_X1 U19291 ( .A(n15850), .ZN(P2_U2840) );
  XOR2_X1 U19292 ( .A(n16318), .B(n15851), .Z(n15860) );
  INV_X1 U19293 ( .A(n16601), .ZN(n16321) );
  AOI21_X1 U19294 ( .B1(n19827), .B2(P2_REIP_REG_14__SCAN_IN), .A(n16423), 
        .ZN(n15852) );
  OAI21_X1 U19295 ( .B1(n19773), .B2(n15853), .A(n15852), .ZN(n15854) );
  AOI21_X1 U19296 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19841), .A(
        n15854), .ZN(n15855) );
  OAI21_X1 U19297 ( .B1(n15856), .B2(n19809), .A(n15855), .ZN(n15858) );
  NOR2_X1 U19298 ( .A1(n16599), .A2(n19833), .ZN(n15857) );
  AOI211_X1 U19299 ( .C1(n19836), .C2(n16321), .A(n15858), .B(n15857), .ZN(
        n15859) );
  OAI21_X1 U19300 ( .B1(n15860), .B2(n19838), .A(n15859), .ZN(P2_U2841) );
  AOI21_X1 U19301 ( .B1(n19827), .B2(P2_REIP_REG_13__SCAN_IN), .A(n16423), 
        .ZN(n15861) );
  OAI21_X1 U19302 ( .B1(n19773), .B2(n15862), .A(n15861), .ZN(n15863) );
  AOI21_X1 U19303 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19841), .A(
        n15863), .ZN(n15864) );
  OAI21_X1 U19304 ( .B1(n15865), .B2(n19809), .A(n15864), .ZN(n15867) );
  NOR2_X1 U19305 ( .A1(n17314), .A2(n16338), .ZN(n15866) );
  AOI211_X1 U19306 ( .C1(n19836), .C2(n16611), .A(n15867), .B(n15866), .ZN(
        n15872) );
  INV_X1 U19307 ( .A(n15868), .ZN(n15869) );
  OAI21_X1 U19308 ( .B1(n15870), .B2(n16338), .A(n15869), .ZN(n15871) );
  OAI211_X1 U19309 ( .C1(n19833), .C2(n16614), .A(n15872), .B(n15871), .ZN(
        P2_U2842) );
  INV_X1 U19310 ( .A(n19765), .ZN(n19762) );
  NOR2_X1 U19311 ( .A1(n19763), .A2(n19762), .ZN(n15873) );
  NOR2_X1 U19312 ( .A1(n19815), .A2(n15873), .ZN(n19764) );
  XOR2_X1 U19313 ( .A(n16348), .B(n19764), .Z(n15884) );
  OAI21_X1 U19314 ( .B1(n15874), .B2(n15875), .A(n14607), .ZN(n16625) );
  AOI21_X1 U19315 ( .B1(n19827), .B2(P2_REIP_REG_12__SCAN_IN), .A(n16423), 
        .ZN(n15876) );
  OAI21_X1 U19316 ( .B1(n19773), .B2(n15877), .A(n15876), .ZN(n15880) );
  NOR2_X1 U19317 ( .A1(n15878), .A2(n19809), .ZN(n15879) );
  AOI211_X1 U19318 ( .C1(n19841), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15880), .B(n15879), .ZN(n15881) );
  OAI21_X1 U19319 ( .B1(n16625), .B2(n19776), .A(n15881), .ZN(n15882) );
  AOI21_X1 U19320 ( .B1(n16628), .B2(n19812), .A(n15882), .ZN(n15883) );
  OAI21_X1 U19321 ( .B1(n15884), .B2(n19838), .A(n15883), .ZN(P2_U2843) );
  NAND2_X1 U19322 ( .A1(n15952), .A2(n15885), .ZN(n15887) );
  INV_X1 U19323 ( .A(n15885), .ZN(n19781) );
  AOI21_X1 U19324 ( .B1(n19781), .B2(n19820), .A(n19842), .ZN(n15886) );
  MUX2_X1 U19325 ( .A(n15887), .B(n15886), .S(n16367), .Z(n15898) );
  AND2_X1 U19326 ( .A1(n15890), .A2(n15889), .ZN(n15891) );
  NOR2_X1 U19327 ( .A1(n15888), .A2(n15891), .ZN(n19858) );
  NAND2_X1 U19328 ( .A1(n15892), .A2(n19829), .ZN(n15895) );
  NOR2_X1 U19329 ( .A1(n19773), .A2(n10531), .ZN(n15893) );
  AOI211_X1 U19330 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19827), .A(n16423), 
        .B(n15893), .ZN(n15894) );
  OAI211_X1 U19331 ( .C1(n19803), .C2(n10418), .A(n15895), .B(n15894), .ZN(
        n15896) );
  AOI21_X1 U19332 ( .B1(n19858), .B2(n19836), .A(n15896), .ZN(n15897) );
  OAI211_X1 U19333 ( .C1(n19833), .C2(n16653), .A(n15898), .B(n15897), .ZN(
        P2_U2845) );
  NOR2_X1 U19334 ( .A1(n19815), .A2(n15899), .ZN(n15900) );
  XOR2_X1 U19335 ( .A(n16394), .B(n15900), .Z(n15909) );
  AOI21_X1 U19336 ( .B1(n19827), .B2(P2_REIP_REG_8__SCAN_IN), .A(n16423), .ZN(
        n15901) );
  OAI21_X1 U19337 ( .B1(n19773), .B2(n15902), .A(n15901), .ZN(n15903) );
  AOI21_X1 U19338 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19841), .A(
        n15903), .ZN(n15904) );
  OAI21_X1 U19339 ( .B1(n15905), .B2(n19809), .A(n15904), .ZN(n15907) );
  NOR2_X1 U19340 ( .A1(n16681), .A2(n19833), .ZN(n15906) );
  AOI211_X1 U19341 ( .C1(n16678), .C2(n19836), .A(n15907), .B(n15906), .ZN(
        n15908) );
  OAI21_X1 U19342 ( .B1(n15909), .B2(n19838), .A(n15908), .ZN(P2_U2847) );
  NAND2_X1 U19343 ( .A1(n15952), .A2(n15910), .ZN(n15913) );
  INV_X1 U19344 ( .A(n15910), .ZN(n15911) );
  AOI21_X1 U19345 ( .B1(n15911), .B2(n19820), .A(n19842), .ZN(n15912) );
  MUX2_X1 U19346 ( .A(n15913), .B(n15912), .S(n16405), .Z(n15920) );
  INV_X1 U19347 ( .A(n16407), .ZN(n16692) );
  NAND2_X1 U19348 ( .A1(n19830), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n15914) );
  OAI211_X1 U19349 ( .C1(n20552), .C2(n19804), .A(n15914), .B(n10176), .ZN(
        n15915) );
  AOI21_X1 U19350 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19841), .A(
        n15915), .ZN(n15916) );
  OAI21_X1 U19351 ( .B1(n15917), .B2(n19809), .A(n15916), .ZN(n15918) );
  AOI21_X1 U19352 ( .B1(n16692), .B2(n19836), .A(n15918), .ZN(n15919) );
  OAI211_X1 U19353 ( .C1(n16689), .C2(n19833), .A(n15920), .B(n15919), .ZN(
        P2_U2848) );
  INV_X1 U19354 ( .A(n15921), .ZN(n19796) );
  AOI21_X1 U19355 ( .B1(n19796), .B2(n19820), .A(n19842), .ZN(n15924) );
  NAND2_X1 U19356 ( .A1(n15952), .A2(n15921), .ZN(n15923) );
  MUX2_X1 U19357 ( .A(n15924), .B(n15923), .S(n15922), .Z(n15931) );
  OAI21_X1 U19358 ( .B1(n19804), .B2(n20550), .A(n10176), .ZN(n15925) );
  AOI21_X1 U19359 ( .B1(P2_EBX_REG_6__SCAN_IN), .B2(n19830), .A(n15925), .ZN(
        n15926) );
  OAI21_X1 U19360 ( .B1(n21556), .B2(n19803), .A(n15926), .ZN(n15928) );
  NOR2_X1 U19361 ( .A1(n16703), .A2(n19776), .ZN(n15927) );
  AOI211_X1 U19362 ( .C1(n19829), .C2(n15929), .A(n15928), .B(n15927), .ZN(
        n15930) );
  OAI211_X1 U19363 ( .C1(n15932), .C2(n19833), .A(n15931), .B(n15930), .ZN(
        P2_U2849) );
  NAND2_X1 U19364 ( .A1(n15952), .A2(n15933), .ZN(n15936) );
  INV_X1 U19365 ( .A(n15933), .ZN(n15934) );
  AOI21_X1 U19366 ( .B1(n15934), .B2(n19820), .A(n19842), .ZN(n15935) );
  MUX2_X1 U19367 ( .A(n15936), .B(n15935), .S(n16451), .Z(n15950) );
  NAND2_X1 U19368 ( .A1(n15939), .A2(n15938), .ZN(n15940) );
  AND2_X1 U19369 ( .A1(n15937), .A2(n15940), .ZN(n20607) );
  NAND2_X1 U19370 ( .A1(n15941), .A2(n19836), .ZN(n15947) );
  AOI22_X1 U19371 ( .A1(n19830), .A2(P2_EBX_REG_3__SCAN_IN), .B1(n19827), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n15946) );
  INV_X1 U19372 ( .A(n15942), .ZN(n15943) );
  NAND2_X1 U19373 ( .A1(n19829), .A2(n15943), .ZN(n15945) );
  NAND2_X1 U19374 ( .A1(n19841), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15944) );
  NAND4_X1 U19375 ( .A1(n15947), .A2(n15946), .A3(n15945), .A4(n15944), .ZN(
        n15948) );
  AOI21_X1 U19376 ( .B1(n19812), .B2(n20607), .A(n15948), .ZN(n15949) );
  OAI211_X1 U19377 ( .C1(n16775), .C2(n19837), .A(n15950), .B(n15949), .ZN(
        P2_U2852) );
  AOI21_X1 U19378 ( .B1(n15966), .B2(n19820), .A(n19842), .ZN(n15955) );
  INV_X1 U19379 ( .A(n15966), .ZN(n15951) );
  NAND2_X1 U19380 ( .A1(n15952), .A2(n15951), .ZN(n15954) );
  MUX2_X1 U19381 ( .A(n15955), .B(n15954), .S(n15953), .Z(n15962) );
  AOI22_X1 U19382 ( .A1(n19830), .A2(P2_EBX_REG_2__SCAN_IN), .B1(n19827), .B2(
        P2_REIP_REG_2__SCAN_IN), .ZN(n15957) );
  NAND2_X1 U19383 ( .A1(n19841), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15956) );
  OAI211_X1 U19384 ( .C1(n19809), .C2(n15958), .A(n15957), .B(n15956), .ZN(
        n15960) );
  NOR2_X1 U19385 ( .A1(n16768), .A2(n19776), .ZN(n15959) );
  AOI211_X1 U19386 ( .C1(n19812), .C2(n19890), .A(n15960), .B(n15959), .ZN(
        n15961) );
  OAI211_X1 U19387 ( .C1(n16799), .C2(n19837), .A(n15962), .B(n15961), .ZN(
        P2_U2853) );
  AND2_X1 U19388 ( .A1(n15964), .A2(n15963), .ZN(n15965) );
  NOR2_X1 U19389 ( .A1(n15966), .A2(n15965), .ZN(n15967) );
  NAND2_X1 U19390 ( .A1(n15968), .A2(n15967), .ZN(n16751) );
  OAI22_X1 U19391 ( .A1(n19809), .A2(n15969), .B1(n19804), .B2(n20542), .ZN(
        n15970) );
  AOI21_X1 U19392 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n19830), .A(n15970), .ZN(
        n15972) );
  NAND2_X1 U19393 ( .A1(n19812), .A2(n19959), .ZN(n15971) );
  OAI211_X1 U19394 ( .C1(n19965), .C2(n19776), .A(n15972), .B(n15971), .ZN(
        n15973) );
  AOI21_X1 U19395 ( .B1(n16797), .B2(n19813), .A(n15973), .ZN(n15975) );
  MUX2_X1 U19396 ( .A(n17314), .B(n19803), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15974) );
  OAI211_X1 U19397 ( .C1(n16751), .C2(n19838), .A(n15975), .B(n15974), .ZN(
        P2_U2854) );
  NOR2_X1 U19398 ( .A1(n15976), .A2(n16065), .ZN(n15977) );
  AOI21_X1 U19399 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16065), .A(n15977), .ZN(
        n15978) );
  OAI21_X1 U19400 ( .B1(n15979), .B2(n19855), .A(n15978), .ZN(P2_U2857) );
  INV_X1 U19401 ( .A(n15980), .ZN(n16073) );
  NAND2_X1 U19402 ( .A1(n15982), .A2(n15981), .ZN(n16072) );
  NAND3_X1 U19403 ( .A1(n16073), .A2(n19863), .A3(n16072), .ZN(n15984) );
  NAND2_X1 U19404 ( .A1(n16065), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15983) );
  OAI211_X1 U19405 ( .C1(n16184), .C2(n16065), .A(n15984), .B(n15983), .ZN(
        P2_U2858) );
  NAND2_X1 U19406 ( .A1(n13269), .A2(n15985), .ZN(n15987) );
  XNOR2_X1 U19407 ( .A(n15987), .B(n15986), .ZN(n16087) );
  NOR2_X1 U19408 ( .A1(n16466), .A2(n16065), .ZN(n15988) );
  AOI21_X1 U19409 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16065), .A(n15988), .ZN(
        n15989) );
  OAI21_X1 U19410 ( .B1(n16087), .B2(n19855), .A(n15989), .ZN(P2_U2859) );
  INV_X1 U19411 ( .A(n16210), .ZN(n15994) );
  NAND2_X1 U19412 ( .A1(n9688), .A2(n19863), .ZN(n15993) );
  NAND2_X1 U19413 ( .A1(n16065), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15992) );
  OAI211_X1 U19414 ( .C1(n15994), .C2(n16065), .A(n15993), .B(n15992), .ZN(
        P2_U2860) );
  NAND2_X1 U19415 ( .A1(n16005), .A2(n16004), .ZN(n16003) );
  NAND2_X1 U19416 ( .A1(n15995), .A2(n16003), .ZN(n16000) );
  NOR2_X1 U19417 ( .A1(n11232), .A2(n15996), .ZN(n15997) );
  XNOR2_X1 U19418 ( .A(n15998), .B(n15997), .ZN(n15999) );
  XNOR2_X1 U19419 ( .A(n16000), .B(n15999), .ZN(n16101) );
  MUX2_X1 U19420 ( .A(n16001), .B(n16481), .S(n19866), .Z(n16002) );
  OAI21_X1 U19421 ( .B1(n16101), .B2(n19855), .A(n16002), .ZN(P2_U2861) );
  OAI21_X1 U19422 ( .B1(n16005), .B2(n16004), .A(n16003), .ZN(n16108) );
  MUX2_X1 U19423 ( .A(n16492), .B(n16006), .S(n16065), .Z(n16007) );
  OAI21_X1 U19424 ( .B1(n19855), .B2(n16108), .A(n16007), .ZN(P2_U2862) );
  AOI21_X1 U19425 ( .B1(n9680), .B2(n16009), .A(n16008), .ZN(n16010) );
  XOR2_X1 U19426 ( .A(n16011), .B(n16010), .Z(n16115) );
  NAND2_X1 U19427 ( .A1(n16505), .A2(n19866), .ZN(n16013) );
  NAND2_X1 U19428 ( .A1(n16065), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16012) );
  OAI211_X1 U19429 ( .C1(n16115), .C2(n19855), .A(n16013), .B(n16012), .ZN(
        P2_U2863) );
  INV_X1 U19430 ( .A(n16517), .ZN(n16019) );
  AOI21_X1 U19431 ( .B1(n16016), .B2(n16015), .A(n16014), .ZN(n16120) );
  NAND2_X1 U19432 ( .A1(n16120), .A2(n19863), .ZN(n16018) );
  NAND2_X1 U19433 ( .A1(n16065), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16017) );
  OAI211_X1 U19434 ( .C1(n16019), .C2(n16065), .A(n16018), .B(n16017), .ZN(
        P2_U2864) );
  NOR2_X1 U19435 ( .A1(n15747), .A2(n16020), .ZN(n16021) );
  OR2_X1 U19436 ( .A1(n15731), .A2(n16021), .ZN(n17304) );
  AOI21_X1 U19437 ( .B1(n16022), .B2(n16024), .A(n9649), .ZN(n16129) );
  AOI22_X1 U19438 ( .A1(n16129), .A2(n19863), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n16065), .ZN(n16023) );
  OAI21_X1 U19439 ( .B1(n17304), .B2(n16065), .A(n16023), .ZN(P2_U2865) );
  INV_X1 U19440 ( .A(n16270), .ZN(n16543) );
  OAI21_X1 U19441 ( .B1(n16031), .B2(n16025), .A(n16024), .ZN(n16026) );
  INV_X1 U19442 ( .A(n16026), .ZN(n16136) );
  AOI22_X1 U19443 ( .A1(n16136), .A2(n19863), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n16065), .ZN(n16027) );
  OAI21_X1 U19444 ( .B1(n16543), .B2(n16065), .A(n16027), .ZN(P2_U2866) );
  INV_X1 U19445 ( .A(n16029), .ZN(n16045) );
  NOR2_X1 U19446 ( .A1(n16028), .A2(n16045), .ZN(n16046) );
  NAND2_X1 U19447 ( .A1(n16046), .A2(n16042), .ZN(n16041) );
  INV_X1 U19448 ( .A(n16030), .ZN(n16038) );
  NOR2_X1 U19449 ( .A1(n16041), .A2(n16038), .ZN(n16037) );
  INV_X1 U19450 ( .A(n16031), .ZN(n16032) );
  OAI21_X1 U19451 ( .B1(n16037), .B2(n16033), .A(n16032), .ZN(n16144) );
  MUX2_X1 U19452 ( .A(n16035), .B(n16034), .S(n19866), .Z(n16036) );
  OAI21_X1 U19453 ( .B1(n19855), .B2(n16144), .A(n16036), .ZN(P2_U2867) );
  AOI21_X1 U19454 ( .B1(n16038), .B2(n16041), .A(n16037), .ZN(n16149) );
  NAND2_X1 U19455 ( .A1(n16149), .A2(n19863), .ZN(n16040) );
  NAND2_X1 U19456 ( .A1(n16065), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n16039) );
  OAI211_X1 U19457 ( .C1(n16276), .C2(n16065), .A(n16040), .B(n16039), .ZN(
        P2_U2868) );
  OAI21_X1 U19458 ( .B1(n16046), .B2(n16042), .A(n16041), .ZN(n16155) );
  MUX2_X1 U19459 ( .A(n16558), .B(n16043), .S(n16065), .Z(n16044) );
  OAI21_X1 U19460 ( .B1(n19855), .B2(n16155), .A(n16044), .ZN(P2_U2869) );
  AND2_X1 U19461 ( .A1(n16028), .A2(n16045), .ZN(n16047) );
  OR2_X1 U19462 ( .A1(n16047), .A2(n16046), .ZN(n16165) );
  NAND2_X1 U19463 ( .A1(n16571), .A2(n19866), .ZN(n16049) );
  NAND2_X1 U19464 ( .A1(n16065), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n16048) );
  OAI211_X1 U19465 ( .C1(n16165), .C2(n19855), .A(n16049), .B(n16048), .ZN(
        P2_U2870) );
  XNOR2_X1 U19466 ( .A(n19848), .B(n19847), .ZN(n16052) );
  NOR2_X1 U19467 ( .A1(n16591), .A2(n16065), .ZN(n16050) );
  AOI21_X1 U19468 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(n16065), .A(n16050), .ZN(
        n16051) );
  OAI21_X1 U19469 ( .B1(n16052), .B2(n19855), .A(n16051), .ZN(P2_U2872) );
  NOR2_X1 U19470 ( .A1(n16054), .A2(n16053), .ZN(n19853) );
  NAND2_X1 U19471 ( .A1(n19853), .A2(n19854), .ZN(n19859) );
  INV_X1 U19472 ( .A(n16062), .ZN(n16055) );
  NOR2_X1 U19473 ( .A1(n19859), .A2(n16055), .ZN(n16059) );
  INV_X1 U19474 ( .A(n16056), .ZN(n16057) );
  OAI211_X1 U19475 ( .C1(n16059), .C2(n16058), .A(n19863), .B(n16057), .ZN(
        n16061) );
  NAND2_X1 U19476 ( .A1(n16065), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n16060) );
  OAI211_X1 U19477 ( .C1(n16625), .C2(n16065), .A(n16061), .B(n16060), .ZN(
        P2_U2875) );
  XOR2_X1 U19478 ( .A(n16062), .B(n19859), .Z(n16068) );
  NOR2_X1 U19479 ( .A1(n15888), .A2(n16063), .ZN(n16064) );
  OR2_X1 U19480 ( .A1(n15874), .A2(n16064), .ZN(n19760) );
  MUX2_X1 U19481 ( .A(n19760), .B(n16066), .S(n16065), .Z(n16067) );
  OAI21_X1 U19482 ( .B1(n16068), .B2(n19855), .A(n16067), .ZN(P2_U2876) );
  NAND2_X1 U19483 ( .A1(n16069), .A2(n19899), .ZN(n16071) );
  AOI22_X1 U19484 ( .A1(n19870), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19898), .ZN(n16070) );
  OAI211_X1 U19485 ( .C1(n17456), .C2(n16154), .A(n16071), .B(n16070), .ZN(
        P2_U2888) );
  NAND3_X1 U19486 ( .A1(n16073), .A2(n19903), .A3(n16072), .ZN(n16079) );
  INV_X1 U19487 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16076) );
  AOI22_X1 U19488 ( .A1(n19868), .A2(n16074), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n19898), .ZN(n16075) );
  OAI21_X1 U19489 ( .B1(n16154), .B2(n16076), .A(n16075), .ZN(n16077) );
  AOI21_X1 U19490 ( .B1(n19870), .B2(BUF2_REG_29__SCAN_IN), .A(n16077), .ZN(
        n16078) );
  OAI211_X1 U19491 ( .C1(n16080), .C2(n16168), .A(n16079), .B(n16078), .ZN(
        P2_U2890) );
  NAND2_X1 U19492 ( .A1(n19870), .A2(BUF2_REG_28__SCAN_IN), .ZN(n16084) );
  NAND2_X1 U19493 ( .A1(n19869), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16083) );
  AOI22_X1 U19494 ( .A1(n19868), .A2(n16081), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19898), .ZN(n16082) );
  NAND3_X1 U19495 ( .A1(n16084), .A2(n16083), .A3(n16082), .ZN(n16085) );
  AOI21_X1 U19496 ( .B1(n16461), .B2(n19899), .A(n16085), .ZN(n16086) );
  OAI21_X1 U19497 ( .B1(n16087), .B2(n16164), .A(n16086), .ZN(P2_U2891) );
  NAND2_X1 U19498 ( .A1(n9688), .A2(n19903), .ZN(n16093) );
  NAND2_X1 U19499 ( .A1(n19870), .A2(BUF2_REG_27__SCAN_IN), .ZN(n16091) );
  NAND2_X1 U19500 ( .A1(n19869), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16090) );
  AOI22_X1 U19501 ( .A1(n19868), .A2(n16088), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n19898), .ZN(n16089) );
  AND3_X1 U19502 ( .A1(n16091), .A2(n16090), .A3(n16089), .ZN(n16092) );
  OAI211_X1 U19503 ( .C1(n16094), .C2(n16168), .A(n16093), .B(n16092), .ZN(
        P2_U2892) );
  AOI22_X1 U19504 ( .A1(n19868), .A2(n16095), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19898), .ZN(n16096) );
  OAI21_X1 U19505 ( .B1(n16154), .B2(n16097), .A(n16096), .ZN(n16099) );
  NOR2_X1 U19506 ( .A1(n16473), .A2(n16168), .ZN(n16098) );
  AOI211_X1 U19507 ( .C1(n19870), .C2(BUF2_REG_26__SCAN_IN), .A(n16099), .B(
        n16098), .ZN(n16100) );
  OAI21_X1 U19508 ( .B1(n16101), .B2(n16164), .A(n16100), .ZN(P2_U2893) );
  NAND2_X1 U19509 ( .A1(n19869), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16104) );
  AOI22_X1 U19510 ( .A1(n19868), .A2(n16102), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n19898), .ZN(n16103) );
  NAND2_X1 U19511 ( .A1(n16104), .A2(n16103), .ZN(n16106) );
  NOR2_X1 U19512 ( .A1(n16486), .A2(n16168), .ZN(n16105) );
  AOI211_X1 U19513 ( .C1(n19870), .C2(BUF2_REG_25__SCAN_IN), .A(n16106), .B(
        n16105), .ZN(n16107) );
  OAI21_X1 U19514 ( .B1(n16164), .B2(n16108), .A(n16107), .ZN(P2_U2894) );
  NAND2_X1 U19515 ( .A1(n19869), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16111) );
  AOI22_X1 U19516 ( .A1(n19868), .A2(n16109), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19898), .ZN(n16110) );
  NAND2_X1 U19517 ( .A1(n16111), .A2(n16110), .ZN(n16113) );
  NOR2_X1 U19518 ( .A1(n16497), .A2(n16168), .ZN(n16112) );
  AOI211_X1 U19519 ( .C1(n19870), .C2(BUF2_REG_24__SCAN_IN), .A(n16113), .B(
        n16112), .ZN(n16114) );
  OAI21_X1 U19520 ( .B1(n16164), .B2(n16115), .A(n16114), .ZN(P2_U2895) );
  INV_X1 U19521 ( .A(n19870), .ZN(n16134) );
  INV_X1 U19522 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16118) );
  AOI22_X1 U19523 ( .A1(n19868), .A2(n20026), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n19898), .ZN(n16117) );
  NAND2_X1 U19524 ( .A1(n19869), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16116) );
  OAI211_X1 U19525 ( .C1(n16134), .C2(n16118), .A(n16117), .B(n16116), .ZN(
        n16119) );
  AOI21_X1 U19526 ( .B1(n16120), .B2(n19903), .A(n16119), .ZN(n16121) );
  OAI21_X1 U19527 ( .B1(n16122), .B2(n16168), .A(n16121), .ZN(P2_U2896) );
  OR2_X1 U19528 ( .A1(n15745), .A2(n16123), .ZN(n16124) );
  NAND2_X1 U19529 ( .A1(n16125), .A2(n16124), .ZN(n17303) );
  AOI22_X1 U19530 ( .A1(n19868), .A2(n20016), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19898), .ZN(n16127) );
  NAND2_X1 U19531 ( .A1(n19869), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16126) );
  OAI211_X1 U19532 ( .C1(n16134), .C2(n19134), .A(n16127), .B(n16126), .ZN(
        n16128) );
  AOI21_X1 U19533 ( .B1(n16129), .B2(n19903), .A(n16128), .ZN(n16130) );
  OAI21_X1 U19534 ( .B1(n17303), .B2(n16168), .A(n16130), .ZN(P2_U2897) );
  INV_X1 U19535 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16133) );
  AOI22_X1 U19536 ( .A1(n19868), .A2(n20007), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n19898), .ZN(n16132) );
  NAND2_X1 U19537 ( .A1(n19869), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16131) );
  OAI211_X1 U19538 ( .C1(n16134), .C2(n16133), .A(n16132), .B(n16131), .ZN(
        n16135) );
  AOI21_X1 U19539 ( .B1(n16136), .B2(n19903), .A(n16135), .ZN(n16137) );
  OAI21_X1 U19540 ( .B1(n16138), .B2(n16168), .A(n16137), .ZN(P2_U2898) );
  NAND2_X1 U19541 ( .A1(n16139), .A2(n19899), .ZN(n16143) );
  AOI22_X1 U19542 ( .A1(n19868), .A2(n20003), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19898), .ZN(n16140) );
  OAI21_X1 U19543 ( .B1(n16154), .B2(n17473), .A(n16140), .ZN(n16141) );
  AOI21_X1 U19544 ( .B1(n19870), .B2(BUF2_REG_20__SCAN_IN), .A(n16141), .ZN(
        n16142) );
  OAI211_X1 U19545 ( .C1(n16164), .C2(n16144), .A(n16143), .B(n16142), .ZN(
        P2_U2899) );
  AOI22_X1 U19546 ( .A1(n19868), .A2(n19998), .B1(P2_EAX_REG_19__SCAN_IN), 
        .B2(n19898), .ZN(n16146) );
  NAND2_X1 U19547 ( .A1(n19870), .A2(BUF2_REG_19__SCAN_IN), .ZN(n16145) );
  OAI211_X1 U19548 ( .C1(n16154), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        n16148) );
  AOI21_X1 U19549 ( .B1(n16149), .B2(n19903), .A(n16148), .ZN(n16150) );
  OAI21_X1 U19550 ( .B1(n16151), .B2(n16168), .A(n16150), .ZN(P2_U2900) );
  INV_X1 U19551 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16153) );
  AOI22_X1 U19552 ( .A1(n19868), .A2(n19993), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19898), .ZN(n16152) );
  OAI21_X1 U19553 ( .B1(n16154), .B2(n16153), .A(n16152), .ZN(n16157) );
  NOR2_X1 U19554 ( .A1(n16155), .A2(n16164), .ZN(n16156) );
  AOI211_X1 U19555 ( .C1(n19870), .C2(BUF2_REG_18__SCAN_IN), .A(n16157), .B(
        n16156), .ZN(n16158) );
  OAI21_X1 U19556 ( .B1(n16552), .B2(n16168), .A(n16158), .ZN(P2_U2901) );
  NAND2_X1 U19557 ( .A1(n19898), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n16159) );
  OAI21_X1 U19558 ( .B1(n16160), .B2(n19908), .A(n16159), .ZN(n16161) );
  AOI21_X1 U19559 ( .B1(n19869), .B2(BUF1_REG_17__SCAN_IN), .A(n16161), .ZN(
        n16163) );
  NAND2_X1 U19560 ( .A1(n19870), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16162) );
  OAI211_X1 U19561 ( .C1(n16165), .C2(n16164), .A(n16163), .B(n16162), .ZN(
        n16166) );
  INV_X1 U19562 ( .A(n16166), .ZN(n16167) );
  OAI21_X1 U19563 ( .B1(n16573), .B2(n16168), .A(n16167), .ZN(P2_U2902) );
  XNOR2_X1 U19564 ( .A(n16170), .B(n16171), .ZN(n19793) );
  XNOR2_X1 U19565 ( .A(n16775), .B(n20607), .ZN(n19885) );
  XNOR2_X1 U19566 ( .A(n16798), .B(n19959), .ZN(n19902) );
  NAND2_X1 U19567 ( .A1(n16813), .A2(n19826), .ZN(n19901) );
  NAND2_X1 U19568 ( .A1(n19902), .A2(n19901), .ZN(n19900) );
  OAI21_X1 U19569 ( .B1(n16797), .B2(n19959), .A(n19900), .ZN(n19892) );
  XNOR2_X1 U19570 ( .A(n16799), .B(n19890), .ZN(n19893) );
  NAND2_X1 U19571 ( .A1(n19892), .A2(n19893), .ZN(n19891) );
  OAI21_X1 U19572 ( .B1(n16769), .B2(n19890), .A(n19891), .ZN(n19884) );
  NAND2_X1 U19573 ( .A1(n19885), .A2(n19884), .ZN(n19883) );
  OAI21_X1 U19574 ( .B1(n20610), .B2(n20607), .A(n19883), .ZN(n16174) );
  NAND2_X1 U19575 ( .A1(n15937), .A2(n16172), .ZN(n16173) );
  NAND2_X1 U19576 ( .A1(n16170), .A2(n16173), .ZN(n19811) );
  NAND2_X1 U19577 ( .A1(n16174), .A2(n19811), .ZN(n19878) );
  INV_X1 U19578 ( .A(n16175), .ZN(n16176) );
  NAND2_X1 U19579 ( .A1(n16179), .A2(n16178), .ZN(n19877) );
  INV_X1 U19580 ( .A(n19877), .ZN(n19864) );
  NAND3_X1 U19581 ( .A1(n19878), .A2(n19903), .A3(n19864), .ZN(n16182) );
  AOI22_X1 U19582 ( .A1(n16180), .A2(n20007), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19898), .ZN(n16181) );
  OAI211_X1 U19583 ( .C1(n19793), .C2(n16183), .A(n16182), .B(n16181), .ZN(
        P2_U2914) );
  NOR2_X1 U19584 ( .A1(n16184), .A2(n16455), .ZN(n16189) );
  NAND2_X1 U19585 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16185) );
  OAI211_X1 U19586 ( .C1(n16187), .C2(n16441), .A(n16186), .B(n16185), .ZN(
        n16188) );
  AOI211_X1 U19587 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n11076), .A(
        n16212), .B(n16193), .ZN(n16195) );
  NAND2_X1 U19588 ( .A1(n16196), .A2(n11076), .ZN(n16197) );
  XNOR2_X1 U19589 ( .A(n16197), .B(n16462), .ZN(n16198) );
  NAND2_X1 U19590 ( .A1(n16460), .A2(n16435), .ZN(n16204) );
  NAND2_X1 U19591 ( .A1(n16423), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n16464) );
  OAI21_X1 U19592 ( .B1(n16424), .B2(n16200), .A(n16464), .ZN(n16202) );
  NOR2_X1 U19593 ( .A1(n16466), .A2(n16455), .ZN(n16201) );
  AOI211_X1 U19594 ( .C1(n16452), .C2(n10605), .A(n16202), .B(n16201), .ZN(
        n16203) );
  OAI211_X1 U19595 ( .C1(n16446), .C2(n16469), .A(n16204), .B(n16203), .ZN(
        P2_U2986) );
  NAND2_X1 U19596 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16205) );
  OAI211_X1 U19597 ( .C1(n16207), .C2(n16441), .A(n16206), .B(n16205), .ZN(
        n16209) );
  INV_X1 U19598 ( .A(n16212), .ZN(n16224) );
  NAND2_X1 U19599 ( .A1(n16213), .A2(n16224), .ZN(n16214) );
  XOR2_X1 U19600 ( .A(n16215), .B(n16214), .Z(n16485) );
  NOR2_X1 U19601 ( .A1(n10176), .A2(n20588), .ZN(n16479) );
  AOI21_X1 U19602 ( .B1(n16450), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16479), .ZN(n16220) );
  NAND2_X1 U19603 ( .A1(n16218), .A2(n16452), .ZN(n16219) );
  OAI211_X1 U19604 ( .C1(n16481), .C2(n16455), .A(n16220), .B(n16219), .ZN(
        n16221) );
  AOI21_X1 U19605 ( .B1(n16484), .B2(n16457), .A(n16221), .ZN(n16222) );
  OAI21_X1 U19606 ( .B1(n16485), .B2(n16459), .A(n16222), .ZN(P2_U2988) );
  NAND2_X1 U19607 ( .A1(n16224), .A2(n16223), .ZN(n16226) );
  XOR2_X1 U19608 ( .A(n16226), .B(n16225), .Z(n16496) );
  NAND2_X1 U19609 ( .A1(n16235), .A2(n16227), .ZN(n16228) );
  NOR2_X1 U19610 ( .A1(n10176), .A2(n20586), .ZN(n16489) );
  NOR2_X1 U19611 ( .A1(n16229), .A2(n16441), .ZN(n16230) );
  AOI211_X1 U19612 ( .C1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n16450), .A(
        n16489), .B(n16230), .ZN(n16231) );
  OAI21_X1 U19613 ( .B1(n16492), .B2(n16455), .A(n16231), .ZN(n16232) );
  OAI21_X1 U19614 ( .B1(n16496), .B2(n16459), .A(n16233), .ZN(P2_U2989) );
  NAND2_X1 U19615 ( .A1(n16236), .A2(n16452), .ZN(n16237) );
  NAND2_X1 U19616 ( .A1(n16423), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16500) );
  OAI211_X1 U19617 ( .C1(n16238), .C2(n16424), .A(n16237), .B(n16500), .ZN(
        n16242) );
  XNOR2_X1 U19618 ( .A(n16239), .B(n16501), .ZN(n16240) );
  XNOR2_X1 U19619 ( .A(n16243), .B(n16244), .ZN(n16521) );
  NAND2_X1 U19620 ( .A1(n16423), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16511) );
  NAND2_X1 U19621 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16245) );
  OAI211_X1 U19622 ( .C1(n16246), .C2(n16441), .A(n16511), .B(n16245), .ZN(
        n16247) );
  AOI21_X1 U19623 ( .B1(n16517), .B2(n16443), .A(n16247), .ZN(n16248) );
  OAI211_X1 U19624 ( .C1(n16521), .C2(n16459), .A(n16249), .B(n16248), .ZN(
        P2_U2991) );
  OAI21_X1 U19625 ( .B1(n9946), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16250), .ZN(n16535) );
  NAND2_X1 U19626 ( .A1(n16253), .A2(n16252), .ZN(n16254) );
  XNOR2_X1 U19627 ( .A(n16251), .B(n16254), .ZN(n16533) );
  AND2_X1 U19628 ( .A1(n16423), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16525) );
  AOI21_X1 U19629 ( .B1(n16450), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16525), .ZN(n16256) );
  NAND2_X1 U19630 ( .A1(n17310), .A2(n16452), .ZN(n16255) );
  OAI211_X1 U19631 ( .C1(n17304), .C2(n16455), .A(n16256), .B(n16255), .ZN(
        n16257) );
  AOI21_X1 U19632 ( .B1(n16435), .B2(n16533), .A(n16257), .ZN(n16258) );
  OAI21_X1 U19633 ( .B1(n16535), .B2(n16446), .A(n16258), .ZN(P2_U2992) );
  NAND2_X1 U19634 ( .A1(n16260), .A2(n16259), .ZN(n16264) );
  NAND2_X1 U19635 ( .A1(n16262), .A2(n16261), .ZN(n16263) );
  XNOR2_X1 U19636 ( .A(n16264), .B(n16263), .ZN(n16549) );
  NAND2_X1 U19637 ( .A1(n16423), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16540) );
  NAND2_X1 U19638 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16265) );
  OAI211_X1 U19639 ( .C1(n16266), .C2(n16441), .A(n16540), .B(n16265), .ZN(
        n16269) );
  OAI21_X1 U19640 ( .B1(n16549), .B2(n16459), .A(n16271), .ZN(P2_U2993) );
  AOI21_X1 U19641 ( .B1(n16450), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16272), .ZN(n16275) );
  NAND2_X1 U19642 ( .A1(n16273), .A2(n16452), .ZN(n16274) );
  OAI211_X1 U19643 ( .C1(n16276), .C2(n16455), .A(n16275), .B(n16274), .ZN(
        n16277) );
  OAI21_X1 U19644 ( .B1(n16279), .B2(n16459), .A(n16278), .ZN(P2_U2995) );
  NAND2_X1 U19645 ( .A1(n16282), .A2(n16281), .ZN(n16283) );
  XNOR2_X1 U19646 ( .A(n16284), .B(n16283), .ZN(n16550) );
  NAND2_X1 U19647 ( .A1(n16550), .A2(n16435), .ZN(n16290) );
  NAND2_X1 U19648 ( .A1(n16423), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16557) );
  OAI21_X1 U19649 ( .B1(n16424), .B2(n16285), .A(n16557), .ZN(n16287) );
  NOR2_X1 U19650 ( .A1(n16558), .A2(n16455), .ZN(n16286) );
  AOI211_X1 U19651 ( .C1(n16452), .C2(n16288), .A(n16287), .B(n16286), .ZN(
        n16289) );
  XOR2_X1 U19652 ( .A(n16292), .B(n16291), .Z(n16575) );
  INV_X1 U19653 ( .A(n16575), .ZN(n16300) );
  AND2_X1 U19654 ( .A1(n16423), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16570) );
  AOI21_X1 U19655 ( .B1(n16450), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16570), .ZN(n16293) );
  OAI21_X1 U19656 ( .B1(n16441), .B2(n16294), .A(n16293), .ZN(n16298) );
  AND2_X1 U19657 ( .A1(n16295), .A2(n16566), .ZN(n16296) );
  OAI21_X1 U19658 ( .B1(n16300), .B2(n16459), .A(n16299), .ZN(P2_U2997) );
  INV_X1 U19659 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20570) );
  NOR2_X1 U19660 ( .A1(n10176), .A2(n20570), .ZN(n16580) );
  AOI21_X1 U19661 ( .B1(n16450), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16580), .ZN(n16301) );
  OAI21_X1 U19662 ( .B1(n16441), .B2(n16302), .A(n16301), .ZN(n16305) );
  NAND2_X1 U19663 ( .A1(n16307), .A2(n16306), .ZN(n16309) );
  XOR2_X1 U19664 ( .A(n16309), .B(n16308), .Z(n16597) );
  AOI21_X1 U19665 ( .B1(n16568), .B2(n16317), .A(n16310), .ZN(n16587) );
  NAND2_X1 U19666 ( .A1(n16587), .A2(n16457), .ZN(n16316) );
  INV_X1 U19667 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16311) );
  NAND2_X1 U19668 ( .A1(n16423), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16590) );
  OAI21_X1 U19669 ( .B1(n16424), .B2(n16311), .A(n16590), .ZN(n16313) );
  NOR2_X1 U19670 ( .A1(n16591), .A2(n16455), .ZN(n16312) );
  AOI211_X1 U19671 ( .C1(n16314), .C2(n16452), .A(n16313), .B(n16312), .ZN(
        n16315) );
  OAI211_X1 U19672 ( .C1(n16597), .C2(n16459), .A(n16316), .B(n16315), .ZN(
        P2_U2999) );
  NOR2_X1 U19673 ( .A1(n16354), .A2(n16615), .ZN(n16335) );
  OAI21_X1 U19674 ( .B1(n16335), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16317), .ZN(n16609) );
  NOR2_X1 U19675 ( .A1(n16441), .A2(n16318), .ZN(n16320) );
  NAND2_X1 U19676 ( .A1(n16423), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n16600) );
  OAI21_X1 U19677 ( .B1(n16424), .B2(n10413), .A(n16600), .ZN(n16319) );
  AOI211_X1 U19678 ( .C1(n16321), .C2(n16443), .A(n16320), .B(n16319), .ZN(
        n16327) );
  NAND2_X1 U19679 ( .A1(n16323), .A2(n16322), .ZN(n16325) );
  XOR2_X1 U19680 ( .A(n16325), .B(n16324), .Z(n16606) );
  NAND2_X1 U19681 ( .A1(n16606), .A2(n16435), .ZN(n16326) );
  OAI211_X1 U19682 ( .C1(n16609), .C2(n16446), .A(n16327), .B(n16326), .ZN(
        P2_U3000) );
  INV_X1 U19683 ( .A(n16369), .ZN(n16328) );
  NOR2_X1 U19684 ( .A1(n9636), .A2(n16328), .ZN(n16356) );
  NAND2_X1 U19685 ( .A1(n16356), .A2(n16360), .ZN(n16343) );
  NAND3_X1 U19686 ( .A1(n16343), .A2(n16342), .A3(n16345), .ZN(n16329) );
  NAND2_X1 U19687 ( .A1(n16329), .A2(n16344), .ZN(n16333) );
  NAND2_X1 U19688 ( .A1(n16331), .A2(n16330), .ZN(n16332) );
  XNOR2_X1 U19689 ( .A(n16333), .B(n16332), .ZN(n16624) );
  INV_X1 U19690 ( .A(n16354), .ZN(n16334) );
  AOI21_X1 U19691 ( .B1(n16334), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16336) );
  NOR2_X1 U19692 ( .A1(n16336), .A2(n16335), .ZN(n16610) );
  NAND2_X1 U19693 ( .A1(n16610), .A2(n16457), .ZN(n16341) );
  NAND2_X1 U19694 ( .A1(n16423), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16612) );
  NAND2_X1 U19695 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16337) );
  OAI211_X1 U19696 ( .C1(n16441), .C2(n16338), .A(n16612), .B(n16337), .ZN(
        n16339) );
  AOI21_X1 U19697 ( .B1(n16611), .B2(n16443), .A(n16339), .ZN(n16340) );
  OAI211_X1 U19698 ( .C1(n16459), .C2(n16624), .A(n16341), .B(n16340), .ZN(
        P2_U3001) );
  XNOR2_X1 U19699 ( .A(n16354), .B(n16632), .ZN(n16637) );
  NAND2_X1 U19700 ( .A1(n16343), .A2(n16342), .ZN(n16347) );
  NAND2_X1 U19701 ( .A1(n16345), .A2(n16344), .ZN(n16346) );
  XNOR2_X1 U19702 ( .A(n16347), .B(n16346), .ZN(n16635) );
  NOR2_X1 U19703 ( .A1(n10176), .A2(n20562), .ZN(n16627) );
  NOR2_X1 U19704 ( .A1(n16441), .A2(n16348), .ZN(n16349) );
  AOI211_X1 U19705 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n16450), .A(
        n16627), .B(n16349), .ZN(n16350) );
  OAI21_X1 U19706 ( .B1(n16625), .B2(n16455), .A(n16350), .ZN(n16351) );
  AOI21_X1 U19707 ( .B1(n16635), .B2(n16435), .A(n16351), .ZN(n16352) );
  OAI21_X1 U19708 ( .B1(n16637), .B2(n16446), .A(n16352), .ZN(P2_U3002) );
  OAI21_X1 U19709 ( .B1(n16353), .B2(n16658), .A(n16640), .ZN(n16355) );
  NAND2_X1 U19710 ( .A1(n16355), .A2(n16354), .ZN(n16650) );
  INV_X1 U19711 ( .A(n16356), .ZN(n16358) );
  NAND2_X1 U19712 ( .A1(n16358), .A2(n16357), .ZN(n16362) );
  NAND2_X1 U19713 ( .A1(n16360), .A2(n16359), .ZN(n16361) );
  XNOR2_X1 U19714 ( .A(n16362), .B(n16361), .ZN(n16648) );
  NOR2_X1 U19715 ( .A1(n19760), .A2(n16455), .ZN(n16365) );
  NAND2_X1 U19716 ( .A1(n16423), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n16642) );
  NAND2_X1 U19717 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16363) );
  OAI211_X1 U19718 ( .C1(n16441), .C2(n19765), .A(n16642), .B(n16363), .ZN(
        n16364) );
  AOI211_X1 U19719 ( .C1(n16648), .C2(n16435), .A(n16365), .B(n16364), .ZN(
        n16366) );
  OAI21_X1 U19720 ( .B1(n16650), .B2(n16446), .A(n16366), .ZN(P2_U3003) );
  XNOR2_X1 U19721 ( .A(n16353), .B(n16658), .ZN(n16663) );
  NAND2_X1 U19722 ( .A1(n16452), .A2(n16367), .ZN(n16368) );
  NAND2_X1 U19723 ( .A1(n16423), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n16652) );
  OAI211_X1 U19724 ( .C1(n10418), .C2(n16424), .A(n16368), .B(n16652), .ZN(
        n16374) );
  NAND2_X1 U19725 ( .A1(n16370), .A2(n16369), .ZN(n16372) );
  NAND2_X1 U19726 ( .A1(n9636), .A2(n16376), .ZN(n16371) );
  XOR2_X1 U19727 ( .A(n16372), .B(n16371), .Z(n16651) );
  NOR2_X1 U19728 ( .A1(n16651), .A2(n16459), .ZN(n16373) );
  AOI211_X1 U19729 ( .C1(n16443), .C2(n19858), .A(n16374), .B(n16373), .ZN(
        n16375) );
  OAI21_X1 U19730 ( .B1(n16446), .B2(n16663), .A(n16375), .ZN(P2_U3004) );
  NAND2_X1 U19731 ( .A1(n16377), .A2(n16376), .ZN(n16378) );
  XOR2_X1 U19732 ( .A(n16378), .B(n9711), .Z(n16675) );
  NAND2_X1 U19733 ( .A1(n16379), .A2(n16638), .ZN(n16664) );
  NAND3_X1 U19734 ( .A1(n16664), .A2(n16457), .A3(n16353), .ZN(n16383) );
  NOR2_X1 U19735 ( .A1(n10176), .A2(n20556), .ZN(n16666) );
  AOI21_X1 U19736 ( .B1(n16450), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16666), .ZN(n16380) );
  OAI21_X1 U19737 ( .B1(n16441), .B2(n19779), .A(n16380), .ZN(n16381) );
  AOI21_X1 U19738 ( .B1(n16667), .B2(n16443), .A(n16381), .ZN(n16382) );
  OAI211_X1 U19739 ( .C1(n16459), .C2(n16675), .A(n16383), .B(n16382), .ZN(
        P2_U3005) );
  XNOR2_X1 U19740 ( .A(n16384), .B(n16704), .ZN(n16410) );
  OAI21_X1 U19741 ( .B1(n16410), .B2(n16411), .A(n16386), .ZN(n16402) );
  AOI21_X1 U19742 ( .B1(n16402), .B2(n16399), .A(n11016), .ZN(n16390) );
  NAND2_X1 U19743 ( .A1(n16388), .A2(n16387), .ZN(n16389) );
  XNOR2_X1 U19744 ( .A(n16390), .B(n16389), .ZN(n16688) );
  OR2_X1 U19745 ( .A1(n16391), .A2(n9652), .ZN(n16676) );
  NAND3_X1 U19746 ( .A1(n16676), .A2(n16457), .A3(n16392), .ZN(n16397) );
  NAND2_X1 U19747 ( .A1(n16423), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16679) );
  NAND2_X1 U19748 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16393) );
  OAI211_X1 U19749 ( .C1(n16441), .C2(n16394), .A(n16679), .B(n16393), .ZN(
        n16395) );
  AOI21_X1 U19750 ( .B1(n16678), .B2(n16443), .A(n16395), .ZN(n16396) );
  OAI211_X1 U19751 ( .C1(n16688), .C2(n16459), .A(n16397), .B(n16396), .ZN(
        P2_U3006) );
  NAND2_X1 U19752 ( .A1(n16400), .A2(n16399), .ZN(n16401) );
  XNOR2_X1 U19753 ( .A(n16402), .B(n16401), .ZN(n16697) );
  NOR2_X1 U19754 ( .A1(n10176), .A2(n20552), .ZN(n16691) );
  NOR2_X1 U19755 ( .A1(n16424), .A2(n16403), .ZN(n16404) );
  AOI211_X1 U19756 ( .C1(n16405), .C2(n16452), .A(n16691), .B(n16404), .ZN(
        n16406) );
  OAI21_X1 U19757 ( .B1(n16407), .B2(n16455), .A(n16406), .ZN(n16408) );
  AOI21_X1 U19758 ( .B1(n16697), .B2(n16435), .A(n16408), .ZN(n16409) );
  OAI21_X1 U19759 ( .B1(n16699), .B2(n16446), .A(n16409), .ZN(P2_U3007) );
  XOR2_X1 U19760 ( .A(n16411), .B(n16410), .Z(n16700) );
  NAND2_X1 U19761 ( .A1(n16700), .A2(n16435), .ZN(n16416) );
  NAND2_X1 U19762 ( .A1(n16423), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n16702) );
  OAI21_X1 U19763 ( .B1(n16424), .B2(n21556), .A(n16702), .ZN(n16413) );
  NOR2_X1 U19764 ( .A1(n16703), .A2(n16455), .ZN(n16412) );
  AOI211_X1 U19765 ( .C1(n16414), .C2(n16452), .A(n16413), .B(n16412), .ZN(
        n16415) );
  OAI211_X1 U19766 ( .C1(n16446), .C2(n16711), .A(n16416), .B(n16415), .ZN(
        P2_U3008) );
  XNOR2_X1 U19767 ( .A(n16417), .B(n16418), .ZN(n16722) );
  AOI21_X1 U19768 ( .B1(n10243), .B2(n16420), .A(n16419), .ZN(n16421) );
  AOI21_X1 U19769 ( .B1(n16422), .B2(n10243), .A(n16421), .ZN(n16712) );
  NAND2_X1 U19770 ( .A1(n16712), .A2(n16457), .ZN(n16428) );
  NOR2_X1 U19771 ( .A1(n16441), .A2(n19794), .ZN(n16426) );
  NAND2_X1 U19772 ( .A1(n16423), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n16715) );
  OAI21_X1 U19773 ( .B1(n16424), .B2(n12468), .A(n16715), .ZN(n16425) );
  AOI211_X1 U19774 ( .C1(n19800), .C2(n16443), .A(n16426), .B(n16425), .ZN(
        n16427) );
  OAI211_X1 U19775 ( .C1(n16722), .C2(n16459), .A(n16428), .B(n16427), .ZN(
        P2_U3009) );
  XNOR2_X1 U19776 ( .A(n16429), .B(n16725), .ZN(n16430) );
  XNOR2_X1 U19777 ( .A(n16431), .B(n16430), .ZN(n16732) );
  XNOR2_X1 U19778 ( .A(n16432), .B(n16736), .ZN(n16448) );
  AOI22_X1 U19779 ( .A1(n16448), .A2(n16447), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16432), .ZN(n16434) );
  XNOR2_X1 U19780 ( .A(n19808), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16433) );
  XNOR2_X1 U19781 ( .A(n16434), .B(n16433), .ZN(n16723) );
  NAND2_X1 U19782 ( .A1(n16723), .A2(n16435), .ZN(n16445) );
  OR2_X1 U19783 ( .A1(n16437), .A2(n16436), .ZN(n16438) );
  AND2_X1 U19784 ( .A1(n14373), .A2(n16438), .ZN(n19862) );
  INV_X1 U19785 ( .A(n19816), .ZN(n16440) );
  AOI22_X1 U19786 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n16423), .ZN(n16439) );
  OAI21_X1 U19787 ( .B1(n16441), .B2(n16440), .A(n16439), .ZN(n16442) );
  AOI21_X1 U19788 ( .B1(n19862), .B2(n16443), .A(n16442), .ZN(n16444) );
  OAI211_X1 U19789 ( .C1(n16446), .C2(n16732), .A(n16445), .B(n16444), .ZN(
        P2_U3010) );
  XNOR2_X1 U19790 ( .A(n16448), .B(n16447), .ZN(n16743) );
  AOI22_X1 U19791 ( .A1(n16450), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n16423), .ZN(n16454) );
  NAND2_X1 U19792 ( .A1(n16452), .A2(n16451), .ZN(n16453) );
  OAI211_X1 U19793 ( .C1(n16733), .C2(n16455), .A(n16454), .B(n16453), .ZN(
        n16456) );
  AOI21_X1 U19794 ( .B1(n16740), .B2(n16457), .A(n16456), .ZN(n16458) );
  OAI21_X1 U19795 ( .B1(n16743), .B2(n16459), .A(n16458), .ZN(P2_U3011) );
  INV_X1 U19796 ( .A(n16460), .ZN(n16472) );
  INV_X1 U19797 ( .A(n16470), .ZN(n16471) );
  OAI21_X1 U19798 ( .B1(n16472), .B2(n19974), .A(n16471), .ZN(P2_U3018) );
  NOR2_X1 U19799 ( .A1(n16473), .A2(n19949), .ZN(n16483) );
  INV_X1 U19800 ( .A(n16474), .ZN(n16502) );
  INV_X1 U19801 ( .A(n16475), .ZN(n16476) );
  AOI21_X1 U19802 ( .B1(n16502), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16476), .ZN(n16490) );
  XNOR2_X1 U19803 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16477) );
  NOR2_X1 U19804 ( .A1(n16487), .A2(n16477), .ZN(n16478) );
  AOI211_X1 U19805 ( .C1(n16490), .C2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16479), .B(n16478), .ZN(n16480) );
  OAI21_X1 U19806 ( .B1(n16481), .B2(n19964), .A(n16480), .ZN(n16482) );
  NOR2_X1 U19807 ( .A1(n16486), .A2(n19949), .ZN(n16494) );
  NOR2_X1 U19808 ( .A1(n16487), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16488) );
  AOI211_X1 U19809 ( .C1(n16490), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16489), .B(n16488), .ZN(n16491) );
  OAI21_X1 U19810 ( .B1(n16492), .B2(n19964), .A(n16491), .ZN(n16493) );
  OAI21_X1 U19811 ( .B1(n16496), .B2(n19974), .A(n16495), .ZN(P2_U3021) );
  NOR2_X1 U19812 ( .A1(n16497), .A2(n19949), .ZN(n16504) );
  INV_X1 U19813 ( .A(n16498), .ZN(n16526) );
  NAND3_X1 U19814 ( .A1(n16526), .A2(n16510), .A3(n16501), .ZN(n16499) );
  OAI211_X1 U19815 ( .C1(n16502), .C2(n16501), .A(n16500), .B(n16499), .ZN(
        n16503) );
  AOI211_X1 U19816 ( .C1(n16505), .C2(n19944), .A(n16504), .B(n16503), .ZN(
        n16508) );
  OR2_X1 U19817 ( .A1(n16506), .A2(n19974), .ZN(n16507) );
  OAI211_X1 U19818 ( .C1(n16509), .C2(n19963), .A(n16508), .B(n16507), .ZN(
        P2_U3022) );
  AOI21_X1 U19819 ( .B1(n10013), .B2(n16515), .A(n16510), .ZN(n16513) );
  INV_X1 U19820 ( .A(n16511), .ZN(n16512) );
  AOI21_X1 U19821 ( .B1(n16526), .B2(n16513), .A(n16512), .ZN(n16514) );
  OAI21_X1 U19822 ( .B1(n16528), .B2(n16515), .A(n16514), .ZN(n16516) );
  AOI21_X1 U19823 ( .B1(n16517), .B2(n19944), .A(n16516), .ZN(n16520) );
  NAND2_X1 U19824 ( .A1(n16518), .A2(n19960), .ZN(n16519) );
  OAI211_X1 U19825 ( .C1(n16521), .C2(n19974), .A(n16520), .B(n16519), .ZN(
        n16522) );
  INV_X1 U19826 ( .A(n16524), .ZN(P2_U3023) );
  NOR2_X1 U19827 ( .A1(n17303), .A2(n19949), .ZN(n16532) );
  AOI21_X1 U19828 ( .B1(n16526), .B2(n10013), .A(n16525), .ZN(n16527) );
  OAI21_X1 U19829 ( .B1(n16528), .B2(n10013), .A(n16527), .ZN(n16529) );
  INV_X1 U19830 ( .A(n16529), .ZN(n16530) );
  OAI21_X1 U19831 ( .B1(n17304), .B2(n19964), .A(n16530), .ZN(n16531) );
  AOI211_X1 U19832 ( .C1(n17444), .C2(n16533), .A(n16532), .B(n16531), .ZN(
        n16534) );
  OAI21_X1 U19833 ( .B1(n16535), .B2(n19963), .A(n16534), .ZN(P2_U3024) );
  INV_X1 U19834 ( .A(n16536), .ZN(n16672) );
  AOI21_X1 U19835 ( .B1(n16537), .B2(n9852), .A(n16672), .ZN(n16542) );
  INV_X1 U19836 ( .A(n16537), .ZN(n16538) );
  NAND3_X1 U19837 ( .A1(n16665), .A2(n16538), .A3(n16541), .ZN(n16539) );
  OAI211_X1 U19838 ( .C1(n16542), .C2(n16541), .A(n16540), .B(n16539), .ZN(
        n16545) );
  NOR2_X1 U19839 ( .A1(n16543), .A2(n19964), .ZN(n16544) );
  AOI211_X1 U19840 ( .C1(n16546), .C2(n19960), .A(n16545), .B(n16544), .ZN(
        n16548) );
  INV_X1 U19841 ( .A(n16550), .ZN(n16563) );
  NOR2_X1 U19842 ( .A1(n16552), .A2(n19949), .ZN(n16561) );
  NOR2_X1 U19843 ( .A1(n16554), .A2(n16553), .ZN(n16560) );
  OR3_X1 U19844 ( .A1(n16616), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16555), .ZN(n16556) );
  OAI211_X1 U19845 ( .C1(n16558), .C2(n19964), .A(n16557), .B(n16556), .ZN(
        n16559) );
  OAI21_X1 U19846 ( .B1(n16563), .B2(n19974), .A(n16562), .ZN(P2_U3028) );
  AOI21_X1 U19847 ( .B1(n16585), .B2(n9852), .A(n16579), .ZN(n16578) );
  INV_X1 U19848 ( .A(n16566), .ZN(n16567) );
  OR2_X1 U19849 ( .A1(n16616), .A2(n16567), .ZN(n16592) );
  AOI21_X1 U19850 ( .B1(n16571), .B2(n19944), .A(n16570), .ZN(n16572) );
  AOI21_X1 U19851 ( .B1(n16575), .B2(n17444), .A(n16574), .ZN(n16576) );
  OAI21_X1 U19852 ( .B1(n16578), .B2(n16577), .A(n16576), .ZN(P2_U3029) );
  INV_X1 U19853 ( .A(n16579), .ZN(n16586) );
  AOI21_X1 U19854 ( .B1(n19851), .B2(n19944), .A(n16580), .ZN(n16582) );
  NAND2_X1 U19855 ( .A1(n19871), .A2(n19960), .ZN(n16581) );
  NAND2_X1 U19856 ( .A1(n16587), .A2(n19946), .ZN(n16596) );
  NAND2_X1 U19857 ( .A1(n16588), .A2(n19960), .ZN(n16589) );
  OAI211_X1 U19858 ( .C1(n16591), .C2(n19964), .A(n16590), .B(n16589), .ZN(
        n16594) );
  NOR2_X1 U19859 ( .A1(n16592), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16593) );
  AOI211_X1 U19860 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16605), .A(
        n16594), .B(n16593), .ZN(n16595) );
  OAI211_X1 U19861 ( .C1(n16597), .C2(n19974), .A(n16596), .B(n16595), .ZN(
        P2_U3031) );
  OAI21_X1 U19862 ( .B1(n16616), .B2(n16615), .A(n16598), .ZN(n16604) );
  NOR2_X1 U19863 ( .A1(n16599), .A2(n19949), .ZN(n16603) );
  OAI21_X1 U19864 ( .B1(n16601), .B2(n19964), .A(n16600), .ZN(n16602) );
  AOI211_X1 U19865 ( .C1(n16605), .C2(n16604), .A(n16603), .B(n16602), .ZN(
        n16608) );
  NAND2_X1 U19866 ( .A1(n16606), .A2(n17444), .ZN(n16607) );
  OAI211_X1 U19867 ( .C1(n16609), .C2(n19963), .A(n16608), .B(n16607), .ZN(
        P2_U3032) );
  NAND2_X1 U19868 ( .A1(n16610), .A2(n19946), .ZN(n16623) );
  INV_X1 U19869 ( .A(n16633), .ZN(n16621) );
  NAND2_X1 U19870 ( .A1(n16611), .A2(n19944), .ZN(n16613) );
  OAI211_X1 U19871 ( .C1(n19949), .C2(n16614), .A(n16613), .B(n16612), .ZN(
        n16620) );
  INV_X1 U19872 ( .A(n16615), .ZN(n16617) );
  AOI211_X1 U19873 ( .C1(n16632), .C2(n16618), .A(n16617), .B(n16616), .ZN(
        n16619) );
  AOI211_X1 U19874 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16621), .A(
        n16620), .B(n16619), .ZN(n16622) );
  OAI211_X1 U19875 ( .C1(n16624), .C2(n19974), .A(n16623), .B(n16622), .ZN(
        P2_U3033) );
  NOR2_X1 U19876 ( .A1(n16625), .A2(n19964), .ZN(n16626) );
  AOI211_X1 U19877 ( .C1(n19960), .C2(n16628), .A(n16627), .B(n16626), .ZN(
        n16631) );
  NAND2_X1 U19878 ( .A1(n16629), .A2(n16632), .ZN(n16630) );
  OAI211_X1 U19879 ( .C1(n16633), .C2(n16632), .A(n16631), .B(n16630), .ZN(
        n16634) );
  AOI21_X1 U19880 ( .B1(n16635), .B2(n17444), .A(n16634), .ZN(n16636) );
  OAI21_X1 U19881 ( .B1(n16637), .B2(n19963), .A(n16636), .ZN(P2_U3034) );
  AOI21_X1 U19882 ( .B1(n16638), .B2(n9852), .A(n16672), .ZN(n16659) );
  AND2_X1 U19883 ( .A1(n16658), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16639) );
  NAND2_X1 U19884 ( .A1(n16665), .A2(n16639), .ZN(n16656) );
  AOI21_X1 U19885 ( .B1(n16659), .B2(n16656), .A(n16640), .ZN(n16647) );
  NAND3_X1 U19886 ( .A1(n16665), .A2(n16641), .A3(n16640), .ZN(n16645) );
  OAI21_X1 U19887 ( .B1(n19760), .B2(n19964), .A(n16642), .ZN(n16643) );
  INV_X1 U19888 ( .A(n16643), .ZN(n16644) );
  OAI211_X1 U19889 ( .C1(n19949), .C2(n19755), .A(n16645), .B(n16644), .ZN(
        n16646) );
  AOI211_X1 U19890 ( .C1(n16648), .C2(n17444), .A(n16647), .B(n16646), .ZN(
        n16649) );
  OAI21_X1 U19891 ( .B1(n16650), .B2(n19963), .A(n16649), .ZN(P2_U3035) );
  INV_X1 U19892 ( .A(n16651), .ZN(n16661) );
  INV_X1 U19893 ( .A(n16652), .ZN(n16655) );
  NOR2_X1 U19894 ( .A1(n16653), .A2(n19949), .ZN(n16654) );
  AOI211_X1 U19895 ( .C1(n19858), .C2(n19944), .A(n16655), .B(n16654), .ZN(
        n16657) );
  OAI211_X1 U19896 ( .C1(n16659), .C2(n16658), .A(n16657), .B(n16656), .ZN(
        n16660) );
  AOI21_X1 U19897 ( .B1(n16661), .B2(n17444), .A(n16660), .ZN(n16662) );
  OAI21_X1 U19898 ( .B1(n16663), .B2(n19963), .A(n16662), .ZN(P2_U3036) );
  NAND3_X1 U19899 ( .A1(n16664), .A2(n19946), .A3(n16353), .ZN(n16674) );
  INV_X1 U19900 ( .A(n16665), .ZN(n16670) );
  AOI21_X1 U19901 ( .B1(n16667), .B2(n19944), .A(n16666), .ZN(n16669) );
  NAND2_X1 U19902 ( .A1(n19785), .A2(n19960), .ZN(n16668) );
  OAI211_X1 U19903 ( .C1(n16670), .C2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16669), .B(n16668), .ZN(n16671) );
  AOI21_X1 U19904 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16672), .A(
        n16671), .ZN(n16673) );
  OAI211_X1 U19905 ( .C1(n16675), .C2(n19974), .A(n16674), .B(n16673), .ZN(
        P2_U3037) );
  NAND3_X1 U19906 ( .A1(n16676), .A2(n19946), .A3(n16392), .ZN(n16687) );
  NAND2_X1 U19907 ( .A1(n16678), .A2(n19944), .ZN(n16680) );
  OAI211_X1 U19908 ( .C1(n19949), .C2(n16681), .A(n16680), .B(n16679), .ZN(
        n16685) );
  OAI21_X1 U19909 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16682), .ZN(n16683) );
  NOR2_X1 U19910 ( .A1(n16695), .A2(n16683), .ZN(n16684) );
  AOI211_X1 U19911 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n10182), .A(
        n16685), .B(n16684), .ZN(n16686) );
  OAI211_X1 U19912 ( .C1(n16688), .C2(n19974), .A(n16687), .B(n16686), .ZN(
        P2_U3038) );
  NAND2_X1 U19913 ( .A1(n10182), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16694) );
  NOR2_X1 U19914 ( .A1(n16689), .A2(n19949), .ZN(n16690) );
  AOI211_X1 U19915 ( .C1(n19944), .C2(n16692), .A(n16691), .B(n16690), .ZN(
        n16693) );
  OAI211_X1 U19916 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16695), .A(
        n16694), .B(n16693), .ZN(n16696) );
  AOI21_X1 U19917 ( .B1(n16697), .B2(n17444), .A(n16696), .ZN(n16698) );
  OAI21_X1 U19918 ( .B1(n16699), .B2(n19963), .A(n16698), .ZN(P2_U3039) );
  NAND2_X1 U19919 ( .A1(n16700), .A2(n17444), .ZN(n16710) );
  OAI211_X1 U19920 ( .C1(n16703), .C2(n19964), .A(n16702), .B(n16701), .ZN(
        n16707) );
  NOR2_X1 U19921 ( .A1(n16705), .A2(n16704), .ZN(n16706) );
  AOI211_X1 U19922 ( .C1(n19960), .C2(n16708), .A(n16707), .B(n16706), .ZN(
        n16709) );
  OAI211_X1 U19923 ( .C1(n16711), .C2(n19963), .A(n16710), .B(n16709), .ZN(
        P2_U3040) );
  NAND2_X1 U19924 ( .A1(n16712), .A2(n19946), .ZN(n16721) );
  OAI211_X1 U19925 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n16714), .B(n16713), .ZN(n16718) );
  INV_X1 U19926 ( .A(n16715), .ZN(n16716) );
  AOI21_X1 U19927 ( .B1(n19800), .B2(n19944), .A(n16716), .ZN(n16717) );
  OAI211_X1 U19928 ( .C1(n19793), .C2(n19949), .A(n16718), .B(n16717), .ZN(
        n16719) );
  AOI21_X1 U19929 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16727), .A(
        n16719), .ZN(n16720) );
  OAI211_X1 U19930 ( .C1(n16722), .C2(n19974), .A(n16721), .B(n16720), .ZN(
        P2_U3041) );
  NAND2_X1 U19931 ( .A1(n16723), .A2(n17444), .ZN(n16731) );
  INV_X1 U19932 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20546) );
  OAI22_X1 U19933 ( .A1(n19949), .A2(n19811), .B1(n20546), .B2(n10176), .ZN(
        n16729) );
  INV_X1 U19934 ( .A(n16724), .ZN(n16726) );
  MUX2_X1 U19935 ( .A(n16727), .B(n16726), .S(n16725), .Z(n16728) );
  AOI211_X1 U19936 ( .C1(n19862), .C2(n19944), .A(n16729), .B(n16728), .ZN(
        n16730) );
  OAI211_X1 U19937 ( .C1(n16732), .C2(n19963), .A(n16731), .B(n16730), .ZN(
        P2_U3042) );
  INV_X1 U19938 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20545) );
  OAI22_X1 U19939 ( .A1(n16733), .A2(n19964), .B1(n20545), .B2(n10176), .ZN(
        n16739) );
  NAND2_X1 U19940 ( .A1(n16736), .A2(n9852), .ZN(n16734) );
  OAI22_X1 U19941 ( .A1(n16737), .A2(n16736), .B1(n16735), .B2(n16734), .ZN(
        n16738) );
  AOI211_X1 U19942 ( .C1(n19960), .C2(n20607), .A(n16739), .B(n16738), .ZN(
        n16742) );
  NAND2_X1 U19943 ( .A1(n16740), .A2(n19946), .ZN(n16741) );
  OAI211_X1 U19944 ( .C1(n16743), .C2(n19974), .A(n16742), .B(n16741), .ZN(
        P2_U3043) );
  OAI21_X1 U19945 ( .B1(n16746), .B2(n16745), .A(n16744), .ZN(n16748) );
  NAND2_X1 U19946 ( .A1(n16759), .A2(n10204), .ZN(n16747) );
  OAI211_X1 U19947 ( .C1(n19965), .C2(n16767), .A(n16748), .B(n16747), .ZN(
        n16865) );
  AOI21_X1 U19948 ( .B1(n19839), .B2(n16749), .A(n16877), .ZN(n16770) );
  NAND2_X1 U19949 ( .A1(n19815), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16750) );
  AND2_X1 U19950 ( .A1(n16751), .A2(n16750), .ZN(n16754) );
  AOI222_X1 U19951 ( .A1(n16865), .A2(n19730), .B1(n16770), .B2(n16754), .C1(
        n16883), .C2(n16797), .ZN(n16753) );
  NAND2_X1 U19952 ( .A1(n16773), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16752) );
  OAI21_X1 U19953 ( .B1(n16753), .B2(n16773), .A(n16752), .ZN(P2_U3600) );
  INV_X1 U19954 ( .A(n16754), .ZN(n16771) );
  NAND2_X1 U19955 ( .A1(n16756), .A2(n16755), .ZN(n16763) );
  INV_X1 U19956 ( .A(n16763), .ZN(n16761) );
  NOR2_X1 U19957 ( .A1(n16758), .A2(n16757), .ZN(n16760) );
  AOI22_X1 U19958 ( .A1(n16762), .A2(n16761), .B1(n16760), .B2(n16759), .ZN(
        n16766) );
  NAND2_X1 U19959 ( .A1(n16764), .A2(n16763), .ZN(n16765) );
  OAI211_X1 U19960 ( .C1(n16768), .C2(n16767), .A(n16766), .B(n16765), .ZN(
        n16842) );
  AOI222_X1 U19961 ( .A1(n16771), .A2(n16770), .B1(n16769), .B2(n16883), .C1(
        n16842), .C2(n19730), .ZN(n16774) );
  NAND2_X1 U19962 ( .A1(n16773), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16772) );
  OAI21_X1 U19963 ( .B1(n16774), .B2(n16773), .A(n16772), .ZN(P2_U3599) );
  AND2_X1 U19964 ( .A1(n20627), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n16817) );
  NAND2_X1 U19965 ( .A1(n16817), .A2(n20080), .ZN(n16793) );
  OAI21_X1 U19966 ( .B1(n16782), .B2(n20619), .A(n16814), .ZN(n16781) );
  NOR2_X4 U19967 ( .A1(n20116), .A2(n20079), .ZN(n20097) );
  INV_X1 U19969 ( .A(n20073), .ZN(n16776) );
  AOI21_X1 U19970 ( .B1(n20109), .B2(n16776), .A(n20408), .ZN(n16779) );
  INV_X1 U19971 ( .A(n16777), .ZN(n16821) );
  INV_X1 U19972 ( .A(n20080), .ZN(n16778) );
  NOR2_X1 U19973 ( .A1(n16821), .A2(n16778), .ZN(n16783) );
  NOR3_X1 U19974 ( .A1(n16779), .A2(n16783), .A3(n20614), .ZN(n16780) );
  OAI21_X1 U19975 ( .B1(n16782), .B2(n20071), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16785) );
  INV_X1 U19976 ( .A(n16783), .ZN(n16784) );
  NAND2_X1 U19977 ( .A1(n16785), .A2(n16784), .ZN(n20072) );
  INV_X1 U19978 ( .A(n20461), .ZN(n20406) );
  AOI22_X1 U19979 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16791), .ZN(n20419) );
  INV_X1 U19980 ( .A(n20473), .ZN(n20379) );
  AOI22_X1 U19981 ( .A1(n20097), .A2(n20470), .B1(n20073), .B2(n20379), .ZN(
        n16792) );
  OAI21_X1 U19982 ( .B1(n20406), .B2(n16793), .A(n16792), .ZN(n16794) );
  AOI21_X1 U19983 ( .B1(n20072), .B2(n20462), .A(n16794), .ZN(n16795) );
  OAI21_X1 U19984 ( .B1(n20077), .B2(n16796), .A(n16795), .ZN(P2_U3064) );
  OAI21_X1 U19985 ( .B1(n20177), .B2(n20218), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16800) );
  OR2_X1 U19986 ( .A1(n20111), .A2(n20145), .ZN(n16807) );
  NAND2_X1 U19987 ( .A1(n16800), .A2(n16807), .ZN(n16806) );
  NAND3_X1 U19988 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20618), .ZN(n20200) );
  INV_X1 U19989 ( .A(n20189), .ZN(n16801) );
  NAND2_X1 U19990 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16801), .ZN(n16802) );
  OAI211_X1 U19991 ( .C1(n20189), .C2(n16814), .A(n16809), .B(n20467), .ZN(
        n16804) );
  INV_X1 U19992 ( .A(n16804), .ZN(n16805) );
  INV_X1 U19993 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16812) );
  AOI22_X1 U19994 ( .A1(n20218), .A2(n20470), .B1(n20177), .B2(n20379), .ZN(
        n16811) );
  OAI21_X1 U19995 ( .B1(n16807), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20619), 
        .ZN(n16808) );
  AOI22_X1 U19996 ( .A1(n20190), .A2(n20462), .B1(n20461), .B2(n20189), .ZN(
        n16810) );
  OAI211_X1 U19997 ( .C1(n20180), .C2(n16812), .A(n16811), .B(n16810), .ZN(
        P2_U3096) );
  AND2_X1 U19998 ( .A1(n16860), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16831) );
  AOI221_X1 U19999 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20311), .C1(
        P2_STATEBS16_REG_SCAN_IN), .C2(n20325), .A(n20290), .ZN(n16816) );
  OAI21_X1 U20000 ( .B1(n16819), .B2(n20619), .A(n16814), .ZN(n16815) );
  NOR2_X1 U20001 ( .A1(n16816), .A2(n16815), .ZN(n16818) );
  INV_X1 U20002 ( .A(n20312), .ZN(n16825) );
  AOI22_X1 U20003 ( .A1(n20325), .A2(n20470), .B1(n20311), .B2(n20379), .ZN(
        n16823) );
  INV_X1 U20004 ( .A(n16831), .ZN(n16826) );
  OAI21_X1 U20005 ( .B1(n16819), .B2(n20309), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16820) );
  AOI22_X1 U20006 ( .A1(n20310), .A2(n20462), .B1(n20309), .B2(n20461), .ZN(
        n16822) );
  OAI211_X1 U20007 ( .C1(n16825), .C2(n16824), .A(n16823), .B(n16822), .ZN(
        P2_U3128) );
  NAND2_X1 U20008 ( .A1(n20610), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20466) );
  OAI22_X1 U20009 ( .A1(n20466), .A2(n20079), .B1(n20335), .B2(n16826), .ZN(
        n16830) );
  NAND2_X1 U20010 ( .A1(n16831), .A2(n20078), .ZN(n16835) );
  NAND2_X1 U20011 ( .A1(n16835), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16827) );
  NAND2_X1 U20012 ( .A1(n16835), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16829) );
  NAND4_X1 U20013 ( .A1(n16830), .A2(n20467), .A3(n16834), .A4(n16829), .ZN(
        n20330) );
  INV_X1 U20014 ( .A(n20330), .ZN(n16839) );
  AOI22_X1 U20015 ( .A1(n20340), .A2(n20470), .B1(n20325), .B2(n20379), .ZN(
        n16837) );
  NAND3_X1 U20016 ( .A1(n16831), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        n16814), .ZN(n16832) );
  NAND2_X1 U20017 ( .A1(n16832), .A2(n20619), .ZN(n16833) );
  INV_X1 U20018 ( .A(n16835), .ZN(n20328) );
  AOI22_X1 U20019 ( .A1(n20329), .A2(n20462), .B1(n20461), .B2(n20328), .ZN(
        n16836) );
  OAI211_X1 U20020 ( .C1(n16839), .C2(n16838), .A(n16837), .B(n16836), .ZN(
        P2_U3136) );
  NAND2_X1 U20021 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n16895) );
  INV_X1 U20022 ( .A(n16840), .ZN(n16879) );
  MUX2_X1 U20023 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16841), .S(
        n16863), .Z(n16876) );
  INV_X1 U20024 ( .A(n16842), .ZN(n16843) );
  MUX2_X1 U20025 ( .A(n10958), .B(n16843), .S(n16863), .Z(n16859) );
  INV_X1 U20026 ( .A(n16859), .ZN(n16875) );
  MUX2_X1 U20027 ( .A(n16846), .B(n16845), .S(n16844), .Z(n16850) );
  NAND2_X1 U20028 ( .A1(n16848), .A2(n16847), .ZN(n16849) );
  AND2_X1 U20029 ( .A1(n16850), .A2(n16849), .ZN(n20635) );
  INV_X1 U20030 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n16852) );
  AOI21_X1 U20031 ( .B1(n16853), .B2(n16852), .A(n16851), .ZN(n16854) );
  AOI211_X1 U20032 ( .C1(n16857), .C2(n16856), .A(n16855), .B(n16854), .ZN(
        n16858) );
  OAI211_X1 U20033 ( .C1(n16863), .C2(n17301), .A(n20635), .B(n16858), .ZN(
        n16874) );
  NOR2_X1 U20034 ( .A1(n16859), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16861) );
  AOI22_X1 U20035 ( .A1(n16861), .A2(n16860), .B1(n16876), .B2(n20618), .ZN(
        n16872) );
  INV_X1 U20036 ( .A(n16861), .ZN(n16862) );
  NAND2_X1 U20037 ( .A1(n16862), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16870) );
  INV_X1 U20038 ( .A(n16863), .ZN(n16867) );
  AOI21_X1 U20039 ( .B1(n16868), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16864) );
  NOR2_X1 U20040 ( .A1(n16865), .A2(n16864), .ZN(n16866) );
  AOI211_X1 U20041 ( .C1(n20078), .C2(n16868), .A(n16867), .B(n16866), .ZN(
        n16869) );
  OAI211_X1 U20042 ( .C1(n16876), .C2(n20618), .A(n16870), .B(n16869), .ZN(
        n16871) );
  AOI21_X1 U20043 ( .B1(n16872), .B2(n16871), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16873) );
  AOI211_X1 U20044 ( .C1(n16876), .C2(n16875), .A(n16874), .B(n16873), .ZN(
        n16889) );
  AOI21_X1 U20045 ( .B1(n16889), .B2(n16877), .A(n16902), .ZN(n16878) );
  AOI21_X1 U20046 ( .B1(n16880), .B2(n16879), .A(n16878), .ZN(n16882) );
  INV_X1 U20047 ( .A(n16882), .ZN(n16894) );
  NAND2_X1 U20048 ( .A1(n16882), .A2(n16881), .ZN(n16897) );
  NOR2_X1 U20049 ( .A1(n16883), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16885) );
  OAI22_X1 U20050 ( .A1(n16897), .A2(n16887), .B1(n16885), .B2(n16884), .ZN(
        n16893) );
  NAND2_X1 U20051 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20619), .ZN(n16896) );
  OAI21_X1 U20052 ( .B1(n16887), .B2(n16896), .A(n16886), .ZN(n16891) );
  NOR2_X1 U20053 ( .A1(n16889), .A2(n16888), .ZN(n16890) );
  AOI211_X1 U20054 ( .C1(n16904), .C2(n20629), .A(n16891), .B(n16890), .ZN(
        n16892) );
  OAI211_X1 U20055 ( .C1(n16895), .C2(n16894), .A(n16893), .B(n16892), .ZN(
        P2_U3176) );
  INV_X1 U20056 ( .A(n16897), .ZN(n16903) );
  INV_X1 U20057 ( .A(n16896), .ZN(n19729) );
  OAI211_X1 U20058 ( .C1(n16903), .C2(n19729), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n20532), .ZN(n16901) );
  NOR3_X1 U20059 ( .A1(n20532), .A2(n16902), .A3(n17296), .ZN(n16898) );
  OAI21_X1 U20060 ( .B1(n16899), .B2(n16898), .A(n16897), .ZN(n16900) );
  NAND3_X1 U20061 ( .A1(n16901), .A2(n19838), .A3(n16900), .ZN(P2_U3177) );
  OAI21_X1 U20062 ( .B1(n16903), .B2(n16902), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n16906) );
  INV_X1 U20063 ( .A(n16904), .ZN(n16905) );
  NAND2_X1 U20064 ( .A1(n16906), .A2(n16905), .ZN(P2_U3593) );
  NAND2_X1 U20065 ( .A1(n19543), .A2(n16907), .ZN(n16908) );
  OR2_X2 U20066 ( .A1(n17547), .A2(n18494), .ZN(n18813) );
  OR2_X2 U20067 ( .A1(n17547), .A2(n19709), .ZN(n18817) );
  INV_X2 U20068 ( .A(n18602), .ZN(n18716) );
  NOR2_X4 U20069 ( .A1(n19390), .A2(n19252), .ZN(n16915) );
  AOI21_X1 U20070 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16914), .A(
        n16915), .ZN(n18598) );
  INV_X1 U20071 ( .A(n18598), .ZN(n16999) );
  NAND2_X1 U20072 ( .A1(n16916), .A2(n16999), .ZN(n16935) );
  XNOR2_X1 U20073 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16913) );
  NOR2_X2 U20074 ( .A1(n18769), .A2(n18790), .ZN(n18820) );
  AND2_X2 U20075 ( .A1(n18820), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18675) );
  AOI21_X1 U20076 ( .B1(n18675), .B2(n17843), .A(n16911), .ZN(n16912) );
  OAI21_X1 U20077 ( .B1(n16935), .B2(n16913), .A(n16912), .ZN(n16919) );
  NOR2_X1 U20078 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18595), .ZN(
        n16943) );
  OR2_X1 U20079 ( .A1(n19206), .A2(n16916), .ZN(n16946) );
  OAI211_X1 U20080 ( .C1(n16917), .C2(n18672), .A(n18810), .B(n16946), .ZN(
        n16942) );
  NOR2_X1 U20081 ( .A1(n16943), .A2(n16942), .ZN(n16931) );
  INV_X1 U20082 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17572) );
  NOR2_X1 U20083 ( .A1(n16931), .A2(n17572), .ZN(n16918) );
  AOI211_X1 U20084 ( .C1(n18716), .C2(n16920), .A(n16919), .B(n16918), .ZN(
        n16921) );
  OAI211_X1 U20085 ( .C1(n16923), .C2(n18813), .A(n16922), .B(n16921), .ZN(
        P3_U2799) );
  OAI21_X1 U20086 ( .B1(n16925), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16924), .ZN(n17081) );
  INV_X1 U20087 ( .A(n17071), .ZN(n17077) );
  OR2_X1 U20088 ( .A1(n16926), .A2(n17098), .ZN(n17076) );
  OR2_X1 U20089 ( .A1(n17076), .A2(n18817), .ZN(n16941) );
  OAI21_X1 U20090 ( .B1(n17077), .B2(n18813), .A(n16941), .ZN(n16951) );
  NAND2_X1 U20091 ( .A1(n18972), .A2(n18780), .ZN(n16928) );
  NAND2_X1 U20092 ( .A1(n18716), .A2(n18713), .ZN(n16927) );
  NOR2_X1 U20093 ( .A1(n18588), .A2(n17097), .ZN(n18546) );
  INV_X1 U20094 ( .A(n18546), .ZN(n16930) );
  NOR3_X1 U20095 ( .A1(n16930), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16929), .ZN(n16937) );
  INV_X1 U20096 ( .A(n16931), .ZN(n16932) );
  NAND2_X1 U20097 ( .A1(n16932), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16934) );
  AND2_X1 U20098 ( .A1(n18905), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17072) );
  AOI21_X1 U20099 ( .B1(n18675), .B2(n17566), .A(n17072), .ZN(n16933) );
  OAI211_X1 U20100 ( .C1(n16935), .C2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16934), .B(n16933), .ZN(n16936) );
  AOI211_X1 U20101 ( .C1(n16951), .C2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16937), .B(n16936), .ZN(n16938) );
  OAI21_X1 U20102 ( .B1(n17081), .B2(n18641), .A(n16938), .ZN(P3_U2800) );
  NAND2_X1 U20103 ( .A1(n16956), .A2(n16939), .ZN(n16940) );
  XNOR2_X1 U20104 ( .A(n16940), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17094) );
  INV_X1 U20105 ( .A(n16941), .ZN(n16950) );
  NAND2_X1 U20106 ( .A1(n16958), .A2(n16947), .ZN(n17068) );
  INV_X1 U20107 ( .A(n17068), .ZN(n17099) );
  AOI22_X1 U20108 ( .A1(n18905), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16942), .ZN(n16945) );
  OAI21_X1 U20109 ( .B1(n16943), .B2(n18675), .A(n17576), .ZN(n16944) );
  OAI211_X1 U20110 ( .C1(n16946), .C2(n9797), .A(n16945), .B(n16944), .ZN(
        n16949) );
  INV_X1 U20111 ( .A(n16947), .ZN(n17103) );
  NOR4_X1 U20112 ( .A1(n17077), .A2(n17118), .A3(n17103), .A4(n18813), .ZN(
        n16948) );
  AOI211_X1 U20113 ( .C1(n16950), .C2(n17099), .A(n16949), .B(n16948), .ZN(
        n16953) );
  NAND2_X1 U20114 ( .A1(n16951), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16952) );
  OAI211_X1 U20115 ( .C1(n17094), .C2(n18641), .A(n16953), .B(n16952), .ZN(
        P3_U2801) );
  NAND2_X1 U20116 ( .A1(n18694), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16954) );
  NAND2_X1 U20117 ( .A1(n16955), .A2(n16954), .ZN(n17108) );
  NAND2_X1 U20118 ( .A1(n16957), .A2(n16956), .ZN(n16971) );
  OAI22_X1 U20119 ( .A1(n18813), .A2(n16959), .B1(n18602), .B2(n16958), .ZN(
        n16979) );
  OR2_X1 U20120 ( .A1(n18830), .A2(n16979), .ZN(n18545) );
  OAI211_X1 U20121 ( .C1(n18780), .C2(n18716), .A(n18545), .B(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16970) );
  INV_X1 U20122 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16960) );
  NAND3_X1 U20123 ( .A1(n18546), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16960), .ZN(n16969) );
  INV_X1 U20124 ( .A(n18672), .ZN(n18552) );
  AOI22_X1 U20125 ( .A1(n11500), .A2(n18790), .B1(n16961), .B2(n18552), .ZN(
        n16962) );
  AND2_X1 U20126 ( .A1(n18810), .A2(n16962), .ZN(n16977) );
  OAI21_X1 U20127 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18595), .A(
        n16977), .ZN(n18539) );
  AOI22_X1 U20128 ( .A1(n18905), .A2(P3_REIP_REG_28__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18539), .ZN(n16965) );
  NOR2_X1 U20129 ( .A1(n18598), .A2(n11500), .ZN(n18544) );
  OAI211_X1 U20130 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n18544), .B(n16963), .ZN(n16964) );
  OAI211_X1 U20131 ( .C1(n18686), .C2(n16966), .A(n16965), .B(n16964), .ZN(
        n16967) );
  INV_X1 U20132 ( .A(n16967), .ZN(n16968) );
  NAND4_X1 U20133 ( .A1(n16971), .A2(n16970), .A3(n16969), .A4(n16968), .ZN(
        P3_U2802) );
  XNOR2_X1 U20134 ( .A(n16972), .B(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17129) );
  AOI21_X1 U20135 ( .B1(n16973), .B2(n16915), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16976) );
  INV_X1 U20136 ( .A(n18595), .ZN(n16974) );
  OAI21_X1 U20137 ( .B1(n18675), .B2(n16974), .A(n17610), .ZN(n16975) );
  NAND2_X1 U20138 ( .A1(n18905), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17123) );
  OAI211_X1 U20139 ( .C1(n16977), .C2(n16976), .A(n16975), .B(n17123), .ZN(
        n16978) );
  AOI221_X1 U20140 ( .B1(n16980), .B2(n17124), .C1(n16979), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n16978), .ZN(n16981) );
  OAI21_X1 U20141 ( .B1(n18641), .B2(n17129), .A(n16981), .ZN(P3_U2804) );
  AND2_X1 U20142 ( .A1(n18694), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18615) );
  NOR2_X1 U20143 ( .A1(n18649), .A2(n18615), .ZN(n16982) );
  XOR2_X1 U20144 ( .A(n16982), .B(n18614), .Z(n17143) );
  NAND2_X1 U20145 ( .A1(n18713), .A2(n13551), .ZN(n17132) );
  NAND2_X1 U20146 ( .A1(n18716), .A2(n17132), .ZN(n18699) );
  OAI21_X1 U20147 ( .B1(n18937), .B2(n18813), .A(n18699), .ZN(n18633) );
  INV_X1 U20148 ( .A(n18633), .ZN(n18683) );
  OAI21_X1 U20149 ( .B1(n17131), .B2(n18684), .A(n18683), .ZN(n18663) );
  INV_X1 U20150 ( .A(n17131), .ZN(n16983) );
  NOR2_X1 U20151 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16983), .ZN(
        n17139) );
  INV_X1 U20152 ( .A(n17139), .ZN(n16988) );
  NOR2_X1 U20153 ( .A1(n18598), .A2(n11504), .ZN(n18643) );
  INV_X1 U20154 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16986) );
  AOI21_X1 U20155 ( .B1(n18790), .B2(n11504), .A(n18769), .ZN(n18658) );
  OAI21_X1 U20156 ( .B1(n16984), .B2(n18672), .A(n18658), .ZN(n18647) );
  NAND2_X1 U20157 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16984), .ZN(
        n17689) );
  OAI21_X1 U20158 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16984), .A(
        n17689), .ZN(n17698) );
  NAND2_X1 U20159 ( .A1(n18905), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17141) );
  OAI21_X1 U20160 ( .B1(n18686), .B2(n17698), .A(n17141), .ZN(n16985) );
  AOI221_X1 U20161 ( .B1(n18643), .B2(n16986), .C1(n18647), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n16985), .ZN(n16987) );
  OAI21_X1 U20162 ( .B1(n18684), .B2(n16988), .A(n16987), .ZN(n16989) );
  AOI21_X1 U20163 ( .B1(n18663), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16989), .ZN(n16990) );
  OAI21_X1 U20164 ( .B1(n18641), .B2(n17143), .A(n16990), .ZN(P3_U2812) );
  NOR2_X1 U20165 ( .A1(n13637), .A2(n18575), .ZN(n17031) );
  NAND2_X1 U20166 ( .A1(n17031), .A2(n18977), .ZN(n17003) );
  NOR2_X1 U20167 ( .A1(n17047), .A2(n18694), .ZN(n18722) );
  INV_X1 U20168 ( .A(n18722), .ZN(n16992) );
  NOR2_X1 U20169 ( .A1(n16992), .A2(n16991), .ZN(n17023) );
  NAND2_X1 U20170 ( .A1(n17023), .A2(n17029), .ZN(n18710) );
  AOI22_X1 U20171 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17003), .B1(
        n18710), .B2(n18969), .ZN(n16993) );
  XOR2_X1 U20172 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n16993), .Z(
        n18951) );
  INV_X1 U20173 ( .A(n17026), .ZN(n18725) );
  NAND2_X1 U20174 ( .A1(n18939), .A2(n18940), .ZN(n18961) );
  NOR2_X1 U20175 ( .A1(n13637), .A2(n16994), .ZN(n18953) );
  OAI22_X1 U20176 ( .A1(n10223), .A2(n18813), .B1(n18953), .B2(n18602), .ZN(
        n17012) );
  NAND2_X1 U20177 ( .A1(n17012), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16998) );
  INV_X1 U20178 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17762) );
  INV_X1 U20179 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17009) );
  NAND2_X1 U20180 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17743), .ZN(
        n17018) );
  NOR2_X1 U20181 ( .A1(n17009), .A2(n17018), .ZN(n17005) );
  INV_X1 U20182 ( .A(n17005), .ZN(n17759) );
  NOR2_X1 U20183 ( .A1(n17744), .A2(n17018), .ZN(n17746) );
  AOI21_X1 U20184 ( .B1(n17762), .B2(n17759), .A(n17746), .ZN(n17757) );
  INV_X1 U20185 ( .A(n18790), .ZN(n17051) );
  OAI21_X1 U20186 ( .B1(n17743), .B2(n17051), .A(n18672), .ZN(n16995) );
  AOI21_X1 U20187 ( .B1(n17018), .B2(n16995), .A(n18769), .ZN(n17008) );
  INV_X1 U20188 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19642) );
  OAI22_X1 U20189 ( .A1(n17008), .A2(n17762), .B1(n18992), .B2(n19642), .ZN(
        n16996) );
  AOI21_X1 U20190 ( .B1(n18675), .B2(n17757), .A(n16996), .ZN(n16997) );
  OAI211_X1 U20191 ( .C1(n18725), .C2(n18961), .A(n16998), .B(n16997), .ZN(
        n17001) );
  NAND2_X1 U20192 ( .A1(n17743), .A2(n16999), .ZN(n18676) );
  AOI211_X1 U20193 ( .C1(n17009), .C2(n17762), .A(n18703), .B(n18676), .ZN(
        n17000) );
  AOI211_X1 U20194 ( .C1(n18951), .C2(n18728), .A(n17001), .B(n17000), .ZN(
        n17002) );
  INV_X1 U20195 ( .A(n17002), .ZN(P3_U2817) );
  NAND2_X1 U20196 ( .A1(n17003), .A2(n18710), .ZN(n17004) );
  XOR2_X1 U20197 ( .A(n17004), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18965) );
  INV_X1 U20198 ( .A(n18965), .ZN(n17014) );
  AOI21_X1 U20199 ( .B1(n17009), .B2(n17018), .A(n17005), .ZN(n17772) );
  INV_X1 U20200 ( .A(n17772), .ZN(n17007) );
  NAND2_X1 U20201 ( .A1(n18977), .A2(n18969), .ZN(n17006) );
  OAI22_X1 U20202 ( .A1(n18686), .A2(n17007), .B1(n18725), .B2(n17006), .ZN(
        n17011) );
  NAND2_X1 U20203 ( .A1(n18905), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18967) );
  OAI221_X1 U20204 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18676), .C1(
        n17009), .C2(n17008), .A(n18967), .ZN(n17010) );
  AOI211_X1 U20205 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17012), .A(
        n17011), .B(n17010), .ZN(n17013) );
  OAI21_X1 U20206 ( .B1(n18641), .B2(n17014), .A(n17013), .ZN(P3_U2818) );
  NAND2_X1 U20207 ( .A1(n18716), .A2(n13637), .ZN(n17048) );
  OR2_X1 U20208 ( .A1(n18813), .A2(n18972), .ZN(n17015) );
  AND2_X1 U20209 ( .A1(n17048), .A2(n17015), .ZN(n17037) );
  OAI21_X1 U20210 ( .B1(n18725), .B2(n18976), .A(n17037), .ZN(n18727) );
  INV_X1 U20211 ( .A(n18727), .ZN(n17030) );
  NAND2_X1 U20212 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17016), .ZN(
        n17842) );
  INV_X1 U20213 ( .A(n17842), .ZN(n17832) );
  NAND2_X1 U20214 ( .A1(n17017), .A2(n17832), .ZN(n17794) );
  INV_X1 U20215 ( .A(n17018), .ZN(n17019) );
  AOI21_X1 U20216 ( .B1(n17793), .B2(n17794), .A(n17019), .ZN(n17785) );
  OR2_X2 U20217 ( .A1(n18675), .A2(n16974), .ZN(n18808) );
  INV_X1 U20218 ( .A(n17033), .ZN(n17806) );
  NOR3_X1 U20219 ( .A1(n19206), .A2(n17020), .A3(n17846), .ZN(n18754) );
  NAND2_X1 U20220 ( .A1(n17806), .A2(n18754), .ZN(n17036) );
  NOR2_X1 U20221 ( .A1(n17035), .A2(n17036), .ZN(n18730) );
  NAND2_X1 U20222 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18730), .ZN(
        n18729) );
  AND2_X1 U20223 ( .A1(n16915), .A2(n17743), .ZN(n18702) );
  AOI211_X1 U20224 ( .C1(n18729), .C2(n17793), .A(n18820), .B(n18702), .ZN(
        n17022) );
  INV_X1 U20225 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19638) );
  NOR2_X1 U20226 ( .A1(n18992), .A2(n19638), .ZN(n17021) );
  AOI211_X1 U20227 ( .C1(n17785), .C2(n18808), .A(n17022), .B(n17021), .ZN(
        n17028) );
  NAND2_X1 U20228 ( .A1(n18976), .A2(n17029), .ZN(n18982) );
  INV_X1 U20229 ( .A(n18982), .ZN(n17025) );
  INV_X1 U20230 ( .A(n17031), .ZN(n18708) );
  NOR2_X1 U20231 ( .A1(n18708), .A2(n19000), .ZN(n18721) );
  AOI21_X1 U20232 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18721), .A(
        n17023), .ZN(n17024) );
  XOR2_X1 U20233 ( .A(n17029), .B(n17024), .Z(n18970) );
  AOI22_X1 U20234 ( .A1(n17026), .A2(n17025), .B1(n18728), .B2(n18970), .ZN(
        n17027) );
  OAI211_X1 U20235 ( .C1(n17030), .C2(n17029), .A(n17028), .B(n17027), .ZN(
        P3_U2819) );
  NOR2_X1 U20236 ( .A1(n18722), .A2(n17031), .ZN(n17032) );
  XNOR2_X1 U20237 ( .A(n17032), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18996) );
  INV_X1 U20238 ( .A(n18996), .ZN(n17042) );
  NOR2_X1 U20239 ( .A1(n17033), .A2(n17842), .ZN(n17046) );
  NAND2_X1 U20240 ( .A1(n17034), .A2(n17832), .ZN(n17796) );
  OAI21_X1 U20241 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17046), .A(
        n17796), .ZN(n17812) );
  INV_X1 U20242 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19634) );
  OAI22_X1 U20243 ( .A1(n18822), .A2(n17812), .B1(n18992), .B2(n19634), .ZN(
        n17040) );
  AOI211_X1 U20244 ( .C1(n17036), .C2(n17035), .A(n18820), .B(n18730), .ZN(
        n17039) );
  OAI22_X1 U20245 ( .A1(n18725), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n17037), .B2(n19000), .ZN(n17038) );
  NOR3_X1 U20246 ( .A1(n17040), .A2(n17039), .A3(n17038), .ZN(n17041) );
  OAI21_X1 U20247 ( .B1(n17042), .B2(n18641), .A(n17041), .ZN(P3_U2821) );
  OR2_X1 U20248 ( .A1(n18691), .A2(n18713), .ZN(n17045) );
  NAND2_X1 U20249 ( .A1(n17043), .A2(n18694), .ZN(n17044) );
  NAND2_X1 U20250 ( .A1(n17045), .A2(n17044), .ZN(n19013) );
  INV_X1 U20251 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17054) );
  NAND2_X1 U20252 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17832), .ZN(
        n17831) );
  AOI21_X1 U20253 ( .B1(n17054), .B2(n17831), .A(n17046), .ZN(n17821) );
  INV_X1 U20254 ( .A(n17047), .ZN(n19010) );
  NOR2_X1 U20255 ( .A1(n17048), .A2(n19010), .ZN(n17059) );
  OAI21_X1 U20256 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17050), .A(
        n17049), .ZN(n19016) );
  OAI21_X1 U20257 ( .B1(n17051), .B2(n17016), .A(n18810), .ZN(n18734) );
  INV_X1 U20258 ( .A(n18734), .ZN(n17055) );
  AOI21_X1 U20259 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17016), .A(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17052) );
  OR3_X1 U20260 ( .A1(n19206), .A2(n17806), .A3(n17052), .ZN(n17053) );
  NAND2_X1 U20261 ( .A1(n18905), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n19018) );
  OAI211_X1 U20262 ( .C1(n17055), .C2(n17054), .A(n17053), .B(n19018), .ZN(
        n17056) );
  INV_X1 U20263 ( .A(n17056), .ZN(n17057) );
  OAI21_X1 U20264 ( .B1(n19016), .B2(n18813), .A(n17057), .ZN(n17058) );
  AOI211_X1 U20265 ( .C1(n17821), .C2(n18808), .A(n17059), .B(n17058), .ZN(
        n17060) );
  OAI21_X1 U20266 ( .B1(n18641), .B2(n19013), .A(n17060), .ZN(P3_U2822) );
  NAND3_X1 U20267 ( .A1(n19592), .A2(n18672), .A3(n18810), .ZN(n17065) );
  NOR2_X1 U20268 ( .A1(n18813), .A2(n17061), .ZN(n17064) );
  OAI22_X1 U20269 ( .A1(n18817), .A2(n17062), .B1(n18992), .B2(n19696), .ZN(
        n17063) );
  AOI211_X1 U20270 ( .C1(n17065), .C2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n17064), .B(n17063), .ZN(n17066) );
  INV_X1 U20271 ( .A(n17066), .ZN(P3_U2830) );
  INV_X1 U20272 ( .A(n18971), .ZN(n18952) );
  OAI22_X1 U20273 ( .A1(n17068), .A2(n18952), .B1(n17103), .B2(n17067), .ZN(
        n17088) );
  NAND3_X1 U20274 ( .A1(n17088), .A2(n19062), .A3(n17069), .ZN(n17070) );
  OAI21_X1 U20275 ( .B1(n17071), .B2(n19095), .A(n17070), .ZN(n17074) );
  AOI21_X1 U20276 ( .B1(n17074), .B2(n17073), .A(n17072), .ZN(n17080) );
  OAI22_X1 U20277 ( .A1(n17077), .A2(n19095), .B1(n17076), .B2(n17075), .ZN(
        n17084) );
  OAI21_X1 U20278 ( .B1(n17084), .B2(n17078), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17079) );
  OAI211_X1 U20279 ( .C1(n17081), .C2(n19012), .A(n17080), .B(n17079), .ZN(
        P3_U2832) );
  INV_X1 U20280 ( .A(n19005), .ZN(n19004) );
  INV_X1 U20281 ( .A(n18978), .ZN(n18983) );
  NAND2_X1 U20282 ( .A1(n18830), .A2(n18983), .ZN(n17082) );
  AND2_X1 U20283 ( .A1(n17083), .A2(n17082), .ZN(n17104) );
  OAI21_X1 U20284 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n19004), .A(
        n17104), .ZN(n17085) );
  AOI211_X1 U20285 ( .C1(n18992), .C2(n17085), .A(n19066), .B(n17084), .ZN(
        n17086) );
  INV_X1 U20286 ( .A(n17086), .ZN(n17092) );
  NOR3_X1 U20287 ( .A1(n17118), .A2(n17103), .A3(n19095), .ZN(n17087) );
  AOI21_X1 U20288 ( .B1(n19062), .B2(n17088), .A(n17087), .ZN(n17090) );
  INV_X1 U20289 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n17089) );
  OAI22_X1 U20290 ( .A1(n17090), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n17089), .B2(n18992), .ZN(n17091) );
  AOI21_X1 U20291 ( .B1(n17092), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17091), .ZN(n17093) );
  OAI21_X1 U20292 ( .B1(n17094), .B2(n19012), .A(n17093), .ZN(P3_U2833) );
  AOI22_X1 U20293 ( .A1(n18972), .A2(n18957), .B1(n18713), .B2(n18971), .ZN(
        n17138) );
  OAI21_X1 U20294 ( .B1(n17138), .B2(n18668), .A(n17095), .ZN(n18863) );
  NAND2_X1 U20295 ( .A1(n18863), .A2(n17096), .ZN(n18857) );
  NOR3_X1 U20296 ( .A1(n18857), .A2(n19082), .A3(n17097), .ZN(n18823) );
  AOI22_X1 U20297 ( .A1(n17101), .A2(n19086), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18823), .ZN(n17114) );
  INV_X1 U20298 ( .A(n19543), .ZN(n17100) );
  NOR3_X1 U20299 ( .A1(n17102), .A2(n17101), .A3(n17100), .ZN(n17107) );
  OAI21_X1 U20300 ( .B1(n17118), .B2(n17103), .A(n18957), .ZN(n17105) );
  NAND3_X1 U20301 ( .A1(n17105), .A2(n17104), .A3(n19090), .ZN(n17106) );
  OAI211_X1 U20302 ( .C1(n17107), .C2(n17106), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18988), .ZN(n17113) );
  NAND2_X1 U20303 ( .A1(n18997), .A2(n17108), .ZN(n17110) );
  INV_X1 U20304 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n17109) );
  OAI22_X1 U20305 ( .A1(n18540), .A2(n17110), .B1(n18992), .B2(n17109), .ZN(
        n17111) );
  INV_X1 U20306 ( .A(n17111), .ZN(n17112) );
  OAI211_X1 U20307 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n17114), .A(
        n17113), .B(n17112), .ZN(P3_U2834) );
  NOR2_X1 U20308 ( .A1(n10220), .A2(n18913), .ZN(n18938) );
  INV_X1 U20309 ( .A(n18938), .ZN(n18994) );
  NOR2_X1 U20310 ( .A1(n18668), .A2(n18994), .ZN(n18919) );
  NAND2_X1 U20311 ( .A1(n17131), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18620) );
  INV_X1 U20312 ( .A(n18620), .ZN(n18872) );
  AOI21_X1 U20313 ( .B1(n18919), .B2(n18872), .A(n18991), .ZN(n18869) );
  NOR2_X1 U20314 ( .A1(n17115), .A2(n18869), .ZN(n18847) );
  OAI21_X1 U20315 ( .B1(n17135), .B2(n17116), .A(n18847), .ZN(n18833) );
  INV_X1 U20316 ( .A(n18825), .ZN(n17127) );
  NAND2_X1 U20317 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17122) );
  NAND3_X1 U20318 ( .A1(n19062), .A2(n17121), .A3(n18863), .ZN(n18855) );
  OAI22_X1 U20319 ( .A1(n17124), .A2(n19082), .B1(n17122), .B2(n18855), .ZN(
        n17126) );
  OAI21_X1 U20320 ( .B1(n19090), .B2(n17124), .A(n17123), .ZN(n17125) );
  AOI21_X1 U20321 ( .B1(n17127), .B2(n17126), .A(n17125), .ZN(n17128) );
  OAI21_X1 U20322 ( .B1(n19012), .B2(n17129), .A(n17128), .ZN(P3_U2836) );
  NAND3_X1 U20323 ( .A1(n18866), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17130), .ZN(n17134) );
  NOR2_X1 U20324 ( .A1(n18957), .A2(n18971), .ZN(n18975) );
  AOI22_X1 U20325 ( .A1(n17131), .A2(n18870), .B1(n18975), .B2(n19546), .ZN(
        n17133) );
  INV_X1 U20326 ( .A(n18957), .ZN(n19545) );
  NAND2_X1 U20327 ( .A1(n17132), .A2(n18971), .ZN(n18930) );
  AOI211_X1 U20328 ( .C1(n19075), .C2(n17134), .A(n17133), .B(n18920), .ZN(
        n18911) );
  AOI221_X1 U20329 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18911), 
        .C1(n17135), .C2(n18911), .A(n18905), .ZN(n17140) );
  INV_X1 U20330 ( .A(n19002), .ZN(n17136) );
  OAI22_X1 U20331 ( .A1(n17136), .A2(n19546), .B1(n19074), .B2(n19003), .ZN(
        n19063) );
  NAND2_X1 U20332 ( .A1(n17137), .A2(n19063), .ZN(n18926) );
  NAND2_X1 U20333 ( .A1(n17138), .A2(n18926), .ZN(n18962) );
  NAND2_X1 U20334 ( .A1(n19062), .A2(n18962), .ZN(n19001) );
  NOR2_X1 U20335 ( .A1(n18668), .A2(n19001), .ZN(n18921) );
  AOI22_X1 U20336 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17140), .B1(
        n18921), .B2(n17139), .ZN(n17142) );
  OAI211_X1 U20337 ( .C1(n17143), .C2(n19012), .A(n17142), .B(n17141), .ZN(
        P3_U2844) );
  INV_X1 U20338 ( .A(n17144), .ZN(n17145) );
  NAND2_X1 U20339 ( .A1(n17145), .A2(n17154), .ZN(n17921) );
  OAI22_X1 U20340 ( .A1(n17147), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n17146), .B2(n17921), .ZN(n19562) );
  INV_X1 U20341 ( .A(n19578), .ZN(n17175) );
  NOR2_X1 U20342 ( .A1(n19592), .A2(n10220), .ZN(n17172) );
  OAI22_X1 U20343 ( .A1(n17148), .A2(n21541), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17170) );
  NAND2_X1 U20344 ( .A1(n17172), .A2(n17170), .ZN(n17149) );
  OAI211_X1 U20345 ( .C1(n17921), .C2(n17175), .A(n17174), .B(n17149), .ZN(
        n17150) );
  AOI21_X1 U20346 ( .B1(n19562), .B2(n17540), .A(n17150), .ZN(n17151) );
  AOI21_X1 U20347 ( .B1(n17178), .B2(n17152), .A(n17151), .ZN(P3_U3289) );
  AND2_X1 U20348 ( .A1(n17153), .A2(n17152), .ZN(n17155) );
  OAI21_X1 U20349 ( .B1(n17156), .B2(n17155), .A(n17154), .ZN(n17161) );
  NAND2_X1 U20350 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18973), .ZN(
        n17158) );
  NAND2_X1 U20351 ( .A1(n17158), .A2(n17157), .ZN(n17159) );
  NAND2_X1 U20352 ( .A1(n17159), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17160) );
  MUX2_X1 U20353 ( .A(n17161), .B(n17160), .S(n9940), .Z(n17169) );
  OAI21_X1 U20354 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n17162), .ZN(n17166) );
  NAND2_X1 U20355 ( .A1(n17164), .A2(n17163), .ZN(n17899) );
  INV_X1 U20356 ( .A(n17899), .ZN(n17165) );
  OAI22_X1 U20357 ( .A1(n19538), .A2(n17166), .B1(n17165), .B2(n19546), .ZN(
        n17167) );
  INV_X1 U20358 ( .A(n17167), .ZN(n17168) );
  NAND2_X1 U20359 ( .A1(n17169), .A2(n17168), .ZN(n19555) );
  INV_X1 U20360 ( .A(n17170), .ZN(n17171) );
  NAND2_X1 U20361 ( .A1(n17172), .A2(n17171), .ZN(n17173) );
  OAI211_X1 U20362 ( .C1(n17899), .C2(n17175), .A(n17174), .B(n17173), .ZN(
        n17176) );
  AOI21_X1 U20363 ( .B1(n19555), .B2(n17540), .A(n17176), .ZN(n17177) );
  AOI21_X1 U20364 ( .B1(n17178), .B2(n9940), .A(n17177), .ZN(P3_U3288) );
  INV_X1 U20365 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17935) );
  INV_X1 U20366 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n18123) );
  INV_X1 U20367 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18157) );
  INV_X1 U20368 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17898) );
  INV_X1 U20369 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18282) );
  NOR2_X1 U20370 ( .A1(n18288), .A2(n18282), .ZN(n18278) );
  INV_X1 U20371 ( .A(n18278), .ZN(n17920) );
  NOR2_X1 U20372 ( .A1(n17898), .A2(n17920), .ZN(n18268) );
  NAND2_X1 U20373 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18173), .ZN(n18153) );
  INV_X1 U20374 ( .A(n17989), .ZN(n17992) );
  NAND2_X1 U20375 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17992), .ZN(n17277) );
  INV_X1 U20376 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17937) );
  AOI22_X1 U20377 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18089), .B1(
        n18192), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17181) );
  OAI21_X1 U20378 ( .B1(n17954), .B2(n17182), .A(n17181), .ZN(n17183) );
  AOI21_X1 U20379 ( .B1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n11603), .A(
        n17183), .ZN(n17186) );
  AOI22_X1 U20380 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20381 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17184) );
  NAND3_X1 U20382 ( .A1(n17186), .A2(n17185), .A3(n17184), .ZN(n17192) );
  AOI22_X1 U20383 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U20384 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20385 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20386 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17187) );
  NAND4_X1 U20387 ( .A1(n17190), .A2(n17189), .A3(n17188), .A4(n17187), .ZN(
        n17191) );
  NOR2_X1 U20388 ( .A1(n17192), .A2(n17191), .ZN(n17990) );
  INV_X1 U20389 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U20390 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17194) );
  NAND2_X1 U20391 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n17193) );
  OAI211_X1 U20392 ( .C1(n17195), .C2(n18216), .A(n17194), .B(n17193), .ZN(
        n17196) );
  INV_X1 U20393 ( .A(n17196), .ZN(n17199) );
  AOI22_X1 U20394 ( .A1(n18235), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U20395 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17197) );
  NAND3_X1 U20396 ( .A1(n17199), .A2(n17198), .A3(n17197), .ZN(n17205) );
  AOI22_X1 U20397 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20398 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20399 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U20400 ( .A1(n11604), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17200) );
  NAND4_X1 U20401 ( .A1(n17203), .A2(n17202), .A3(n17201), .A4(n17200), .ZN(
        n17204) );
  NOR2_X1 U20402 ( .A1(n17205), .A2(n17204), .ZN(n17998) );
  INV_X1 U20403 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18108) );
  INV_X1 U20404 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17206) );
  INV_X1 U20405 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18106) );
  INV_X1 U20406 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17209) );
  OAI22_X1 U20407 ( .A1(n11598), .A2(n18106), .B1(n11548), .B2(n17209), .ZN(
        n17210) );
  AOI211_X1 U20408 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17211), .B(n17210), .ZN(n17213) );
  AOI22_X1 U20409 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17212) );
  OAI211_X1 U20410 ( .C1(n18216), .C2(n18108), .A(n17213), .B(n17212), .ZN(
        n17219) );
  AOI22_X1 U20411 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20412 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20413 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U20414 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17214) );
  NAND4_X1 U20415 ( .A1(n17217), .A2(n17216), .A3(n17215), .A4(n17214), .ZN(
        n17218) );
  OR2_X1 U20416 ( .A1(n17219), .A2(n17218), .ZN(n18002) );
  INV_X1 U20417 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17221) );
  INV_X1 U20418 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17220) );
  INV_X1 U20419 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18130) );
  OAI22_X1 U20420 ( .A1(n11598), .A2(n18130), .B1(n11548), .B2(n17961), .ZN(
        n17222) );
  AOI211_X1 U20421 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n17223), .B(n17222), .ZN(n17225) );
  AOI22_X1 U20422 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17224) );
  OAI211_X1 U20423 ( .C1(n18216), .C2(n17226), .A(n17225), .B(n17224), .ZN(
        n17232) );
  AOI22_X1 U20424 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20425 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20426 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20427 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17227) );
  NAND4_X1 U20428 ( .A1(n17230), .A2(n17229), .A3(n17228), .A4(n17227), .ZN(
        n17231) );
  OR2_X1 U20429 ( .A1(n17232), .A2(n17231), .ZN(n18003) );
  NAND2_X1 U20430 ( .A1(n18002), .A2(n18003), .ZN(n18001) );
  NOR2_X1 U20431 ( .A1(n17998), .A2(n18001), .ZN(n17995) );
  INV_X1 U20432 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17239) );
  INV_X1 U20433 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18201) );
  INV_X1 U20434 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18076) );
  INV_X1 U20435 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17234) );
  OAI22_X1 U20436 ( .A1(n11598), .A2(n18076), .B1(n11548), .B2(n17234), .ZN(
        n17235) );
  AOI211_X1 U20437 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17236), .B(n17235), .ZN(n17238) );
  AOI22_X1 U20438 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17237) );
  OAI211_X1 U20439 ( .C1(n18251), .C2(n17239), .A(n17238), .B(n17237), .ZN(
        n17245) );
  AOI22_X1 U20440 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17243) );
  AOI22_X1 U20441 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20442 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20443 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17240) );
  NAND4_X1 U20444 ( .A1(n17243), .A2(n17242), .A3(n17241), .A4(n17240), .ZN(
        n17244) );
  OR2_X1 U20445 ( .A1(n17245), .A2(n17244), .ZN(n17994) );
  NAND2_X1 U20446 ( .A1(n17995), .A2(n17994), .ZN(n17993) );
  NOR2_X1 U20447 ( .A1(n17990), .A2(n17993), .ZN(n17987) );
  INV_X1 U20448 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17255) );
  INV_X1 U20449 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17247) );
  INV_X1 U20450 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17246) );
  INV_X1 U20451 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17249) );
  INV_X1 U20452 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17248) );
  OAI22_X1 U20453 ( .A1(n11598), .A2(n17249), .B1(n11548), .B2(n17248), .ZN(
        n17250) );
  AOI211_X1 U20454 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17251), .B(n17250), .ZN(n17254) );
  AOI22_X1 U20455 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17253) );
  OAI211_X1 U20456 ( .C1(n18251), .C2(n17255), .A(n17254), .B(n17253), .ZN(
        n17261) );
  AOI22_X1 U20457 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U20458 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20459 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U20460 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17256) );
  NAND4_X1 U20461 ( .A1(n17259), .A2(n17258), .A3(n17257), .A4(n17256), .ZN(
        n17260) );
  OR2_X1 U20462 ( .A1(n17261), .A2(n17260), .ZN(n17986) );
  NAND2_X1 U20463 ( .A1(n17987), .A2(n17986), .ZN(n17985) );
  INV_X1 U20464 ( .A(n17985), .ZN(n17978) );
  INV_X1 U20465 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18023) );
  INV_X1 U20466 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17262) );
  INV_X1 U20467 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18021) );
  INV_X1 U20468 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17264) );
  OAI22_X1 U20469 ( .A1(n11598), .A2(n18021), .B1(n11548), .B2(n17264), .ZN(
        n17265) );
  AOI211_X1 U20470 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n17266), .B(n17265), .ZN(n17268) );
  INV_X1 U20471 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21462) );
  AOI22_X1 U20472 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17267) );
  OAI211_X1 U20473 ( .C1(n18251), .C2(n18023), .A(n17268), .B(n17267), .ZN(
        n17275) );
  AOI22_X1 U20474 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U20475 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17272) );
  AOI22_X1 U20476 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20477 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17270) );
  NAND4_X1 U20478 ( .A1(n17273), .A2(n17272), .A3(n17271), .A4(n17270), .ZN(
        n17274) );
  OR2_X1 U20479 ( .A1(n17275), .A2(n17274), .ZN(n17979) );
  XOR2_X1 U20480 ( .A(n17978), .B(n17979), .Z(n18307) );
  AOI22_X1 U20481 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17983), .B1(n18286), 
        .B2(n18307), .ZN(n17276) );
  OAI21_X1 U20482 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17277), .A(n17276), .ZN(
        P3_U2675) );
  INV_X1 U20483 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18022) );
  AOI22_X1 U20484 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17278), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17279) );
  OAI21_X1 U20485 ( .B1(n17954), .B2(n18022), .A(n17279), .ZN(n17280) );
  AOI21_X1 U20486 ( .B1(n11603), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n17280), .ZN(n17284) );
  AOI22_X1 U20487 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20488 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17282) );
  NAND3_X1 U20489 ( .A1(n17284), .A2(n17283), .A3(n17282), .ZN(n17290) );
  AOI22_X1 U20490 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U20491 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20492 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20493 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17285) );
  NAND4_X1 U20494 ( .A1(n17288), .A2(n17287), .A3(n17286), .A4(n17285), .ZN(
        n17289) );
  NOR2_X1 U20495 ( .A1(n17290), .A2(n17289), .ZN(n18388) );
  OAI211_X1 U20496 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n18173), .A(n18153), .B(
        n18270), .ZN(n17291) );
  OAI21_X1 U20497 ( .B1(n18388), .B2(n18270), .A(n17291), .ZN(P3_U2690) );
  NAND2_X1 U20498 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19251) );
  AOI221_X1 U20499 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19251), .C1(n17293), 
        .C2(n19251), .A(n17292), .ZN(n19102) );
  NOR2_X1 U20500 ( .A1(n17294), .A2(n11652), .ZN(n17295) );
  OAI21_X1 U20501 ( .B1(n17295), .B2(n19450), .A(n19103), .ZN(n19100) );
  AOI22_X1 U20502 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19102), .B1(
        n19100), .B2(n19568), .ZN(P3_U2865) );
  NAND2_X1 U20503 ( .A1(n17302), .A2(n17299), .ZN(n17300) );
  OAI21_X1 U20504 ( .B1(n17302), .B2(n17301), .A(n17300), .ZN(P2_U3595) );
  OAI22_X1 U20505 ( .A1(n17304), .A2(n19776), .B1(n19833), .B2(n17303), .ZN(
        n17305) );
  INV_X1 U20506 ( .A(n17305), .ZN(n17319) );
  INV_X1 U20507 ( .A(n17306), .ZN(n17317) );
  INV_X1 U20508 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20509 ( .A1(n19830), .A2(P2_EBX_REG_22__SCAN_IN), .B1(n19827), 
        .B2(P2_REIP_REG_22__SCAN_IN), .ZN(n17307) );
  OAI21_X1 U20510 ( .B1(n19803), .B2(n17308), .A(n17307), .ZN(n17316) );
  INV_X1 U20511 ( .A(n17309), .ZN(n17312) );
  INV_X1 U20512 ( .A(n17310), .ZN(n17311) );
  OAI21_X1 U20513 ( .B1(n17312), .B2(n17311), .A(n19820), .ZN(n17313) );
  AOI21_X1 U20514 ( .B1(n17314), .B2(n17313), .A(n15734), .ZN(n17315) );
  AOI211_X1 U20515 ( .C1(n19829), .C2(n17317), .A(n17316), .B(n17315), .ZN(
        n17318) );
  NAND2_X1 U20516 ( .A1(n17319), .A2(n17318), .ZN(P2_U2833) );
  INV_X1 U20517 ( .A(n17320), .ZN(n17331) );
  INV_X1 U20518 ( .A(n17321), .ZN(n17322) );
  OAI211_X1 U20519 ( .C1(n12593), .C2(n17323), .A(n17322), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17329) );
  INV_X1 U20520 ( .A(n17329), .ZN(n17327) );
  INV_X1 U20521 ( .A(n17324), .ZN(n17326) );
  OAI22_X1 U20522 ( .A1(n17327), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n17326), .B2(n17325), .ZN(n17328) );
  OAI21_X1 U20523 ( .B1(n17329), .B2(n21432), .A(n17328), .ZN(n17330) );
  AOI222_X1 U20524 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17331), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17330), .C1(n17331), 
        .C2(n17330), .ZN(n17332) );
  OR2_X1 U20525 ( .A1(n17332), .A2(n21132), .ZN(n17333) );
  AOI22_X1 U20526 ( .A1(n17334), .A2(n17333), .B1(n17332), .B2(n21132), .ZN(
        n17341) );
  OR2_X1 U20527 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n17338) );
  INV_X1 U20528 ( .A(n17335), .ZN(n17337) );
  AOI211_X1 U20529 ( .C1(n17339), .C2(n17338), .A(n17337), .B(n17336), .ZN(
        n17340) );
  OAI21_X1 U20530 ( .B1(n17341), .B2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n17340), .ZN(n17342) );
  NOR3_X1 U20531 ( .A1(n17344), .A2(n17343), .A3(n17342), .ZN(n17356) );
  INV_X1 U20532 ( .A(n17356), .ZN(n17350) );
  NAND4_X1 U20533 ( .A1(n12451), .A2(n20828), .A3(n17346), .A4(n17345), .ZN(
        n17349) );
  OAI21_X1 U20534 ( .B1(n17347), .B2(n21404), .A(n17355), .ZN(n17348) );
  NAND2_X1 U20535 ( .A1(n17349), .A2(n17348), .ZN(n17435) );
  AOI21_X1 U20536 ( .B1(n17352), .B2(n12586), .A(n17351), .ZN(n17354) );
  OAI211_X1 U20537 ( .C1(n17356), .C2(n17355), .A(n17354), .B(n17353), .ZN(
        n17357) );
  NOR2_X1 U20538 ( .A1(n17439), .A2(n17357), .ZN(n17362) );
  NAND2_X1 U20539 ( .A1(n17359), .A2(n17358), .ZN(n17360) );
  NAND2_X1 U20540 ( .A1(n10287), .A2(n17360), .ZN(n17361) );
  OAI22_X1 U20541 ( .A1(n17362), .A2(n10287), .B1(n17439), .B2(n17361), .ZN(
        P1_U3161) );
  INV_X1 U20542 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17534) );
  NOR2_X1 U20543 ( .A1(n20772), .A2(n17534), .ZN(P1_U2905) );
  NOR2_X1 U20544 ( .A1(n17363), .A2(n20626), .ZN(P2_U3047) );
  AOI22_X1 U20545 ( .A1(n17370), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n17416), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17369) );
  XNOR2_X1 U20546 ( .A(n17364), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17365) );
  XNOR2_X1 U20547 ( .A(n17366), .B(n17365), .ZN(n17412) );
  INV_X1 U20548 ( .A(n17367), .ZN(n20686) );
  AOI22_X1 U20549 ( .A1(n17412), .A2(n17382), .B1(n20686), .B2(n17381), .ZN(
        n17368) );
  OAI211_X1 U20550 ( .C1(n17377), .C2(n20680), .A(n17369), .B(n17368), .ZN(
        P1_U2992) );
  AOI22_X1 U20551 ( .A1(n17370), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n17416), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17376) );
  NAND2_X1 U20552 ( .A1(n17372), .A2(n17371), .ZN(n17373) );
  XNOR2_X1 U20553 ( .A(n17374), .B(n17373), .ZN(n17417) );
  AOI22_X1 U20554 ( .A1(n20697), .A2(n17381), .B1(n17417), .B2(n17382), .ZN(
        n17375) );
  OAI211_X1 U20555 ( .C1(n17377), .C2(n20691), .A(n17376), .B(n17375), .ZN(
        P1_U2993) );
  INV_X1 U20556 ( .A(n20712), .ZN(n17380) );
  AOI222_X1 U20557 ( .A1(n17430), .A2(n17382), .B1(n17381), .B2(n20709), .C1(
        n17380), .C2(n17379), .ZN(n17384) );
  NOR2_X1 U20558 ( .A1(n20716), .A2(n20692), .ZN(n17423) );
  INV_X1 U20559 ( .A(n17423), .ZN(n17383) );
  OAI211_X1 U20560 ( .C1(n20701), .C2(n17385), .A(n17384), .B(n17383), .ZN(
        P1_U2994) );
  NOR2_X1 U20561 ( .A1(n17387), .A2(n17386), .ZN(n17395) );
  INV_X1 U20562 ( .A(n17388), .ZN(n17389) );
  OAI21_X1 U20563 ( .B1(n17391), .B2(n17390), .A(n17389), .ZN(n17392) );
  AOI221_X1 U20564 ( .B1(n17395), .B2(n17394), .C1(n17393), .C2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n17392), .ZN(n17396) );
  OAI21_X1 U20565 ( .B1(n17398), .B2(n17397), .A(n17396), .ZN(P1_U3017) );
  OR2_X1 U20566 ( .A1(n17400), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17426) );
  AOI221_X1 U20567 ( .B1(n17402), .B2(n17401), .C1(n17400), .C2(n17401), .A(
        n17399), .ZN(n17432) );
  OAI21_X1 U20568 ( .B1(n17403), .B2(n17426), .A(n17432), .ZN(n17418) );
  AOI21_X1 U20569 ( .B1(n17408), .B2(n17404), .A(n17418), .ZN(n17415) );
  INV_X1 U20570 ( .A(n17405), .ZN(n17406) );
  AOI222_X1 U20571 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n17416), .B1(n17424), 
        .B2(n17407), .C1(n17429), .C2(n17406), .ZN(n17410) );
  NOR2_X1 U20572 ( .A1(n17421), .A2(n17408), .ZN(n17411) );
  OAI221_X1 U20573 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n12130), .C2(n15294), .A(
        n17411), .ZN(n17409) );
  OAI211_X1 U20574 ( .C1(n17415), .C2(n12130), .A(n17410), .B(n17409), .ZN(
        P1_U3023) );
  AOI22_X1 U20575 ( .A1(n20678), .A2(n17424), .B1(n17416), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U20576 ( .A1(n17412), .A2(n17429), .B1(n15294), .B2(n17411), .ZN(
        n17413) );
  OAI211_X1 U20577 ( .C1(n17415), .C2(n15294), .A(n17414), .B(n17413), .ZN(
        P1_U3024) );
  AOI22_X1 U20578 ( .A1(n17424), .A2(n20689), .B1(n17416), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20579 ( .A1(n17418), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n17429), .B2(n17417), .ZN(n17419) );
  OAI211_X1 U20580 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n17421), .A(
        n17420), .B(n17419), .ZN(P1_U3025) );
  INV_X1 U20581 ( .A(n17422), .ZN(n17427) );
  AOI21_X1 U20582 ( .B1(n20707), .B2(n17424), .A(n17423), .ZN(n17425) );
  OAI21_X1 U20583 ( .B1(n17427), .B2(n17426), .A(n17425), .ZN(n17428) );
  AOI21_X1 U20584 ( .B1(n17430), .B2(n17429), .A(n17428), .ZN(n17431) );
  OAI21_X1 U20585 ( .B1(n17432), .B2(n21471), .A(n17431), .ZN(P1_U3026) );
  NAND4_X1 U20586 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n12586), .A4(n21404), .ZN(n17433) );
  NAND2_X1 U20587 ( .A1(n17434), .A2(n17433), .ZN(n21358) );
  OAI21_X1 U20588 ( .B1(n17436), .B2(n21358), .A(n17435), .ZN(n17437) );
  OAI221_X1 U20589 ( .B1(n21399), .B2(n21197), .C1(n21399), .C2(n21404), .A(
        n17437), .ZN(n17438) );
  AOI221_X1 U20590 ( .B1(n17439), .B2(n21357), .C1(n10287), .C2(n21357), .A(
        n17438), .ZN(P1_U3162) );
  NOR2_X1 U20591 ( .A1(n17439), .A2(n10287), .ZN(n17441) );
  OAI21_X1 U20592 ( .B1(n17441), .B2(n21197), .A(n17440), .ZN(P1_U3466) );
  INV_X1 U20593 ( .A(n17442), .ZN(n17443) );
  AOI22_X1 U20594 ( .A1(n17444), .A2(n17443), .B1(n19960), .B2(n19826), .ZN(
        n17452) );
  OAI22_X1 U20595 ( .A1(n17446), .A2(n19941), .B1(n19964), .B2(n17445), .ZN(
        n17450) );
  OAI21_X1 U20596 ( .B1(n19963), .B2(n17448), .A(n17447), .ZN(n17449) );
  NOR2_X1 U20597 ( .A1(n17450), .A2(n17449), .ZN(n17451) );
  OAI211_X1 U20598 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19970), .A(
        n17452), .B(n17451), .ZN(P2_U3046) );
  NOR3_X1 U20599 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17454) );
  NOR4_X1 U20600 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17453) );
  NAND4_X1 U20601 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17454), .A3(n17453), .A4(
        U215), .ZN(U213) );
  INV_X1 U20602 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19909) );
  OAI222_X1 U20603 ( .A1(U212), .A2(n19909), .B1(n17503), .B2(n17456), .C1(
        U214), .C2(n17534), .ZN(U216) );
  INV_X1 U20604 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20012) );
  AOI22_X1 U20605 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n17501), .ZN(n17457) );
  OAI21_X1 U20606 ( .B1(n20012), .B2(n17503), .A(n17457), .ZN(U217) );
  AOI22_X1 U20607 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17501), .ZN(n17458) );
  OAI21_X1 U20608 ( .B1(n16076), .B2(n17503), .A(n17458), .ZN(U218) );
  AOI22_X1 U20609 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17501), .ZN(n17459) );
  OAI21_X1 U20610 ( .B1(n17460), .B2(n17503), .A(n17459), .ZN(U219) );
  INV_X1 U20611 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U20612 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17501), .ZN(n17461) );
  OAI21_X1 U20613 ( .B1(n17462), .B2(n17503), .A(n17461), .ZN(U220) );
  AOI22_X1 U20614 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17501), .ZN(n17463) );
  OAI21_X1 U20615 ( .B1(n16097), .B2(n17503), .A(n17463), .ZN(U221) );
  AOI22_X1 U20616 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17501), .ZN(n17464) );
  OAI21_X1 U20617 ( .B1(n15131), .B2(n17503), .A(n17464), .ZN(U222) );
  INV_X1 U20618 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U20619 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17501), .ZN(n17465) );
  OAI21_X1 U20620 ( .B1(n17466), .B2(n17503), .A(n17465), .ZN(U223) );
  INV_X1 U20621 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20622 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17501), .ZN(n17467) );
  OAI21_X1 U20623 ( .B1(n17468), .B2(n17503), .A(n17467), .ZN(U224) );
  AOI222_X1 U20624 ( .A1(n17498), .A2(P1_DATAO_REG_22__SCAN_IN), .B1(n17499), 
        .B2(BUF1_REG_22__SCAN_IN), .C1(n17501), .C2(P2_DATAO_REG_22__SCAN_IN), 
        .ZN(n17469) );
  INV_X1 U20625 ( .A(n17469), .ZN(U225) );
  INV_X1 U20626 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17471) );
  AOI22_X1 U20627 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17501), .ZN(n17470) );
  OAI21_X1 U20628 ( .B1(n17471), .B2(n17503), .A(n17470), .ZN(U226) );
  AOI22_X1 U20629 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17501), .ZN(n17472) );
  OAI21_X1 U20630 ( .B1(n17473), .B2(n17503), .A(n17472), .ZN(U227) );
  AOI22_X1 U20631 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17501), .ZN(n17474) );
  OAI21_X1 U20632 ( .B1(n16147), .B2(n17503), .A(n17474), .ZN(U228) );
  AOI22_X1 U20633 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17501), .ZN(n17475) );
  OAI21_X1 U20634 ( .B1(n16153), .B2(n17503), .A(n17475), .ZN(U229) );
  INV_X1 U20635 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U20636 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17501), .ZN(n17476) );
  OAI21_X1 U20637 ( .B1(n17477), .B2(n17503), .A(n17476), .ZN(U230) );
  INV_X1 U20638 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17479) );
  AOI22_X1 U20639 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17501), .ZN(n17478) );
  OAI21_X1 U20640 ( .B1(n17479), .B2(n17503), .A(n17478), .ZN(U231) );
  INV_X1 U20641 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n21494) );
  AOI22_X1 U20642 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n17498), .ZN(n17480) );
  OAI21_X1 U20643 ( .B1(n21494), .B2(U212), .A(n17480), .ZN(U232) );
  INV_X1 U20644 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U20645 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n17498), .ZN(n17481) );
  OAI21_X1 U20646 ( .B1(n17482), .B2(U212), .A(n17481), .ZN(U233) );
  INV_X1 U20647 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n17515) );
  AOI22_X1 U20648 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n17498), .ZN(n17483) );
  OAI21_X1 U20649 ( .B1(n17515), .B2(U212), .A(n17483), .ZN(U234) );
  INV_X1 U20650 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n21465) );
  AOI22_X1 U20651 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n17498), .ZN(n17484) );
  OAI21_X1 U20652 ( .B1(n21465), .B2(U212), .A(n17484), .ZN(U235) );
  INV_X1 U20653 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n21483) );
  AOI22_X1 U20654 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17498), .ZN(n17485) );
  OAI21_X1 U20655 ( .B1(n21483), .B2(U212), .A(n17485), .ZN(U236) );
  INV_X1 U20656 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17487) );
  AOI22_X1 U20657 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17501), .ZN(n17486) );
  OAI21_X1 U20658 ( .B1(n17487), .B2(n17503), .A(n17486), .ZN(U237) );
  INV_X1 U20659 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U20660 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n17498), .ZN(n17488) );
  OAI21_X1 U20661 ( .B1(n17513), .B2(U212), .A(n17488), .ZN(U238) );
  INV_X1 U20662 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n21466) );
  AOI22_X1 U20663 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n17499), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17501), .ZN(n17489) );
  OAI21_X1 U20664 ( .B1(n21466), .B2(U214), .A(n17489), .ZN(U239) );
  INV_X1 U20665 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17511) );
  AOI22_X1 U20666 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17498), .ZN(n17490) );
  OAI21_X1 U20667 ( .B1(n17511), .B2(U212), .A(n17490), .ZN(U240) );
  INV_X1 U20668 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U20669 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17501), .ZN(n17491) );
  OAI21_X1 U20670 ( .B1(n17492), .B2(n17503), .A(n17491), .ZN(U241) );
  INV_X1 U20671 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n20771) );
  INV_X1 U20672 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n17493) );
  INV_X1 U20673 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n21477) );
  OAI222_X1 U20674 ( .A1(U214), .A2(n20771), .B1(n17503), .B2(n17493), .C1(
        U212), .C2(n21477), .ZN(U242) );
  INV_X1 U20675 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17495) );
  AOI22_X1 U20676 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17501), .ZN(n17494) );
  OAI21_X1 U20677 ( .B1(n17495), .B2(n17503), .A(n17494), .ZN(U243) );
  INV_X1 U20678 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17508) );
  AOI22_X1 U20679 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17498), .ZN(n17496) );
  OAI21_X1 U20680 ( .B1(n17508), .B2(U212), .A(n17496), .ZN(U244) );
  INV_X1 U20681 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U20682 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n17498), .ZN(n17497) );
  OAI21_X1 U20683 ( .B1(n17507), .B2(U212), .A(n17497), .ZN(U245) );
  INV_X1 U20684 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n17506) );
  AOI22_X1 U20685 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17499), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17498), .ZN(n17500) );
  OAI21_X1 U20686 ( .B1(n17506), .B2(U212), .A(n17500), .ZN(U246) );
  INV_X1 U20687 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n17504) );
  AOI22_X1 U20688 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n17498), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n17501), .ZN(n17502) );
  OAI21_X1 U20689 ( .B1(n17504), .B2(n17503), .A(n17502), .ZN(U247) );
  OAI22_X1 U20690 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n17532), .ZN(n17505) );
  INV_X1 U20691 ( .A(n17505), .ZN(U251) );
  INV_X1 U20692 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n19112) );
  AOI22_X1 U20693 ( .A1(n17532), .A2(n17506), .B1(n19112), .B2(U215), .ZN(U252) );
  AOI22_X1 U20694 ( .A1(n17532), .A2(n17507), .B1(n19116), .B2(U215), .ZN(U253) );
  INV_X1 U20695 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19121) );
  AOI22_X1 U20696 ( .A1(n17532), .A2(n17508), .B1(n19121), .B2(U215), .ZN(U254) );
  OAI22_X1 U20697 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17532), .ZN(n17509) );
  INV_X1 U20698 ( .A(n17509), .ZN(U255) );
  INV_X1 U20699 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19130) );
  AOI22_X1 U20700 ( .A1(n17532), .A2(n21477), .B1(n19130), .B2(U215), .ZN(U256) );
  OAI22_X1 U20701 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n17532), .ZN(n17510) );
  INV_X1 U20702 ( .A(n17510), .ZN(U257) );
  AOI22_X1 U20703 ( .A1(n17532), .A2(n17511), .B1(n14047), .B2(U215), .ZN(U258) );
  OAI22_X1 U20704 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17532), .ZN(n17512) );
  INV_X1 U20705 ( .A(n17512), .ZN(U259) );
  AOI22_X1 U20706 ( .A1(n17532), .A2(n17513), .B1(n14028), .B2(U215), .ZN(U260) );
  OAI22_X1 U20707 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17532), .ZN(n17514) );
  INV_X1 U20708 ( .A(n17514), .ZN(U261) );
  AOI22_X1 U20709 ( .A1(n17532), .A2(n21483), .B1(n14034), .B2(U215), .ZN(U262) );
  AOI22_X1 U20710 ( .A1(n17532), .A2(n21465), .B1(n14024), .B2(U215), .ZN(U263) );
  AOI22_X1 U20711 ( .A1(n17532), .A2(n17515), .B1(n14014), .B2(U215), .ZN(U264) );
  OAI22_X1 U20712 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17532), .ZN(n17516) );
  INV_X1 U20713 ( .A(n17516), .ZN(U265) );
  OAI22_X1 U20714 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17532), .ZN(n17517) );
  INV_X1 U20715 ( .A(n17517), .ZN(U266) );
  OAI22_X1 U20716 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17532), .ZN(n17518) );
  INV_X1 U20717 ( .A(n17518), .ZN(U267) );
  OAI22_X1 U20718 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17532), .ZN(n17519) );
  INV_X1 U20719 ( .A(n17519), .ZN(U268) );
  OAI22_X1 U20720 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17532), .ZN(n17520) );
  INV_X1 U20721 ( .A(n17520), .ZN(U269) );
  OAI22_X1 U20722 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17532), .ZN(n17521) );
  INV_X1 U20723 ( .A(n17521), .ZN(U270) );
  OAI22_X1 U20724 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17532), .ZN(n17522) );
  INV_X1 U20725 ( .A(n17522), .ZN(U271) );
  OAI22_X1 U20726 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17532), .ZN(n17523) );
  INV_X1 U20727 ( .A(n17523), .ZN(U272) );
  INV_X1 U20728 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n21524) );
  AOI22_X1 U20729 ( .A1(n17532), .A2(n21524), .B1(n19134), .B2(U215), .ZN(U273) );
  OAI22_X1 U20730 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17532), .ZN(n17524) );
  INV_X1 U20731 ( .A(n17524), .ZN(U274) );
  OAI22_X1 U20732 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17532), .ZN(n17525) );
  INV_X1 U20733 ( .A(n17525), .ZN(U275) );
  OAI22_X1 U20734 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17532), .ZN(n17526) );
  INV_X1 U20735 ( .A(n17526), .ZN(U276) );
  OAI22_X1 U20736 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17532), .ZN(n17527) );
  INV_X1 U20737 ( .A(n17527), .ZN(U277) );
  OAI22_X1 U20738 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17532), .ZN(n17528) );
  INV_X1 U20739 ( .A(n17528), .ZN(U278) );
  OAI22_X1 U20740 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17532), .ZN(n17529) );
  INV_X1 U20741 ( .A(n17529), .ZN(U279) );
  OAI22_X1 U20742 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17532), .ZN(n17530) );
  INV_X1 U20743 ( .A(n17530), .ZN(U280) );
  OAI22_X1 U20744 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17532), .ZN(n17531) );
  INV_X1 U20745 ( .A(n17531), .ZN(U281) );
  INV_X1 U20746 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18298) );
  AOI22_X1 U20747 ( .A1(n17532), .A2(n19909), .B1(n18298), .B2(U215), .ZN(U282) );
  INV_X1 U20748 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17533) );
  AOI222_X1 U20749 ( .A1(n17534), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19909), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17533), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17535) );
  INV_X2 U20750 ( .A(n17537), .ZN(n17536) );
  INV_X1 U20751 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19637) );
  INV_X1 U20752 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20559) );
  AOI22_X1 U20753 ( .A1(n17536), .A2(n19637), .B1(n20559), .B2(n17537), .ZN(
        U347) );
  INV_X1 U20754 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19635) );
  INV_X1 U20755 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20557) );
  AOI22_X1 U20756 ( .A1(n17536), .A2(n19635), .B1(n20557), .B2(n17537), .ZN(
        U348) );
  INV_X1 U20757 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19632) );
  INV_X1 U20758 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20555) );
  AOI22_X1 U20759 ( .A1(n17536), .A2(n19632), .B1(n20555), .B2(n17537), .ZN(
        U349) );
  INV_X1 U20760 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19631) );
  INV_X1 U20761 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20553) );
  AOI22_X1 U20762 ( .A1(n17536), .A2(n19631), .B1(n20553), .B2(n17537), .ZN(
        U350) );
  INV_X1 U20763 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19629) );
  INV_X1 U20764 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20551) );
  AOI22_X1 U20765 ( .A1(n17536), .A2(n19629), .B1(n20551), .B2(n17537), .ZN(
        U351) );
  INV_X1 U20766 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19627) );
  INV_X1 U20767 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20549) );
  AOI22_X1 U20768 ( .A1(n17536), .A2(n19627), .B1(n20549), .B2(n17537), .ZN(
        U352) );
  INV_X1 U20769 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19625) );
  INV_X1 U20770 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20547) );
  AOI22_X1 U20771 ( .A1(n17536), .A2(n19625), .B1(n20547), .B2(n17537), .ZN(
        U353) );
  INV_X1 U20772 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19623) );
  AOI22_X1 U20773 ( .A1(n17536), .A2(n19623), .B1(n20544), .B2(n17537), .ZN(
        U354) );
  INV_X1 U20774 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19676) );
  INV_X1 U20775 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20598) );
  AOI22_X1 U20776 ( .A1(n17536), .A2(n19676), .B1(n20598), .B2(n17537), .ZN(
        U355) );
  INV_X1 U20777 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19673) );
  INV_X1 U20778 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20595) );
  AOI22_X1 U20779 ( .A1(n17536), .A2(n19673), .B1(n20595), .B2(n17537), .ZN(
        U356) );
  INV_X1 U20780 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19672) );
  INV_X1 U20781 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20593) );
  AOI22_X1 U20782 ( .A1(n17536), .A2(n19672), .B1(n20593), .B2(n17537), .ZN(
        U357) );
  INV_X1 U20783 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19671) );
  INV_X1 U20784 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20590) );
  AOI22_X1 U20785 ( .A1(n17536), .A2(n19671), .B1(n20590), .B2(n17537), .ZN(
        U358) );
  INV_X1 U20786 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19669) );
  INV_X1 U20787 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20589) );
  AOI22_X1 U20788 ( .A1(n17536), .A2(n19669), .B1(n20589), .B2(n17537), .ZN(
        U359) );
  INV_X1 U20789 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19667) );
  INV_X1 U20790 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20587) );
  AOI22_X1 U20791 ( .A1(n17536), .A2(n19667), .B1(n20587), .B2(n17537), .ZN(
        U360) );
  INV_X1 U20792 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19665) );
  INV_X1 U20793 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20585) );
  AOI22_X1 U20794 ( .A1(n17536), .A2(n19665), .B1(n20585), .B2(n17537), .ZN(
        U361) );
  INV_X1 U20795 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19662) );
  INV_X1 U20796 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20583) );
  AOI22_X1 U20797 ( .A1(n17536), .A2(n19662), .B1(n20583), .B2(n17537), .ZN(
        U362) );
  INV_X1 U20798 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19661) );
  INV_X1 U20799 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20581) );
  AOI22_X1 U20800 ( .A1(n17536), .A2(n19661), .B1(n20581), .B2(n17537), .ZN(
        U363) );
  INV_X1 U20801 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19659) );
  INV_X1 U20802 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20580) );
  AOI22_X1 U20803 ( .A1(n17536), .A2(n19659), .B1(n20580), .B2(n17537), .ZN(
        U364) );
  INV_X1 U20804 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19621) );
  INV_X1 U20805 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20543) );
  AOI22_X1 U20806 ( .A1(n17536), .A2(n19621), .B1(n20543), .B2(n17537), .ZN(
        U365) );
  INV_X1 U20807 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19656) );
  INV_X1 U20808 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20578) );
  AOI22_X1 U20809 ( .A1(n17536), .A2(n19656), .B1(n20578), .B2(n17537), .ZN(
        U366) );
  INV_X1 U20810 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19655) );
  INV_X1 U20811 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20576) );
  AOI22_X1 U20812 ( .A1(n17536), .A2(n19655), .B1(n20576), .B2(n17537), .ZN(
        U367) );
  INV_X1 U20813 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19653) );
  INV_X1 U20814 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20574) );
  AOI22_X1 U20815 ( .A1(n17536), .A2(n19653), .B1(n20574), .B2(n17537), .ZN(
        U368) );
  INV_X1 U20816 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19651) );
  INV_X1 U20817 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n21463) );
  AOI22_X1 U20818 ( .A1(n17536), .A2(n19651), .B1(n21463), .B2(n17537), .ZN(
        U369) );
  INV_X1 U20819 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19649) );
  INV_X1 U20820 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20571) );
  AOI22_X1 U20821 ( .A1(n17536), .A2(n19649), .B1(n20571), .B2(n17537), .ZN(
        U370) );
  INV_X1 U20822 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19647) );
  INV_X1 U20823 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20569) );
  AOI22_X1 U20824 ( .A1(n17535), .A2(n19647), .B1(n20569), .B2(n17537), .ZN(
        U371) );
  INV_X1 U20825 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19644) );
  INV_X1 U20826 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20567) );
  AOI22_X1 U20827 ( .A1(n17535), .A2(n19644), .B1(n20567), .B2(n17537), .ZN(
        U372) );
  INV_X1 U20828 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19643) );
  INV_X1 U20829 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20565) );
  AOI22_X1 U20830 ( .A1(n17535), .A2(n19643), .B1(n20565), .B2(n17537), .ZN(
        U373) );
  INV_X1 U20831 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19641) );
  INV_X1 U20832 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20563) );
  AOI22_X1 U20833 ( .A1(n17535), .A2(n19641), .B1(n20563), .B2(n17537), .ZN(
        U374) );
  INV_X1 U20834 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19639) );
  INV_X1 U20835 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20561) );
  AOI22_X1 U20836 ( .A1(n17536), .A2(n19639), .B1(n20561), .B2(n17537), .ZN(
        U375) );
  INV_X1 U20837 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19619) );
  INV_X1 U20838 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20541) );
  AOI22_X1 U20839 ( .A1(n17536), .A2(n19619), .B1(n20541), .B2(n17537), .ZN(
        U376) );
  NAND3_X1 U20840 ( .A1(n19618), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n17538) );
  NAND2_X1 U20841 ( .A1(n19615), .A2(n19607), .ZN(n19603) );
  NAND2_X1 U20842 ( .A1(n17538), .A2(n19603), .ZN(n19687) );
  AOI21_X1 U20843 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19687), .ZN(n17539) );
  INV_X1 U20844 ( .A(n17539), .ZN(P3_U2633) );
  AOI21_X1 U20845 ( .B1(n18493), .B2(n17546), .A(n18492), .ZN(n17542) );
  INV_X1 U20846 ( .A(P3_CODEFETCH_REG_SCAN_IN), .ZN(n21557) );
  NAND2_X1 U20847 ( .A1(n17540), .A2(n19582), .ZN(n17541) );
  OAI22_X1 U20848 ( .A1(n17542), .A2(n21557), .B1(n19591), .B2(n17541), .ZN(
        P3_U2634) );
  AOI21_X1 U20849 ( .B1(n19615), .B2(n19618), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17543) );
  AOI22_X1 U20850 ( .A1(n19682), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17543), 
        .B2(n19717), .ZN(P3_U2635) );
  OAI21_X1 U20851 ( .B1(n17544), .B2(BS16), .A(n19687), .ZN(n19685) );
  OAI21_X1 U20852 ( .B1(n19687), .B2(n21509), .A(n19685), .ZN(P3_U2636) );
  AOI211_X1 U20853 ( .C1(n18493), .C2(n17546), .A(n17545), .B(n19541), .ZN(
        n19548) );
  NOR2_X1 U20854 ( .A1(n19548), .A2(n19588), .ZN(n19700) );
  OAI21_X1 U20855 ( .B1(n19700), .B2(n19097), .A(n17547), .ZN(P3_U2637) );
  NOR4_X1 U20856 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n17551) );
  NOR4_X1 U20857 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17550) );
  NOR4_X1 U20858 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17549) );
  NOR4_X1 U20859 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17548) );
  NAND4_X1 U20860 ( .A1(n17551), .A2(n17550), .A3(n17549), .A4(n17548), .ZN(
        n17557) );
  NOR4_X1 U20861 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17555) );
  AOI211_X1 U20862 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_3__SCAN_IN), .B(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17554) );
  NOR4_X1 U20863 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n17553) );
  NOR4_X1 U20864 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n17552) );
  NAND4_X1 U20865 ( .A1(n17555), .A2(n17554), .A3(n17553), .A4(n17552), .ZN(
        n17556) );
  NOR2_X1 U20866 ( .A1(n17557), .A2(n17556), .ZN(n19694) );
  INV_X1 U20867 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17559) );
  NOR3_X1 U20868 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17560) );
  OAI21_X1 U20869 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17560), .A(n19694), .ZN(
        n17558) );
  OAI21_X1 U20870 ( .B1(n19694), .B2(n17559), .A(n17558), .ZN(P3_U2638) );
  INV_X1 U20871 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n21537) );
  INV_X1 U20872 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19686) );
  AOI21_X1 U20873 ( .B1(n21537), .B2(n19686), .A(n17560), .ZN(n17562) );
  INV_X1 U20874 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17561) );
  INV_X1 U20875 ( .A(n19694), .ZN(n19697) );
  AOI22_X1 U20876 ( .A1(n19694), .A2(n17562), .B1(n17561), .B2(n19697), .ZN(
        P3_U2639) );
  NOR3_X1 U20877 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19677), .A3(n17563), 
        .ZN(n17564) );
  AOI21_X1 U20878 ( .B1(n17916), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17564), .ZN(
        n17571) );
  INV_X1 U20879 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17944) );
  NAND2_X1 U20880 ( .A1(n17843), .A2(n19598), .ZN(n17919) );
  INV_X1 U20881 ( .A(n17567), .ZN(n17568) );
  INV_X1 U20882 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19675) );
  AOI21_X1 U20883 ( .B1(n17578), .B2(n17568), .A(n19675), .ZN(n17569) );
  NOR2_X1 U20884 ( .A1(n17586), .A2(n17982), .ZN(n17584) );
  INV_X1 U20885 ( .A(n17573), .ZN(n17574) );
  AOI211_X1 U20886 ( .C1(n17576), .C2(n17575), .A(n17574), .B(n17879), .ZN(
        n17580) );
  OAI22_X1 U20887 ( .A1(n17578), .A2(n17089), .B1(n17577), .B2(n17918), .ZN(
        n17579) );
  NAND3_X1 U20888 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n17585), .A3(n17089), 
        .ZN(n17581) );
  OAI211_X1 U20889 ( .C1(n17584), .C2(n17583), .A(n17582), .B(n17581), .ZN(
        P3_U2642) );
  INV_X1 U20890 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17595) );
  AOI22_X1 U20891 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17916), .B1(n17585), 
        .B2(n17109), .ZN(n17594) );
  INV_X1 U20892 ( .A(n17606), .ZN(n17599) );
  OAI21_X1 U20893 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n17605), .A(n17599), 
        .ZN(n17592) );
  AOI211_X1 U20894 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17602), .A(n17586), .B(
        n17928), .ZN(n17591) );
  AOI211_X1 U20895 ( .C1(n17589), .C2(n17588), .A(n17587), .B(n17879), .ZN(
        n17590) );
  AOI211_X1 U20896 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17592), .A(n17591), 
        .B(n17590), .ZN(n17593) );
  OAI211_X1 U20897 ( .C1(n17595), .C2(n17918), .A(n17594), .B(n17593), .ZN(
        P3_U2643) );
  INV_X1 U20898 ( .A(n17596), .ZN(n17597) );
  AOI211_X1 U20899 ( .C1(n18538), .C2(n17598), .A(n17597), .B(n17879), .ZN(
        n17601) );
  OAI22_X1 U20900 ( .A1(n18543), .A2(n17918), .B1(n19670), .B2(n17599), .ZN(
        n17600) );
  AOI211_X1 U20901 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n17916), .A(n17601), .B(
        n17600), .ZN(n17604) );
  OAI211_X1 U20902 ( .C1(n17608), .C2(n17936), .A(n17887), .B(n17602), .ZN(
        n17603) );
  OAI211_X1 U20903 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17605), .A(n17604), 
        .B(n17603), .ZN(P3_U2644) );
  AOI22_X1 U20904 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17910), .B1(
        n17916), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17615) );
  OAI21_X1 U20905 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n17607), .A(n17606), 
        .ZN(n17614) );
  AOI211_X1 U20906 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17622), .A(n17608), .B(
        n17928), .ZN(n17612) );
  AOI211_X1 U20907 ( .C1(n17610), .C2(n9724), .A(n17609), .B(n17879), .ZN(
        n17611) );
  NOR2_X1 U20908 ( .A1(n17612), .A2(n17611), .ZN(n17613) );
  NAND3_X1 U20909 ( .A1(n17615), .A2(n17614), .A3(n17613), .ZN(P3_U2645) );
  AOI22_X1 U20910 ( .A1(n17915), .A2(n19664), .B1(n17930), .B2(n17629), .ZN(
        n17626) );
  AOI211_X1 U20911 ( .C1(n17618), .C2(n17617), .A(n17616), .B(n17879), .ZN(
        n17621) );
  OAI22_X1 U20912 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17619), .B1(n17623), 
        .B2(n17929), .ZN(n17620) );
  AOI211_X1 U20913 ( .C1(n17910), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17621), .B(n17620), .ZN(n17625) );
  OAI211_X1 U20914 ( .C1(n17630), .C2(n17623), .A(n17887), .B(n17622), .ZN(
        n17624) );
  OAI211_X1 U20915 ( .C1(n17626), .C2(n19666), .A(n17625), .B(n17624), .ZN(
        P3_U2646) );
  NOR2_X1 U20916 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17906), .ZN(n17627) );
  AOI22_X1 U20917 ( .A1(n17916), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17628), 
        .B2(n17627), .ZN(n17636) );
  AND2_X1 U20918 ( .A1(n17930), .A2(n17629), .ZN(n17643) );
  AOI211_X1 U20919 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17644), .A(n17630), .B(
        n17928), .ZN(n17634) );
  INV_X1 U20920 ( .A(n17631), .ZN(n17632) );
  AOI211_X1 U20921 ( .C1(n17643), .C2(P3_REIP_REG_24__SCAN_IN), .A(n17634), 
        .B(n17633), .ZN(n17635) );
  OAI211_X1 U20922 ( .C1(n18568), .C2(n17918), .A(n17636), .B(n17635), .ZN(
        P3_U2647) );
  OAI21_X1 U20923 ( .B1(n17906), .B2(n17637), .A(n19663), .ZN(n17642) );
  AOI211_X1 U20924 ( .C1(n18579), .C2(n17639), .A(n17638), .B(n17879), .ZN(
        n17641) );
  OAI22_X1 U20925 ( .A1(n18583), .A2(n17918), .B1(n17929), .B2(n17645), .ZN(
        n17640) );
  AOI211_X1 U20926 ( .C1(n17643), .C2(n17642), .A(n17641), .B(n17640), .ZN(
        n17647) );
  OAI211_X1 U20927 ( .C1(n17653), .C2(n17645), .A(n17887), .B(n17644), .ZN(
        n17646) );
  NAND2_X1 U20928 ( .A1(n17647), .A2(n17646), .ZN(P3_U2648) );
  NOR2_X1 U20929 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17906), .ZN(n17648) );
  AOI22_X1 U20930 ( .A1(n17916), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n17649), 
        .B2(n17648), .ZN(n17661) );
  NOR2_X1 U20931 ( .A1(n17924), .A2(n17651), .ZN(n17750) );
  NOR2_X1 U20932 ( .A1(n17650), .A2(n17750), .ZN(n17752) );
  AOI21_X1 U20933 ( .B1(n17652), .B2(n17930), .A(n17752), .ZN(n17681) );
  INV_X1 U20934 ( .A(n17726), .ZN(n17682) );
  OR3_X1 U20935 ( .A1(n17652), .A2(n17682), .A3(P3_REIP_REG_21__SCAN_IN), .ZN(
        n17666) );
  NAND2_X1 U20936 ( .A1(n17681), .A2(n17666), .ZN(n17659) );
  AOI211_X1 U20937 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17669), .A(n17653), .B(
        n17928), .ZN(n17658) );
  INV_X1 U20938 ( .A(n17654), .ZN(n17655) );
  AOI211_X1 U20939 ( .C1(n18596), .C2(n17656), .A(n17655), .B(n17879), .ZN(
        n17657) );
  AOI211_X1 U20940 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17659), .A(n17658), 
        .B(n17657), .ZN(n17660) );
  OAI211_X1 U20941 ( .C1(n17662), .C2(n17918), .A(n17661), .B(n17660), .ZN(
        P3_U2649) );
  AOI211_X1 U20942 ( .C1(n17665), .C2(n17664), .A(n17663), .B(n17879), .ZN(
        n17668) );
  OAI21_X1 U20943 ( .B1(n18037), .B2(n17929), .A(n17666), .ZN(n17667) );
  AOI211_X1 U20944 ( .C1(n17910), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n17668), .B(n17667), .ZN(n17671) );
  OAI211_X1 U20945 ( .C1(n17672), .C2(n18037), .A(n17887), .B(n17669), .ZN(
        n17670) );
  OAI211_X1 U20946 ( .C1(n17681), .C2(n19658), .A(n17671), .B(n17670), .ZN(
        P3_U2650) );
  INV_X1 U20947 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19657) );
  AOI22_X1 U20948 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17910), .B1(
        n17916), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n17680) );
  NOR2_X1 U20949 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17682), .ZN(n17677) );
  AOI211_X1 U20950 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17684), .A(n17672), .B(
        n17928), .ZN(n17676) );
  AOI211_X1 U20951 ( .C1(n18639), .C2(n17674), .A(n17673), .B(n17879), .ZN(
        n17675) );
  AOI211_X1 U20952 ( .C1(n17678), .C2(n17677), .A(n17676), .B(n17675), .ZN(
        n17679) );
  OAI211_X1 U20953 ( .C1(n17681), .C2(n19657), .A(n17680), .B(n17679), .ZN(
        P3_U2651) );
  NAND2_X1 U20954 ( .A1(n17695), .A2(n17750), .ZN(n17714) );
  OAI21_X1 U20955 ( .B1(n19652), .B2(n17714), .A(n17930), .ZN(n17705) );
  NOR4_X1 U20956 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n19652), .A3(n17683), 
        .A4(n17682), .ZN(n17688) );
  OAI211_X1 U20957 ( .C1(n17700), .C2(n17686), .A(n17887), .B(n17684), .ZN(
        n17685) );
  OAI211_X1 U20958 ( .C1(n17929), .C2(n17686), .A(n18992), .B(n17685), .ZN(
        n17687) );
  AOI211_X1 U20959 ( .C1(n17910), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n17688), .B(n17687), .ZN(n17694) );
  INV_X1 U20960 ( .A(n17719), .ZN(n17732) );
  OAI21_X1 U20961 ( .B1(n17732), .B2(n17689), .A(n17843), .ZN(n17699) );
  INV_X1 U20962 ( .A(n17689), .ZN(n17691) );
  OAI21_X1 U20963 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17691), .A(
        n17690), .ZN(n18645) );
  AOI21_X1 U20964 ( .B1(n17699), .B2(n18645), .A(n17879), .ZN(n17692) );
  OAI21_X1 U20965 ( .B1(n17699), .B2(n18645), .A(n17692), .ZN(n17693) );
  OAI211_X1 U20966 ( .C1(n19654), .C2(n17705), .A(n17694), .B(n17693), .ZN(
        P3_U2652) );
  AOI21_X1 U20967 ( .B1(n17695), .B2(n17726), .A(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n17706) );
  AOI21_X1 U20968 ( .B1(n17916), .B2(P3_EBX_REG_18__SCAN_IN), .A(n18905), .ZN(
        n17704) );
  NAND2_X1 U20969 ( .A1(n19598), .A2(n17882), .ZN(n17913) );
  INV_X1 U20970 ( .A(n11504), .ZN(n17696) );
  INV_X1 U20971 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17917) );
  NAND2_X1 U20972 ( .A1(n17917), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17905) );
  INV_X1 U20973 ( .A(n17905), .ZN(n17742) );
  OAI221_X1 U20974 ( .B1(n17698), .B2(n17696), .C1(n17698), .C2(n17742), .A(
        n19598), .ZN(n17697) );
  AOI22_X1 U20975 ( .A1(n17699), .A2(n17698), .B1(n17913), .B2(n17697), .ZN(
        n17702) );
  AOI211_X1 U20976 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17709), .A(n17700), .B(
        n17928), .ZN(n17701) );
  AOI211_X1 U20977 ( .C1(n17910), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17702), .B(n17701), .ZN(n17703) );
  OAI211_X1 U20978 ( .C1(n17706), .C2(n17705), .A(n17704), .B(n17703), .ZN(
        P3_U2653) );
  AOI21_X1 U20979 ( .B1(n18656), .B2(n17742), .A(n17882), .ZN(n17708) );
  INV_X1 U20980 ( .A(n18673), .ZN(n17745) );
  NOR2_X1 U20981 ( .A1(n18678), .A2(n17745), .ZN(n17718) );
  OAI21_X1 U20982 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17718), .A(
        n17707), .ZN(n18667) );
  XOR2_X1 U20983 ( .A(n17708), .B(n18667), .Z(n17717) );
  AOI22_X1 U20984 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17910), .B1(
        n17916), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n17713) );
  OAI211_X1 U20985 ( .C1(n17721), .C2(n17710), .A(n17887), .B(n17709), .ZN(
        n17712) );
  NAND4_X1 U20986 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n17726), .A4(n19650), .ZN(n17711) );
  AND4_X1 U20987 ( .A1(n17713), .A2(n18988), .A3(n17712), .A4(n17711), .ZN(
        n17716) );
  NAND3_X1 U20988 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17930), .A3(n17714), 
        .ZN(n17715) );
  OAI211_X1 U20989 ( .C1(n17879), .C2(n17717), .A(n17716), .B(n17715), .ZN(
        P3_U2654) );
  INV_X1 U20990 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17723) );
  AOI21_X1 U20991 ( .B1(n17723), .B2(n17731), .A(n17718), .ZN(n18674) );
  NOR2_X1 U20992 ( .A1(n17719), .A2(n17882), .ZN(n17720) );
  XNOR2_X1 U20993 ( .A(n18674), .B(n17720), .ZN(n17730) );
  AOI211_X1 U20994 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17737), .A(n17721), .B(
        n17928), .ZN(n17725) );
  NAND3_X1 U20995 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n17726), .A3(n19648), 
        .ZN(n17722) );
  OAI211_X1 U20996 ( .C1(n17723), .C2(n17918), .A(n18992), .B(n17722), .ZN(
        n17724) );
  AOI211_X1 U20997 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17916), .A(n17725), .B(
        n17724), .ZN(n17729) );
  NAND2_X1 U20998 ( .A1(n19646), .A2(n17726), .ZN(n17740) );
  INV_X1 U20999 ( .A(n17740), .ZN(n17727) );
  OAI21_X1 U21000 ( .B1(n17752), .B2(n17727), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n17728) );
  OAI211_X1 U21001 ( .C1(n17730), .C2(n17879), .A(n17729), .B(n17728), .ZN(
        P3_U2655) );
  OAI21_X1 U21002 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18673), .A(
        n17731), .ZN(n18685) );
  OAI21_X1 U21003 ( .B1(n17882), .B2(n17917), .A(n19598), .ZN(n17927) );
  AOI211_X1 U21004 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17913), .A(
        n18685), .B(n17927), .ZN(n17736) );
  NAND2_X1 U21005 ( .A1(n17732), .A2(n18685), .ZN(n17734) );
  AOI22_X1 U21006 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17910), .B1(
        n17916), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n17733) );
  OAI21_X1 U21007 ( .B1(n17919), .B2(n17734), .A(n17733), .ZN(n17735) );
  AOI211_X1 U21008 ( .C1(n17752), .C2(P3_REIP_REG_15__SCAN_IN), .A(n17736), 
        .B(n17735), .ZN(n17741) );
  OAI211_X1 U21009 ( .C1(n17747), .C2(n17738), .A(n17887), .B(n17737), .ZN(
        n17739) );
  NAND4_X1 U21010 ( .A1(n17741), .A2(n18988), .A3(n17740), .A4(n17739), .ZN(
        P3_U2656) );
  AOI21_X1 U21011 ( .B1(n17743), .B2(n17742), .A(n17882), .ZN(n17771) );
  AOI21_X1 U21012 ( .B1(n17843), .B2(n17744), .A(n17771), .ZN(n17756) );
  OAI21_X1 U21013 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17746), .A(
        n17745), .ZN(n18704) );
  XNOR2_X1 U21014 ( .A(n17756), .B(n18704), .ZN(n17755) );
  AOI211_X1 U21015 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17760), .A(n17747), .B(
        n17928), .ZN(n17748) );
  AOI21_X1 U21016 ( .B1(n17910), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17748), .ZN(n17754) );
  NAND3_X1 U21017 ( .A1(n17915), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n17763), 
        .ZN(n17749) );
  OAI22_X1 U21018 ( .A1(n17750), .A2(n17749), .B1(n17929), .B2(n18157), .ZN(
        n17751) );
  AOI211_X1 U21019 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n17752), .A(n18905), 
        .B(n17751), .ZN(n17753) );
  OAI211_X1 U21020 ( .C1(n17879), .C2(n17755), .A(n17754), .B(n17753), .ZN(
        P3_U2657) );
  AOI21_X1 U21021 ( .B1(n17915), .B2(n17775), .A(n17924), .ZN(n17787) );
  NAND2_X1 U21022 ( .A1(n17915), .A2(n19640), .ZN(n17774) );
  NOR3_X1 U21023 ( .A1(n17757), .A2(n17756), .A3(n17879), .ZN(n17769) );
  INV_X1 U21024 ( .A(n17757), .ZN(n17758) );
  AOI211_X1 U21025 ( .C1(n17843), .C2(n17759), .A(n17758), .B(n17927), .ZN(
        n17768) );
  OAI211_X1 U21026 ( .C1(n17773), .C2(n17764), .A(n17887), .B(n17760), .ZN(
        n17761) );
  OAI211_X1 U21027 ( .C1(n17762), .C2(n17918), .A(n18988), .B(n17761), .ZN(
        n17767) );
  NAND2_X1 U21028 ( .A1(n17915), .A2(n17763), .ZN(n17765) );
  OAI22_X1 U21029 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17765), .B1(n17929), 
        .B2(n17764), .ZN(n17766) );
  NOR4_X1 U21030 ( .A1(n17769), .A2(n17768), .A3(n17767), .A4(n17766), .ZN(
        n17770) );
  OAI221_X1 U21031 ( .B1(n19642), .B2(n17787), .C1(n19642), .C2(n17774), .A(
        n17770), .ZN(P3_U2658) );
  AOI22_X1 U21032 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17910), .B1(
        n17916), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n17780) );
  XOR2_X1 U21033 ( .A(n17772), .B(n17771), .Z(n17778) );
  AOI211_X1 U21034 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17790), .A(n17773), .B(
        n17928), .ZN(n17777) );
  OAI21_X1 U21035 ( .B1(n17775), .B2(n17774), .A(n18992), .ZN(n17776) );
  AOI211_X1 U21036 ( .C1(n17778), .C2(n19598), .A(n17777), .B(n17776), .ZN(
        n17779) );
  OAI211_X1 U21037 ( .C1(n19640), .C2(n17787), .A(n17780), .B(n17779), .ZN(
        P3_U2659) );
  INV_X1 U21038 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19636) );
  NOR2_X1 U21039 ( .A1(n19636), .A2(n19634), .ZN(n17782) );
  INV_X1 U21040 ( .A(n17781), .ZN(n17822) );
  NOR2_X1 U21041 ( .A1(n17906), .A2(n17822), .ZN(n17799) );
  AOI21_X1 U21042 ( .B1(n17782), .B2(n17799), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17788) );
  OAI21_X1 U21043 ( .B1(n17783), .B2(n17905), .A(n17843), .ZN(n17784) );
  XOR2_X1 U21044 ( .A(n17785), .B(n17784), .Z(n17786) );
  OAI22_X1 U21045 ( .A1(n17788), .A2(n17787), .B1(n17879), .B2(n17786), .ZN(
        n17789) );
  AOI211_X1 U21046 ( .C1(n17916), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18905), .B(
        n17789), .ZN(n17792) );
  OAI211_X1 U21047 ( .C1(n17797), .C2(n18188), .A(n17887), .B(n17790), .ZN(
        n17791) );
  OAI211_X1 U21048 ( .C1(n17918), .C2(n17793), .A(n17792), .B(n17791), .ZN(
        P3_U2660) );
  INV_X1 U21049 ( .A(n17796), .ZN(n17795) );
  OAI21_X1 U21050 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17795), .A(
        n17794), .ZN(n18719) );
  OAI21_X1 U21051 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17796), .A(
        n17843), .ZN(n17807) );
  XNOR2_X1 U21052 ( .A(n18719), .B(n17807), .ZN(n17805) );
  AOI22_X1 U21053 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17910), .B1(
        n17916), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n17804) );
  AOI21_X1 U21054 ( .B1(n17915), .B2(n17822), .A(n17924), .ZN(n17829) );
  NAND2_X1 U21055 ( .A1(n17799), .A2(n19634), .ZN(n17810) );
  AOI21_X1 U21056 ( .B1(n17829), .B2(n17810), .A(n19636), .ZN(n17802) );
  AOI211_X1 U21057 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17798), .A(n17797), .B(
        n17928), .ZN(n17801) );
  AND3_X1 U21058 ( .A1(n19636), .A2(P3_REIP_REG_9__SCAN_IN), .A3(n17799), .ZN(
        n17800) );
  NOR4_X1 U21059 ( .A1(n18905), .A2(n17802), .A3(n17801), .A4(n17800), .ZN(
        n17803) );
  OAI211_X1 U21060 ( .C1(n17879), .C2(n17805), .A(n17804), .B(n17803), .ZN(
        P3_U2661) );
  NOR2_X1 U21061 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17842), .ZN(
        n17830) );
  AOI21_X1 U21062 ( .B1(n17806), .B2(n17830), .A(n17812), .ZN(n17808) );
  NOR3_X1 U21063 ( .A1(n17808), .A2(n17807), .A3(n17879), .ZN(n17809) );
  AOI211_X1 U21064 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17910), .A(
        n18905), .B(n17809), .ZN(n17817) );
  NOR2_X1 U21065 ( .A1(n17811), .A2(n17928), .ZN(n17819) );
  INV_X1 U21066 ( .A(n17810), .ZN(n17815) );
  AOI21_X1 U21067 ( .B1(n17887), .B2(n17811), .A(n17916), .ZN(n17813) );
  OAI22_X1 U21068 ( .A1(n18231), .A2(n17813), .B1(n17812), .B2(n17913), .ZN(
        n17814) );
  AOI211_X1 U21069 ( .C1(n17819), .C2(n18231), .A(n17815), .B(n17814), .ZN(
        n17816) );
  OAI211_X1 U21070 ( .C1(n17829), .C2(n19634), .A(n17817), .B(n17816), .ZN(
        P3_U2662) );
  NAND2_X1 U21071 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17834), .ZN(n17818) );
  AOI22_X1 U21072 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17910), .B1(
        n17819), .B2(n17818), .ZN(n17828) );
  AOI21_X1 U21073 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17830), .A(
        n17882), .ZN(n17820) );
  XOR2_X1 U21074 ( .A(n17821), .B(n17820), .Z(n17826) );
  INV_X1 U21075 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n18256) );
  NAND2_X1 U21076 ( .A1(n17915), .A2(n17822), .ZN(n17823) );
  OAI22_X1 U21077 ( .A1(n17929), .A2(n18256), .B1(n17824), .B2(n17823), .ZN(
        n17825) );
  AOI211_X1 U21078 ( .C1(n19598), .C2(n17826), .A(n18905), .B(n17825), .ZN(
        n17827) );
  OAI211_X1 U21079 ( .C1(n17829), .C2(n19633), .A(n17828), .B(n17827), .ZN(
        P3_U2663) );
  INV_X1 U21080 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18735) );
  NOR2_X1 U21081 ( .A1(n17830), .A2(n17882), .ZN(n17847) );
  OAI21_X1 U21082 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17832), .A(
        n17831), .ZN(n18745) );
  XNOR2_X1 U21083 ( .A(n17847), .B(n18745), .ZN(n17838) );
  AOI21_X1 U21084 ( .B1(n17915), .B2(n17833), .A(n17924), .ZN(n17860) );
  INV_X1 U21085 ( .A(n17833), .ZN(n17857) );
  NAND3_X1 U21086 ( .A1(n17915), .A2(n17857), .A3(n19628), .ZN(n17845) );
  INV_X1 U21087 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19630) );
  AOI21_X1 U21088 ( .B1(n17860), .B2(n17845), .A(n19630), .ZN(n17837) );
  OAI211_X1 U21089 ( .C1(n17844), .C2(n18255), .A(n17887), .B(n17834), .ZN(
        n17835) );
  OAI211_X1 U21090 ( .C1(n17929), .C2(n18255), .A(n18992), .B(n17835), .ZN(
        n17836) );
  AOI211_X1 U21091 ( .C1(n17838), .C2(n19598), .A(n17837), .B(n17836), .ZN(
        n17841) );
  NAND3_X1 U21092 ( .A1(n17915), .A2(n17839), .A3(n19630), .ZN(n17840) );
  OAI211_X1 U21093 ( .C1(n17918), .C2(n18735), .A(n17841), .B(n17840), .ZN(
        P3_U2664) );
  NOR2_X1 U21094 ( .A1(n18821), .A2(n17020), .ZN(n17855) );
  OAI21_X1 U21095 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17855), .A(
        n17842), .ZN(n18752) );
  AOI211_X1 U21096 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n17843), .A(
        n18752), .B(n17927), .ZN(n17853) );
  AOI211_X1 U21097 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17863), .A(n17844), .B(
        n17928), .ZN(n17852) );
  OAI211_X1 U21098 ( .C1(n17846), .C2(n17918), .A(n18992), .B(n17845), .ZN(
        n17851) );
  INV_X1 U21099 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17849) );
  NAND3_X1 U21100 ( .A1(n19598), .A2(n17847), .A3(n18752), .ZN(n17848) );
  OAI21_X1 U21101 ( .B1(n17849), .B2(n17929), .A(n17848), .ZN(n17850) );
  NOR4_X1 U21102 ( .A1(n17853), .A2(n17852), .A3(n17851), .A4(n17850), .ZN(
        n17854) );
  OAI21_X1 U21103 ( .B1(n17860), .B2(n19628), .A(n17854), .ZN(P3_U2665) );
  AND2_X1 U21104 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18762), .ZN(
        n17867) );
  INV_X1 U21105 ( .A(n17855), .ZN(n17856) );
  OAI21_X1 U21106 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17867), .A(
        n17856), .ZN(n18763) );
  AOI21_X1 U21107 ( .B1(n17867), .B2(n17917), .A(n17882), .ZN(n17870) );
  XNOR2_X1 U21108 ( .A(n18763), .B(n17870), .ZN(n17862) );
  INV_X1 U21109 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19626) );
  NOR2_X1 U21110 ( .A1(n17857), .A2(n17906), .ZN(n17858) );
  AOI22_X1 U21111 ( .A1(n17916), .A2(P3_EBX_REG_5__SCAN_IN), .B1(n17871), .B2(
        n17858), .ZN(n17859) );
  OAI211_X1 U21112 ( .C1(n17860), .C2(n19626), .A(n17859), .B(n18992), .ZN(
        n17861) );
  AOI21_X1 U21113 ( .B1(n17862), .B2(n19598), .A(n17861), .ZN(n17865) );
  OAI211_X1 U21114 ( .C1(n17873), .C2(n18158), .A(n17887), .B(n17863), .ZN(
        n17864) );
  OAI211_X1 U21115 ( .C1(n17918), .C2(n10369), .A(n17865), .B(n17864), .ZN(
        P3_U2666) );
  OR2_X1 U21116 ( .A1(n18821), .A2(n17866), .ZN(n17881) );
  AOI21_X1 U21117 ( .B1(n18783), .B2(n17881), .A(n17867), .ZN(n18779) );
  INV_X1 U21118 ( .A(n18779), .ZN(n17869) );
  NOR3_X1 U21119 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17866), .A3(
        n17905), .ZN(n17868) );
  AOI221_X1 U21120 ( .B1(n17870), .B2(n17869), .C1(n17882), .C2(n18779), .A(
        n17868), .ZN(n17880) );
  AOI211_X1 U21121 ( .C1(n19624), .C2(n17892), .A(n17871), .B(n17906), .ZN(
        n17872) );
  AOI21_X1 U21122 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17916), .A(n17872), .ZN(
        n17878) );
  AOI211_X1 U21123 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17886), .A(n17873), .B(
        n17928), .ZN(n17876) );
  INV_X1 U21124 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19551) );
  NOR2_X1 U21125 ( .A1(n18432), .A2(n19720), .ZN(n17884) );
  AOI21_X1 U21126 ( .B1(n11548), .B2(n19551), .A(n19723), .ZN(n17875) );
  OAI22_X1 U21127 ( .A1(n18783), .A2(n17918), .B1(n19624), .B2(n17932), .ZN(
        n17874) );
  NOR4_X1 U21128 ( .A1(n18905), .A2(n17876), .A3(n17875), .A4(n17874), .ZN(
        n17877) );
  OAI211_X1 U21129 ( .C1(n17880), .C2(n17879), .A(n17878), .B(n17877), .ZN(
        P3_U2667) );
  INV_X1 U21130 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21512) );
  NAND2_X1 U21131 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17903) );
  INV_X1 U21132 ( .A(n17903), .ZN(n17895) );
  OAI21_X1 U21133 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17895), .A(
        n17881), .ZN(n18793) );
  AOI21_X1 U21134 ( .B1(n17895), .B2(n17917), .A(n17882), .ZN(n17883) );
  XNOR2_X1 U21135 ( .A(n18793), .B(n17883), .ZN(n17891) );
  AOI22_X1 U21136 ( .A1(n17924), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n17885), 
        .B2(n17884), .ZN(n17889) );
  OAI211_X1 U21137 ( .C1(n17896), .C2(n18269), .A(n17887), .B(n17886), .ZN(
        n17888) );
  OAI211_X1 U21138 ( .C1(n18269), .C2(n17929), .A(n17889), .B(n17888), .ZN(
        n17890) );
  AOI21_X1 U21139 ( .B1(n17891), .B2(n19598), .A(n17890), .ZN(n17894) );
  INV_X1 U21140 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19620) );
  NOR2_X1 U21141 ( .A1(n21537), .A2(n19620), .ZN(n17907) );
  OAI211_X1 U21142 ( .C1(P3_REIP_REG_3__SCAN_IN), .C2(n17907), .A(n17915), .B(
        n17892), .ZN(n17893) );
  OAI211_X1 U21143 ( .C1(n17918), .C2(n21512), .A(n17894), .B(n17893), .ZN(
        P3_U2668) );
  INV_X1 U21144 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18811) );
  AOI21_X1 U21145 ( .B1(n18821), .B2(n18811), .A(n17895), .ZN(n18807) );
  INV_X1 U21146 ( .A(n18807), .ZN(n17914) );
  NAND2_X1 U21147 ( .A1(n18288), .A2(n18282), .ZN(n17897) );
  AOI211_X1 U21148 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17897), .A(n17896), .B(
        n17928), .ZN(n17902) );
  OAI22_X1 U21149 ( .A1(n17929), .A2(n17898), .B1(n19620), .B2(n17932), .ZN(
        n17901) );
  NOR2_X1 U21150 ( .A1(n17899), .A2(n19723), .ZN(n17900) );
  NOR3_X1 U21151 ( .A1(n17902), .A2(n17901), .A3(n17900), .ZN(n17912) );
  NOR2_X1 U21152 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17903), .ZN(
        n17904) );
  AOI211_X1 U21153 ( .C1(n18807), .C2(n17905), .A(n17904), .B(n17919), .ZN(
        n17909) );
  AOI211_X1 U21154 ( .C1(n21537), .C2(n19620), .A(n17907), .B(n17906), .ZN(
        n17908) );
  AOI211_X1 U21155 ( .C1(n17910), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17909), .B(n17908), .ZN(n17911) );
  OAI211_X1 U21156 ( .C1(n17914), .C2(n17913), .A(n17912), .B(n17911), .ZN(
        P3_U2669) );
  AOI22_X1 U21157 ( .A1(n17916), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n17915), .B2(
        n21537), .ZN(n17926) );
  AOI221_X1 U21158 ( .B1(n17919), .B2(n17918), .C1(n17917), .C2(n17918), .A(
        n18821), .ZN(n17923) );
  OAI21_X1 U21159 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17920), .ZN(n18283) );
  OAI22_X1 U21160 ( .A1(n17928), .A2(n18283), .B1(n19723), .B2(n17921), .ZN(
        n17922) );
  AOI211_X1 U21161 ( .C1(n17924), .C2(P3_REIP_REG_1__SCAN_IN), .A(n17923), .B(
        n17922), .ZN(n17925) );
  OAI211_X1 U21162 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17927), .A(
        n17926), .B(n17925), .ZN(P3_U2670) );
  NAND2_X1 U21163 ( .A1(n17929), .A2(n17928), .ZN(n17931) );
  AOI22_X1 U21164 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17931), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17930), .ZN(n17934) );
  NAND3_X1 U21165 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19719), .A3(
        n17932), .ZN(n17933) );
  OAI211_X1 U21166 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n19723), .A(
        n17934), .B(n17933), .ZN(P3_U2671) );
  NOR4_X1 U21167 ( .A1(n17937), .A2(n17936), .A3(n17935), .A4(n18037), .ZN(
        n17940) );
  NAND2_X1 U21168 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .ZN(n17938) );
  NOR4_X1 U21169 ( .A1(n17982), .A2(n10149), .A3(n18069), .A4(n17938), .ZN(
        n17939) );
  NAND4_X1 U21170 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17940), .A4(n17939), .ZN(n17943) );
  NOR2_X1 U21171 ( .A1(n17944), .A2(n17943), .ZN(n17977) );
  NAND2_X1 U21172 ( .A1(n18270), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17942) );
  NAND2_X1 U21173 ( .A1(n17977), .A2(n19140), .ZN(n17941) );
  OAI22_X1 U21174 ( .A1(n17977), .A2(n17942), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17941), .ZN(P3_U2672) );
  NAND2_X1 U21175 ( .A1(n17944), .A2(n17943), .ZN(n17945) );
  NAND2_X1 U21176 ( .A1(n17945), .A2(n18270), .ZN(n17976) );
  AOI22_X1 U21177 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17949) );
  AOI22_X1 U21178 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17948) );
  AOI22_X1 U21179 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17947) );
  AOI22_X1 U21180 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17946) );
  NAND4_X1 U21181 ( .A1(n17949), .A2(n17948), .A3(n17947), .A4(n17946), .ZN(
        n17958) );
  INV_X1 U21182 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18012) );
  INV_X1 U21183 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17951) );
  INV_X1 U21184 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17950) );
  OAI22_X1 U21185 ( .A1(n18198), .A2(n18013), .B1(n18200), .B2(n10130), .ZN(
        n17952) );
  AOI211_X1 U21186 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17953), .B(n17952), .ZN(n17956) );
  AOI22_X1 U21187 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17955) );
  OAI211_X1 U21188 ( .C1(n18251), .C2(n18012), .A(n17956), .B(n17955), .ZN(
        n17957) );
  OR2_X1 U21189 ( .A1(n17958), .A2(n17957), .ZN(n17980) );
  NAND3_X1 U21190 ( .A1(n17979), .A2(n17978), .A3(n17980), .ZN(n17975) );
  AOI22_X1 U21191 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17960) );
  NAND2_X1 U21192 ( .A1(n13434), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n17959) );
  OAI211_X1 U21193 ( .C1(n17961), .C2(n18216), .A(n17960), .B(n17959), .ZN(
        n17967) );
  INV_X1 U21194 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18132) );
  OAI22_X1 U21195 ( .A1(n18198), .A2(n17962), .B1(n18196), .B2(n18132), .ZN(
        n17966) );
  INV_X1 U21196 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17964) );
  OAI22_X1 U21197 ( .A1(n18202), .A2(n17964), .B1(n18200), .B2(n17963), .ZN(
        n17965) );
  OR3_X1 U21198 ( .A1(n17967), .A2(n17966), .A3(n17965), .ZN(n17973) );
  AOI22_X1 U21199 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17971) );
  AOI22_X1 U21200 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18192), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17970) );
  AOI22_X1 U21201 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17969) );
  AOI22_X1 U21202 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17968) );
  NAND4_X1 U21203 ( .A1(n17971), .A2(n17970), .A3(n17969), .A4(n17968), .ZN(
        n17972) );
  NOR2_X1 U21204 ( .A1(n17973), .A2(n17972), .ZN(n17974) );
  XNOR2_X1 U21205 ( .A(n17975), .B(n17974), .ZN(n18299) );
  OAI22_X1 U21206 ( .A1(n17977), .A2(n17976), .B1(n18299), .B2(n18270), .ZN(
        P3_U2673) );
  NAND2_X1 U21207 ( .A1(n17979), .A2(n17978), .ZN(n17981) );
  XOR2_X1 U21208 ( .A(n17981), .B(n17980), .Z(n18306) );
  OAI21_X1 U21209 ( .B1(n18270), .B2(n18306), .A(n17984), .ZN(P3_U2674) );
  OAI21_X1 U21210 ( .B1(n17987), .B2(n17986), .A(n17985), .ZN(n18315) );
  NAND3_X1 U21211 ( .A1(n17989), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18270), 
        .ZN(n17988) );
  OAI221_X1 U21212 ( .B1(n17989), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18270), 
        .C2(n18315), .A(n17988), .ZN(P3_U2676) );
  AOI21_X1 U21213 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18270), .A(n17997), .ZN(
        n17991) );
  XNOR2_X1 U21214 ( .A(n17990), .B(n17993), .ZN(n18319) );
  OAI22_X1 U21215 ( .A1(n17992), .A2(n17991), .B1(n18270), .B2(n18319), .ZN(
        P3_U2677) );
  AOI21_X1 U21216 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18270), .A(n18000), .ZN(
        n17996) );
  OAI21_X1 U21217 ( .B1(n17995), .B2(n17994), .A(n17993), .ZN(n18323) );
  OAI22_X1 U21218 ( .A1(n17997), .A2(n17996), .B1(n18270), .B2(n18323), .ZN(
        P3_U2678) );
  AOI21_X1 U21219 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18270), .A(n9735), .ZN(
        n17999) );
  XNOR2_X1 U21220 ( .A(n17998), .B(n18001), .ZN(n18329) );
  OAI22_X1 U21221 ( .A1(n18000), .A2(n17999), .B1(n18270), .B2(n18329), .ZN(
        P3_U2679) );
  AOI22_X1 U21222 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n18270), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n18005), .ZN(n18004) );
  OAI21_X1 U21223 ( .B1(n18003), .B2(n18002), .A(n18001), .ZN(n18335) );
  OAI22_X1 U21224 ( .A1(n9735), .A2(n18004), .B1(n18270), .B2(n18335), .ZN(
        P3_U2680) );
  AOI22_X1 U21225 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18009) );
  AOI22_X1 U21226 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18008) );
  AOI22_X1 U21227 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18007) );
  AOI22_X1 U21228 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18006) );
  NAND4_X1 U21229 ( .A1(n18009), .A2(n18008), .A3(n18007), .A4(n18006), .ZN(
        n18019) );
  INV_X1 U21230 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18140) );
  INV_X1 U21231 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18011) );
  INV_X1 U21232 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18010) );
  OAI22_X1 U21233 ( .A1(n18079), .A2(n18013), .B1(n11548), .B2(n18012), .ZN(
        n18014) );
  AOI211_X1 U21234 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n18015), .B(n18014), .ZN(n18017) );
  AOI22_X1 U21235 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18016) );
  OAI211_X1 U21236 ( .C1(n18251), .C2(n18140), .A(n18017), .B(n18016), .ZN(
        n18018) );
  NOR2_X1 U21237 ( .A1(n18019), .A2(n18018), .ZN(n18338) );
  NAND3_X1 U21238 ( .A1(n10151), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n18270), 
        .ZN(n18020) );
  OAI221_X1 U21239 ( .B1(n10151), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n18270), 
        .C2(n18338), .A(n18020), .ZN(P3_U2681) );
  OAI21_X1 U21240 ( .B1(n10149), .B2(n18069), .A(n18270), .ZN(n18054) );
  INV_X1 U21241 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18029) );
  INV_X1 U21242 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18024) );
  OAI22_X1 U21243 ( .A1(n11598), .A2(n18024), .B1(n11548), .B2(n18023), .ZN(
        n18025) );
  AOI211_X1 U21244 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n18026), .B(n18025), .ZN(n18028) );
  AOI22_X1 U21245 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18027) );
  OAI211_X1 U21246 ( .C1(n18216), .C2(n18029), .A(n18028), .B(n18027), .ZN(
        n18035) );
  AOI22_X1 U21247 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18033) );
  AOI22_X1 U21248 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18032) );
  AOI22_X1 U21249 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18031) );
  AOI22_X1 U21250 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18030) );
  NAND4_X1 U21251 ( .A1(n18033), .A2(n18032), .A3(n18031), .A4(n18030), .ZN(
        n18034) );
  OR2_X1 U21252 ( .A1(n18035), .A2(n18034), .ZN(n18343) );
  NAND2_X1 U21253 ( .A1(n18286), .A2(n18343), .ZN(n18036) );
  OAI221_X1 U21254 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18038), .C1(n18037), 
        .C2(n18054), .A(n18036), .ZN(P3_U2682) );
  INV_X1 U21255 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18041) );
  NAND2_X1 U21256 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n18040) );
  NAND2_X1 U21257 ( .A1(n11604), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n18039) );
  OAI211_X1 U21258 ( .C1(n18216), .C2(n18041), .A(n18040), .B(n18039), .ZN(
        n18042) );
  INV_X1 U21259 ( .A(n18042), .ZN(n18046) );
  AOI22_X1 U21260 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18045) );
  AOI22_X1 U21261 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18044) );
  NAND2_X1 U21262 ( .A1(n17252), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n18043) );
  NAND4_X1 U21263 ( .A1(n18046), .A2(n18045), .A3(n18044), .A4(n18043), .ZN(
        n18052) );
  AOI22_X1 U21264 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17269), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18050) );
  AOI22_X1 U21265 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18049) );
  AOI22_X1 U21266 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18048) );
  AOI22_X1 U21267 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18047) );
  NAND4_X1 U21268 ( .A1(n18050), .A2(n18049), .A3(n18048), .A4(n18047), .ZN(
        n18051) );
  NOR2_X1 U21269 ( .A1(n18052), .A2(n18051), .ZN(n18347) );
  NOR2_X1 U21270 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18053), .ZN(n18055) );
  OAI22_X1 U21271 ( .A1(n18347), .A2(n18270), .B1(n18055), .B2(n18054), .ZN(
        P3_U2683) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n9589), .B1(
        n18192), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18056) );
  OAI21_X1 U21273 ( .B1(n17954), .B2(n18057), .A(n18056), .ZN(n18058) );
  AOI21_X1 U21274 ( .B1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n11603), .A(
        n18058), .ZN(n18061) );
  AOI22_X1 U21275 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18060) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n9593), .B1(
        n18219), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18059) );
  NAND3_X1 U21277 ( .A1(n18061), .A2(n18060), .A3(n18059), .ZN(n18068) );
  AOI22_X1 U21278 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18066) );
  AOI22_X1 U21279 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18065) );
  AOI22_X1 U21280 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18064) );
  AOI22_X1 U21281 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18063) );
  NAND4_X1 U21282 ( .A1(n18066), .A2(n18065), .A3(n18064), .A4(n18063), .ZN(
        n18067) );
  NOR2_X1 U21283 ( .A1(n18068), .A2(n18067), .ZN(n18356) );
  OAI21_X1 U21284 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18088), .A(n18069), .ZN(
        n18070) );
  AOI22_X1 U21285 ( .A1(n18286), .A2(n18356), .B1(n18070), .B2(n18270), .ZN(
        P3_U2684) );
  OAI21_X1 U21286 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n18071), .A(n18270), .ZN(
        n18087) );
  AOI22_X1 U21287 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18075) );
  AOI22_X1 U21288 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U21289 ( .A1(n11607), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18073) );
  AOI22_X1 U21290 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18072) );
  NAND4_X1 U21291 ( .A1(n18075), .A2(n18074), .A3(n18073), .A4(n18072), .ZN(
        n18086) );
  INV_X1 U21292 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18084) );
  INV_X1 U21293 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18077) );
  INV_X1 U21294 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18078) );
  OAI22_X1 U21295 ( .A1(n18079), .A2(n18195), .B1(n18200), .B2(n18078), .ZN(
        n18080) );
  AOI211_X1 U21296 ( .C1(n18244), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n18081), .B(n18080), .ZN(n18083) );
  AOI22_X1 U21297 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18082) );
  OAI211_X1 U21298 ( .C1(n18216), .C2(n18084), .A(n18083), .B(n18082), .ZN(
        n18085) );
  NOR2_X1 U21299 ( .A1(n18086), .A2(n18085), .ZN(n18361) );
  OAI22_X1 U21300 ( .A1(n18088), .A2(n18087), .B1(n18361), .B2(n18270), .ZN(
        P3_U2685) );
  INV_X1 U21301 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18092) );
  AOI22_X1 U21302 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18091) );
  NAND2_X1 U21303 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n18090) );
  OAI211_X1 U21304 ( .C1(n18092), .C2(n18216), .A(n18091), .B(n18090), .ZN(
        n18093) );
  INV_X1 U21305 ( .A(n18093), .ZN(n18096) );
  AOI22_X1 U21306 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18095) );
  AOI22_X1 U21307 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18094) );
  NAND3_X1 U21308 ( .A1(n18096), .A2(n18095), .A3(n18094), .ZN(n18102) );
  AOI22_X1 U21309 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18244), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18100) );
  AOI22_X1 U21310 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18099) );
  AOI22_X1 U21311 ( .A1(n11607), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18219), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18098) );
  AOI22_X1 U21312 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18097) );
  NAND4_X1 U21313 ( .A1(n18100), .A2(n18099), .A3(n18098), .A4(n18097), .ZN(
        n18101) );
  NOR2_X1 U21314 ( .A1(n18102), .A2(n18101), .ZN(n18366) );
  OAI21_X1 U21315 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18104), .A(n18103), .ZN(
        n18105) );
  AOI22_X1 U21316 ( .A1(n18286), .A2(n18366), .B1(n18105), .B2(n18270), .ZN(
        P3_U2686) );
  NAND2_X1 U21317 ( .A1(n18270), .A2(n18120), .ZN(n18136) );
  INV_X1 U21318 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18247) );
  OAI22_X1 U21319 ( .A1(n11598), .A2(n18247), .B1(n11548), .B2(n18108), .ZN(
        n18109) );
  AOI211_X1 U21320 ( .C1(n18244), .C2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n18110), .B(n18109), .ZN(n18112) );
  AOI22_X1 U21321 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18111) );
  OAI211_X1 U21322 ( .C1(n18216), .C2(n18113), .A(n18112), .B(n18111), .ZN(
        n18119) );
  AOI22_X1 U21323 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18117) );
  AOI22_X1 U21324 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18116) );
  AOI22_X1 U21325 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18115) );
  AOI22_X1 U21326 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18114) );
  NAND4_X1 U21327 ( .A1(n18117), .A2(n18116), .A3(n18115), .A4(n18114), .ZN(
        n18118) );
  OR2_X1 U21328 ( .A1(n18119), .A2(n18118), .ZN(n18367) );
  NOR3_X1 U21329 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18277), .A3(n18120), .ZN(
        n18121) );
  AOI21_X1 U21330 ( .B1(n18286), .B2(n18367), .A(n18121), .ZN(n18122) );
  OAI21_X1 U21331 ( .B1(n18123), .B2(n18136), .A(n18122), .ZN(P3_U2687) );
  AOI22_X1 U21332 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18174), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18127) );
  AOI22_X1 U21333 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18126) );
  AOI22_X1 U21334 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18125) );
  AOI22_X1 U21335 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18124) );
  NAND4_X1 U21336 ( .A1(n18127), .A2(n18126), .A3(n18125), .A4(n18124), .ZN(
        n18134) );
  AOI22_X1 U21337 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18129) );
  AOI22_X1 U21338 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18128) );
  AOI22_X1 U21339 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18131) );
  OAI211_X1 U21340 ( .C1(n18216), .C2(n18132), .A(n9794), .B(n18131), .ZN(
        n18133) );
  NOR2_X1 U21341 ( .A1(n18134), .A2(n18133), .ZN(n18378) );
  NOR2_X1 U21342 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n18135), .ZN(n18137) );
  OAI22_X1 U21343 ( .A1(n18378), .A2(n18270), .B1(n18137), .B2(n18136), .ZN(
        P3_U2688) );
  NAND2_X1 U21344 ( .A1(n18270), .A2(n18153), .ZN(n18156) );
  INV_X1 U21345 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18146) );
  INV_X1 U21346 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18139) );
  INV_X1 U21347 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18138) );
  OAI22_X1 U21348 ( .A1(n11598), .A2(n18141), .B1(n11548), .B2(n18140), .ZN(
        n18142) );
  AOI211_X1 U21349 ( .C1(n17252), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n18143), .B(n18142), .ZN(n18145) );
  AOI22_X1 U21350 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18144) );
  OAI211_X1 U21351 ( .C1(n18216), .C2(n18146), .A(n18145), .B(n18144), .ZN(
        n18152) );
  AOI22_X1 U21352 ( .A1(n18248), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18150) );
  AOI22_X1 U21353 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18149) );
  AOI22_X1 U21354 ( .A1(n18219), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18148) );
  AOI22_X1 U21355 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18147) );
  NAND4_X1 U21356 ( .A1(n18150), .A2(n18149), .A3(n18148), .A4(n18147), .ZN(
        n18151) );
  OR2_X1 U21357 ( .A1(n18152), .A2(n18151), .ZN(n18381) );
  NOR3_X1 U21358 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18277), .A3(n18153), .ZN(
        n18154) );
  AOI21_X1 U21359 ( .B1(n18286), .B2(n18381), .A(n18154), .ZN(n18155) );
  OAI21_X1 U21360 ( .B1(n18157), .B2(n18156), .A(n18155), .ZN(P3_U2689) );
  NOR2_X1 U21361 ( .A1(n18158), .A2(n18264), .ZN(n18267) );
  NAND2_X1 U21362 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18267), .ZN(n18262) );
  NOR2_X1 U21363 ( .A1(n18255), .A2(n18262), .ZN(n18254) );
  NAND2_X1 U21364 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18254), .ZN(n18230) );
  NAND2_X1 U21365 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18234), .ZN(n18212) );
  NOR2_X1 U21366 ( .A1(n18188), .A2(n18212), .ZN(n18191) );
  OAI21_X1 U21367 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n18191), .A(n18270), .ZN(
        n18172) );
  AOI22_X1 U21368 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18160) );
  NAND2_X1 U21369 ( .A1(n11603), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n18159) );
  OAI211_X1 U21370 ( .C1(n18161), .C2(n18196), .A(n18160), .B(n18159), .ZN(
        n18162) );
  INV_X1 U21371 ( .A(n18162), .ZN(n18165) );
  AOI22_X1 U21372 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18164) );
  AOI22_X1 U21373 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18219), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18163) );
  NAND3_X1 U21374 ( .A1(n18165), .A2(n18164), .A3(n18163), .ZN(n18171) );
  AOI22_X1 U21375 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18169) );
  AOI22_X1 U21376 ( .A1(n17269), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18168) );
  AOI22_X1 U21377 ( .A1(n11607), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18167) );
  AOI22_X1 U21378 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18166) );
  NAND4_X1 U21379 ( .A1(n18169), .A2(n18168), .A3(n18167), .A4(n18166), .ZN(
        n18170) );
  NOR2_X1 U21380 ( .A1(n18171), .A2(n18170), .ZN(n18392) );
  OAI22_X1 U21381 ( .A1(n18173), .A2(n18172), .B1(n18392), .B2(n18270), .ZN(
        P3_U2691) );
  INV_X1 U21382 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18177) );
  AOI22_X1 U21383 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18176) );
  NAND2_X1 U21384 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n18175) );
  OAI211_X1 U21385 ( .C1(n18216), .C2(n18177), .A(n18176), .B(n18175), .ZN(
        n18178) );
  INV_X1 U21386 ( .A(n18178), .ZN(n18181) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18219), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18180) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n17281), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18179) );
  NAND3_X1 U21389 ( .A1(n18181), .A2(n18180), .A3(n18179), .ZN(n18187) );
  AOI22_X1 U21390 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18185) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n9589), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18184) );
  AOI22_X1 U21392 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18183) );
  AOI22_X1 U21393 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18182) );
  NAND4_X1 U21394 ( .A1(n18185), .A2(n18184), .A3(n18183), .A4(n18182), .ZN(
        n18186) );
  NOR2_X1 U21395 ( .A1(n18187), .A2(n18186), .ZN(n18395) );
  AOI21_X1 U21396 ( .B1(n18188), .B2(n18212), .A(n18286), .ZN(n18189) );
  INV_X1 U21397 ( .A(n18189), .ZN(n18190) );
  OAI22_X1 U21398 ( .A1(n18395), .A2(n18270), .B1(n18191), .B2(n18190), .ZN(
        P3_U2692) );
  INV_X1 U21399 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18281) );
  AOI22_X1 U21400 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18194) );
  NAND2_X1 U21401 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n18193) );
  OAI211_X1 U21402 ( .C1(n18281), .C2(n18216), .A(n18194), .B(n18193), .ZN(
        n18205) );
  INV_X1 U21403 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18197) );
  OAI22_X1 U21404 ( .A1(n18198), .A2(n18197), .B1(n18196), .B2(n18195), .ZN(
        n18204) );
  INV_X1 U21405 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18199) );
  OAI22_X1 U21406 ( .A1(n18202), .A2(n18201), .B1(n18200), .B2(n18199), .ZN(
        n18203) );
  OR3_X1 U21407 ( .A1(n18205), .A2(n18204), .A3(n18203), .ZN(n18211) );
  AOI22_X1 U21408 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18209) );
  AOI22_X1 U21409 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18208) );
  AOI22_X1 U21410 ( .A1(n11607), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18207) );
  AOI22_X1 U21411 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18206) );
  NAND4_X1 U21412 ( .A1(n18209), .A2(n18208), .A3(n18207), .A4(n18206), .ZN(
        n18210) );
  NOR2_X1 U21413 ( .A1(n18211), .A2(n18210), .ZN(n18402) );
  OAI21_X1 U21414 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18234), .A(n18212), .ZN(
        n18213) );
  AOI22_X1 U21415 ( .A1(n18286), .A2(n18402), .B1(n18213), .B2(n18270), .ZN(
        P3_U2693) );
  INV_X1 U21416 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18217) );
  AOI22_X1 U21417 ( .A1(n18089), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18215) );
  NAND2_X1 U21418 ( .A1(n11605), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n18214) );
  OAI211_X1 U21419 ( .C1(n18217), .C2(n18216), .A(n18215), .B(n18214), .ZN(
        n18218) );
  INV_X1 U21420 ( .A(n18218), .ZN(n18222) );
  AOI22_X1 U21421 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18221) );
  AOI22_X1 U21422 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18219), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18220) );
  NAND3_X1 U21423 ( .A1(n18222), .A2(n18221), .A3(n18220), .ZN(n18229) );
  AOI22_X1 U21424 ( .A1(n18223), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17252), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18227) );
  AOI22_X1 U21425 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18192), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18226) );
  AOI22_X1 U21426 ( .A1(n18174), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18238), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18225) );
  AOI22_X1 U21427 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18224) );
  NAND4_X1 U21428 ( .A1(n18227), .A2(n18226), .A3(n18225), .A4(n18224), .ZN(
        n18228) );
  NOR2_X1 U21429 ( .A1(n18229), .A2(n18228), .ZN(n18404) );
  AOI21_X1 U21430 ( .B1(n18231), .B2(n18230), .A(n18286), .ZN(n18232) );
  INV_X1 U21431 ( .A(n18232), .ZN(n18233) );
  OAI22_X1 U21432 ( .A1(n18404), .A2(n18270), .B1(n18234), .B2(n18233), .ZN(
        P3_U2694) );
  AOI22_X1 U21433 ( .A1(n11607), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18235), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18242) );
  AOI22_X1 U21434 ( .A1(n18237), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18236), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18241) );
  AOI22_X1 U21435 ( .A1(n18192), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17208), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18240) );
  AOI22_X1 U21436 ( .A1(n18238), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13434), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18239) );
  NAND4_X1 U21437 ( .A1(n18242), .A2(n18241), .A3(n18240), .A4(n18239), .ZN(
        n18253) );
  INV_X1 U21438 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18250) );
  AOI22_X1 U21439 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9589), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18246) );
  AOI22_X1 U21440 ( .A1(n18244), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18243), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18245) );
  AOI22_X1 U21441 ( .A1(n17281), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18249) );
  OAI211_X1 U21442 ( .C1(n18251), .C2(n18250), .A(n9795), .B(n18249), .ZN(
        n18252) );
  NOR2_X1 U21443 ( .A1(n18253), .A2(n18252), .ZN(n18407) );
  NOR2_X1 U21444 ( .A1(n18286), .A2(n18254), .ZN(n18259) );
  NOR3_X1 U21445 ( .A1(n18277), .A2(n18255), .A3(n18262), .ZN(n18257) );
  AOI22_X1 U21446 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18259), .B1(n18257), .B2(
        n18256), .ZN(n18258) );
  OAI21_X1 U21447 ( .B1(n18407), .B2(n18270), .A(n18258), .ZN(P3_U2695) );
  INV_X1 U21448 ( .A(n18262), .ZN(n18260) );
  OAI21_X1 U21449 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18260), .A(n18259), .ZN(
        n18261) );
  OAI21_X1 U21450 ( .B1(n18270), .B2(n18132), .A(n18261), .ZN(P3_U2696) );
  OAI21_X1 U21451 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18267), .A(n18262), .ZN(
        n18263) );
  AOI22_X1 U21452 ( .A1(n18286), .A2(n18146), .B1(n18263), .B2(n18270), .ZN(
        P3_U2697) );
  INV_X1 U21453 ( .A(n18264), .ZN(n18273) );
  OAI21_X1 U21454 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18273), .A(n18270), .ZN(
        n18266) );
  INV_X1 U21455 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18265) );
  OAI22_X1 U21456 ( .A1(n18267), .A2(n18266), .B1(n18265), .B2(n18270), .ZN(
        P3_U2698) );
  NAND2_X1 U21457 ( .A1(n19140), .A2(n18289), .ZN(n18284) );
  INV_X1 U21458 ( .A(n18284), .ZN(n18285) );
  NAND2_X1 U21459 ( .A1(n18268), .A2(n18285), .ZN(n18274) );
  NOR2_X1 U21460 ( .A1(n18269), .A2(n18274), .ZN(n18276) );
  AOI21_X1 U21461 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18270), .A(n18276), .ZN(
        n18272) );
  INV_X1 U21462 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18271) );
  OAI22_X1 U21463 ( .A1(n18273), .A2(n18272), .B1(n18271), .B2(n18270), .ZN(
        P3_U2699) );
  INV_X1 U21464 ( .A(n18274), .ZN(n18279) );
  AOI21_X1 U21465 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18270), .A(n18279), .ZN(
        n18275) );
  OAI22_X1 U21466 ( .A1(n18276), .A2(n18275), .B1(n18177), .B2(n18270), .ZN(
        P3_U2700) );
  AOI221_X1 U21467 ( .B1(n18278), .B2(n18289), .C1(n18277), .C2(n18289), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n18280) );
  AOI211_X1 U21468 ( .C1(n18286), .C2(n18281), .A(n18280), .B(n18279), .ZN(
        P3_U2701) );
  OAI222_X1 U21469 ( .A1(n18284), .A2(n18283), .B1(n18282), .B2(n18289), .C1(
        n18217), .C2(n18270), .ZN(P3_U2702) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18286), .B1(
        n18285), .B2(n18288), .ZN(n18287) );
  OAI21_X1 U21471 ( .B1(n18289), .B2(n18288), .A(n18287), .ZN(P3_U2703) );
  INV_X1 U21472 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18438) );
  INV_X1 U21473 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18443) );
  INV_X1 U21474 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18445) );
  INV_X1 U21475 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18458) );
  NAND4_X1 U21476 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n18292)
         );
  NAND4_X1 U21477 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_5__SCAN_IN), .ZN(n18291) );
  INV_X1 U21478 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18484) );
  INV_X1 U21479 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18486) );
  NOR4_X1 U21480 ( .A1(n18484), .A2(n18486), .A3(n18515), .A4(n18491), .ZN(
        n18380) );
  NAND4_X1 U21481 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18380), .A3(
        P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n18290) );
  NOR4_X2 U21482 ( .A1(n18293), .A2(n18292), .A3(n18291), .A4(n18290), .ZN(
        n18383) );
  NAND2_X1 U21483 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n18383), .ZN(n18375) );
  NOR2_X2 U21484 ( .A1(n18458), .A2(n18375), .ZN(n18369) );
  INV_X1 U21485 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18497) );
  NAND3_X1 U21486 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .ZN(n18336) );
  NOR3_X1 U21487 ( .A1(n21491), .A2(n18497), .A3(n18336), .ZN(n18340) );
  NAND3_X1 U21488 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18369), .A3(n18340), 
        .ZN(n18331) );
  NOR2_X2 U21489 ( .A1(n18445), .A2(n18331), .ZN(n18330) );
  NAND2_X1 U21490 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18311), .ZN(n18308) );
  NOR2_X1 U21491 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n18302), .ZN(n18296) );
  AOI22_X1 U21492 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18296), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18295), .ZN(n18297) );
  OAI21_X1 U21493 ( .B1(n18298), .B2(n18337), .A(n18297), .ZN(P3_U2704) );
  INV_X1 U21494 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18512) );
  NAND2_X1 U21495 ( .A1(n19131), .A2(n18370), .ZN(n18374) );
  INV_X1 U21496 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n20014) );
  OAI22_X1 U21497 ( .A1(n18299), .A2(n18427), .B1(n20014), .B2(n18337), .ZN(
        n18300) );
  AOI21_X1 U21498 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18362), .A(n18300), .ZN(
        n18301) );
  OAI221_X1 U21499 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18302), .C1(n18512), 
        .C2(n9699), .A(n18301), .ZN(P3_U2705) );
  AOI22_X1 U21500 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18362), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18368), .ZN(n18305) );
  OAI211_X1 U21501 ( .C1(n18303), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18425), .B(
        n18302), .ZN(n18304) );
  OAI211_X1 U21502 ( .C1(n18427), .C2(n18306), .A(n18305), .B(n18304), .ZN(
        P3_U2706) );
  AOI22_X1 U21503 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18362), .B1(n18307), .B2(
        n18382), .ZN(n18310) );
  OAI211_X1 U21504 ( .C1(n18311), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18425), .B(
        n18308), .ZN(n18309) );
  OAI211_X1 U21505 ( .C1(n18337), .C2(n19125), .A(n18310), .B(n18309), .ZN(
        P3_U2707) );
  AOI22_X1 U21506 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18362), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18368), .ZN(n18314) );
  AOI211_X1 U21507 ( .C1(n18438), .C2(n18316), .A(n18311), .B(n18370), .ZN(
        n18312) );
  INV_X1 U21508 ( .A(n18312), .ZN(n18313) );
  OAI211_X1 U21509 ( .C1(n18427), .C2(n18315), .A(n18314), .B(n18313), .ZN(
        P3_U2708) );
  AOI22_X1 U21510 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18362), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18368), .ZN(n18318) );
  OAI211_X1 U21511 ( .C1(n9639), .C2(P3_EAX_REG_26__SCAN_IN), .A(n18425), .B(
        n18316), .ZN(n18317) );
  OAI211_X1 U21512 ( .C1(n18319), .C2(n18427), .A(n18318), .B(n18317), .ZN(
        P3_U2709) );
  AOI22_X1 U21513 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18362), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18368), .ZN(n18322) );
  AOI211_X1 U21514 ( .C1(n18441), .C2(n18325), .A(n9639), .B(n18370), .ZN(
        n18320) );
  INV_X1 U21515 ( .A(n18320), .ZN(n18321) );
  OAI211_X1 U21516 ( .C1(n18323), .C2(n18427), .A(n18322), .B(n18321), .ZN(
        P3_U2710) );
  AOI22_X1 U21517 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18362), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18368), .ZN(n18328) );
  OAI21_X1 U21518 ( .B1(n18443), .B2(n18370), .A(n18324), .ZN(n18326) );
  NAND2_X1 U21519 ( .A1(n18326), .A2(n18325), .ZN(n18327) );
  OAI211_X1 U21520 ( .C1(n18329), .C2(n18427), .A(n18328), .B(n18327), .ZN(
        P3_U2711) );
  AOI211_X1 U21521 ( .C1(n18445), .C2(n18331), .A(n18370), .B(n18330), .ZN(
        n18332) );
  AOI21_X1 U21522 ( .B1(n18368), .B2(BUF2_REG_23__SCAN_IN), .A(n18332), .ZN(
        n18334) );
  NAND2_X1 U21523 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18362), .ZN(n18333) );
  OAI211_X1 U21524 ( .C1(n18335), .C2(n18427), .A(n18334), .B(n18333), .ZN(
        P3_U2712) );
  NAND3_X1 U21525 ( .A1(n19140), .A2(n18369), .A3(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n18363) );
  NOR2_X1 U21526 ( .A1(n18336), .A2(n18363), .ZN(n18352) );
  NOR2_X1 U21527 ( .A1(n18370), .A2(n18352), .ZN(n18349) );
  AND2_X1 U21528 ( .A1(n21491), .A2(n18352), .ZN(n18344) );
  OAI22_X1 U21529 ( .A1(n18338), .A2(n18427), .B1(n19134), .B2(n18337), .ZN(
        n18339) );
  AOI221_X1 U21530 ( .B1(n18349), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n18344), 
        .C2(P3_EAX_REG_22__SCAN_IN), .A(n18339), .ZN(n18342) );
  INV_X1 U21531 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18447) );
  NAND4_X1 U21532 ( .A1(n19140), .A2(n18369), .A3(n18340), .A4(n18447), .ZN(
        n18341) );
  OAI211_X1 U21533 ( .C1(n18374), .C2(n14001), .A(n18342), .B(n18341), .ZN(
        P3_U2713) );
  AOI22_X1 U21534 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18368), .B1(n18382), .B2(
        n18343), .ZN(n18346) );
  AOI21_X1 U21535 ( .B1(n18349), .B2(P3_EAX_REG_21__SCAN_IN), .A(n18344), .ZN(
        n18345) );
  OAI211_X1 U21536 ( .C1(n19130), .C2(n18374), .A(n18346), .B(n18345), .ZN(
        P3_U2714) );
  INV_X1 U21537 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18454) );
  NOR2_X1 U21538 ( .A1(n18454), .A2(n18363), .ZN(n18357) );
  NAND2_X1 U21539 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18357), .ZN(n18353) );
  INV_X1 U21540 ( .A(n18347), .ZN(n18348) );
  AOI22_X1 U21541 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18362), .B1(n18382), .B2(
        n18348), .ZN(n18351) );
  AOI22_X1 U21542 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18368), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n18349), .ZN(n18350) );
  OAI211_X1 U21543 ( .C1(n18352), .C2(n18353), .A(n18351), .B(n18350), .ZN(
        P3_U2715) );
  AOI22_X1 U21544 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18362), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18368), .ZN(n18355) );
  OAI211_X1 U21545 ( .C1(n18357), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18425), .B(
        n18353), .ZN(n18354) );
  OAI211_X1 U21546 ( .C1(n18356), .C2(n18427), .A(n18355), .B(n18354), .ZN(
        P3_U2716) );
  AOI22_X1 U21547 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18362), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18368), .ZN(n18360) );
  AOI211_X1 U21548 ( .C1(n18454), .C2(n18363), .A(n18357), .B(n18370), .ZN(
        n18358) );
  INV_X1 U21549 ( .A(n18358), .ZN(n18359) );
  OAI211_X1 U21550 ( .C1(n18361), .C2(n18427), .A(n18360), .B(n18359), .ZN(
        P3_U2717) );
  AOI22_X1 U21551 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18362), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18368), .ZN(n18365) );
  OAI211_X1 U21552 ( .C1(n18369), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18425), .B(
        n18363), .ZN(n18364) );
  OAI211_X1 U21553 ( .C1(n18366), .C2(n18427), .A(n18365), .B(n18364), .ZN(
        P3_U2718) );
  AOI22_X1 U21554 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n18368), .B1(n18382), .B2(
        n18367), .ZN(n18373) );
  AOI211_X1 U21555 ( .C1(n18458), .C2(n18375), .A(n18370), .B(n18369), .ZN(
        n18371) );
  INV_X1 U21556 ( .A(n18371), .ZN(n18372) );
  OAI211_X1 U21557 ( .C1(n18374), .C2(n19105), .A(n18373), .B(n18372), .ZN(
        P3_U2719) );
  OAI211_X1 U21558 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n18383), .A(n18425), .B(
        n18375), .ZN(n18377) );
  NAND2_X1 U21559 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18398), .ZN(n18376) );
  OAI211_X1 U21560 ( .C1(n18378), .C2(n18427), .A(n18377), .B(n18376), .ZN(
        P3_U2720) );
  INV_X1 U21561 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18465) );
  INV_X1 U21562 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18471) );
  INV_X1 U21563 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18475) );
  NAND2_X1 U21564 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18420), .ZN(n18410) );
  NAND2_X1 U21565 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18413), .ZN(n18403) );
  NOR2_X2 U21566 ( .A1(n18471), .A2(n18403), .ZN(n18406) );
  NAND3_X1 U21567 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(n18406), .ZN(n18391) );
  NAND2_X1 U21568 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18394), .ZN(n18387) );
  AOI22_X1 U21569 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18398), .B1(n18382), .B2(
        n18381), .ZN(n18386) );
  INV_X1 U21570 ( .A(n18383), .ZN(n18384) );
  NAND3_X1 U21571 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18425), .A3(n18384), 
        .ZN(n18385) );
  OAI211_X1 U21572 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n18387), .A(n18386), .B(
        n18385), .ZN(P3_U2721) );
  INV_X1 U21573 ( .A(n18387), .ZN(n18390) );
  AOI21_X1 U21574 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18425), .A(n18394), .ZN(
        n18389) );
  OAI222_X1 U21575 ( .A1(n18430), .A2(n14014), .B1(n18390), .B2(n18389), .C1(
        n18427), .C2(n18388), .ZN(P3_U2722) );
  INV_X1 U21576 ( .A(n18391), .ZN(n18397) );
  AOI21_X1 U21577 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18425), .A(n18397), .ZN(
        n18393) );
  OAI222_X1 U21578 ( .A1(n18430), .A2(n14024), .B1(n18394), .B2(n18393), .C1(
        n18427), .C2(n18392), .ZN(P3_U2723) );
  AOI22_X1 U21579 ( .A1(n18406), .A2(P3_EAX_REG_10__SCAN_IN), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n18425), .ZN(n18396) );
  OAI222_X1 U21580 ( .A1(n18430), .A2(n14034), .B1(n18397), .B2(n18396), .C1(
        n18427), .C2(n18395), .ZN(P3_U2724) );
  NAND2_X1 U21581 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18398), .ZN(n18401) );
  NAND2_X1 U21582 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18406), .ZN(n18399) );
  OAI211_X1 U21583 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n18406), .A(n18425), .B(
        n18399), .ZN(n18400) );
  OAI211_X1 U21584 ( .C1(n18402), .C2(n18427), .A(n18401), .B(n18400), .ZN(
        P3_U2725) );
  INV_X1 U21585 ( .A(n18403), .ZN(n18409) );
  AOI21_X1 U21586 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18425), .A(n18409), .ZN(
        n18405) );
  OAI222_X1 U21587 ( .A1(n18430), .A2(n14028), .B1(n18406), .B2(n18405), .C1(
        n18427), .C2(n18404), .ZN(P3_U2726) );
  AOI21_X1 U21588 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n18425), .A(n18413), .ZN(
        n18408) );
  OAI222_X1 U21589 ( .A1(n18430), .A2(n14031), .B1(n18409), .B2(n18408), .C1(
        n18427), .C2(n18407), .ZN(P3_U2727) );
  INV_X1 U21590 ( .A(n18410), .ZN(n18416) );
  AOI21_X1 U21591 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18425), .A(n18416), .ZN(
        n18412) );
  OAI222_X1 U21592 ( .A1(n18430), .A2(n14047), .B1(n18413), .B2(n18412), .C1(
        n18427), .C2(n18411), .ZN(P3_U2728) );
  AOI21_X1 U21593 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18425), .A(n18420), .ZN(
        n18415) );
  OAI222_X1 U21594 ( .A1(n14001), .A2(n18430), .B1(n18416), .B2(n18415), .C1(
        n18427), .C2(n18414), .ZN(P3_U2729) );
  INV_X1 U21595 ( .A(n18417), .ZN(n18423) );
  AOI21_X1 U21596 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18425), .A(n18423), .ZN(
        n18419) );
  OAI222_X1 U21597 ( .A1(n19130), .A2(n18430), .B1(n18420), .B2(n18419), .C1(
        n18427), .C2(n18418), .ZN(P3_U2730) );
  INV_X1 U21598 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19126) );
  AOI21_X1 U21599 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18425), .A(n18429), .ZN(
        n18422) );
  OAI222_X1 U21600 ( .A1(n19126), .A2(n18430), .B1(n18423), .B2(n18422), .C1(
        n18427), .C2(n18421), .ZN(P3_U2731) );
  AOI21_X1 U21601 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18425), .A(n18424), .ZN(
        n18428) );
  OAI222_X1 U21602 ( .A1(n19121), .A2(n18430), .B1(n18429), .B2(n18428), .C1(
        n18427), .C2(n18426), .ZN(P3_U2732) );
  NOR2_X4 U21603 ( .A1(n18488), .A2(n18460), .ZN(n18476) );
  AND2_X1 U21604 ( .A1(n18476), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AOI22_X1 U21605 ( .A1(n18488), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18433) );
  OAI21_X1 U21606 ( .B1(n18512), .B2(n18457), .A(n18433), .ZN(P3_U2737) );
  AOI22_X1 U21607 ( .A1(n18488), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18434) );
  OAI21_X1 U21608 ( .B1(n10299), .B2(n18457), .A(n18434), .ZN(P3_U2738) );
  INV_X1 U21609 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18436) );
  AOI22_X1 U21610 ( .A1(n18488), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18435) );
  OAI21_X1 U21611 ( .B1(n18436), .B2(n18457), .A(n18435), .ZN(P3_U2739) );
  AOI22_X1 U21612 ( .A1(n18488), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18437) );
  OAI21_X1 U21613 ( .B1(n18438), .B2(n18457), .A(n18437), .ZN(P3_U2740) );
  AOI22_X1 U21614 ( .A1(n18488), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18439) );
  OAI21_X1 U21615 ( .B1(n10306), .B2(n18457), .A(n18439), .ZN(P3_U2741) );
  AOI22_X1 U21616 ( .A1(n18488), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18440) );
  OAI21_X1 U21617 ( .B1(n18441), .B2(n18457), .A(n18440), .ZN(P3_U2742) );
  AOI22_X1 U21618 ( .A1(n18488), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18442) );
  OAI21_X1 U21619 ( .B1(n18443), .B2(n18457), .A(n18442), .ZN(P3_U2743) );
  AOI22_X1 U21620 ( .A1(n18488), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18444) );
  OAI21_X1 U21621 ( .B1(n18445), .B2(n18457), .A(n18444), .ZN(P3_U2744) );
  AOI22_X1 U21622 ( .A1(n18488), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18446) );
  OAI21_X1 U21623 ( .B1(n18447), .B2(n18457), .A(n18446), .ZN(P3_U2745) );
  AOI22_X1 U21624 ( .A1(n18488), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18448) );
  OAI21_X1 U21625 ( .B1(n21491), .B2(n18457), .A(n18448), .ZN(P3_U2746) );
  INV_X1 U21626 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18450) );
  AOI22_X1 U21627 ( .A1(n18488), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18449) );
  OAI21_X1 U21628 ( .B1(n18450), .B2(n18457), .A(n18449), .ZN(P3_U2747) );
  INV_X1 U21629 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18452) );
  AOI22_X1 U21630 ( .A1(n18488), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18451) );
  OAI21_X1 U21631 ( .B1(n18452), .B2(n18457), .A(n18451), .ZN(P3_U2748) );
  AOI22_X1 U21632 ( .A1(n18488), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18453) );
  OAI21_X1 U21633 ( .B1(n18454), .B2(n18457), .A(n18453), .ZN(P3_U2749) );
  AOI22_X1 U21634 ( .A1(n18488), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18455) );
  OAI21_X1 U21635 ( .B1(n18497), .B2(n18457), .A(n18455), .ZN(P3_U2750) );
  AOI22_X1 U21636 ( .A1(n18488), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18456) );
  OAI21_X1 U21637 ( .B1(n18458), .B2(n18457), .A(n18456), .ZN(P3_U2751) );
  INV_X1 U21638 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18537) );
  AOI22_X1 U21639 ( .A1(n18488), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18459) );
  OAI21_X1 U21640 ( .B1(n18537), .B2(n18490), .A(n18459), .ZN(P3_U2752) );
  INV_X1 U21641 ( .A(P3_LWORD_REG_14__SCAN_IN), .ZN(n21453) );
  AOI22_X1 U21642 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18460), .B1(n18476), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18461) );
  OAI21_X1 U21643 ( .B1(n21453), .B2(n19704), .A(n18461), .ZN(P3_U2753) );
  INV_X1 U21644 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18463) );
  AOI22_X1 U21645 ( .A1(n18488), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18462) );
  OAI21_X1 U21646 ( .B1(n18463), .B2(n18490), .A(n18462), .ZN(P3_U2754) );
  AOI22_X1 U21647 ( .A1(n18488), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18464) );
  OAI21_X1 U21648 ( .B1(n18465), .B2(n18490), .A(n18464), .ZN(P3_U2755) );
  INV_X1 U21649 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18467) );
  AOI22_X1 U21650 ( .A1(n18488), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18466) );
  OAI21_X1 U21651 ( .B1(n18467), .B2(n18490), .A(n18466), .ZN(P3_U2756) );
  INV_X1 U21652 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18469) );
  AOI22_X1 U21653 ( .A1(n18488), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18468) );
  OAI21_X1 U21654 ( .B1(n18469), .B2(n18490), .A(n18468), .ZN(P3_U2757) );
  AOI22_X1 U21655 ( .A1(n18488), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18470) );
  OAI21_X1 U21656 ( .B1(n18471), .B2(n18490), .A(n18470), .ZN(P3_U2758) );
  INV_X1 U21657 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18473) );
  AOI22_X1 U21658 ( .A1(n18488), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18472) );
  OAI21_X1 U21659 ( .B1(n18473), .B2(n18490), .A(n18472), .ZN(P3_U2759) );
  AOI22_X1 U21660 ( .A1(n18488), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18474) );
  OAI21_X1 U21661 ( .B1(n18475), .B2(n18490), .A(n18474), .ZN(P3_U2760) );
  INV_X1 U21662 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18478) );
  AOI22_X1 U21663 ( .A1(n18488), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18477) );
  OAI21_X1 U21664 ( .B1(n18478), .B2(n18490), .A(n18477), .ZN(P3_U2761) );
  AOI22_X1 U21665 ( .A1(n18488), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18479) );
  OAI21_X1 U21666 ( .B1(n18480), .B2(n18490), .A(n18479), .ZN(P3_U2762) );
  INV_X1 U21667 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18482) );
  AOI22_X1 U21668 ( .A1(n18488), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18481) );
  OAI21_X1 U21669 ( .B1(n18482), .B2(n18490), .A(n18481), .ZN(P3_U2763) );
  AOI22_X1 U21670 ( .A1(n18488), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18483) );
  OAI21_X1 U21671 ( .B1(n18484), .B2(n18490), .A(n18483), .ZN(P3_U2764) );
  AOI22_X1 U21672 ( .A1(n18488), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18485) );
  OAI21_X1 U21673 ( .B1(n18486), .B2(n18490), .A(n18485), .ZN(P3_U2765) );
  AOI22_X1 U21674 ( .A1(n18488), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18487) );
  OAI21_X1 U21675 ( .B1(n18515), .B2(n18490), .A(n18487), .ZN(P3_U2766) );
  AOI22_X1 U21676 ( .A1(n18488), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18476), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18489) );
  OAI21_X1 U21677 ( .B1(n18491), .B2(n18490), .A(n18489), .ZN(P3_U2767) );
  AOI22_X1 U21678 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18530), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18533), .ZN(n18495) );
  OAI21_X1 U21679 ( .B1(n19105), .B2(n18529), .A(n18495), .ZN(P3_U2768) );
  AOI22_X1 U21680 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18534), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18533), .ZN(n18496) );
  OAI21_X1 U21681 ( .B1(n18497), .B2(n18536), .A(n18496), .ZN(P3_U2769) );
  AOI22_X1 U21682 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18530), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18533), .ZN(n18498) );
  OAI21_X1 U21683 ( .B1(n19116), .B2(n18529), .A(n18498), .ZN(P3_U2770) );
  AOI22_X1 U21684 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18530), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18533), .ZN(n18499) );
  OAI21_X1 U21685 ( .B1(n19121), .B2(n18529), .A(n18499), .ZN(P3_U2771) );
  AOI22_X1 U21686 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18530), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18533), .ZN(n18500) );
  OAI21_X1 U21687 ( .B1(n19126), .B2(n18529), .A(n18500), .ZN(P3_U2772) );
  AOI22_X1 U21688 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18530), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18533), .ZN(n18501) );
  OAI21_X1 U21689 ( .B1(n19130), .B2(n18529), .A(n18501), .ZN(P3_U2773) );
  AOI22_X1 U21690 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18530), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18533), .ZN(n18502) );
  OAI21_X1 U21691 ( .B1(n14001), .B2(n18529), .A(n18502), .ZN(P3_U2774) );
  AOI22_X1 U21692 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18508), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18533), .ZN(n18503) );
  OAI21_X1 U21693 ( .B1(n14047), .B2(n18529), .A(n18503), .ZN(P3_U2775) );
  AOI22_X1 U21694 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18508), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18533), .ZN(n18504) );
  OAI21_X1 U21695 ( .B1(n14031), .B2(n18529), .A(n18504), .ZN(P3_U2776) );
  AOI22_X1 U21696 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18508), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18533), .ZN(n18505) );
  OAI21_X1 U21697 ( .B1(n14028), .B2(n18529), .A(n18505), .ZN(P3_U2777) );
  AOI22_X1 U21698 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18508), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18533), .ZN(n18506) );
  OAI21_X1 U21699 ( .B1(n18525), .B2(n18529), .A(n18506), .ZN(P3_U2778) );
  AOI22_X1 U21700 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n18508), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18533), .ZN(n18507) );
  OAI21_X1 U21701 ( .B1(n14034), .B2(n18529), .A(n18507), .ZN(P3_U2779) );
  AOI22_X1 U21702 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18508), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18533), .ZN(n18509) );
  OAI21_X1 U21703 ( .B1(n14024), .B2(n18529), .A(n18509), .ZN(P3_U2780) );
  AOI22_X1 U21704 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18530), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18533), .ZN(n18510) );
  OAI21_X1 U21705 ( .B1(n14014), .B2(n18529), .A(n18510), .ZN(P3_U2781) );
  AOI22_X1 U21706 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18534), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18533), .ZN(n18511) );
  OAI21_X1 U21707 ( .B1(n18512), .B2(n18536), .A(n18511), .ZN(P3_U2782) );
  AOI22_X1 U21708 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18533), .ZN(n18513) );
  OAI21_X1 U21709 ( .B1(n19105), .B2(n18529), .A(n18513), .ZN(P3_U2783) );
  AOI22_X1 U21710 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18534), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18533), .ZN(n18514) );
  OAI21_X1 U21711 ( .B1(n18515), .B2(n18536), .A(n18514), .ZN(P3_U2784) );
  AOI22_X1 U21712 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18533), .ZN(n18516) );
  OAI21_X1 U21713 ( .B1(n19116), .B2(n18529), .A(n18516), .ZN(P3_U2785) );
  AOI22_X1 U21714 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18533), .ZN(n18517) );
  OAI21_X1 U21715 ( .B1(n19121), .B2(n18529), .A(n18517), .ZN(P3_U2786) );
  AOI22_X1 U21716 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18533), .ZN(n18518) );
  OAI21_X1 U21717 ( .B1(n19126), .B2(n18529), .A(n18518), .ZN(P3_U2787) );
  AOI22_X1 U21718 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18533), .ZN(n18519) );
  OAI21_X1 U21719 ( .B1(n19130), .B2(n18529), .A(n18519), .ZN(P3_U2788) );
  AOI22_X1 U21720 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18533), .ZN(n18520) );
  OAI21_X1 U21721 ( .B1(n14001), .B2(n18529), .A(n18520), .ZN(P3_U2789) );
  AOI22_X1 U21722 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18533), .ZN(n18521) );
  OAI21_X1 U21723 ( .B1(n14047), .B2(n18529), .A(n18521), .ZN(P3_U2790) );
  AOI22_X1 U21724 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18533), .ZN(n18522) );
  OAI21_X1 U21725 ( .B1(n14031), .B2(n18529), .A(n18522), .ZN(P3_U2791) );
  AOI22_X1 U21726 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18533), .ZN(n18523) );
  OAI21_X1 U21727 ( .B1(n14028), .B2(n18529), .A(n18523), .ZN(P3_U2792) );
  AOI22_X1 U21728 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18533), .ZN(n18524) );
  OAI21_X1 U21729 ( .B1(n18525), .B2(n18529), .A(n18524), .ZN(P3_U2793) );
  AOI22_X1 U21730 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18533), .ZN(n18526) );
  OAI21_X1 U21731 ( .B1(n14034), .B2(n18529), .A(n18526), .ZN(P3_U2794) );
  AOI22_X1 U21732 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18533), .ZN(n18527) );
  OAI21_X1 U21733 ( .B1(n14024), .B2(n18529), .A(n18527), .ZN(P3_U2795) );
  AOI22_X1 U21734 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18530), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18533), .ZN(n18528) );
  OAI21_X1 U21735 ( .B1(n14014), .B2(n18529), .A(n18528), .ZN(P3_U2796) );
  AOI22_X1 U21736 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18534), .B1(
        P3_EAX_REG_14__SCAN_IN), .B2(n18530), .ZN(n18531) );
  OAI21_X1 U21737 ( .B1(n18532), .B2(n21453), .A(n18531), .ZN(P3_U2797) );
  AOI22_X1 U21738 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18534), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18533), .ZN(n18535) );
  OAI21_X1 U21739 ( .B1(n18537), .B2(n18536), .A(n18535), .ZN(P3_U2798) );
  AOI22_X1 U21740 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18539), .B1(
        n18675), .B2(n18538), .ZN(n18549) );
  NOR2_X1 U21741 ( .A1(n10448), .A2(n18541), .ZN(n18542) );
  XNOR2_X1 U21742 ( .A(n18542), .B(n18694), .ZN(n18827) );
  AOI22_X1 U21743 ( .A1(n18728), .A2(n18827), .B1(n18544), .B2(n18543), .ZN(
        n18548) );
  OAI21_X1 U21744 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18546), .A(
        n18545), .ZN(n18547) );
  NAND2_X1 U21745 ( .A1(n18905), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18828) );
  NAND4_X1 U21746 ( .A1(n18549), .A2(n18548), .A3(n18547), .A4(n18828), .ZN(
        P3_U2803) );
  XOR2_X1 U21747 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18550), .Z(
        n18836) );
  AND2_X1 U21748 ( .A1(n11501), .A2(n16915), .ZN(n18580) );
  AOI211_X1 U21749 ( .C1(n18552), .C2(n18551), .A(n18769), .B(n18580), .ZN(
        n18584) );
  OAI21_X1 U21750 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18595), .A(
        n18584), .ZN(n18567) );
  NOR2_X1 U21751 ( .A1(n18598), .A2(n11501), .ZN(n18569) );
  OAI211_X1 U21752 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18569), .B(n18553), .ZN(n18554) );
  NAND2_X1 U21753 ( .A1(n18905), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18842) );
  OAI211_X1 U21754 ( .C1(n18686), .C2(n18555), .A(n18554), .B(n18842), .ZN(
        n18556) );
  AOI21_X1 U21755 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18567), .A(
        n18556), .ZN(n18563) );
  XOR2_X1 U21756 ( .A(n18557), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18832) );
  INV_X1 U21757 ( .A(n18558), .ZN(n18559) );
  NAND2_X1 U21758 ( .A1(n18560), .A2(n18559), .ZN(n18561) );
  XNOR2_X1 U21759 ( .A(n18561), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18831) );
  AOI22_X1 U21760 ( .A1(n18780), .A2(n18832), .B1(n18728), .B2(n18831), .ZN(
        n18562) );
  OAI211_X1 U21761 ( .C1(n18602), .C2(n18836), .A(n18563), .B(n18562), .ZN(
        P3_U2805) );
  AOI22_X1 U21762 ( .A1(n18780), .A2(n18845), .B1(n18716), .B2(n18844), .ZN(
        n18587) );
  AOI22_X1 U21763 ( .A1(n18905), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18675), 
        .B2(n18564), .ZN(n18565) );
  INV_X1 U21764 ( .A(n18565), .ZN(n18566) );
  AOI221_X1 U21765 ( .B1(n18569), .B2(n18568), .C1(n18567), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18566), .ZN(n18574) );
  OAI21_X1 U21766 ( .B1(n9748), .B2(n18854), .A(n18570), .ZN(n18851) );
  NOR3_X1 U21767 ( .A1(n18684), .A2(n18571), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18572) );
  AOI21_X1 U21768 ( .B1(n18728), .B2(n18851), .A(n18572), .ZN(n18573) );
  OAI211_X1 U21769 ( .C1(n18587), .C2(n18854), .A(n18574), .B(n18573), .ZN(
        P3_U2806) );
  INV_X1 U21770 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18623) );
  AND2_X1 U21771 ( .A1(n18618), .A2(n18623), .ZN(n18590) );
  NAND2_X1 U21772 ( .A1(n18575), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18576) );
  OAI211_X1 U21773 ( .C1(n18577), .C2(n18590), .A(n18625), .B(n18576), .ZN(
        n18578) );
  XNOR2_X1 U21774 ( .A(n18578), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18860) );
  AOI22_X1 U21775 ( .A1(n18581), .A2(n18580), .B1(n18579), .B2(n18808), .ZN(
        n18582) );
  NAND2_X1 U21776 ( .A1(n18905), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18861) );
  OAI211_X1 U21777 ( .C1(n18584), .C2(n18583), .A(n18582), .B(n18861), .ZN(
        n18585) );
  AOI21_X1 U21778 ( .B1(n18728), .B2(n18860), .A(n18585), .ZN(n18586) );
  OAI221_X1 U21779 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18588), 
        .C1(n18856), .C2(n18587), .A(n18586), .ZN(P3_U2807) );
  INV_X1 U21780 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18589) );
  NOR3_X1 U21781 ( .A1(n18617), .A2(n18875), .A3(n18589), .ZN(n18591) );
  OAI21_X1 U21782 ( .B1(n18591), .B2(n18590), .A(n18625), .ZN(n18592) );
  XOR2_X1 U21783 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18592), .Z(
        n18882) );
  OAI21_X1 U21784 ( .B1(n18593), .B2(n18672), .A(n18810), .ZN(n18594) );
  AOI21_X1 U21785 ( .B1(n18790), .B2(n18597), .A(n18594), .ZN(n18632) );
  OAI21_X1 U21786 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18595), .A(
        n18632), .ZN(n18611) );
  INV_X1 U21787 ( .A(n18596), .ZN(n18601) );
  NAND2_X1 U21788 ( .A1(n18905), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18880) );
  NOR2_X1 U21789 ( .A1(n18598), .A2(n18597), .ZN(n18613) );
  OAI211_X1 U21790 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18613), .B(n18599), .ZN(n18600) );
  OAI211_X1 U21791 ( .C1(n18601), .C2(n18686), .A(n18880), .B(n18600), .ZN(
        n18607) );
  NOR2_X1 U21792 ( .A1(n18875), .A2(n18620), .ZN(n18873) );
  INV_X1 U21793 ( .A(n18873), .ZN(n18603) );
  NOR2_X1 U21794 ( .A1(n18684), .A2(n18603), .ZN(n18605) );
  NAND2_X1 U21795 ( .A1(n18813), .A2(n18602), .ZN(n18634) );
  AOI21_X1 U21796 ( .B1(n18634), .B2(n18603), .A(n18633), .ZN(n18624) );
  INV_X1 U21797 ( .A(n18624), .ZN(n18604) );
  MUX2_X1 U21798 ( .A(n18605), .B(n18604), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n18606) );
  AOI211_X1 U21799 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n18611), .A(
        n18607), .B(n18606), .ZN(n18608) );
  OAI21_X1 U21800 ( .B1(n18641), .B2(n18882), .A(n18608), .ZN(P3_U2808) );
  INV_X1 U21801 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18612) );
  OAI22_X1 U21802 ( .A1(n18992), .A2(n19658), .B1(n18686), .B2(n18609), .ZN(
        n18610) );
  AOI221_X1 U21803 ( .B1(n18613), .B2(n18612), .C1(n18611), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18610), .ZN(n18622) );
  INV_X1 U21804 ( .A(n18614), .ZN(n18650) );
  INV_X1 U21805 ( .A(n18615), .ZN(n18616) );
  NOR2_X1 U21806 ( .A1(n18617), .A2(n18616), .ZN(n18648) );
  AOI22_X1 U21807 ( .A1(n18650), .A2(n18618), .B1(n18884), .B2(n18648), .ZN(
        n18619) );
  XNOR2_X1 U21808 ( .A(n18619), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18889) );
  AND2_X1 U21809 ( .A1(n18623), .A2(n18884), .ZN(n18887) );
  NOR2_X1 U21810 ( .A1(n18684), .A2(n18620), .ZN(n18652) );
  AOI22_X1 U21811 ( .A1(n18728), .A2(n18889), .B1(n18887), .B2(n18652), .ZN(
        n18621) );
  OAI211_X1 U21812 ( .C1(n18624), .C2(n18623), .A(n18622), .B(n18621), .ZN(
        P3_U2809) );
  INV_X1 U21813 ( .A(n18625), .ZN(n18627) );
  OAI22_X1 U21814 ( .A1(n18648), .A2(n18895), .B1(n18649), .B2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18626) );
  NOR2_X1 U21815 ( .A1(n18627), .A2(n18626), .ZN(n18628) );
  XOR2_X1 U21816 ( .A(n18629), .B(n18628), .Z(n18899) );
  AOI21_X1 U21817 ( .B1(n16915), .B2(n18630), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18631) );
  NAND2_X1 U21818 ( .A1(n18905), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18898) );
  OAI21_X1 U21819 ( .B1(n18632), .B2(n18631), .A(n18898), .ZN(n18638) );
  NAND2_X1 U21820 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18872), .ZN(
        n18865) );
  NOR2_X1 U21821 ( .A1(n18684), .A2(n18865), .ZN(n18636) );
  AOI21_X1 U21822 ( .B1(n18634), .B2(n18865), .A(n18633), .ZN(n18655) );
  INV_X1 U21823 ( .A(n18655), .ZN(n18635) );
  MUX2_X1 U21824 ( .A(n18636), .B(n18635), .S(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n18637) );
  AOI211_X1 U21825 ( .C1(n18639), .C2(n18808), .A(n18638), .B(n18637), .ZN(
        n18640) );
  OAI21_X1 U21826 ( .B1(n18641), .B2(n18899), .A(n18640), .ZN(P3_U2810) );
  OAI211_X1 U21827 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18643), .B(n18642), .ZN(n18644) );
  NAND2_X1 U21828 ( .A1(n18905), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18902) );
  OAI211_X1 U21829 ( .C1(n18686), .C2(n18645), .A(n18644), .B(n18902), .ZN(
        n18646) );
  AOI21_X1 U21830 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18647), .A(
        n18646), .ZN(n18654) );
  AOI21_X1 U21831 ( .B1(n18650), .B2(n18649), .A(n18648), .ZN(n18651) );
  XOR2_X1 U21832 ( .A(n18895), .B(n18651), .Z(n18900) );
  AOI22_X1 U21833 ( .A1(n18728), .A2(n18900), .B1(n18652), .B2(n18895), .ZN(
        n18653) );
  OAI211_X1 U21834 ( .C1(n18655), .C2(n18895), .A(n18654), .B(n18653), .ZN(
        P3_U2811) );
  AOI21_X1 U21835 ( .B1(n18656), .B2(n16915), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18657) );
  OR2_X1 U21836 ( .A1(n18658), .A2(n18657), .ZN(n18661) );
  XNOR2_X1 U21837 ( .A(n18659), .B(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18906) );
  NAND2_X1 U21838 ( .A1(n18906), .A2(n18728), .ZN(n18660) );
  OAI211_X1 U21839 ( .C1(n19650), .C2(n18988), .A(n18661), .B(n18660), .ZN(
        n18662) );
  INV_X1 U21840 ( .A(n18662), .ZN(n18666) );
  OAI221_X1 U21841 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18664), .A(n18663), .ZN(
        n18665) );
  OAI211_X1 U21842 ( .C1(n18822), .C2(n18667), .A(n18666), .B(n18665), .ZN(
        P3_U2813) );
  OAI22_X1 U21843 ( .A1(n18669), .A2(n18694), .B1(n18708), .B2(n18668), .ZN(
        n18670) );
  XOR2_X1 U21844 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n18670), .Z(
        n18922) );
  AOI21_X1 U21845 ( .B1(n18790), .B2(n18671), .A(n18769), .ZN(n18706) );
  OAI21_X1 U21846 ( .B1(n18673), .B2(n18672), .A(n18706), .ZN(n18688) );
  AOI22_X1 U21847 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18688), .B1(
        n18675), .B2(n18674), .ZN(n18680) );
  NAND2_X1 U21848 ( .A1(n18703), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18677) );
  NOR2_X1 U21849 ( .A1(n18677), .A2(n18676), .ZN(n18690) );
  OAI211_X1 U21850 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18690), .B(n18678), .ZN(n18679) );
  OAI211_X1 U21851 ( .C1(n19648), .C2(n18992), .A(n18680), .B(n18679), .ZN(
        n18681) );
  AOI21_X1 U21852 ( .B1(n18728), .B2(n18922), .A(n18681), .ZN(n18682) );
  OAI221_X1 U21853 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18684), 
        .C1(n10082), .C2(n18683), .A(n18682), .ZN(P3_U2814) );
  NOR2_X1 U21854 ( .A1(n13637), .A2(n18917), .ZN(n18714) );
  NOR2_X1 U21855 ( .A1(n18714), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18931) );
  INV_X1 U21856 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18689) );
  OAI22_X1 U21857 ( .A1(n18992), .A2(n19646), .B1(n18686), .B2(n18685), .ZN(
        n18687) );
  AOI221_X1 U21858 ( .B1(n18690), .B2(n18689), .C1(n18688), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18687), .ZN(n18698) );
  NAND3_X1 U21859 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n18977), .ZN(n18692) );
  OAI22_X1 U21860 ( .A1(n18710), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n18692), .B2(n18691), .ZN(n18693) );
  OAI221_X1 U21861 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n10228), 
        .C1(n18969), .C2(n18694), .A(n18693), .ZN(n18695) );
  XOR2_X1 U21862 ( .A(n18912), .B(n18695), .Z(n18932) );
  NOR2_X1 U21863 ( .A1(n18937), .A2(n18813), .ZN(n18696) );
  NAND2_X1 U21864 ( .A1(n18700), .A2(n18912), .ZN(n18925) );
  AOI22_X1 U21865 ( .A1(n18728), .A2(n18932), .B1(n18696), .B2(n18925), .ZN(
        n18697) );
  OAI211_X1 U21866 ( .C1(n18931), .C2(n18699), .A(n18698), .B(n18697), .ZN(
        P3_U2815) );
  OAI21_X1 U21867 ( .B1(n18701), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18700), .ZN(n18950) );
  AOI21_X1 U21868 ( .B1(n18703), .B2(n18702), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18705) );
  OAI22_X1 U21869 ( .A1(n18706), .A2(n18705), .B1(n18822), .B2(n18704), .ZN(
        n18707) );
  AOI21_X1 U21870 ( .B1(n18905), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18707), 
        .ZN(n18718) );
  NAND2_X1 U21871 ( .A1(n18969), .A2(n18940), .ZN(n18709) );
  OAI22_X1 U21872 ( .A1(n18710), .A2(n18709), .B1(n18927), .B2(n18708), .ZN(
        n18711) );
  XOR2_X1 U21873 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18711), .Z(
        n18946) );
  AOI21_X1 U21874 ( .B1(n18713), .B2(n18712), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18715) );
  NOR2_X1 U21875 ( .A1(n18715), .A2(n18714), .ZN(n18942) );
  AOI22_X1 U21876 ( .A1(n18946), .A2(n18728), .B1(n18716), .B2(n18942), .ZN(
        n18717) );
  OAI211_X1 U21877 ( .C1(n18813), .C2(n18950), .A(n18718), .B(n18717), .ZN(
        P3_U2816) );
  INV_X1 U21878 ( .A(n18719), .ZN(n18720) );
  AOI22_X1 U21879 ( .A1(n18905), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18720), 
        .B2(n18808), .ZN(n18733) );
  AOI21_X1 U21880 ( .B1(n18722), .B2(n19000), .A(n18721), .ZN(n18723) );
  XOR2_X1 U21881 ( .A(n18724), .B(n18723), .Z(n18986) );
  OAI21_X1 U21882 ( .B1(n18725), .B2(n19000), .A(n18724), .ZN(n18726) );
  AOI22_X1 U21883 ( .A1(n18728), .A2(n18986), .B1(n18727), .B2(n18726), .ZN(
        n18732) );
  INV_X1 U21884 ( .A(n18820), .ZN(n18761) );
  OAI211_X1 U21885 ( .C1(n18730), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18761), .B(n18729), .ZN(n18731) );
  NAND3_X1 U21886 ( .A1(n18733), .A2(n18732), .A3(n18731), .ZN(P3_U2820) );
  NOR2_X1 U21887 ( .A1(n18992), .A2(n19630), .ZN(n19023) );
  AOI221_X1 U21888 ( .B1(n18754), .B2(n18735), .C1(n18734), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n19023), .ZN(n18744) );
  AOI21_X1 U21889 ( .B1(n18738), .B2(n18737), .A(n18736), .ZN(n18739) );
  XOR2_X1 U21890 ( .A(n18739), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n19025) );
  INV_X1 U21891 ( .A(n18817), .ZN(n18796) );
  OAI21_X1 U21892 ( .B1(n18741), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18740), .ZN(n18742) );
  INV_X1 U21893 ( .A(n18742), .ZN(n19024) );
  AOI22_X1 U21894 ( .A1(n18780), .A2(n19025), .B1(n18796), .B2(n19024), .ZN(
        n18743) );
  OAI211_X1 U21895 ( .C1(n18822), .C2(n18745), .A(n18744), .B(n18743), .ZN(
        P3_U2823) );
  OAI21_X1 U21896 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18747), .A(
        n18746), .ZN(n19031) );
  OR2_X1 U21897 ( .A1(n18749), .A2(n18748), .ZN(n18750) );
  AND2_X1 U21898 ( .A1(n18751), .A2(n18750), .ZN(n19033) );
  NOR2_X1 U21899 ( .A1(n19206), .A2(n17020), .ZN(n18765) );
  AOI21_X1 U21900 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18761), .A(
        n18765), .ZN(n18753) );
  OAI22_X1 U21901 ( .A1(n18754), .A2(n18753), .B1(n18822), .B2(n18752), .ZN(
        n18755) );
  AOI21_X1 U21902 ( .B1(n18796), .B2(n19033), .A(n18755), .ZN(n18756) );
  NAND2_X1 U21903 ( .A1(n18905), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n19039) );
  OAI211_X1 U21904 ( .C1(n18813), .C2(n19031), .A(n18756), .B(n19039), .ZN(
        P3_U2824) );
  OAI21_X1 U21905 ( .B1(n18759), .B2(n18758), .A(n18757), .ZN(n19051) );
  XNOR2_X1 U21906 ( .A(n18760), .B(n10273), .ZN(n19046) );
  NAND2_X1 U21907 ( .A1(n18905), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n19049) );
  INV_X1 U21908 ( .A(n19049), .ZN(n18767) );
  OAI221_X1 U21909 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18762), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18810), .A(n18761), .ZN(n18764) );
  OAI22_X1 U21910 ( .A1(n18765), .A2(n18764), .B1(n18822), .B2(n18763), .ZN(
        n18766) );
  AOI211_X1 U21911 ( .C1(n18796), .C2(n19046), .A(n18767), .B(n18766), .ZN(
        n18768) );
  OAI21_X1 U21912 ( .B1(n18813), .B2(n19051), .A(n18768), .ZN(P3_U2825) );
  AOI21_X1 U21913 ( .B1(n18790), .B2(n17866), .A(n18769), .ZN(n18789) );
  OAI21_X1 U21914 ( .B1(n18772), .B2(n18771), .A(n18770), .ZN(n18773) );
  INV_X1 U21915 ( .A(n18773), .ZN(n19053) );
  NOR3_X1 U21916 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17866), .A3(
        n19206), .ZN(n18774) );
  NOR2_X1 U21917 ( .A1(n18988), .A2(n19624), .ZN(n19052) );
  AOI211_X1 U21918 ( .C1(n18796), .C2(n19053), .A(n18774), .B(n19052), .ZN(
        n18782) );
  AOI21_X1 U21919 ( .B1(n18777), .B2(n18776), .A(n18775), .ZN(n18778) );
  XOR2_X1 U21920 ( .A(n18778), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n19056) );
  AOI22_X1 U21921 ( .A1(n18780), .A2(n19056), .B1(n18779), .B2(n18808), .ZN(
        n18781) );
  OAI211_X1 U21922 ( .C1(n18789), .C2(n18783), .A(n18782), .B(n18781), .ZN(
        P3_U2826) );
  OAI21_X1 U21923 ( .B1(n18786), .B2(n18785), .A(n18784), .ZN(n19073) );
  INV_X1 U21924 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18787) );
  XNOR2_X1 U21925 ( .A(n18788), .B(n18787), .ZN(n19065) );
  NOR2_X1 U21926 ( .A1(n18789), .A2(n21512), .ZN(n18795) );
  NAND2_X1 U21927 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18810), .ZN(
        n18792) );
  NAND2_X1 U21928 ( .A1(n18790), .A2(n17866), .ZN(n18791) );
  OAI22_X1 U21929 ( .A1(n18822), .A2(n18793), .B1(n18792), .B2(n18791), .ZN(
        n18794) );
  AOI211_X1 U21930 ( .C1(n18796), .C2(n19065), .A(n18795), .B(n18794), .ZN(
        n18798) );
  AND2_X1 U21931 ( .A1(n18905), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19064) );
  INV_X1 U21932 ( .A(n19064), .ZN(n18797) );
  OAI211_X1 U21933 ( .C1(n18813), .C2(n19073), .A(n18798), .B(n18797), .ZN(
        P3_U2827) );
  OAI21_X1 U21934 ( .B1(n18801), .B2(n18800), .A(n18799), .ZN(n19094) );
  NOR2_X1 U21935 ( .A1(n18813), .A2(n19094), .ZN(n18806) );
  OAI21_X1 U21936 ( .B1(n18804), .B2(n18803), .A(n18802), .ZN(n19084) );
  NAND2_X1 U21937 ( .A1(n18905), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n19087) );
  OAI21_X1 U21938 ( .B1(n18817), .B2(n19084), .A(n19087), .ZN(n18805) );
  AOI211_X1 U21939 ( .C1(n18808), .C2(n18807), .A(n18806), .B(n18805), .ZN(
        n18809) );
  OAI221_X1 U21940 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19206), .C1(
        n18811), .C2(n18810), .A(n18809), .ZN(P3_U2828) );
  OR2_X1 U21941 ( .A1(n18813), .A2(n18812), .ZN(n18815) );
  OAI211_X1 U21942 ( .C1(n18817), .C2(n18816), .A(n18815), .B(n18814), .ZN(
        n18818) );
  INV_X1 U21943 ( .A(n18818), .ZN(n18819) );
  OAI221_X1 U21944 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18822), .C1(
        n18821), .C2(n18820), .A(n18819), .ZN(P3_U2829) );
  AOI21_X1 U21945 ( .B1(n19062), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18823), .ZN(n18824) );
  AOI21_X1 U21946 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18825), .A(
        n18824), .ZN(n18826) );
  AOI21_X1 U21947 ( .B1(n18827), .B2(n18997), .A(n18826), .ZN(n18829) );
  OAI211_X1 U21948 ( .C1(n19090), .C2(n18830), .A(n18829), .B(n18828), .ZN(
        P3_U2835) );
  AOI22_X1 U21949 ( .A1(n19057), .A2(n18832), .B1(n18997), .B2(n18831), .ZN(
        n18843) );
  AOI211_X1 U21950 ( .C1(n18916), .C2(n18835), .A(n18834), .B(n18833), .ZN(
        n18837) );
  OAI22_X1 U21951 ( .A1(n18837), .A2(n10442), .B1(n18952), .B2(n18836), .ZN(
        n18839) );
  OAI221_X1 U21952 ( .B1(n18839), .B2(n18838), .C1(n18839), .C2(n10442), .A(
        n19062), .ZN(n18841) );
  NAND2_X1 U21953 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19066), .ZN(
        n18840) );
  NAND4_X1 U21954 ( .A1(n18843), .A2(n18842), .A3(n18841), .A4(n18840), .ZN(
        P3_U2837) );
  AOI22_X1 U21955 ( .A1(n18957), .A2(n18845), .B1(n18971), .B2(n18844), .ZN(
        n18846) );
  NAND3_X1 U21956 ( .A1(n18847), .A2(n18846), .A3(n19090), .ZN(n18850) );
  NOR3_X1 U21957 ( .A1(n18850), .A2(n18856), .A3(n18848), .ZN(n18849) );
  NOR2_X1 U21958 ( .A1(n18849), .A2(n18905), .ZN(n18859) );
  OAI21_X1 U21959 ( .B1(n19005), .B2(n18850), .A(n18859), .ZN(n18853) );
  AOI22_X1 U21960 ( .A1(n18851), .A2(n18997), .B1(n18905), .B2(
        P3_REIP_REG_24__SCAN_IN), .ZN(n18852) );
  OAI221_X1 U21961 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18855), 
        .C1(n18854), .C2(n18853), .A(n18852), .ZN(P3_U2838) );
  OAI21_X1 U21962 ( .B1(n19066), .B2(n18857), .A(n18856), .ZN(n18858) );
  AOI22_X1 U21963 ( .A1(n18997), .A2(n18860), .B1(n18859), .B2(n18858), .ZN(
        n18862) );
  NAND2_X1 U21964 ( .A1(n18862), .A2(n18861), .ZN(P3_U2839) );
  INV_X1 U21965 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18864) );
  NAND3_X1 U21966 ( .A1(n19062), .A2(n18872), .A3(n18863), .ZN(n18904) );
  OAI22_X1 U21967 ( .A1(n18864), .A2(n19082), .B1(n18875), .B2(n18904), .ZN(
        n18879) );
  INV_X1 U21968 ( .A(n18865), .ZN(n18892) );
  AOI21_X1 U21969 ( .B1(n18866), .B2(n18892), .A(n18877), .ZN(n18868) );
  OAI211_X1 U21970 ( .C1(n18872), .C2(n19546), .A(n18871), .B(n18870), .ZN(
        n18883) );
  OAI22_X1 U21971 ( .A1(n18877), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18975), .B2(n18873), .ZN(n18886) );
  AOI211_X1 U21972 ( .C1(n18875), .C2(n18874), .A(n18883), .B(n18886), .ZN(
        n18876) );
  OAI211_X1 U21973 ( .C1(n18877), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18876), .ZN(n18878) );
  AOI22_X1 U21974 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19066), .B1(
        n18879), .B2(n18878), .ZN(n18881) );
  OAI211_X1 U21975 ( .C1(n19012), .C2(n18882), .A(n18881), .B(n18880), .ZN(
        P3_U2840) );
  OAI21_X1 U21976 ( .B1(n18884), .B2(n18894), .A(n18893), .ZN(n18885) );
  OAI21_X1 U21977 ( .B1(n18886), .B2(n18885), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18891) );
  INV_X1 U21978 ( .A(n18904), .ZN(n18888) );
  AOI22_X1 U21979 ( .A1(n18997), .A2(n18889), .B1(n18888), .B2(n18887), .ZN(
        n18890) );
  OAI221_X1 U21980 ( .B1(n18905), .B2(n18891), .C1(n18988), .C2(n19658), .A(
        n18890), .ZN(P3_U2841) );
  NOR3_X1 U21981 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18894), .A3(
        n19582), .ZN(n18897) );
  NOR3_X1 U21982 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18895), .A3(
        n18904), .ZN(n18896) );
  AOI22_X1 U21983 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18901), .B1(
        n18997), .B2(n18900), .ZN(n18903) );
  OAI211_X1 U21984 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18904), .A(
        n18903), .B(n18902), .ZN(P3_U2843) );
  NAND2_X1 U21985 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18992), .ZN(
        n18910) );
  AOI22_X1 U21986 ( .A1(n18906), .A2(n18997), .B1(n18905), .B2(
        P3_REIP_REG_17__SCAN_IN), .ZN(n18909) );
  INV_X1 U21987 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18907) );
  NAND3_X1 U21988 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18921), .A3(
        n18907), .ZN(n18908) );
  OAI211_X1 U21989 ( .C1(n18911), .C2(n18910), .A(n18909), .B(n18908), .ZN(
        P3_U2845) );
  NOR2_X1 U21990 ( .A1(n18973), .A2(n18912), .ZN(n18918) );
  AOI22_X1 U21991 ( .A1(n18916), .A2(n18915), .B1(n18914), .B2(n18913), .ZN(
        n18990) );
  NAND2_X1 U21992 ( .A1(n18983), .A2(n18917), .ZN(n18944) );
  OAI211_X1 U21993 ( .C1(n18919), .C2(n18918), .A(n18990), .B(n18944), .ZN(
        n18928) );
  OAI221_X1 U21994 ( .B1(n18920), .B2(n19005), .C1(n18920), .C2(n18928), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18924) );
  AOI22_X1 U21995 ( .A1(n18997), .A2(n18922), .B1(n18921), .B2(n10082), .ZN(
        n18923) );
  OAI221_X1 U21996 ( .B1(n18905), .B2(n18924), .C1(n18988), .C2(n19648), .A(
        n18923), .ZN(P3_U2846) );
  NAND2_X1 U21997 ( .A1(n19057), .A2(n18925), .ZN(n18936) );
  AOI22_X1 U21998 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19066), .B1(
        n18905), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18935) );
  NOR2_X1 U21999 ( .A1(n18927), .A2(n18926), .ZN(n18941) );
  OAI221_X1 U22000 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18941), .A(n18928), .ZN(
        n18929) );
  OAI21_X1 U22001 ( .B1(n18931), .B2(n18930), .A(n18929), .ZN(n18933) );
  AOI22_X1 U22002 ( .A1(n19062), .A2(n18933), .B1(n18997), .B2(n18932), .ZN(
        n18934) );
  OAI211_X1 U22003 ( .C1(n18937), .C2(n18936), .A(n18935), .B(n18934), .ZN(
        P3_U2847) );
  AOI22_X1 U22004 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19066), .B1(
        n18905), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n18949) );
  AOI22_X1 U22005 ( .A1(n18991), .A2(n18990), .B1(n18939), .B2(n18938), .ZN(
        n18955) );
  AOI21_X1 U22006 ( .B1(n18973), .B2(n18940), .A(n18955), .ZN(n18945) );
  AOI22_X1 U22007 ( .A1(n18942), .A2(n18971), .B1(n18941), .B2(n10228), .ZN(
        n18943) );
  OAI221_X1 U22008 ( .B1(n10228), .B2(n18945), .C1(n10228), .C2(n18944), .A(
        n18943), .ZN(n18947) );
  AOI22_X1 U22009 ( .A1(n19062), .A2(n18947), .B1(n18997), .B2(n18946), .ZN(
        n18948) );
  OAI211_X1 U22010 ( .C1(n19095), .C2(n18950), .A(n18949), .B(n18948), .ZN(
        P3_U2848) );
  AOI22_X1 U22011 ( .A1(n18905), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18997), 
        .B2(n18951), .ZN(n18960) );
  OAI22_X1 U22012 ( .A1(n18953), .A2(n18952), .B1(n18978), .B2(n18977), .ZN(
        n18954) );
  AOI211_X1 U22013 ( .C1(n18957), .C2(n18956), .A(n18955), .B(n18954), .ZN(
        n18964) );
  OAI211_X1 U22014 ( .C1(n18978), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n19062), .B(n18964), .ZN(n18958) );
  NAND3_X1 U22015 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18988), .A3(
        n18958), .ZN(n18959) );
  OAI211_X1 U22016 ( .C1(n18961), .C2(n19001), .A(n18960), .B(n18959), .ZN(
        P3_U2849) );
  NAND3_X1 U22017 ( .A1(n18977), .A2(n18962), .A3(n18969), .ZN(n18963) );
  OAI21_X1 U22018 ( .B1(n18964), .B2(n18969), .A(n18963), .ZN(n18966) );
  AOI22_X1 U22019 ( .A1(n19062), .A2(n18966), .B1(n18997), .B2(n18965), .ZN(
        n18968) );
  OAI211_X1 U22020 ( .C1(n19090), .C2(n18969), .A(n18968), .B(n18967), .ZN(
        P3_U2850) );
  AOI22_X1 U22021 ( .A1(n18905), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18997), 
        .B2(n18970), .ZN(n18981) );
  NAND2_X1 U22022 ( .A1(n13637), .A2(n18971), .ZN(n19009) );
  OAI211_X1 U22023 ( .C1(n18972), .C2(n19545), .A(n19062), .B(n19009), .ZN(
        n18995) );
  AOI221_X1 U22024 ( .B1(n19000), .B2(n18973), .C1(n18994), .C2(n18973), .A(
        n18995), .ZN(n18974) );
  OAI211_X1 U22025 ( .C1(n18976), .C2(n18975), .A(n18990), .B(n18974), .ZN(
        n18984) );
  OAI22_X1 U22026 ( .A1(n18978), .A2(n18977), .B1(n18991), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18979) );
  OAI211_X1 U22027 ( .C1(n18984), .C2(n18979), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18988), .ZN(n18980) );
  OAI211_X1 U22028 ( .C1(n18982), .C2(n19001), .A(n18981), .B(n18980), .ZN(
        P3_U2851) );
  OAI221_X1 U22029 ( .B1(n18984), .B2(n18983), .C1(n18984), .C2(n19000), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18989) );
  NOR3_X1 U22030 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n19000), .A3(
        n19001), .ZN(n18985) );
  AOI21_X1 U22031 ( .B1(n18997), .B2(n18986), .A(n18985), .ZN(n18987) );
  OAI221_X1 U22032 ( .B1(n18905), .B2(n18989), .C1(n18988), .C2(n19636), .A(
        n18987), .ZN(P3_U2852) );
  NAND2_X1 U22033 ( .A1(n18991), .A2(n18990), .ZN(n18993) );
  OAI221_X1 U22034 ( .B1(n18995), .B2(n18994), .C1(n18995), .C2(n18993), .A(
        n18992), .ZN(n18999) );
  AOI22_X1 U22035 ( .A1(n18905), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18997), 
        .B2(n18996), .ZN(n18998) );
  OAI221_X1 U22036 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19001), .C1(
        n19000), .C2(n18999), .A(n18998), .ZN(P3_U2853) );
  INV_X1 U22037 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n19020) );
  NOR2_X1 U22038 ( .A1(n19546), .A2(n19002), .ZN(n19079) );
  AOI211_X1 U22039 ( .C1(n19075), .C2(n19003), .A(n19079), .B(n19076), .ZN(
        n19054) );
  OAI211_X1 U22040 ( .C1(n19004), .C2(n19022), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n19054), .ZN(n19021) );
  NAND3_X1 U22041 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19005), .A3(
        n19021), .ZN(n19008) );
  NAND3_X1 U22042 ( .A1(n19006), .A2(n19020), .A3(n19063), .ZN(n19007) );
  OAI211_X1 U22043 ( .C1(n19010), .C2(n19009), .A(n19008), .B(n19007), .ZN(
        n19011) );
  NAND2_X1 U22044 ( .A1(n19011), .A2(n19062), .ZN(n19015) );
  OR2_X1 U22045 ( .A1(n19013), .A2(n19012), .ZN(n19014) );
  OAI211_X1 U22046 ( .C1(n19016), .C2(n19095), .A(n19015), .B(n19014), .ZN(
        n19017) );
  INV_X1 U22047 ( .A(n19017), .ZN(n19019) );
  OAI211_X1 U22048 ( .C1(n19090), .C2(n19020), .A(n19019), .B(n19018), .ZN(
        P3_U2854) );
  OAI221_X1 U22049 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n19022), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n19063), .A(n19021), .ZN(
        n19028) );
  AOI21_X1 U22050 ( .B1(n19066), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n19023), .ZN(n19027) );
  AOI22_X1 U22051 ( .A1(n19025), .A2(n19057), .B1(n19086), .B2(n19024), .ZN(
        n19026) );
  OAI211_X1 U22052 ( .C1(n19082), .C2(n19028), .A(n19027), .B(n19026), .ZN(
        P3_U2855) );
  OAI21_X1 U22053 ( .B1(n19054), .B2(n19082), .A(n19090), .ZN(n19029) );
  AOI21_X1 U22054 ( .B1(n19030), .B2(n19036), .A(n19029), .ZN(n19043) );
  NAND3_X1 U22055 ( .A1(n19062), .A2(n19041), .A3(n19063), .ZN(n19037) );
  INV_X1 U22056 ( .A(n19031), .ZN(n19032) );
  NAND2_X1 U22057 ( .A1(n19057), .A2(n19032), .ZN(n19035) );
  NAND2_X1 U22058 ( .A1(n19086), .A2(n19033), .ZN(n19034) );
  OAI211_X1 U22059 ( .C1(n19037), .C2(n19036), .A(n19035), .B(n19034), .ZN(
        n19038) );
  INV_X1 U22060 ( .A(n19038), .ZN(n19040) );
  OAI211_X1 U22061 ( .C1(n19043), .C2(n19041), .A(n19040), .B(n19039), .ZN(
        P3_U2856) );
  NAND3_X1 U22062 ( .A1(n19062), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n19063), .ZN(n19061) );
  NOR2_X1 U22063 ( .A1(n19042), .A2(n19061), .ZN(n19045) );
  INV_X1 U22064 ( .A(n19043), .ZN(n19044) );
  MUX2_X1 U22065 ( .A(n19045), .B(n19044), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n19048) );
  AND2_X1 U22066 ( .A1(n19086), .A2(n19046), .ZN(n19047) );
  NOR2_X1 U22067 ( .A1(n19048), .A2(n19047), .ZN(n19050) );
  OAI211_X1 U22068 ( .C1(n19051), .C2(n19095), .A(n19050), .B(n19049), .ZN(
        P3_U2857) );
  AOI21_X1 U22069 ( .B1(n19086), .B2(n19053), .A(n19052), .ZN(n19060) );
  AND2_X1 U22070 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19054), .ZN(
        n19070) );
  OAI21_X1 U22071 ( .B1(n19070), .B2(n19055), .A(n19090), .ZN(n19058) );
  AOI22_X1 U22072 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n19058), .B1(
        n19057), .B2(n19056), .ZN(n19059) );
  OAI211_X1 U22073 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n19061), .A(
        n19060), .B(n19059), .ZN(P3_U2858) );
  OAI21_X1 U22074 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19063), .A(
        n19062), .ZN(n19069) );
  AOI21_X1 U22075 ( .B1(n19086), .B2(n19065), .A(n19064), .ZN(n19068) );
  NAND2_X1 U22076 ( .A1(n19066), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19067) );
  OAI211_X1 U22077 ( .C1(n19070), .C2(n19069), .A(n19068), .B(n19067), .ZN(
        n19071) );
  INV_X1 U22078 ( .A(n19071), .ZN(n19072) );
  OAI21_X1 U22079 ( .B1(n19095), .B2(n19073), .A(n19072), .ZN(P3_U2859) );
  NOR2_X1 U22080 ( .A1(n21541), .A2(n19074), .ZN(n19081) );
  NAND2_X1 U22081 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19078) );
  OAI21_X1 U22082 ( .B1(n19076), .B2(n21541), .A(n19075), .ZN(n19077) );
  OAI21_X1 U22083 ( .B1(n19078), .B2(n19546), .A(n19077), .ZN(n19080) );
  AOI221_X1 U22084 ( .B1(n19081), .B2(n19089), .C1(n19080), .C2(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n19079), .ZN(n19083) );
  NOR2_X1 U22085 ( .A1(n19083), .A2(n19082), .ZN(n19092) );
  INV_X1 U22086 ( .A(n19084), .ZN(n19085) );
  NAND2_X1 U22087 ( .A1(n19086), .A2(n19085), .ZN(n19088) );
  OAI211_X1 U22088 ( .C1(n19090), .C2(n19089), .A(n19088), .B(n19087), .ZN(
        n19091) );
  NOR2_X1 U22089 ( .A1(n19092), .A2(n19091), .ZN(n19093) );
  OAI21_X1 U22090 ( .B1(n19095), .B2(n19094), .A(n19093), .ZN(P3_U2860) );
  AOI21_X1 U22091 ( .B1(n19098), .B2(n19097), .A(n19096), .ZN(n19583) );
  OAI21_X1 U22092 ( .B1(n19583), .B2(n19144), .A(n19103), .ZN(n19099) );
  OAI221_X1 U22093 ( .B1(n11653), .B2(n19702), .C1(n11653), .C2(n19103), .A(
        n19099), .ZN(P3_U2863) );
  INV_X1 U22094 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19570) );
  NAND2_X1 U22095 ( .A1(n19568), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19363) );
  INV_X1 U22096 ( .A(n19363), .ZN(n19320) );
  INV_X1 U22097 ( .A(n19229), .ZN(n19276) );
  NOR2_X1 U22098 ( .A1(n19320), .A2(n19276), .ZN(n19101) );
  OAI22_X1 U22099 ( .A1(n19102), .A2(n19570), .B1(n19101), .B2(n19100), .ZN(
        P3_U2866) );
  NOR2_X1 U22100 ( .A1(n19571), .A2(n19103), .ZN(P3_U2867) );
  NAND2_X1 U22101 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19419) );
  INV_X1 U22102 ( .A(n19419), .ZN(n19421) );
  NOR2_X1 U22103 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n11653), .ZN(
        n19319) );
  NAND2_X1 U22104 ( .A1(n19421), .A2(n19319), .ZN(n19520) );
  NAND2_X1 U22105 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n16915), .ZN(n19455) );
  NOR2_X1 U22106 ( .A1(n19570), .A2(n19251), .ZN(n19482) );
  NAND2_X1 U22107 ( .A1(n11653), .A2(n19482), .ZN(n19462) );
  INV_X1 U22108 ( .A(n19462), .ZN(n19474) );
  INV_X1 U22109 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19104) );
  NOR2_X2 U22110 ( .A1(n19206), .A2(n19104), .ZN(n19484) );
  NOR2_X2 U22111 ( .A1(n19252), .A2(n19105), .ZN(n19479) );
  NOR2_X1 U22112 ( .A1(n11652), .A2(n11653), .ZN(n19558) );
  NAND2_X1 U22113 ( .A1(n19558), .A2(n19421), .ZN(n19494) );
  NOR2_X1 U22114 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19388) );
  NAND2_X1 U22115 ( .A1(n19388), .A2(n19185), .ZN(n19205) );
  NAND2_X1 U22116 ( .A1(n19494), .A2(n19205), .ZN(n19164) );
  AND2_X1 U22117 ( .A1(n19478), .A2(n19164), .ZN(n19138) );
  AOI22_X1 U22118 ( .A1(n19474), .A2(n19484), .B1(n19479), .B2(n19138), .ZN(
        n19110) );
  NAND2_X1 U22119 ( .A1(n19520), .A2(n19462), .ZN(n19451) );
  AOI21_X1 U22120 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n19252), .ZN(n19448) );
  AOI22_X1 U22121 ( .A1(n16915), .A2(n19451), .B1(n19448), .B2(n19164), .ZN(
        n19141) );
  NAND2_X1 U22122 ( .A1(n19107), .A2(n19106), .ZN(n19139) );
  NOR2_X1 U22123 ( .A1(n19108), .A2(n19139), .ZN(n19452) );
  AOI22_X1 U22124 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19141), .B1(
        n19198), .B2(n19452), .ZN(n19109) );
  OAI211_X1 U22125 ( .C1(n19520), .C2(n19455), .A(n19110), .B(n19109), .ZN(
        P3_U2868) );
  NAND2_X1 U22126 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n16915), .ZN(n19428) );
  INV_X1 U22127 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19111) );
  NOR2_X2 U22128 ( .A1(n19206), .A2(n19111), .ZN(n19490) );
  NOR2_X2 U22129 ( .A1(n19252), .A2(n19112), .ZN(n19488) );
  AOI22_X1 U22130 ( .A1(n19474), .A2(n19490), .B1(n19138), .B2(n19488), .ZN(
        n19114) );
  AOI22_X1 U22131 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19141), .B1(
        n19198), .B2(n19425), .ZN(n19113) );
  OAI211_X1 U22132 ( .C1(n19520), .C2(n19428), .A(n19114), .B(n19113), .ZN(
        P3_U2869) );
  NAND2_X1 U22133 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n16915), .ZN(n19500) );
  INV_X1 U22134 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n19115) );
  NOR2_X2 U22135 ( .A1(n19206), .A2(n19115), .ZN(n19496) );
  NOR2_X2 U22136 ( .A1(n19252), .A2(n19116), .ZN(n19495) );
  AOI22_X1 U22137 ( .A1(n19474), .A2(n19496), .B1(n19138), .B2(n19495), .ZN(
        n19119) );
  AOI22_X1 U22138 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19141), .B1(
        n19198), .B2(n19497), .ZN(n19118) );
  OAI211_X1 U22139 ( .C1(n19520), .C2(n19500), .A(n19119), .B(n19118), .ZN(
        P3_U2870) );
  INV_X1 U22140 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19120) );
  NOR2_X1 U22141 ( .A1(n19206), .A2(n19120), .ZN(n19502) );
  INV_X1 U22142 ( .A(n19502), .ZN(n19434) );
  INV_X1 U22143 ( .A(n19520), .ZN(n19530) );
  NAND2_X1 U22144 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n16915), .ZN(n19506) );
  INV_X1 U22145 ( .A(n19506), .ZN(n19431) );
  NOR2_X2 U22146 ( .A1(n19252), .A2(n19121), .ZN(n19501) );
  AOI22_X1 U22147 ( .A1(n19530), .A2(n19431), .B1(n19138), .B2(n19501), .ZN(
        n19124) );
  NOR2_X2 U22148 ( .A1(n19122), .A2(n19139), .ZN(n19503) );
  AOI22_X1 U22149 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19141), .B1(
        n19198), .B2(n19503), .ZN(n19123) );
  OAI211_X1 U22150 ( .C1(n19462), .C2(n19434), .A(n19124), .B(n19123), .ZN(
        P3_U2871) );
  NOR2_X1 U22151 ( .A1(n19125), .A2(n19206), .ZN(n19508) );
  NAND2_X1 U22152 ( .A1(n16915), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19512) );
  INV_X1 U22153 ( .A(n19512), .ZN(n19374) );
  NOR2_X2 U22154 ( .A1(n19252), .A2(n19126), .ZN(n19507) );
  AOI22_X1 U22155 ( .A1(n19474), .A2(n19374), .B1(n19138), .B2(n19507), .ZN(
        n19129) );
  NOR2_X2 U22156 ( .A1(n19127), .A2(n19139), .ZN(n19509) );
  AOI22_X1 U22157 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19141), .B1(
        n19198), .B2(n19509), .ZN(n19128) );
  OAI211_X1 U22158 ( .C1(n19520), .C2(n19377), .A(n19129), .B(n19128), .ZN(
        P3_U2872) );
  NOR2_X1 U22159 ( .A1(n19206), .A2(n16133), .ZN(n19404) );
  NAND2_X1 U22160 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n16915), .ZN(n19408) );
  INV_X1 U22161 ( .A(n19408), .ZN(n19515) );
  NOR2_X2 U22162 ( .A1(n19252), .A2(n19130), .ZN(n19513) );
  AOI22_X1 U22163 ( .A1(n19530), .A2(n19515), .B1(n19138), .B2(n19513), .ZN(
        n19133) );
  NOR2_X2 U22164 ( .A1(n19131), .A2(n19139), .ZN(n19516) );
  AOI22_X1 U22165 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19141), .B1(
        n19198), .B2(n19516), .ZN(n19132) );
  OAI211_X1 U22166 ( .C1(n19462), .C2(n19519), .A(n19133), .B(n19132), .ZN(
        P3_U2873) );
  NOR2_X1 U22167 ( .A1(n19206), .A2(n19134), .ZN(n19522) );
  NAND2_X1 U22168 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n16915), .ZN(n19526) );
  INV_X1 U22169 ( .A(n19526), .ZN(n19409) );
  NOR2_X2 U22170 ( .A1(n19252), .A2(n14001), .ZN(n19521) );
  AOI22_X1 U22171 ( .A1(n19530), .A2(n19409), .B1(n19138), .B2(n19521), .ZN(
        n19137) );
  NOR2_X2 U22172 ( .A1(n19135), .A2(n19139), .ZN(n19523) );
  AOI22_X1 U22173 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19141), .B1(
        n19198), .B2(n19523), .ZN(n19136) );
  OAI211_X1 U22174 ( .C1(n19462), .C2(n19412), .A(n19137), .B(n19136), .ZN(
        P3_U2874) );
  NAND2_X1 U22175 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n16915), .ZN(n19447) );
  NAND2_X1 U22176 ( .A1(n16915), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19537) );
  INV_X1 U22177 ( .A(n19537), .ZN(n19443) );
  NOR2_X2 U22178 ( .A1(n14047), .A2(n19252), .ZN(n19528) );
  AOI22_X1 U22179 ( .A1(n19530), .A2(n19443), .B1(n19138), .B2(n19528), .ZN(
        n19143) );
  NOR2_X2 U22180 ( .A1(n19140), .A2(n19139), .ZN(n19531) );
  AOI22_X1 U22181 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19141), .B1(
        n19198), .B2(n19531), .ZN(n19142) );
  OAI211_X1 U22182 ( .C1(n19462), .C2(n19447), .A(n19143), .B(n19142), .ZN(
        P3_U2875) );
  NAND2_X1 U22183 ( .A1(n19319), .A2(n19185), .ZN(n19223) );
  INV_X1 U22184 ( .A(n19455), .ZN(n19480) );
  INV_X1 U22185 ( .A(n19185), .ZN(n19163) );
  NAND2_X1 U22186 ( .A1(n11652), .A2(n19478), .ZN(n19418) );
  NOR2_X1 U22187 ( .A1(n19163), .A2(n19418), .ZN(n19159) );
  AOI22_X1 U22188 ( .A1(n19474), .A2(n19480), .B1(n19479), .B2(n19159), .ZN(
        n19146) );
  NOR2_X1 U22189 ( .A1(n19252), .A2(n19144), .ZN(n19481) );
  INV_X1 U22190 ( .A(n19481), .ZN(n19184) );
  NOR2_X1 U22191 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19184), .ZN(
        n19420) );
  AOI22_X1 U22192 ( .A1(n16915), .A2(n19482), .B1(n19185), .B2(n19420), .ZN(
        n19160) );
  INV_X1 U22193 ( .A(n19494), .ZN(n19532) );
  AOI22_X1 U22194 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19160), .B1(
        n19532), .B2(n19484), .ZN(n19145) );
  OAI211_X1 U22195 ( .C1(n19487), .C2(n19223), .A(n19146), .B(n19145), .ZN(
        P3_U2876) );
  INV_X1 U22196 ( .A(n19425), .ZN(n19493) );
  INV_X1 U22197 ( .A(n19428), .ZN(n19489) );
  AOI22_X1 U22198 ( .A1(n19474), .A2(n19489), .B1(n19488), .B2(n19159), .ZN(
        n19148) );
  AOI22_X1 U22199 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19160), .B1(
        n19532), .B2(n19490), .ZN(n19147) );
  OAI211_X1 U22200 ( .C1(n19493), .C2(n19223), .A(n19148), .B(n19147), .ZN(
        P3_U2877) );
  AOI22_X1 U22201 ( .A1(n19532), .A2(n19496), .B1(n19495), .B2(n19159), .ZN(
        n19150) );
  AOI22_X1 U22202 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19160), .B1(
        n19497), .B2(n19225), .ZN(n19149) );
  OAI211_X1 U22203 ( .C1(n19462), .C2(n19500), .A(n19150), .B(n19149), .ZN(
        P3_U2878) );
  AOI22_X1 U22204 ( .A1(n19474), .A2(n19431), .B1(n19501), .B2(n19159), .ZN(
        n19152) );
  AOI22_X1 U22205 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19160), .B1(
        n19503), .B2(n19225), .ZN(n19151) );
  OAI211_X1 U22206 ( .C1(n19494), .C2(n19434), .A(n19152), .B(n19151), .ZN(
        P3_U2879) );
  AOI22_X1 U22207 ( .A1(n19532), .A2(n19374), .B1(n19507), .B2(n19159), .ZN(
        n19154) );
  AOI22_X1 U22208 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19160), .B1(
        n19509), .B2(n19225), .ZN(n19153) );
  OAI211_X1 U22209 ( .C1(n19462), .C2(n19377), .A(n19154), .B(n19153), .ZN(
        P3_U2880) );
  AOI22_X1 U22210 ( .A1(n19474), .A2(n19515), .B1(n19513), .B2(n19159), .ZN(
        n19156) );
  AOI22_X1 U22211 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19160), .B1(
        n19516), .B2(n19225), .ZN(n19155) );
  OAI211_X1 U22212 ( .C1(n19494), .C2(n19519), .A(n19156), .B(n19155), .ZN(
        P3_U2881) );
  AOI22_X1 U22213 ( .A1(n19474), .A2(n19409), .B1(n19521), .B2(n19159), .ZN(
        n19158) );
  AOI22_X1 U22214 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19160), .B1(
        n19523), .B2(n19225), .ZN(n19157) );
  OAI211_X1 U22215 ( .C1(n19494), .C2(n19412), .A(n19158), .B(n19157), .ZN(
        P3_U2882) );
  INV_X1 U22216 ( .A(n19447), .ZN(n19529) );
  AOI22_X1 U22217 ( .A1(n19532), .A2(n19529), .B1(n19528), .B2(n19159), .ZN(
        n19162) );
  AOI22_X1 U22218 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19160), .B1(
        n19531), .B2(n19225), .ZN(n19161) );
  OAI211_X1 U22219 ( .C1(n19462), .C2(n19537), .A(n19162), .B(n19161), .ZN(
        P3_U2883) );
  NOR2_X1 U22220 ( .A1(n11652), .A2(n19163), .ZN(n19230) );
  NAND2_X1 U22221 ( .A1(n19230), .A2(n11653), .ZN(n19250) );
  INV_X1 U22222 ( .A(n19478), .ZN(n19595) );
  NAND2_X1 U22223 ( .A1(n19223), .A2(n19250), .ZN(n19165) );
  INV_X1 U22224 ( .A(n19165), .ZN(n19207) );
  NOR2_X1 U22225 ( .A1(n19595), .A2(n19207), .ZN(n19180) );
  AOI22_X1 U22226 ( .A1(n19532), .A2(n19480), .B1(n19479), .B2(n19180), .ZN(
        n19167) );
  OAI221_X1 U22227 ( .B1(n19165), .B2(n19450), .C1(n19165), .C2(n19164), .A(
        n19448), .ZN(n19181) );
  AOI22_X1 U22228 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19181), .B1(
        n19198), .B2(n19484), .ZN(n19166) );
  OAI211_X1 U22229 ( .C1(n19487), .C2(n19250), .A(n19167), .B(n19166), .ZN(
        P3_U2884) );
  AOI22_X1 U22230 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19181), .B1(
        n19488), .B2(n19180), .ZN(n19169) );
  AOI22_X1 U22231 ( .A1(n19198), .A2(n19490), .B1(n19425), .B2(n19243), .ZN(
        n19168) );
  OAI211_X1 U22232 ( .C1(n19494), .C2(n19428), .A(n19169), .B(n19168), .ZN(
        P3_U2885) );
  AOI22_X1 U22233 ( .A1(n19532), .A2(n19458), .B1(n19495), .B2(n19180), .ZN(
        n19171) );
  AOI22_X1 U22234 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19181), .B1(
        n19198), .B2(n19496), .ZN(n19170) );
  OAI211_X1 U22235 ( .C1(n19461), .C2(n19250), .A(n19171), .B(n19170), .ZN(
        P3_U2886) );
  AOI22_X1 U22236 ( .A1(n19198), .A2(n19502), .B1(n19501), .B2(n19180), .ZN(
        n19173) );
  AOI22_X1 U22237 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19181), .B1(
        n19503), .B2(n19243), .ZN(n19172) );
  OAI211_X1 U22238 ( .C1(n19494), .C2(n19506), .A(n19173), .B(n19172), .ZN(
        P3_U2887) );
  AOI22_X1 U22239 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19181), .B1(
        n19507), .B2(n19180), .ZN(n19175) );
  AOI22_X1 U22240 ( .A1(n19198), .A2(n19374), .B1(n19509), .B2(n19243), .ZN(
        n19174) );
  OAI211_X1 U22241 ( .C1(n19494), .C2(n19377), .A(n19175), .B(n19174), .ZN(
        P3_U2888) );
  AOI22_X1 U22242 ( .A1(n19532), .A2(n19515), .B1(n19513), .B2(n19180), .ZN(
        n19177) );
  AOI22_X1 U22243 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19181), .B1(
        n19516), .B2(n19243), .ZN(n19176) );
  OAI211_X1 U22244 ( .C1(n19205), .C2(n19519), .A(n19177), .B(n19176), .ZN(
        P3_U2889) );
  AOI22_X1 U22245 ( .A1(n19532), .A2(n19409), .B1(n19521), .B2(n19180), .ZN(
        n19179) );
  AOI22_X1 U22246 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19181), .B1(
        n19523), .B2(n19243), .ZN(n19178) );
  OAI211_X1 U22247 ( .C1(n19205), .C2(n19412), .A(n19179), .B(n19178), .ZN(
        P3_U2890) );
  AOI22_X1 U22248 ( .A1(n19532), .A2(n19443), .B1(n19528), .B2(n19180), .ZN(
        n19183) );
  AOI22_X1 U22249 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19181), .B1(
        n19531), .B2(n19243), .ZN(n19182) );
  OAI211_X1 U22250 ( .C1(n19205), .C2(n19447), .A(n19183), .B(n19182), .ZN(
        P3_U2891) );
  AND2_X1 U22251 ( .A1(n19478), .A2(n19230), .ZN(n19201) );
  AOI22_X1 U22252 ( .A1(n19484), .A2(n19225), .B1(n19479), .B2(n19201), .ZN(
        n19187) );
  AOI21_X1 U22253 ( .B1(n11652), .B2(n19390), .A(n19184), .ZN(n19275) );
  NAND2_X1 U22254 ( .A1(n19185), .A2(n19275), .ZN(n19202) );
  NAND2_X1 U22255 ( .A1(n19558), .A2(n19185), .ZN(n19274) );
  INV_X1 U22256 ( .A(n19274), .ZN(n19263) );
  AOI22_X1 U22257 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19202), .B1(
        n19452), .B2(n19263), .ZN(n19186) );
  OAI211_X1 U22258 ( .C1(n19205), .C2(n19455), .A(n19187), .B(n19186), .ZN(
        P3_U2892) );
  AOI22_X1 U22259 ( .A1(n19198), .A2(n19489), .B1(n19488), .B2(n19201), .ZN(
        n19189) );
  AOI22_X1 U22260 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19202), .B1(
        n19490), .B2(n19225), .ZN(n19188) );
  OAI211_X1 U22261 ( .C1(n19493), .C2(n19274), .A(n19189), .B(n19188), .ZN(
        P3_U2893) );
  AOI22_X1 U22262 ( .A1(n19496), .A2(n19225), .B1(n19495), .B2(n19201), .ZN(
        n19191) );
  AOI22_X1 U22263 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19202), .B1(
        n19497), .B2(n19263), .ZN(n19190) );
  OAI211_X1 U22264 ( .C1(n19205), .C2(n19500), .A(n19191), .B(n19190), .ZN(
        P3_U2894) );
  AOI22_X1 U22265 ( .A1(n19198), .A2(n19431), .B1(n19501), .B2(n19201), .ZN(
        n19193) );
  AOI22_X1 U22266 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19202), .B1(
        n19503), .B2(n19263), .ZN(n19192) );
  OAI211_X1 U22267 ( .C1(n19434), .C2(n19223), .A(n19193), .B(n19192), .ZN(
        P3_U2895) );
  AOI22_X1 U22268 ( .A1(n19198), .A2(n19508), .B1(n19507), .B2(n19201), .ZN(
        n19195) );
  AOI22_X1 U22269 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19202), .B1(
        n19509), .B2(n19263), .ZN(n19194) );
  OAI211_X1 U22270 ( .C1(n19512), .C2(n19223), .A(n19195), .B(n19194), .ZN(
        P3_U2896) );
  AOI22_X1 U22271 ( .A1(n19198), .A2(n19515), .B1(n19513), .B2(n19201), .ZN(
        n19197) );
  AOI22_X1 U22272 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19202), .B1(
        n19516), .B2(n19263), .ZN(n19196) );
  OAI211_X1 U22273 ( .C1(n19519), .C2(n19223), .A(n19197), .B(n19196), .ZN(
        P3_U2897) );
  AOI22_X1 U22274 ( .A1(n19198), .A2(n19409), .B1(n19521), .B2(n19201), .ZN(
        n19200) );
  AOI22_X1 U22275 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19202), .B1(
        n19523), .B2(n19263), .ZN(n19199) );
  OAI211_X1 U22276 ( .C1(n19412), .C2(n19223), .A(n19200), .B(n19199), .ZN(
        P3_U2898) );
  AOI22_X1 U22277 ( .A1(n19529), .A2(n19225), .B1(n19528), .B2(n19201), .ZN(
        n19204) );
  AOI22_X1 U22278 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19202), .B1(
        n19531), .B2(n19263), .ZN(n19203) );
  OAI211_X1 U22279 ( .C1(n19205), .C2(n19537), .A(n19204), .B(n19203), .ZN(
        P3_U2899) );
  INV_X1 U22280 ( .A(n19388), .ZN(n19563) );
  NOR2_X2 U22281 ( .A1(n19563), .A2(n19229), .ZN(n19289) );
  NOR2_X1 U22282 ( .A1(n19263), .A2(n19289), .ZN(n19253) );
  NOR2_X1 U22283 ( .A1(n19595), .A2(n19253), .ZN(n19224) );
  AOI22_X1 U22284 ( .A1(n19480), .A2(n19225), .B1(n19479), .B2(n19224), .ZN(
        n19210) );
  OAI22_X1 U22285 ( .A1(n19207), .A2(n19206), .B1(n19253), .B2(n19252), .ZN(
        n19208) );
  OAI21_X1 U22286 ( .B1(n19289), .B2(n19690), .A(n19208), .ZN(n19226) );
  AOI22_X1 U22287 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19226), .B1(
        n19484), .B2(n19243), .ZN(n19209) );
  OAI211_X1 U22288 ( .C1(n19487), .C2(n19296), .A(n19210), .B(n19209), .ZN(
        P3_U2900) );
  AOI22_X1 U22289 ( .A1(n19489), .A2(n19225), .B1(n19488), .B2(n19224), .ZN(
        n19212) );
  AOI22_X1 U22290 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19226), .B1(
        n19490), .B2(n19243), .ZN(n19211) );
  OAI211_X1 U22291 ( .C1(n19493), .C2(n19296), .A(n19212), .B(n19211), .ZN(
        P3_U2901) );
  AOI22_X1 U22292 ( .A1(n19458), .A2(n19225), .B1(n19495), .B2(n19224), .ZN(
        n19214) );
  AOI22_X1 U22293 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19226), .B1(
        n19496), .B2(n19243), .ZN(n19213) );
  OAI211_X1 U22294 ( .C1(n19461), .C2(n19296), .A(n19214), .B(n19213), .ZN(
        P3_U2902) );
  AOI22_X1 U22295 ( .A1(n19502), .A2(n19243), .B1(n19501), .B2(n19224), .ZN(
        n19216) );
  AOI22_X1 U22296 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19226), .B1(
        n19503), .B2(n19289), .ZN(n19215) );
  OAI211_X1 U22297 ( .C1(n19506), .C2(n19223), .A(n19216), .B(n19215), .ZN(
        P3_U2903) );
  AOI22_X1 U22298 ( .A1(n19374), .A2(n19243), .B1(n19507), .B2(n19224), .ZN(
        n19218) );
  AOI22_X1 U22299 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19226), .B1(
        n19509), .B2(n19289), .ZN(n19217) );
  OAI211_X1 U22300 ( .C1(n19377), .C2(n19223), .A(n19218), .B(n19217), .ZN(
        P3_U2904) );
  AOI22_X1 U22301 ( .A1(n19404), .A2(n19243), .B1(n19513), .B2(n19224), .ZN(
        n19220) );
  AOI22_X1 U22302 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19226), .B1(
        n19516), .B2(n19289), .ZN(n19219) );
  OAI211_X1 U22303 ( .C1(n19408), .C2(n19223), .A(n19220), .B(n19219), .ZN(
        P3_U2905) );
  AOI22_X1 U22304 ( .A1(n19522), .A2(n19243), .B1(n19521), .B2(n19224), .ZN(
        n19222) );
  AOI22_X1 U22305 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19226), .B1(
        n19523), .B2(n19289), .ZN(n19221) );
  OAI211_X1 U22306 ( .C1(n19526), .C2(n19223), .A(n19222), .B(n19221), .ZN(
        P3_U2906) );
  AOI22_X1 U22307 ( .A1(n19443), .A2(n19225), .B1(n19528), .B2(n19224), .ZN(
        n19228) );
  AOI22_X1 U22308 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19226), .B1(
        n19531), .B2(n19289), .ZN(n19227) );
  OAI211_X1 U22309 ( .C1(n19447), .C2(n19250), .A(n19228), .B(n19227), .ZN(
        P3_U2907) );
  NAND2_X1 U22310 ( .A1(n19276), .A2(n19319), .ZN(n19313) );
  NOR2_X1 U22311 ( .A1(n19229), .A2(n19418), .ZN(n19246) );
  AOI22_X1 U22312 ( .A1(n19480), .A2(n19243), .B1(n19479), .B2(n19246), .ZN(
        n19232) );
  AOI22_X1 U22313 ( .A1(n16915), .A2(n19230), .B1(n19276), .B2(n19420), .ZN(
        n19247) );
  AOI22_X1 U22314 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19247), .B1(
        n19484), .B2(n19263), .ZN(n19231) );
  OAI211_X1 U22315 ( .C1(n19487), .C2(n19313), .A(n19232), .B(n19231), .ZN(
        P3_U2908) );
  AOI22_X1 U22316 ( .A1(n19490), .A2(n19263), .B1(n19488), .B2(n19246), .ZN(
        n19234) );
  AOI22_X1 U22317 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19247), .B1(
        n19489), .B2(n19243), .ZN(n19233) );
  OAI211_X1 U22318 ( .C1(n19493), .C2(n19313), .A(n19234), .B(n19233), .ZN(
        P3_U2909) );
  AOI22_X1 U22319 ( .A1(n19496), .A2(n19263), .B1(n19495), .B2(n19246), .ZN(
        n19236) );
  AOI22_X1 U22320 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19247), .B1(
        n19458), .B2(n19243), .ZN(n19235) );
  OAI211_X1 U22321 ( .C1(n19461), .C2(n19313), .A(n19236), .B(n19235), .ZN(
        P3_U2910) );
  AOI22_X1 U22322 ( .A1(n19502), .A2(n19263), .B1(n19501), .B2(n19246), .ZN(
        n19238) );
  INV_X1 U22323 ( .A(n19313), .ZN(n19315) );
  AOI22_X1 U22324 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19247), .B1(
        n19503), .B2(n19315), .ZN(n19237) );
  OAI211_X1 U22325 ( .C1(n19506), .C2(n19250), .A(n19238), .B(n19237), .ZN(
        P3_U2911) );
  AOI22_X1 U22326 ( .A1(n19374), .A2(n19263), .B1(n19507), .B2(n19246), .ZN(
        n19240) );
  AOI22_X1 U22327 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19247), .B1(
        n19509), .B2(n19315), .ZN(n19239) );
  OAI211_X1 U22328 ( .C1(n19377), .C2(n19250), .A(n19240), .B(n19239), .ZN(
        P3_U2912) );
  AOI22_X1 U22329 ( .A1(n19515), .A2(n19243), .B1(n19513), .B2(n19246), .ZN(
        n19242) );
  AOI22_X1 U22330 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19247), .B1(
        n19516), .B2(n19315), .ZN(n19241) );
  OAI211_X1 U22331 ( .C1(n19519), .C2(n19274), .A(n19242), .B(n19241), .ZN(
        P3_U2913) );
  AOI22_X1 U22332 ( .A1(n19409), .A2(n19243), .B1(n19521), .B2(n19246), .ZN(
        n19245) );
  AOI22_X1 U22333 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19247), .B1(
        n19523), .B2(n19315), .ZN(n19244) );
  OAI211_X1 U22334 ( .C1(n19412), .C2(n19274), .A(n19245), .B(n19244), .ZN(
        P3_U2914) );
  AOI22_X1 U22335 ( .A1(n19529), .A2(n19263), .B1(n19528), .B2(n19246), .ZN(
        n19249) );
  AOI22_X1 U22336 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19247), .B1(
        n19531), .B2(n19315), .ZN(n19248) );
  OAI211_X1 U22337 ( .C1(n19537), .C2(n19250), .A(n19249), .B(n19248), .ZN(
        P3_U2915) );
  NOR2_X1 U22338 ( .A1(n19251), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19321) );
  NAND2_X1 U22339 ( .A1(n11653), .A2(n19321), .ZN(n19340) );
  NOR2_X1 U22340 ( .A1(n19315), .A2(n19328), .ZN(n19297) );
  NOR2_X1 U22341 ( .A1(n19595), .A2(n19297), .ZN(n19270) );
  AOI22_X1 U22342 ( .A1(n19484), .A2(n19289), .B1(n19479), .B2(n19270), .ZN(
        n19256) );
  INV_X1 U22343 ( .A(n19252), .ZN(n19393) );
  OAI21_X1 U22344 ( .B1(n19253), .B2(n19390), .A(n19297), .ZN(n19254) );
  OAI211_X1 U22345 ( .C1(n19328), .C2(n19690), .A(n19393), .B(n19254), .ZN(
        n19271) );
  AOI22_X1 U22346 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19271), .B1(
        n19452), .B2(n19328), .ZN(n19255) );
  OAI211_X1 U22347 ( .C1(n19455), .C2(n19274), .A(n19256), .B(n19255), .ZN(
        P3_U2916) );
  AOI22_X1 U22348 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19271), .B1(
        n19488), .B2(n19270), .ZN(n19258) );
  AOI22_X1 U22349 ( .A1(n19425), .A2(n19328), .B1(n19490), .B2(n19289), .ZN(
        n19257) );
  OAI211_X1 U22350 ( .C1(n19428), .C2(n19274), .A(n19258), .B(n19257), .ZN(
        P3_U2917) );
  AOI22_X1 U22351 ( .A1(n19458), .A2(n19263), .B1(n19495), .B2(n19270), .ZN(
        n19260) );
  AOI22_X1 U22352 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19271), .B1(
        n19496), .B2(n19289), .ZN(n19259) );
  OAI211_X1 U22353 ( .C1(n19461), .C2(n19340), .A(n19260), .B(n19259), .ZN(
        P3_U2918) );
  AOI22_X1 U22354 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19271), .B1(
        n19501), .B2(n19270), .ZN(n19262) );
  AOI22_X1 U22355 ( .A1(n19502), .A2(n19289), .B1(n19503), .B2(n19328), .ZN(
        n19261) );
  OAI211_X1 U22356 ( .C1(n19506), .C2(n19274), .A(n19262), .B(n19261), .ZN(
        P3_U2919) );
  AOI22_X1 U22357 ( .A1(n19508), .A2(n19263), .B1(n19507), .B2(n19270), .ZN(
        n19265) );
  AOI22_X1 U22358 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19271), .B1(
        n19509), .B2(n19328), .ZN(n19264) );
  OAI211_X1 U22359 ( .C1(n19512), .C2(n19296), .A(n19265), .B(n19264), .ZN(
        P3_U2920) );
  AOI22_X1 U22360 ( .A1(n19404), .A2(n19289), .B1(n19513), .B2(n19270), .ZN(
        n19267) );
  AOI22_X1 U22361 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19271), .B1(
        n19516), .B2(n19328), .ZN(n19266) );
  OAI211_X1 U22362 ( .C1(n19408), .C2(n19274), .A(n19267), .B(n19266), .ZN(
        P3_U2921) );
  AOI22_X1 U22363 ( .A1(n19522), .A2(n19289), .B1(n19521), .B2(n19270), .ZN(
        n19269) );
  AOI22_X1 U22364 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19271), .B1(
        n19523), .B2(n19328), .ZN(n19268) );
  OAI211_X1 U22365 ( .C1(n19526), .C2(n19274), .A(n19269), .B(n19268), .ZN(
        P3_U2922) );
  AOI22_X1 U22366 ( .A1(n19529), .A2(n19289), .B1(n19528), .B2(n19270), .ZN(
        n19273) );
  AOI22_X1 U22367 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19271), .B1(
        n19531), .B2(n19328), .ZN(n19272) );
  OAI211_X1 U22368 ( .C1(n19537), .C2(n19274), .A(n19273), .B(n19272), .ZN(
        P3_U2923) );
  AND2_X1 U22369 ( .A1(n19478), .A2(n19321), .ZN(n19292) );
  AOI22_X1 U22370 ( .A1(n19484), .A2(n19315), .B1(n19479), .B2(n19292), .ZN(
        n19278) );
  NAND2_X1 U22371 ( .A1(n19276), .A2(n19275), .ZN(n19293) );
  NAND2_X1 U22372 ( .A1(n19558), .A2(n19276), .ZN(n19362) );
  AOI22_X1 U22373 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19293), .B1(
        n19452), .B2(n19355), .ZN(n19277) );
  OAI211_X1 U22374 ( .C1(n19455), .C2(n19296), .A(n19278), .B(n19277), .ZN(
        P3_U2924) );
  AOI22_X1 U22375 ( .A1(n19490), .A2(n19315), .B1(n19488), .B2(n19292), .ZN(
        n19280) );
  AOI22_X1 U22376 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19293), .B1(
        n19425), .B2(n19355), .ZN(n19279) );
  OAI211_X1 U22377 ( .C1(n19428), .C2(n19296), .A(n19280), .B(n19279), .ZN(
        P3_U2925) );
  AOI22_X1 U22378 ( .A1(n19458), .A2(n19289), .B1(n19495), .B2(n19292), .ZN(
        n19282) );
  AOI22_X1 U22379 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19293), .B1(
        n19496), .B2(n19315), .ZN(n19281) );
  OAI211_X1 U22380 ( .C1(n19461), .C2(n19362), .A(n19282), .B(n19281), .ZN(
        P3_U2926) );
  AOI22_X1 U22381 ( .A1(n19502), .A2(n19315), .B1(n19501), .B2(n19292), .ZN(
        n19284) );
  AOI22_X1 U22382 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19293), .B1(
        n19503), .B2(n19355), .ZN(n19283) );
  OAI211_X1 U22383 ( .C1(n19506), .C2(n19296), .A(n19284), .B(n19283), .ZN(
        P3_U2927) );
  AOI22_X1 U22384 ( .A1(n19374), .A2(n19315), .B1(n19507), .B2(n19292), .ZN(
        n19286) );
  AOI22_X1 U22385 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19293), .B1(
        n19509), .B2(n19355), .ZN(n19285) );
  OAI211_X1 U22386 ( .C1(n19377), .C2(n19296), .A(n19286), .B(n19285), .ZN(
        P3_U2928) );
  AOI22_X1 U22387 ( .A1(n19515), .A2(n19289), .B1(n19513), .B2(n19292), .ZN(
        n19288) );
  AOI22_X1 U22388 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19293), .B1(
        n19516), .B2(n19355), .ZN(n19287) );
  OAI211_X1 U22389 ( .C1(n19519), .C2(n19313), .A(n19288), .B(n19287), .ZN(
        P3_U2929) );
  AOI22_X1 U22390 ( .A1(n19409), .A2(n19289), .B1(n19521), .B2(n19292), .ZN(
        n19291) );
  AOI22_X1 U22391 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19293), .B1(
        n19523), .B2(n19355), .ZN(n19290) );
  OAI211_X1 U22392 ( .C1(n19412), .C2(n19313), .A(n19291), .B(n19290), .ZN(
        P3_U2930) );
  AOI22_X1 U22393 ( .A1(n19529), .A2(n19315), .B1(n19528), .B2(n19292), .ZN(
        n19295) );
  AOI22_X1 U22394 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19293), .B1(
        n19531), .B2(n19355), .ZN(n19294) );
  OAI211_X1 U22395 ( .C1(n19537), .C2(n19296), .A(n19295), .B(n19294), .ZN(
        P3_U2931) );
  NOR2_X2 U22396 ( .A1(n19563), .A2(n19363), .ZN(n19384) );
  INV_X1 U22397 ( .A(n19384), .ZN(n19380) );
  NOR2_X1 U22398 ( .A1(n19355), .A2(n19384), .ZN(n19341) );
  NOR2_X1 U22399 ( .A1(n19595), .A2(n19341), .ZN(n19314) );
  AOI22_X1 U22400 ( .A1(n19480), .A2(n19315), .B1(n19479), .B2(n19314), .ZN(
        n19300) );
  OAI21_X1 U22401 ( .B1(n19297), .B2(n19390), .A(n19341), .ZN(n19298) );
  OAI211_X1 U22402 ( .C1(n19384), .C2(n19690), .A(n19393), .B(n19298), .ZN(
        n19316) );
  AOI22_X1 U22403 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19316), .B1(
        n19484), .B2(n19328), .ZN(n19299) );
  OAI211_X1 U22404 ( .C1(n19487), .C2(n19380), .A(n19300), .B(n19299), .ZN(
        P3_U2932) );
  AOI22_X1 U22405 ( .A1(n19489), .A2(n19315), .B1(n19488), .B2(n19314), .ZN(
        n19302) );
  AOI22_X1 U22406 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19316), .B1(
        n19490), .B2(n19328), .ZN(n19301) );
  OAI211_X1 U22407 ( .C1(n19493), .C2(n19380), .A(n19302), .B(n19301), .ZN(
        P3_U2933) );
  AOI22_X1 U22408 ( .A1(n19496), .A2(n19328), .B1(n19495), .B2(n19314), .ZN(
        n19304) );
  AOI22_X1 U22409 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19316), .B1(
        n19497), .B2(n19384), .ZN(n19303) );
  OAI211_X1 U22410 ( .C1(n19500), .C2(n19313), .A(n19304), .B(n19303), .ZN(
        P3_U2934) );
  AOI22_X1 U22411 ( .A1(n19502), .A2(n19328), .B1(n19501), .B2(n19314), .ZN(
        n19306) );
  AOI22_X1 U22412 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19316), .B1(
        n19503), .B2(n19384), .ZN(n19305) );
  OAI211_X1 U22413 ( .C1(n19506), .C2(n19313), .A(n19306), .B(n19305), .ZN(
        P3_U2935) );
  AOI22_X1 U22414 ( .A1(n19508), .A2(n19315), .B1(n19507), .B2(n19314), .ZN(
        n19308) );
  AOI22_X1 U22415 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19316), .B1(
        n19509), .B2(n19384), .ZN(n19307) );
  OAI211_X1 U22416 ( .C1(n19512), .C2(n19340), .A(n19308), .B(n19307), .ZN(
        P3_U2936) );
  AOI22_X1 U22417 ( .A1(n19404), .A2(n19328), .B1(n19513), .B2(n19314), .ZN(
        n19310) );
  AOI22_X1 U22418 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19316), .B1(
        n19516), .B2(n19384), .ZN(n19309) );
  OAI211_X1 U22419 ( .C1(n19408), .C2(n19313), .A(n19310), .B(n19309), .ZN(
        P3_U2937) );
  AOI22_X1 U22420 ( .A1(n19522), .A2(n19328), .B1(n19521), .B2(n19314), .ZN(
        n19312) );
  AOI22_X1 U22421 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19316), .B1(
        n19523), .B2(n19384), .ZN(n19311) );
  OAI211_X1 U22422 ( .C1(n19526), .C2(n19313), .A(n19312), .B(n19311), .ZN(
        P3_U2938) );
  AOI22_X1 U22423 ( .A1(n19443), .A2(n19315), .B1(n19528), .B2(n19314), .ZN(
        n19318) );
  AOI22_X1 U22424 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19316), .B1(
        n19531), .B2(n19384), .ZN(n19317) );
  OAI211_X1 U22425 ( .C1(n19447), .C2(n19340), .A(n19318), .B(n19317), .ZN(
        P3_U2939) );
  NAND2_X1 U22426 ( .A1(n19320), .A2(n19319), .ZN(n19407) );
  NOR2_X1 U22427 ( .A1(n19363), .A2(n19418), .ZN(n19365) );
  AOI22_X1 U22428 ( .A1(n19484), .A2(n19355), .B1(n19479), .B2(n19365), .ZN(
        n19323) );
  AOI22_X1 U22429 ( .A1(n16915), .A2(n19321), .B1(n19320), .B2(n19420), .ZN(
        n19337) );
  AOI22_X1 U22430 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19337), .B1(
        n19480), .B2(n19328), .ZN(n19322) );
  OAI211_X1 U22431 ( .C1(n19487), .C2(n19407), .A(n19323), .B(n19322), .ZN(
        P3_U2940) );
  AOI22_X1 U22432 ( .A1(n19489), .A2(n19328), .B1(n19488), .B2(n19365), .ZN(
        n19325) );
  AOI22_X1 U22433 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19337), .B1(
        n19490), .B2(n19355), .ZN(n19324) );
  OAI211_X1 U22434 ( .C1(n19493), .C2(n19407), .A(n19325), .B(n19324), .ZN(
        P3_U2941) );
  AOI22_X1 U22435 ( .A1(n19458), .A2(n19328), .B1(n19495), .B2(n19365), .ZN(
        n19327) );
  AOI22_X1 U22436 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19337), .B1(
        n19496), .B2(n19355), .ZN(n19326) );
  OAI211_X1 U22437 ( .C1(n19461), .C2(n19407), .A(n19327), .B(n19326), .ZN(
        P3_U2942) );
  AOI22_X1 U22438 ( .A1(n19501), .A2(n19365), .B1(n19431), .B2(n19328), .ZN(
        n19330) );
  AOI22_X1 U22439 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19337), .B1(
        n19503), .B2(n19414), .ZN(n19329) );
  OAI211_X1 U22440 ( .C1(n19434), .C2(n19362), .A(n19330), .B(n19329), .ZN(
        P3_U2943) );
  AOI22_X1 U22441 ( .A1(n19374), .A2(n19355), .B1(n19507), .B2(n19365), .ZN(
        n19332) );
  AOI22_X1 U22442 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19337), .B1(
        n19509), .B2(n19414), .ZN(n19331) );
  OAI211_X1 U22443 ( .C1(n19377), .C2(n19340), .A(n19332), .B(n19331), .ZN(
        P3_U2944) );
  AOI22_X1 U22444 ( .A1(n19404), .A2(n19355), .B1(n19513), .B2(n19365), .ZN(
        n19334) );
  AOI22_X1 U22445 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19337), .B1(
        n19516), .B2(n19414), .ZN(n19333) );
  OAI211_X1 U22446 ( .C1(n19408), .C2(n19340), .A(n19334), .B(n19333), .ZN(
        P3_U2945) );
  AOI22_X1 U22447 ( .A1(n19522), .A2(n19355), .B1(n19521), .B2(n19365), .ZN(
        n19336) );
  AOI22_X1 U22448 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19337), .B1(
        n19523), .B2(n19414), .ZN(n19335) );
  OAI211_X1 U22449 ( .C1(n19526), .C2(n19340), .A(n19336), .B(n19335), .ZN(
        P3_U2946) );
  AOI22_X1 U22450 ( .A1(n19529), .A2(n19355), .B1(n19528), .B2(n19365), .ZN(
        n19339) );
  AOI22_X1 U22451 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19337), .B1(
        n19531), .B2(n19414), .ZN(n19338) );
  OAI211_X1 U22452 ( .C1(n19537), .C2(n19340), .A(n19339), .B(n19338), .ZN(
        P3_U2947) );
  NOR2_X1 U22453 ( .A1(n11652), .A2(n19363), .ZN(n19422) );
  NAND2_X1 U22454 ( .A1(n11653), .A2(n19422), .ZN(n19441) );
  INV_X1 U22455 ( .A(n19441), .ZN(n19442) );
  NOR2_X1 U22456 ( .A1(n19414), .A2(n19442), .ZN(n19391) );
  NOR2_X1 U22457 ( .A1(n19595), .A2(n19391), .ZN(n19358) );
  AOI22_X1 U22458 ( .A1(n19484), .A2(n19384), .B1(n19479), .B2(n19358), .ZN(
        n19344) );
  OAI21_X1 U22459 ( .B1(n19341), .B2(n19390), .A(n19391), .ZN(n19342) );
  OAI211_X1 U22460 ( .C1(n19442), .C2(n19690), .A(n19393), .B(n19342), .ZN(
        n19359) );
  AOI22_X1 U22461 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19359), .B1(
        n19452), .B2(n19442), .ZN(n19343) );
  OAI211_X1 U22462 ( .C1(n19455), .C2(n19362), .A(n19344), .B(n19343), .ZN(
        P3_U2948) );
  AOI22_X1 U22463 ( .A1(n19490), .A2(n19384), .B1(n19488), .B2(n19358), .ZN(
        n19346) );
  AOI22_X1 U22464 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19359), .B1(
        n19425), .B2(n19442), .ZN(n19345) );
  OAI211_X1 U22465 ( .C1(n19428), .C2(n19362), .A(n19346), .B(n19345), .ZN(
        P3_U2949) );
  AOI22_X1 U22466 ( .A1(n19458), .A2(n19355), .B1(n19495), .B2(n19358), .ZN(
        n19348) );
  AOI22_X1 U22467 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19359), .B1(
        n19496), .B2(n19384), .ZN(n19347) );
  OAI211_X1 U22468 ( .C1(n19461), .C2(n19441), .A(n19348), .B(n19347), .ZN(
        P3_U2950) );
  AOI22_X1 U22469 ( .A1(n19502), .A2(n19384), .B1(n19501), .B2(n19358), .ZN(
        n19350) );
  AOI22_X1 U22470 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19359), .B1(
        n19503), .B2(n19442), .ZN(n19349) );
  OAI211_X1 U22471 ( .C1(n19506), .C2(n19362), .A(n19350), .B(n19349), .ZN(
        P3_U2951) );
  AOI22_X1 U22472 ( .A1(n19508), .A2(n19355), .B1(n19507), .B2(n19358), .ZN(
        n19352) );
  AOI22_X1 U22473 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19359), .B1(
        n19509), .B2(n19442), .ZN(n19351) );
  OAI211_X1 U22474 ( .C1(n19512), .C2(n19380), .A(n19352), .B(n19351), .ZN(
        P3_U2952) );
  AOI22_X1 U22475 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19359), .B1(
        n19513), .B2(n19358), .ZN(n19354) );
  AOI22_X1 U22476 ( .A1(n19404), .A2(n19384), .B1(n19516), .B2(n19442), .ZN(
        n19353) );
  OAI211_X1 U22477 ( .C1(n19408), .C2(n19362), .A(n19354), .B(n19353), .ZN(
        P3_U2953) );
  AOI22_X1 U22478 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19359), .B1(
        n19521), .B2(n19358), .ZN(n19357) );
  AOI22_X1 U22479 ( .A1(n19523), .A2(n19442), .B1(n19409), .B2(n19355), .ZN(
        n19356) );
  OAI211_X1 U22480 ( .C1(n19412), .C2(n19380), .A(n19357), .B(n19356), .ZN(
        P3_U2954) );
  AOI22_X1 U22481 ( .A1(n19529), .A2(n19384), .B1(n19528), .B2(n19358), .ZN(
        n19361) );
  AOI22_X1 U22482 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19359), .B1(
        n19531), .B2(n19442), .ZN(n19360) );
  OAI211_X1 U22483 ( .C1(n19537), .C2(n19362), .A(n19361), .B(n19360), .ZN(
        P3_U2955) );
  INV_X1 U22484 ( .A(n19558), .ZN(n19364) );
  NOR2_X2 U22485 ( .A1(n19364), .A2(n19363), .ZN(n19467) );
  INV_X1 U22486 ( .A(n19467), .ZN(n19477) );
  AND2_X1 U22487 ( .A1(n19478), .A2(n19422), .ZN(n19383) );
  AOI22_X1 U22488 ( .A1(n19480), .A2(n19384), .B1(n19479), .B2(n19383), .ZN(
        n19367) );
  AOI22_X1 U22489 ( .A1(n16915), .A2(n19365), .B1(n19481), .B2(n19422), .ZN(
        n19385) );
  AOI22_X1 U22490 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19385), .B1(
        n19484), .B2(n19414), .ZN(n19366) );
  OAI211_X1 U22491 ( .C1(n19487), .C2(n19477), .A(n19367), .B(n19366), .ZN(
        P3_U2956) );
  AOI22_X1 U22492 ( .A1(n19490), .A2(n19414), .B1(n19488), .B2(n19383), .ZN(
        n19369) );
  AOI22_X1 U22493 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19385), .B1(
        n19489), .B2(n19384), .ZN(n19368) );
  OAI211_X1 U22494 ( .C1(n19493), .C2(n19477), .A(n19369), .B(n19368), .ZN(
        P3_U2957) );
  AOI22_X1 U22495 ( .A1(n19496), .A2(n19414), .B1(n19495), .B2(n19383), .ZN(
        n19371) );
  AOI22_X1 U22496 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19385), .B1(
        n19458), .B2(n19384), .ZN(n19370) );
  OAI211_X1 U22497 ( .C1(n19461), .C2(n19477), .A(n19371), .B(n19370), .ZN(
        P3_U2958) );
  AOI22_X1 U22498 ( .A1(n19501), .A2(n19383), .B1(n19431), .B2(n19384), .ZN(
        n19373) );
  AOI22_X1 U22499 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19385), .B1(
        n19503), .B2(n19467), .ZN(n19372) );
  OAI211_X1 U22500 ( .C1(n19434), .C2(n19407), .A(n19373), .B(n19372), .ZN(
        P3_U2959) );
  AOI22_X1 U22501 ( .A1(n19374), .A2(n19414), .B1(n19507), .B2(n19383), .ZN(
        n19376) );
  AOI22_X1 U22502 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19385), .B1(
        n19509), .B2(n19467), .ZN(n19375) );
  OAI211_X1 U22503 ( .C1(n19377), .C2(n19380), .A(n19376), .B(n19375), .ZN(
        P3_U2960) );
  AOI22_X1 U22504 ( .A1(n19404), .A2(n19414), .B1(n19513), .B2(n19383), .ZN(
        n19379) );
  AOI22_X1 U22505 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19385), .B1(
        n19516), .B2(n19467), .ZN(n19378) );
  OAI211_X1 U22506 ( .C1(n19408), .C2(n19380), .A(n19379), .B(n19378), .ZN(
        P3_U2961) );
  AOI22_X1 U22507 ( .A1(n19409), .A2(n19384), .B1(n19521), .B2(n19383), .ZN(
        n19382) );
  AOI22_X1 U22508 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19385), .B1(
        n19523), .B2(n19467), .ZN(n19381) );
  OAI211_X1 U22509 ( .C1(n19412), .C2(n19407), .A(n19382), .B(n19381), .ZN(
        P3_U2962) );
  AOI22_X1 U22510 ( .A1(n19443), .A2(n19384), .B1(n19528), .B2(n19383), .ZN(
        n19387) );
  AOI22_X1 U22511 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19385), .B1(
        n19531), .B2(n19467), .ZN(n19386) );
  OAI211_X1 U22512 ( .C1(n19447), .C2(n19407), .A(n19387), .B(n19386), .ZN(
        P3_U2963) );
  NAND2_X1 U22513 ( .A1(n19388), .A2(n19421), .ZN(n19536) );
  NAND2_X1 U22514 ( .A1(n19477), .A2(n19536), .ZN(n19449) );
  INV_X1 U22515 ( .A(n19449), .ZN(n19389) );
  NOR2_X1 U22516 ( .A1(n19595), .A2(n19389), .ZN(n19413) );
  AOI22_X1 U22517 ( .A1(n19484), .A2(n19442), .B1(n19479), .B2(n19413), .ZN(
        n19395) );
  INV_X1 U22518 ( .A(n19536), .ZN(n19514) );
  OAI21_X1 U22519 ( .B1(n19391), .B2(n19390), .A(n19389), .ZN(n19392) );
  OAI211_X1 U22520 ( .C1(n19514), .C2(n19690), .A(n19393), .B(n19392), .ZN(
        n19415) );
  AOI22_X1 U22521 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19415), .B1(
        n19452), .B2(n19514), .ZN(n19394) );
  OAI211_X1 U22522 ( .C1(n19455), .C2(n19407), .A(n19395), .B(n19394), .ZN(
        P3_U2964) );
  AOI22_X1 U22523 ( .A1(n19490), .A2(n19442), .B1(n19488), .B2(n19413), .ZN(
        n19397) );
  AOI22_X1 U22524 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19415), .B1(
        n19425), .B2(n19514), .ZN(n19396) );
  OAI211_X1 U22525 ( .C1(n19428), .C2(n19407), .A(n19397), .B(n19396), .ZN(
        P3_U2965) );
  AOI22_X1 U22526 ( .A1(n19458), .A2(n19414), .B1(n19495), .B2(n19413), .ZN(
        n19399) );
  AOI22_X1 U22527 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19415), .B1(
        n19496), .B2(n19442), .ZN(n19398) );
  OAI211_X1 U22528 ( .C1(n19461), .C2(n19536), .A(n19399), .B(n19398), .ZN(
        P3_U2966) );
  AOI22_X1 U22529 ( .A1(n19502), .A2(n19442), .B1(n19501), .B2(n19413), .ZN(
        n19401) );
  AOI22_X1 U22530 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19415), .B1(
        n19503), .B2(n19514), .ZN(n19400) );
  OAI211_X1 U22531 ( .C1(n19506), .C2(n19407), .A(n19401), .B(n19400), .ZN(
        P3_U2967) );
  AOI22_X1 U22532 ( .A1(n19508), .A2(n19414), .B1(n19507), .B2(n19413), .ZN(
        n19403) );
  AOI22_X1 U22533 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19415), .B1(
        n19509), .B2(n19514), .ZN(n19402) );
  OAI211_X1 U22534 ( .C1(n19512), .C2(n19441), .A(n19403), .B(n19402), .ZN(
        P3_U2968) );
  AOI22_X1 U22535 ( .A1(n19404), .A2(n19442), .B1(n19513), .B2(n19413), .ZN(
        n19406) );
  AOI22_X1 U22536 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19415), .B1(
        n19516), .B2(n19514), .ZN(n19405) );
  OAI211_X1 U22537 ( .C1(n19408), .C2(n19407), .A(n19406), .B(n19405), .ZN(
        P3_U2969) );
  AOI22_X1 U22538 ( .A1(n19409), .A2(n19414), .B1(n19521), .B2(n19413), .ZN(
        n19411) );
  AOI22_X1 U22539 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19415), .B1(
        n19523), .B2(n19514), .ZN(n19410) );
  OAI211_X1 U22540 ( .C1(n19412), .C2(n19441), .A(n19411), .B(n19410), .ZN(
        P3_U2970) );
  AOI22_X1 U22541 ( .A1(n19443), .A2(n19414), .B1(n19528), .B2(n19413), .ZN(
        n19417) );
  AOI22_X1 U22542 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19415), .B1(
        n19531), .B2(n19514), .ZN(n19416) );
  OAI211_X1 U22543 ( .C1(n19447), .C2(n19441), .A(n19417), .B(n19416), .ZN(
        P3_U2971) );
  NOR2_X1 U22544 ( .A1(n19419), .A2(n19418), .ZN(n19483) );
  AOI22_X1 U22545 ( .A1(n19480), .A2(n19442), .B1(n19479), .B2(n19483), .ZN(
        n19424) );
  AOI22_X1 U22546 ( .A1(n16915), .A2(n19422), .B1(n19421), .B2(n19420), .ZN(
        n19444) );
  AOI22_X1 U22547 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19444), .B1(
        n19484), .B2(n19467), .ZN(n19423) );
  OAI211_X1 U22548 ( .C1(n19520), .C2(n19487), .A(n19424), .B(n19423), .ZN(
        P3_U2972) );
  AOI22_X1 U22549 ( .A1(n19490), .A2(n19467), .B1(n19488), .B2(n19483), .ZN(
        n19427) );
  AOI22_X1 U22550 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19444), .B1(
        n19530), .B2(n19425), .ZN(n19426) );
  OAI211_X1 U22551 ( .C1(n19428), .C2(n19441), .A(n19427), .B(n19426), .ZN(
        P3_U2973) );
  AOI22_X1 U22552 ( .A1(n19496), .A2(n19467), .B1(n19495), .B2(n19483), .ZN(
        n19430) );
  AOI22_X1 U22553 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19444), .B1(
        n19530), .B2(n19497), .ZN(n19429) );
  OAI211_X1 U22554 ( .C1(n19500), .C2(n19441), .A(n19430), .B(n19429), .ZN(
        P3_U2974) );
  AOI22_X1 U22555 ( .A1(n19501), .A2(n19483), .B1(n19431), .B2(n19442), .ZN(
        n19433) );
  AOI22_X1 U22556 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19444), .B1(
        n19530), .B2(n19503), .ZN(n19432) );
  OAI211_X1 U22557 ( .C1(n19434), .C2(n19477), .A(n19433), .B(n19432), .ZN(
        P3_U2975) );
  AOI22_X1 U22558 ( .A1(n19508), .A2(n19442), .B1(n19507), .B2(n19483), .ZN(
        n19436) );
  AOI22_X1 U22559 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19444), .B1(
        n19530), .B2(n19509), .ZN(n19435) );
  OAI211_X1 U22560 ( .C1(n19512), .C2(n19477), .A(n19436), .B(n19435), .ZN(
        P3_U2976) );
  AOI22_X1 U22561 ( .A1(n19515), .A2(n19442), .B1(n19513), .B2(n19483), .ZN(
        n19438) );
  AOI22_X1 U22562 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19444), .B1(
        n19530), .B2(n19516), .ZN(n19437) );
  OAI211_X1 U22563 ( .C1(n19519), .C2(n19477), .A(n19438), .B(n19437), .ZN(
        P3_U2977) );
  AOI22_X1 U22564 ( .A1(n19522), .A2(n19467), .B1(n19521), .B2(n19483), .ZN(
        n19440) );
  AOI22_X1 U22565 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19444), .B1(
        n19530), .B2(n19523), .ZN(n19439) );
  OAI211_X1 U22566 ( .C1(n19526), .C2(n19441), .A(n19440), .B(n19439), .ZN(
        P3_U2978) );
  AOI22_X1 U22567 ( .A1(n19443), .A2(n19442), .B1(n19528), .B2(n19483), .ZN(
        n19446) );
  AOI22_X1 U22568 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19444), .B1(
        n19530), .B2(n19531), .ZN(n19445) );
  OAI211_X1 U22569 ( .C1(n19447), .C2(n19477), .A(n19446), .B(n19445), .ZN(
        P3_U2979) );
  OAI221_X1 U22570 ( .B1(n19451), .B2(n19450), .C1(n19451), .C2(n19449), .A(
        n19448), .ZN(n19473) );
  AND2_X1 U22571 ( .A1(n19478), .A2(n19451), .ZN(n19472) );
  AOI22_X1 U22572 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19473), .B1(
        n19479), .B2(n19472), .ZN(n19454) );
  AOI22_X1 U22573 ( .A1(n19474), .A2(n19452), .B1(n19484), .B2(n19514), .ZN(
        n19453) );
  OAI211_X1 U22574 ( .C1(n19455), .C2(n19477), .A(n19454), .B(n19453), .ZN(
        P3_U2980) );
  AOI22_X1 U22575 ( .A1(n19489), .A2(n19467), .B1(n19488), .B2(n19472), .ZN(
        n19457) );
  AOI22_X1 U22576 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19473), .B1(
        n19490), .B2(n19514), .ZN(n19456) );
  OAI211_X1 U22577 ( .C1(n19462), .C2(n19493), .A(n19457), .B(n19456), .ZN(
        P3_U2981) );
  AOI22_X1 U22578 ( .A1(n19458), .A2(n19467), .B1(n19495), .B2(n19472), .ZN(
        n19460) );
  AOI22_X1 U22579 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19473), .B1(
        n19496), .B2(n19514), .ZN(n19459) );
  OAI211_X1 U22580 ( .C1(n19462), .C2(n19461), .A(n19460), .B(n19459), .ZN(
        P3_U2982) );
  AOI22_X1 U22581 ( .A1(n19502), .A2(n19514), .B1(n19501), .B2(n19472), .ZN(
        n19464) );
  AOI22_X1 U22582 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19473), .B1(
        n19474), .B2(n19503), .ZN(n19463) );
  OAI211_X1 U22583 ( .C1(n19506), .C2(n19477), .A(n19464), .B(n19463), .ZN(
        P3_U2983) );
  AOI22_X1 U22584 ( .A1(n19508), .A2(n19467), .B1(n19507), .B2(n19472), .ZN(
        n19466) );
  AOI22_X1 U22585 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19473), .B1(
        n19474), .B2(n19509), .ZN(n19465) );
  OAI211_X1 U22586 ( .C1(n19512), .C2(n19536), .A(n19466), .B(n19465), .ZN(
        P3_U2984) );
  AOI22_X1 U22587 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19473), .B1(
        n19513), .B2(n19472), .ZN(n19469) );
  AOI22_X1 U22588 ( .A1(n19474), .A2(n19516), .B1(n19515), .B2(n19467), .ZN(
        n19468) );
  OAI211_X1 U22589 ( .C1(n19519), .C2(n19536), .A(n19469), .B(n19468), .ZN(
        P3_U2985) );
  AOI22_X1 U22590 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19473), .B1(
        n19521), .B2(n19472), .ZN(n19471) );
  AOI22_X1 U22591 ( .A1(n19474), .A2(n19523), .B1(n19522), .B2(n19514), .ZN(
        n19470) );
  OAI211_X1 U22592 ( .C1(n19526), .C2(n19477), .A(n19471), .B(n19470), .ZN(
        P3_U2986) );
  AOI22_X1 U22593 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19473), .B1(
        n19528), .B2(n19472), .ZN(n19476) );
  AOI22_X1 U22594 ( .A1(n19474), .A2(n19531), .B1(n19529), .B2(n19514), .ZN(
        n19475) );
  OAI211_X1 U22595 ( .C1(n19537), .C2(n19477), .A(n19476), .B(n19475), .ZN(
        P3_U2987) );
  AND2_X1 U22596 ( .A1(n19478), .A2(n19482), .ZN(n19527) );
  AOI22_X1 U22597 ( .A1(n19480), .A2(n19514), .B1(n19479), .B2(n19527), .ZN(
        n19486) );
  AOI22_X1 U22598 ( .A1(n16915), .A2(n19483), .B1(n19482), .B2(n19481), .ZN(
        n19533) );
  AOI22_X1 U22599 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19533), .B1(
        n19530), .B2(n19484), .ZN(n19485) );
  OAI211_X1 U22600 ( .C1(n19494), .C2(n19487), .A(n19486), .B(n19485), .ZN(
        P3_U2988) );
  AOI22_X1 U22601 ( .A1(n19489), .A2(n19514), .B1(n19488), .B2(n19527), .ZN(
        n19492) );
  AOI22_X1 U22602 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19533), .B1(
        n19530), .B2(n19490), .ZN(n19491) );
  OAI211_X1 U22603 ( .C1(n19494), .C2(n19493), .A(n19492), .B(n19491), .ZN(
        P3_U2989) );
  AOI22_X1 U22604 ( .A1(n19530), .A2(n19496), .B1(n19495), .B2(n19527), .ZN(
        n19499) );
  AOI22_X1 U22605 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19497), .ZN(n19498) );
  OAI211_X1 U22606 ( .C1(n19500), .C2(n19536), .A(n19499), .B(n19498), .ZN(
        P3_U2990) );
  AOI22_X1 U22607 ( .A1(n19530), .A2(n19502), .B1(n19501), .B2(n19527), .ZN(
        n19505) );
  AOI22_X1 U22608 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19503), .ZN(n19504) );
  OAI211_X1 U22609 ( .C1(n19506), .C2(n19536), .A(n19505), .B(n19504), .ZN(
        P3_U2991) );
  AOI22_X1 U22610 ( .A1(n19508), .A2(n19514), .B1(n19507), .B2(n19527), .ZN(
        n19511) );
  AOI22_X1 U22611 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19509), .ZN(n19510) );
  OAI211_X1 U22612 ( .C1(n19520), .C2(n19512), .A(n19511), .B(n19510), .ZN(
        P3_U2992) );
  AOI22_X1 U22613 ( .A1(n19515), .A2(n19514), .B1(n19513), .B2(n19527), .ZN(
        n19518) );
  AOI22_X1 U22614 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19516), .ZN(n19517) );
  OAI211_X1 U22615 ( .C1(n19520), .C2(n19519), .A(n19518), .B(n19517), .ZN(
        P3_U2993) );
  AOI22_X1 U22616 ( .A1(n19530), .A2(n19522), .B1(n19521), .B2(n19527), .ZN(
        n19525) );
  AOI22_X1 U22617 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19523), .ZN(n19524) );
  OAI211_X1 U22618 ( .C1(n19526), .C2(n19536), .A(n19525), .B(n19524), .ZN(
        P3_U2994) );
  AOI22_X1 U22619 ( .A1(n19530), .A2(n19529), .B1(n19528), .B2(n19527), .ZN(
        n19535) );
  AOI22_X1 U22620 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19533), .B1(
        n19532), .B2(n19531), .ZN(n19534) );
  OAI211_X1 U22621 ( .C1(n19537), .C2(n19536), .A(n19535), .B(n19534), .ZN(
        P3_U2995) );
  NAND2_X1 U22622 ( .A1(n19539), .A2(n19538), .ZN(n19540) );
  AOI22_X1 U22623 ( .A1(n19543), .A2(n19542), .B1(n19541), .B2(n19540), .ZN(
        n19544) );
  OAI221_X1 U22624 ( .B1(n19547), .B2(n19546), .C1(n19547), .C2(n19545), .A(
        n19544), .ZN(n19701) );
  OAI21_X1 U22625 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19548), .ZN(n19549) );
  OAI211_X1 U22626 ( .C1(n19557), .C2(n19551), .A(n19550), .B(n19549), .ZN(
        n19576) );
  NAND2_X1 U22627 ( .A1(n19557), .A2(n19552), .ZN(n19553) );
  AOI22_X1 U22628 ( .A1(n19557), .A2(n19554), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19553), .ZN(n19574) );
  INV_X1 U22629 ( .A(n19555), .ZN(n19556) );
  INV_X1 U22630 ( .A(n19557), .ZN(n19566) );
  AOI22_X1 U22631 ( .A1(n19557), .A2(n19556), .B1(n19566), .B2(n9940), .ZN(
        n19569) );
  NAND2_X1 U22632 ( .A1(n19559), .A2(n19558), .ZN(n19561) );
  INV_X1 U22633 ( .A(n19559), .ZN(n19560) );
  AOI22_X1 U22634 ( .A1(n19562), .A2(n19561), .B1(n11652), .B2(n19560), .ZN(
        n19565) );
  NAND2_X1 U22635 ( .A1(n19569), .A2(n19568), .ZN(n19564) );
  OAI211_X1 U22636 ( .C1(n19566), .C2(n19565), .A(n19564), .B(n19563), .ZN(
        n19567) );
  OAI211_X1 U22637 ( .C1(n19568), .C2(n19569), .A(n19567), .B(n19571), .ZN(
        n19573) );
  AOI21_X1 U22638 ( .B1(n19571), .B2(n19570), .A(n19569), .ZN(n19572) );
  AOI222_X1 U22639 ( .A1(n19574), .A2(n19573), .B1(n19574), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19573), .C2(n19572), .ZN(
        n19575) );
  NOR4_X1 U22640 ( .A1(n19577), .A2(n19701), .A3(n19576), .A4(n19575), .ZN(
        n19589) );
  AOI22_X1 U22641 ( .A1(n19578), .A2(n19712), .B1(n19705), .B2(n18488), .ZN(
        n19579) );
  INV_X1 U22642 ( .A(n19579), .ZN(n19585) );
  OAI211_X1 U22643 ( .C1(n19581), .C2(n19580), .A(n19703), .B(n19589), .ZN(
        n19689) );
  NAND2_X1 U22644 ( .A1(n19705), .A2(n19582), .ZN(n19590) );
  NAND2_X1 U22645 ( .A1(n19689), .A2(n19590), .ZN(n19593) );
  NOR2_X1 U22646 ( .A1(n19583), .A2(n19593), .ZN(n19584) );
  MUX2_X1 U22647 ( .A(n19585), .B(n19584), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19587) );
  OAI211_X1 U22648 ( .C1(n19589), .C2(n19588), .A(n19587), .B(n19586), .ZN(
        P3_U2996) );
  NOR2_X1 U22649 ( .A1(n19710), .A2(n19704), .ZN(n19597) );
  NOR3_X1 U22650 ( .A1(n19592), .A2(n19591), .A3(n19590), .ZN(n19600) );
  NOR3_X1 U22651 ( .A1(n19595), .A2(n19594), .A3(n19593), .ZN(n19596) );
  OR4_X1 U22652 ( .A1(n19598), .A2(n19597), .A3(n19600), .A4(n19596), .ZN(
        P3_U2997) );
  NOR4_X1 U22653 ( .A1(n19712), .A2(n19601), .A3(n19600), .A4(n19599), .ZN(
        P3_U2998) );
  AND2_X1 U22654 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19602), .ZN(
        P3_U2999) );
  AND2_X1 U22655 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19602), .ZN(
        P3_U3000) );
  AND2_X1 U22656 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19602), .ZN(
        P3_U3001) );
  AND2_X1 U22657 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19602), .ZN(
        P3_U3002) );
  AND2_X1 U22658 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19602), .ZN(
        P3_U3003) );
  AND2_X1 U22659 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19602), .ZN(
        P3_U3004) );
  AND2_X1 U22660 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19602), .ZN(
        P3_U3005) );
  AND2_X1 U22661 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19602), .ZN(
        P3_U3006) );
  AND2_X1 U22662 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19602), .ZN(
        P3_U3007) );
  AND2_X1 U22663 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19602), .ZN(
        P3_U3008) );
  AND2_X1 U22664 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19602), .ZN(
        P3_U3009) );
  AND2_X1 U22665 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19602), .ZN(
        P3_U3010) );
  AND2_X1 U22666 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19602), .ZN(
        P3_U3011) );
  AND2_X1 U22667 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19602), .ZN(
        P3_U3012) );
  AND2_X1 U22668 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19602), .ZN(
        P3_U3013) );
  AND2_X1 U22669 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19602), .ZN(
        P3_U3014) );
  AND2_X1 U22670 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19602), .ZN(
        P3_U3015) );
  AND2_X1 U22671 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19602), .ZN(
        P3_U3016) );
  AND2_X1 U22672 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19602), .ZN(
        P3_U3017) );
  AND2_X1 U22673 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19602), .ZN(
        P3_U3018) );
  AND2_X1 U22674 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19602), .ZN(
        P3_U3019) );
  AND2_X1 U22675 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19602), .ZN(
        P3_U3020) );
  INV_X1 U22676 ( .A(P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21468) );
  NOR2_X1 U22677 ( .A1(n21468), .A2(n19687), .ZN(P3_U3021) );
  AND2_X1 U22678 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19602), .ZN(P3_U3022) );
  AND2_X1 U22679 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19602), .ZN(P3_U3023) );
  AND2_X1 U22680 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19602), .ZN(P3_U3024) );
  AND2_X1 U22681 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19602), .ZN(P3_U3025) );
  AND2_X1 U22682 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19602), .ZN(P3_U3026) );
  INV_X1 U22683 ( .A(P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21446) );
  NOR2_X1 U22684 ( .A1(n21446), .A2(n19687), .ZN(P3_U3027) );
  AND2_X1 U22685 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19602), .ZN(P3_U3028) );
  NOR2_X1 U22686 ( .A1(n19618), .A2(n21363), .ZN(n19613) );
  INV_X1 U22687 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19606) );
  AOI211_X1 U22688 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n19613), .B(
        n19606), .ZN(n19605) );
  AOI21_X1 U22689 ( .B1(n19705), .B2(P3_STATE_REG_1__SCAN_IN), .A(n19615), 
        .ZN(n19617) );
  OAI21_X1 U22690 ( .B1(n21362), .B2(n19603), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19616) );
  INV_X1 U22691 ( .A(n19616), .ZN(n19604) );
  OAI22_X1 U22692 ( .A1(n19682), .A2(n19605), .B1(n19617), .B2(n19604), .ZN(
        P3_U3029) );
  NOR2_X1 U22693 ( .A1(n19613), .A2(n19606), .ZN(n19609) );
  NOR2_X1 U22694 ( .A1(n19607), .A2(n21363), .ZN(n19608) );
  AOI22_X1 U22695 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19609), .B1(n19608), 
        .B2(n19618), .ZN(n19610) );
  NAND2_X1 U22696 ( .A1(n19705), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19611) );
  NAND3_X1 U22697 ( .A1(n19610), .A2(n19708), .A3(n19611), .ZN(P3_U3030) );
  OAI22_X1 U22698 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19611), .ZN(n19612) );
  OAI22_X1 U22699 ( .A1(n19613), .A2(n19612), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19614) );
  OAI22_X1 U22700 ( .A1(n19617), .A2(n19616), .B1(n19615), .B2(n19614), .ZN(
        P3_U3031) );
  NAND2_X2 U22701 ( .A1(n19682), .A2(n19618), .ZN(n19674) );
  OAI222_X1 U22702 ( .A1(n21537), .A2(n19678), .B1(n19619), .B2(n19682), .C1(
        n19620), .C2(n19674), .ZN(P3_U3032) );
  INV_X1 U22703 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19622) );
  OAI222_X1 U22704 ( .A1(n19674), .A2(n19622), .B1(n19621), .B2(n19682), .C1(
        n19620), .C2(n19678), .ZN(P3_U3033) );
  OAI222_X1 U22705 ( .A1(n19674), .A2(n19624), .B1(n19623), .B2(n19682), .C1(
        n19622), .C2(n19678), .ZN(P3_U3034) );
  OAI222_X1 U22706 ( .A1(n19674), .A2(n19626), .B1(n19625), .B2(n19682), .C1(
        n19624), .C2(n19678), .ZN(P3_U3035) );
  OAI222_X1 U22707 ( .A1(n19674), .A2(n19628), .B1(n19627), .B2(n19682), .C1(
        n19626), .C2(n19678), .ZN(P3_U3036) );
  OAI222_X1 U22708 ( .A1(n19674), .A2(n19630), .B1(n19629), .B2(n19682), .C1(
        n19628), .C2(n19678), .ZN(P3_U3037) );
  OAI222_X1 U22709 ( .A1(n19674), .A2(n19633), .B1(n19631), .B2(n19682), .C1(
        n19630), .C2(n19678), .ZN(P3_U3038) );
  OAI222_X1 U22710 ( .A1(n19633), .A2(n19678), .B1(n19632), .B2(n19682), .C1(
        n19634), .C2(n19674), .ZN(P3_U3039) );
  OAI222_X1 U22711 ( .A1(n19674), .A2(n19636), .B1(n19635), .B2(n19682), .C1(
        n19634), .C2(n19678), .ZN(P3_U3040) );
  OAI222_X1 U22712 ( .A1(n19674), .A2(n19638), .B1(n19637), .B2(n19682), .C1(
        n19636), .C2(n19678), .ZN(P3_U3041) );
  OAI222_X1 U22713 ( .A1(n19674), .A2(n19640), .B1(n19639), .B2(n19682), .C1(
        n19638), .C2(n19678), .ZN(P3_U3042) );
  OAI222_X1 U22714 ( .A1(n19674), .A2(n19642), .B1(n19641), .B2(n19682), .C1(
        n19640), .C2(n19678), .ZN(P3_U3043) );
  INV_X1 U22715 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19645) );
  OAI222_X1 U22716 ( .A1(n19674), .A2(n19645), .B1(n19643), .B2(n19682), .C1(
        n19642), .C2(n19678), .ZN(P3_U3044) );
  OAI222_X1 U22717 ( .A1(n19645), .A2(n19678), .B1(n19644), .B2(n19682), .C1(
        n19646), .C2(n19674), .ZN(P3_U3045) );
  OAI222_X1 U22718 ( .A1(n19674), .A2(n19648), .B1(n19647), .B2(n19682), .C1(
        n19646), .C2(n19678), .ZN(P3_U3046) );
  OAI222_X1 U22719 ( .A1(n19674), .A2(n19650), .B1(n19649), .B2(n19682), .C1(
        n19648), .C2(n19678), .ZN(P3_U3047) );
  OAI222_X1 U22720 ( .A1(n19674), .A2(n19652), .B1(n19651), .B2(n19682), .C1(
        n19650), .C2(n19678), .ZN(P3_U3048) );
  OAI222_X1 U22721 ( .A1(n19674), .A2(n19654), .B1(n19653), .B2(n19682), .C1(
        n19652), .C2(n19678), .ZN(P3_U3049) );
  OAI222_X1 U22722 ( .A1(n19674), .A2(n19657), .B1(n19655), .B2(n19682), .C1(
        n19654), .C2(n19678), .ZN(P3_U3050) );
  OAI222_X1 U22723 ( .A1(n19657), .A2(n19678), .B1(n19656), .B2(n19682), .C1(
        n19658), .C2(n19674), .ZN(P3_U3051) );
  INV_X1 U22724 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19660) );
  OAI222_X1 U22725 ( .A1(n19674), .A2(n19660), .B1(n19659), .B2(n19682), .C1(
        n19658), .C2(n19678), .ZN(P3_U3052) );
  OAI222_X1 U22726 ( .A1(n19674), .A2(n19663), .B1(n19661), .B2(n19682), .C1(
        n19660), .C2(n19678), .ZN(P3_U3053) );
  OAI222_X1 U22727 ( .A1(n19663), .A2(n19678), .B1(n19662), .B2(n19682), .C1(
        n19664), .C2(n19674), .ZN(P3_U3054) );
  OAI222_X1 U22728 ( .A1(n19674), .A2(n19666), .B1(n19665), .B2(n19682), .C1(
        n19664), .C2(n19678), .ZN(P3_U3055) );
  INV_X1 U22729 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19668) );
  OAI222_X1 U22730 ( .A1(n19674), .A2(n19668), .B1(n19667), .B2(n19682), .C1(
        n19666), .C2(n19678), .ZN(P3_U3056) );
  OAI222_X1 U22731 ( .A1(n19674), .A2(n19670), .B1(n19669), .B2(n19682), .C1(
        n19668), .C2(n19678), .ZN(P3_U3057) );
  OAI222_X1 U22732 ( .A1(n19674), .A2(n17109), .B1(n19671), .B2(n19682), .C1(
        n19670), .C2(n19678), .ZN(P3_U3058) );
  OAI222_X1 U22733 ( .A1(n17109), .A2(n19678), .B1(n19672), .B2(n19682), .C1(
        n17089), .C2(n19674), .ZN(P3_U3059) );
  OAI222_X1 U22734 ( .A1(n19674), .A2(n19677), .B1(n19673), .B2(n19682), .C1(
        n17089), .C2(n19678), .ZN(P3_U3060) );
  OAI222_X1 U22735 ( .A1(n19678), .A2(n19677), .B1(n19676), .B2(n19682), .C1(
        n19675), .C2(n19674), .ZN(P3_U3061) );
  OAI22_X1 U22736 ( .A1(n19717), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19682), .ZN(n19679) );
  INV_X1 U22737 ( .A(n19679), .ZN(P3_U3274) );
  OAI22_X1 U22738 ( .A1(n19717), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19682), .ZN(n19680) );
  INV_X1 U22739 ( .A(n19680), .ZN(P3_U3275) );
  OAI22_X1 U22740 ( .A1(n19717), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19682), .ZN(n19681) );
  INV_X1 U22741 ( .A(n19681), .ZN(P3_U3276) );
  OAI22_X1 U22742 ( .A1(n19717), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19682), .ZN(n19683) );
  INV_X1 U22743 ( .A(n19683), .ZN(P3_U3277) );
  OAI21_X1 U22744 ( .B1(n19687), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19685), 
        .ZN(n19684) );
  INV_X1 U22745 ( .A(n19684), .ZN(P3_U3280) );
  OAI21_X1 U22746 ( .B1(n19687), .B2(n19686), .A(n19685), .ZN(P3_U3281) );
  OAI221_X1 U22747 ( .B1(n19690), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19690), 
        .C2(n19689), .A(n19688), .ZN(P3_U3282) );
  AOI21_X1 U22748 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19691) );
  AOI22_X1 U22749 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19691), .B2(n21537), .ZN(n19693) );
  INV_X1 U22750 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19692) );
  AOI22_X1 U22751 ( .A1(n19694), .A2(n19693), .B1(n19692), .B2(n19697), .ZN(
        P3_U3292) );
  INV_X1 U22752 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19698) );
  NOR2_X1 U22753 ( .A1(n19697), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19695) );
  AOI22_X1 U22754 ( .A1(n19698), .A2(n19697), .B1(n19696), .B2(n19695), .ZN(
        P3_U3293) );
  INV_X1 U22755 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19699) );
  AOI22_X1 U22756 ( .A1(n19682), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19699), 
        .B2(n19717), .ZN(P3_U3294) );
  MUX2_X1 U22757 ( .A(P3_MORE_REG_SCAN_IN), .B(n19701), .S(n19700), .Z(
        P3_U3295) );
  OAI22_X1 U22758 ( .A1(n19705), .A2(n19704), .B1(n19703), .B2(n19702), .ZN(
        n19706) );
  NOR2_X1 U22759 ( .A1(n19707), .A2(n19706), .ZN(n19716) );
  AOI21_X1 U22760 ( .B1(n19709), .B2(n21509), .A(n19708), .ZN(n19711) );
  OAI211_X1 U22761 ( .C1(n19711), .C2(n19721), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19710), .ZN(n19713) );
  AOI21_X1 U22762 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19713), .A(n19712), 
        .ZN(n19715) );
  NAND2_X1 U22763 ( .A1(n19716), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19714) );
  OAI21_X1 U22764 ( .B1(n19716), .B2(n19715), .A(n19714), .ZN(P3_U3296) );
  OAI22_X1 U22765 ( .A1(n19717), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19682), .ZN(n19718) );
  INV_X1 U22766 ( .A(n19718), .ZN(P3_U3297) );
  OAI21_X1 U22767 ( .B1(n19719), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n19720), 
        .ZN(n19724) );
  OAI22_X1 U22768 ( .A1(n19721), .A2(n19720), .B1(n19724), .B2(
        P3_READREQUEST_REG_SCAN_IN), .ZN(n19722) );
  INV_X1 U22769 ( .A(n19722), .ZN(P3_U3298) );
  OAI21_X1 U22770 ( .B1(n19724), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19723), 
        .ZN(n19725) );
  INV_X1 U22771 ( .A(n19725), .ZN(P3_U3299) );
  INV_X1 U22772 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19732) );
  NAND2_X1 U22773 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20540), .ZN(n20530) );
  NAND2_X1 U22774 ( .A1(n19732), .A2(n19726), .ZN(n20527) );
  OAI21_X1 U22775 ( .B1(n19732), .B2(n20530), .A(n20527), .ZN(n20606) );
  AOI21_X1 U22776 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20606), .ZN(n19727) );
  INV_X1 U22777 ( .A(n19727), .ZN(P2_U2815) );
  AOI22_X1 U22778 ( .A1(n19730), .A2(n19729), .B1(n19728), .B2(
        P2_CODEFETCH_REG_SCAN_IN), .ZN(n19731) );
  INV_X1 U22779 ( .A(n19731), .ZN(P2_U2816) );
  NAND2_X1 U22780 ( .A1(n19732), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20638) );
  INV_X2 U22781 ( .A(n20638), .ZN(n20597) );
  INV_X1 U22782 ( .A(n19734), .ZN(n20535) );
  NAND2_X1 U22783 ( .A1(n20535), .A2(n20638), .ZN(n20524) );
  AOI21_X1 U22784 ( .B1(n19732), .B2(n20524), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19733) );
  AOI21_X1 U22785 ( .B1(n20597), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n19733), 
        .ZN(P2_U2817) );
  OAI21_X1 U22786 ( .B1(n19734), .B2(BS16), .A(n20606), .ZN(n20604) );
  OAI21_X1 U22787 ( .B1(n20606), .B2(n20408), .A(n20604), .ZN(P2_U2818) );
  NOR4_X1 U22788 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19738) );
  NOR4_X1 U22789 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19737) );
  NOR4_X1 U22790 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19736) );
  NOR4_X1 U22791 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19735) );
  NAND4_X1 U22792 ( .A1(n19738), .A2(n19737), .A3(n19736), .A4(n19735), .ZN(
        n19744) );
  NOR4_X1 U22793 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19742) );
  AOI211_X1 U22794 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19741) );
  NOR4_X1 U22795 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19740) );
  NOR4_X1 U22796 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19739) );
  NAND4_X1 U22797 ( .A1(n19742), .A2(n19741), .A3(n19740), .A4(n19739), .ZN(
        n19743) );
  NOR2_X1 U22798 ( .A1(n19744), .A2(n19743), .ZN(n19754) );
  INV_X1 U22799 ( .A(n19754), .ZN(n19753) );
  NOR2_X1 U22800 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19753), .ZN(n19747) );
  INV_X1 U22801 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19745) );
  AOI22_X1 U22802 ( .A1(n19747), .A2(n19748), .B1(n19753), .B2(n19745), .ZN(
        P2_U2820) );
  OR3_X1 U22803 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19752) );
  INV_X1 U22804 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19746) );
  AOI22_X1 U22805 ( .A1(n19747), .A2(n19752), .B1(n19753), .B2(n19746), .ZN(
        P2_U2821) );
  INV_X1 U22806 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20605) );
  NAND2_X1 U22807 ( .A1(n19747), .A2(n20605), .ZN(n19751) );
  OAI21_X1 U22808 ( .B1(n19748), .B2(n20542), .A(n19754), .ZN(n19749) );
  OAI21_X1 U22809 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19754), .A(n19749), 
        .ZN(n19750) );
  OAI221_X1 U22810 ( .B1(n19751), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19751), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19750), .ZN(P2_U2822) );
  INV_X1 U22811 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21538) );
  OAI221_X1 U22812 ( .B1(n19754), .B2(n21538), .C1(n19753), .C2(n19752), .A(
        n19751), .ZN(P2_U2823) );
  AOI22_X1 U22813 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19841), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n19830), .ZN(n19770) );
  INV_X1 U22814 ( .A(n19755), .ZN(n19759) );
  AOI21_X1 U22815 ( .B1(n19827), .B2(P2_REIP_REG_11__SCAN_IN), .A(n16423), 
        .ZN(n19756) );
  OAI21_X1 U22816 ( .B1(n19757), .B2(n19809), .A(n19756), .ZN(n19758) );
  AOI21_X1 U22817 ( .B1(n19759), .B2(n19812), .A(n19758), .ZN(n19769) );
  INV_X1 U22818 ( .A(n19760), .ZN(n19761) );
  AOI22_X1 U22819 ( .A1(n19842), .A2(n19762), .B1(n19836), .B2(n19761), .ZN(
        n19768) );
  INV_X1 U22820 ( .A(n19763), .ZN(n19766) );
  OAI211_X1 U22821 ( .C1(n19766), .C2(n19765), .A(n19764), .B(n19820), .ZN(
        n19767) );
  NAND4_X1 U22822 ( .A1(n19770), .A2(n19769), .A3(n19768), .A4(n19767), .ZN(
        P2_U2844) );
  AOI21_X1 U22823 ( .B1(n19827), .B2(P2_REIP_REG_9__SCAN_IN), .A(n16423), .ZN(
        n19771) );
  OAI21_X1 U22824 ( .B1(n19773), .B2(n19772), .A(n19771), .ZN(n19774) );
  AOI21_X1 U22825 ( .B1(n19775), .B2(n19829), .A(n19774), .ZN(n19787) );
  NOR2_X1 U22826 ( .A1(n19777), .A2(n19776), .ZN(n19784) );
  NOR2_X1 U22827 ( .A1(n19778), .A2(n19779), .ZN(n19780) );
  MUX2_X1 U22828 ( .A(n19780), .B(n19779), .S(n19815), .Z(n19782) );
  NOR3_X1 U22829 ( .A1(n19782), .A2(n19781), .A3(n19838), .ZN(n19783) );
  AOI211_X1 U22830 ( .C1(n19785), .C2(n19812), .A(n19784), .B(n19783), .ZN(
        n19786) );
  OAI211_X1 U22831 ( .C1(n19788), .C2(n19803), .A(n19787), .B(n19786), .ZN(
        P2_U2846) );
  AOI21_X1 U22832 ( .B1(n19827), .B2(P2_REIP_REG_5__SCAN_IN), .A(n16423), .ZN(
        n19790) );
  NAND2_X1 U22833 ( .A1(n19830), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n19789) );
  OAI211_X1 U22834 ( .C1(n19791), .C2(n19809), .A(n19790), .B(n19789), .ZN(
        n19792) );
  INV_X1 U22835 ( .A(n19792), .ZN(n19802) );
  NOR2_X1 U22836 ( .A1(n19793), .A2(n19833), .ZN(n19799) );
  NOR2_X1 U22837 ( .A1(n19818), .A2(n19794), .ZN(n19795) );
  MUX2_X1 U22838 ( .A(n19795), .B(n19794), .S(n19815), .Z(n19797) );
  NOR3_X1 U22839 ( .A1(n19797), .A2(n19796), .A3(n19838), .ZN(n19798) );
  AOI211_X1 U22840 ( .C1(n19800), .C2(n19836), .A(n19799), .B(n19798), .ZN(
        n19801) );
  OAI211_X1 U22841 ( .C1(n12468), .C2(n19803), .A(n19802), .B(n19801), .ZN(
        P2_U2850) );
  NAND2_X1 U22842 ( .A1(n19841), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19807) );
  OAI21_X1 U22843 ( .B1(n19804), .B2(n20546), .A(n10176), .ZN(n19805) );
  INV_X1 U22844 ( .A(n19805), .ZN(n19806) );
  OAI211_X1 U22845 ( .C1(n19809), .C2(n19808), .A(n19807), .B(n19806), .ZN(
        n19810) );
  INV_X1 U22846 ( .A(n19810), .ZN(n19825) );
  INV_X1 U22847 ( .A(n19811), .ZN(n19876) );
  AOI22_X1 U22848 ( .A1(n19876), .A2(n19812), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n19830), .ZN(n19824) );
  AOI22_X1 U22849 ( .A1(n19864), .A2(n19813), .B1(n19836), .B2(n19862), .ZN(
        n19823) );
  NAND2_X1 U22850 ( .A1(n19814), .A2(n19816), .ZN(n19817) );
  MUX2_X1 U22851 ( .A(n19817), .B(n19816), .S(n19815), .Z(n19821) );
  INV_X1 U22852 ( .A(n19818), .ZN(n19819) );
  NAND3_X1 U22853 ( .A1(n19821), .A2(n19820), .A3(n19819), .ZN(n19822) );
  NAND4_X1 U22854 ( .A1(n19825), .A2(n19824), .A3(n19823), .A4(n19822), .ZN(
        P2_U2851) );
  INV_X1 U22855 ( .A(n19826), .ZN(n19834) );
  AOI22_X1 U22856 ( .A1(n19829), .A2(n19828), .B1(n19827), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n19832) );
  NAND2_X1 U22857 ( .A1(n19830), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n19831) );
  OAI211_X1 U22858 ( .C1(n19834), .C2(n19833), .A(n19832), .B(n19831), .ZN(
        n19835) );
  OAI22_X1 U22859 ( .A1(n19839), .A2(n19838), .B1(n19837), .B2(n20622), .ZN(
        n19840) );
  INV_X1 U22860 ( .A(n19840), .ZN(n19844) );
  OAI21_X1 U22861 ( .B1(n19842), .B2(n19841), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19843) );
  NAND3_X1 U22862 ( .A1(n19845), .A2(n19844), .A3(n19843), .ZN(P2_U2855) );
  AOI21_X1 U22863 ( .B1(n19848), .B2(n19847), .A(n19846), .ZN(n19850) );
  INV_X1 U22864 ( .A(n16028), .ZN(n19849) );
  NOR2_X1 U22865 ( .A1(n19850), .A2(n19849), .ZN(n19872) );
  AOI22_X1 U22866 ( .A1(n19851), .A2(n19866), .B1(n19863), .B2(n19872), .ZN(
        n19852) );
  OAI21_X1 U22867 ( .B1(n19866), .B2(n15824), .A(n19852), .ZN(P2_U2871) );
  INV_X1 U22868 ( .A(n19853), .ZN(n19857) );
  INV_X1 U22869 ( .A(n19854), .ZN(n19856) );
  AOI21_X1 U22870 ( .B1(n19857), .B2(n19856), .A(n19855), .ZN(n19860) );
  AOI22_X1 U22871 ( .A1(n19860), .A2(n19859), .B1(n19866), .B2(n19858), .ZN(
        n19861) );
  OAI21_X1 U22872 ( .B1(n19866), .B2(n10531), .A(n19861), .ZN(P2_U2877) );
  AOI22_X1 U22873 ( .A1(n19864), .A2(n19863), .B1(n19866), .B2(n19862), .ZN(
        n19865) );
  OAI21_X1 U22874 ( .B1(n19866), .B2(n11121), .A(n19865), .ZN(P2_U2883) );
  AOI22_X1 U22875 ( .A1(n19868), .A2(n19867), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19898), .ZN(n19875) );
  AOI22_X1 U22876 ( .A1(n19870), .A2(BUF2_REG_16__SCAN_IN), .B1(n19869), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U22877 ( .A1(n19903), .A2(n19872), .B1(n19871), .B2(n19899), .ZN(
        n19873) );
  NAND3_X1 U22878 ( .A1(n19875), .A2(n19874), .A3(n19873), .ZN(P2_U2903) );
  AOI22_X1 U22879 ( .A1(n19876), .A2(n19899), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19898), .ZN(n19881) );
  XNOR2_X1 U22880 ( .A(n19878), .B(n19877), .ZN(n19879) );
  NAND2_X1 U22881 ( .A1(n19879), .A2(n19903), .ZN(n19880) );
  OAI211_X1 U22882 ( .C1(n19882), .C2(n19907), .A(n19881), .B(n19880), .ZN(
        P2_U2915) );
  AOI22_X1 U22883 ( .A1(n20607), .A2(n19899), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19898), .ZN(n19888) );
  OAI21_X1 U22884 ( .B1(n19885), .B2(n19884), .A(n19883), .ZN(n19886) );
  NAND2_X1 U22885 ( .A1(n19886), .A2(n19903), .ZN(n19887) );
  OAI211_X1 U22886 ( .C1(n19889), .C2(n19907), .A(n19888), .B(n19887), .ZN(
        P2_U2916) );
  AOI22_X1 U22887 ( .A1(n19899), .A2(n19890), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19898), .ZN(n19896) );
  OAI21_X1 U22888 ( .B1(n19893), .B2(n19892), .A(n19891), .ZN(n19894) );
  NAND2_X1 U22889 ( .A1(n19894), .A2(n19903), .ZN(n19895) );
  OAI211_X1 U22890 ( .C1(n19897), .C2(n19907), .A(n19896), .B(n19895), .ZN(
        P2_U2917) );
  AOI22_X1 U22891 ( .A1(n19899), .A2(n19959), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19898), .ZN(n19906) );
  OAI21_X1 U22892 ( .B1(n19902), .B2(n19901), .A(n19900), .ZN(n19904) );
  NAND2_X1 U22893 ( .A1(n19904), .A2(n19903), .ZN(n19905) );
  OAI211_X1 U22894 ( .C1(n19908), .C2(n19907), .A(n19906), .B(n19905), .ZN(
        P2_U2918) );
  NOR2_X1 U22895 ( .A1(n19930), .A2(n19909), .ZN(P2_U2920) );
  INV_X1 U22896 ( .A(n19910), .ZN(n19911) );
  AOI22_X1 U22897 ( .A1(n19911), .A2(P2_EAX_REG_22__SCAN_IN), .B1(
        P2_UWORD_REG_6__SCAN_IN), .B2(n19927), .ZN(n19912) );
  OAI21_X1 U22898 ( .B1(n21524), .B2(n19930), .A(n19912), .ZN(P2_U2929) );
  AOI22_X1 U22899 ( .A1(P2_EAX_REG_15__SCAN_IN), .A2(n19928), .B1(n19927), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n19913) );
  OAI21_X1 U22900 ( .B1(n21494), .B2(n19930), .A(n19913), .ZN(P2_U2936) );
  AOI22_X1 U22901 ( .A1(n19927), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19914) );
  OAI21_X1 U22902 ( .B1(n19915), .B2(n19938), .A(n19914), .ZN(P2_U2937) );
  AOI22_X1 U22903 ( .A1(n19927), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19916) );
  OAI21_X1 U22904 ( .B1(n14022), .B2(n19938), .A(n19916), .ZN(P2_U2938) );
  AOI22_X1 U22905 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19928), .B1(n19927), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19917) );
  OAI21_X1 U22906 ( .B1(n21465), .B2(n19930), .A(n19917), .ZN(P2_U2939) );
  AOI22_X1 U22907 ( .A1(P2_EAX_REG_11__SCAN_IN), .A2(n19928), .B1(n19927), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n19918) );
  OAI21_X1 U22908 ( .B1(n21483), .B2(n19930), .A(n19918), .ZN(P2_U2940) );
  AOI22_X1 U22909 ( .A1(n19927), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19919) );
  OAI21_X1 U22910 ( .B1(n19920), .B2(n19938), .A(n19919), .ZN(P2_U2941) );
  AOI22_X1 U22911 ( .A1(n19927), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19921) );
  OAI21_X1 U22912 ( .B1(n14076), .B2(n19938), .A(n19921), .ZN(P2_U2942) );
  AOI22_X1 U22913 ( .A1(n19927), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19922) );
  OAI21_X1 U22914 ( .B1(n14070), .B2(n19938), .A(n19922), .ZN(P2_U2943) );
  AOI22_X1 U22915 ( .A1(n19927), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19923) );
  OAI21_X1 U22916 ( .B1(n19924), .B2(n19938), .A(n19923), .ZN(P2_U2944) );
  AOI22_X1 U22917 ( .A1(n19927), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19925) );
  OAI21_X1 U22918 ( .B1(n19926), .B2(n19938), .A(n19925), .ZN(P2_U2945) );
  AOI22_X1 U22919 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19928), .B1(n19927), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n19929) );
  OAI21_X1 U22920 ( .B1(n21477), .B2(n19930), .A(n19929), .ZN(P2_U2946) );
  AOI22_X1 U22921 ( .A1(n19927), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19931) );
  OAI21_X1 U22922 ( .B1(n14008), .B2(n19938), .A(n19931), .ZN(P2_U2947) );
  AOI22_X1 U22923 ( .A1(n19927), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19932) );
  OAI21_X1 U22924 ( .B1(n14012), .B2(n19938), .A(n19932), .ZN(P2_U2948) );
  AOI22_X1 U22925 ( .A1(n19927), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19933) );
  OAI21_X1 U22926 ( .B1(n19934), .B2(n19938), .A(n19933), .ZN(P2_U2949) );
  AOI22_X1 U22927 ( .A1(n19927), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19935) );
  OAI21_X1 U22928 ( .B1(n19936), .B2(n19938), .A(n19935), .ZN(P2_U2950) );
  AOI22_X1 U22929 ( .A1(n19927), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n14475), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19937) );
  OAI21_X1 U22930 ( .B1(n14018), .B2(n19938), .A(n19937), .ZN(P2_U2951) );
  NOR2_X1 U22931 ( .A1(n19940), .A2(n19939), .ZN(n19957) );
  INV_X1 U22932 ( .A(n19957), .ZN(n19955) );
  INV_X1 U22933 ( .A(n19941), .ZN(n19961) );
  NOR2_X1 U22934 ( .A1(n19974), .A2(n19942), .ZN(n19952) );
  AOI22_X1 U22935 ( .A1(n19946), .A2(n19945), .B1(n19944), .B2(n19943), .ZN(
        n19948) );
  OAI211_X1 U22936 ( .C1(n19950), .C2(n19949), .A(n19948), .B(n19947), .ZN(
        n19951) );
  AOI211_X1 U22937 ( .C1(n19961), .C2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n19952), .B(n19951), .ZN(n19953) );
  OAI221_X1 U22938 ( .B1(n19957), .B2(n19956), .C1(n19955), .C2(n19954), .A(
        n19953), .ZN(P2_U3044) );
  OAI21_X1 U22939 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19958), .ZN(n19969) );
  AOI22_X1 U22940 ( .A1(n19961), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19960), .B2(n19959), .ZN(n19968) );
  OAI22_X1 U22941 ( .A1(n19965), .A2(n19964), .B1(n19963), .B2(n19962), .ZN(
        n19966) );
  INV_X1 U22942 ( .A(n19966), .ZN(n19967) );
  OAI211_X1 U22943 ( .C1(n19970), .C2(n19969), .A(n19968), .B(n19967), .ZN(
        n19971) );
  INV_X1 U22944 ( .A(n19971), .ZN(n19973) );
  OAI211_X1 U22945 ( .C1(n19975), .C2(n19974), .A(n19973), .B(n19972), .ZN(
        P2_U3045) );
  OAI21_X1 U22946 ( .B1(n20515), .B2(n20020), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19976) );
  NAND2_X1 U22947 ( .A1(n19976), .A2(n20266), .ZN(n19986) );
  OAI21_X1 U22948 ( .B1(n19978), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20614), 
        .ZN(n19979) );
  OAI21_X1 U22949 ( .B1(n19986), .B2(n20511), .A(n19979), .ZN(n19980) );
  NAND2_X1 U22950 ( .A1(n20080), .A2(n20335), .ZN(n20034) );
  NAND2_X1 U22951 ( .A1(n19980), .A2(n19982), .ZN(n19981) );
  INV_X1 U22952 ( .A(n19982), .ZN(n20024) );
  AOI22_X1 U22953 ( .A1(n20515), .A2(n20379), .B1(n20461), .B2(n20024), .ZN(
        n19988) );
  NOR2_X1 U22954 ( .A1(n20024), .A2(n20511), .ZN(n19985) );
  OAI21_X1 U22955 ( .B1(n19983), .B2(n20024), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19984) );
  AOI22_X1 U22956 ( .A1(n20462), .A2(n20027), .B1(n20020), .B2(n20470), .ZN(
        n19987) );
  OAI211_X1 U22957 ( .C1(n20025), .C2(n13149), .A(n19988), .B(n19987), .ZN(
        P2_U3048) );
  INV_X1 U22958 ( .A(n20479), .ZN(n20382) );
  AOI22_X1 U22959 ( .A1(n20515), .A2(n20382), .B1(n20024), .B2(n20474), .ZN(
        n19991) );
  AOI22_X1 U22960 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16791), .ZN(n20421) );
  AOI22_X1 U22961 ( .A1(n20475), .A2(n20027), .B1(n20020), .B2(n20476), .ZN(
        n19990) );
  OAI211_X1 U22962 ( .C1(n20025), .C2(n13164), .A(n19991), .B(n19990), .ZN(
        P2_U3049) );
  INV_X1 U22963 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19996) );
  INV_X1 U22964 ( .A(n20485), .ZN(n20385) );
  AOI22_X1 U22965 ( .A1(n20515), .A2(n20385), .B1(n20024), .B2(n20480), .ZN(
        n19995) );
  AOI22_X1 U22966 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16791), .ZN(n20426) );
  AOI22_X1 U22967 ( .A1(n20481), .A2(n20027), .B1(n20020), .B2(n20482), .ZN(
        n19994) );
  OAI211_X1 U22968 ( .C1(n20025), .C2(n19996), .A(n19995), .B(n19994), .ZN(
        P2_U3050) );
  AOI22_X2 U22969 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n16791), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20021), .ZN(n20491) );
  INV_X1 U22970 ( .A(n20491), .ZN(n20388) );
  AOI22_X1 U22971 ( .A1(n20515), .A2(n20388), .B1(n20024), .B2(n20486), .ZN(
        n20000) );
  AOI22_X1 U22972 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16791), .ZN(n20434) );
  AOI22_X1 U22973 ( .A1(n20487), .A2(n20027), .B1(n20020), .B2(n20488), .ZN(
        n19999) );
  OAI211_X1 U22974 ( .C1(n20025), .C2(n20001), .A(n20000), .B(n19999), .ZN(
        P2_U3051) );
  AOI22_X1 U22975 ( .A1(n20515), .A2(n20391), .B1(n20024), .B2(n20492), .ZN(
        n20005) );
  AOI22_X1 U22976 ( .A1(n20493), .A2(n20027), .B1(n20020), .B2(n20494), .ZN(
        n20004) );
  OAI211_X1 U22977 ( .C1(n20025), .C2(n13244), .A(n20005), .B(n20004), .ZN(
        P2_U3052) );
  INV_X1 U22978 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n21495) );
  INV_X1 U22979 ( .A(n20021), .ZN(n20011) );
  AOI22_X1 U22980 ( .A1(n20440), .A2(n20515), .B1(n20024), .B2(n20498), .ZN(
        n20009) );
  AOI22_X1 U22981 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16791), .ZN(n20443) );
  AOI22_X1 U22982 ( .A1(n20499), .A2(n20027), .B1(n20020), .B2(n20500), .ZN(
        n20008) );
  OAI211_X1 U22983 ( .C1(n20025), .C2(n20010), .A(n20009), .B(n20008), .ZN(
        P2_U3053) );
  AOI22_X1 U22984 ( .A1(n20446), .A2(n20515), .B1(n20024), .B2(n20504), .ZN(
        n20018) );
  AOI22_X1 U22985 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16791), .ZN(n20449) );
  AOI22_X1 U22986 ( .A1(n20505), .A2(n20027), .B1(n20020), .B2(n20506), .ZN(
        n20017) );
  OAI211_X1 U22987 ( .C1(n20025), .C2(n20019), .A(n20018), .B(n20017), .ZN(
        P2_U3054) );
  AOI22_X2 U22988 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20021), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n16791), .ZN(n20520) );
  INV_X1 U22989 ( .A(n20520), .ZN(n20399) );
  AOI22_X1 U22990 ( .A1(n20515), .A2(n20399), .B1(n20024), .B2(n20510), .ZN(
        n20030) );
  INV_X1 U22991 ( .A(n20025), .ZN(n20028) );
  AOI22_X1 U22992 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20028), .B1(
        n20512), .B2(n20027), .ZN(n20029) );
  OAI211_X1 U22993 ( .C1(n20458), .C2(n20058), .A(n20030), .B(n20029), .ZN(
        P2_U3055) );
  OR2_X1 U22994 ( .A1(n20034), .A2(n20627), .ZN(n20035) );
  NAND2_X1 U22995 ( .A1(n20035), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20031) );
  OAI21_X1 U22996 ( .B1(n20034), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20619), 
        .ZN(n20033) );
  AND2_X1 U22997 ( .A1(n20037), .A2(n20033), .ZN(n20054) );
  AOI22_X1 U22998 ( .A1(n20054), .A2(n20462), .B1(n20461), .B2(n20053), .ZN(
        n20040) );
  NOR2_X1 U22999 ( .A1(n20610), .A2(n20408), .ZN(n20199) );
  INV_X1 U23000 ( .A(n20199), .ZN(n20144) );
  OAI21_X1 U23001 ( .B1(n20144), .B2(n20267), .A(n20034), .ZN(n20038) );
  NAND2_X1 U23002 ( .A1(n20035), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20036) );
  NAND4_X1 U23003 ( .A1(n20038), .A2(n20467), .A3(n20037), .A4(n20036), .ZN(
        n20055) );
  AOI22_X1 U23004 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20055), .B1(
        n20073), .B2(n20470), .ZN(n20039) );
  OAI211_X1 U23005 ( .C1(n20473), .C2(n20058), .A(n20040), .B(n20039), .ZN(
        P2_U3056) );
  AOI22_X1 U23006 ( .A1(n20054), .A2(n20475), .B1(n20474), .B2(n20053), .ZN(
        n20042) );
  AOI22_X1 U23007 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20055), .B1(
        n20073), .B2(n20476), .ZN(n20041) );
  OAI211_X1 U23008 ( .C1(n20479), .C2(n20058), .A(n20042), .B(n20041), .ZN(
        P2_U3057) );
  AOI22_X1 U23009 ( .A1(n20054), .A2(n20481), .B1(n20480), .B2(n20053), .ZN(
        n20044) );
  AOI22_X1 U23010 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20055), .B1(
        n20073), .B2(n20482), .ZN(n20043) );
  OAI211_X1 U23011 ( .C1(n20485), .C2(n20058), .A(n20044), .B(n20043), .ZN(
        P2_U3058) );
  AOI22_X1 U23012 ( .A1(n20054), .A2(n20487), .B1(n20486), .B2(n20053), .ZN(
        n20046) );
  AOI22_X1 U23013 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20055), .B1(
        n20073), .B2(n20488), .ZN(n20045) );
  OAI211_X1 U23014 ( .C1(n20491), .C2(n20058), .A(n20046), .B(n20045), .ZN(
        P2_U3059) );
  AOI22_X1 U23015 ( .A1(n20054), .A2(n20493), .B1(n20492), .B2(n20053), .ZN(
        n20048) );
  AOI22_X1 U23016 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20055), .B1(
        n20073), .B2(n20494), .ZN(n20047) );
  OAI211_X1 U23017 ( .C1(n20497), .C2(n20058), .A(n20048), .B(n20047), .ZN(
        P2_U3060) );
  AOI22_X1 U23018 ( .A1(n20054), .A2(n20499), .B1(n20498), .B2(n20053), .ZN(
        n20050) );
  AOI22_X1 U23019 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20055), .B1(
        n20073), .B2(n20500), .ZN(n20049) );
  OAI211_X1 U23020 ( .C1(n20503), .C2(n20058), .A(n20050), .B(n20049), .ZN(
        P2_U3061) );
  AOI22_X1 U23021 ( .A1(n20054), .A2(n20505), .B1(n20504), .B2(n20053), .ZN(
        n20052) );
  AOI22_X1 U23022 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20055), .B1(
        n20073), .B2(n20506), .ZN(n20051) );
  OAI211_X1 U23023 ( .C1(n20509), .C2(n20058), .A(n20052), .B(n20051), .ZN(
        P2_U3062) );
  AOI22_X1 U23024 ( .A1(n20054), .A2(n20512), .B1(n20510), .B2(n20053), .ZN(
        n20057) );
  AOI22_X1 U23025 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20055), .B1(
        n20073), .B2(n20514), .ZN(n20056) );
  OAI211_X1 U23026 ( .C1(n20520), .C2(n20058), .A(n20057), .B(n20056), .ZN(
        P2_U3063) );
  AOI22_X1 U23027 ( .A1(n20072), .A2(n20475), .B1(n20071), .B2(n20474), .ZN(
        n20060) );
  AOI22_X1 U23028 ( .A1(n20097), .A2(n20476), .B1(n20073), .B2(n20382), .ZN(
        n20059) );
  OAI211_X1 U23029 ( .C1(n20077), .C2(n13162), .A(n20060), .B(n20059), .ZN(
        P2_U3065) );
  AOI22_X1 U23030 ( .A1(n20072), .A2(n20481), .B1(n20071), .B2(n20480), .ZN(
        n20062) );
  AOI22_X1 U23031 ( .A1(n20097), .A2(n20482), .B1(n20073), .B2(n20385), .ZN(
        n20061) );
  OAI211_X1 U23032 ( .C1(n20077), .C2(n13201), .A(n20062), .B(n20061), .ZN(
        P2_U3066) );
  AOI22_X1 U23033 ( .A1(n20072), .A2(n20487), .B1(n20071), .B2(n20486), .ZN(
        n20064) );
  AOI22_X1 U23034 ( .A1(n20097), .A2(n20488), .B1(n20073), .B2(n20388), .ZN(
        n20063) );
  OAI211_X1 U23035 ( .C1(n20077), .C2(n13212), .A(n20064), .B(n20063), .ZN(
        P2_U3067) );
  AOI22_X1 U23036 ( .A1(n20072), .A2(n20493), .B1(n20071), .B2(n20492), .ZN(
        n20066) );
  AOI22_X1 U23037 ( .A1(n20073), .A2(n20391), .B1(n20097), .B2(n20494), .ZN(
        n20065) );
  OAI211_X1 U23038 ( .C1(n20077), .C2(n13241), .A(n20066), .B(n20065), .ZN(
        P2_U3068) );
  AOI22_X1 U23039 ( .A1(n20072), .A2(n20499), .B1(n20071), .B2(n20498), .ZN(
        n20068) );
  AOI22_X1 U23040 ( .A1(n20097), .A2(n20500), .B1(n20073), .B2(n20440), .ZN(
        n20067) );
  OAI211_X1 U23041 ( .C1(n20077), .C2(n13270), .A(n20068), .B(n20067), .ZN(
        P2_U3069) );
  AOI22_X1 U23042 ( .A1(n20072), .A2(n20505), .B1(n20071), .B2(n20504), .ZN(
        n20070) );
  AOI22_X1 U23043 ( .A1(n20097), .A2(n20506), .B1(n20073), .B2(n20446), .ZN(
        n20069) );
  OAI211_X1 U23044 ( .C1(n20077), .C2(n13297), .A(n20070), .B(n20069), .ZN(
        P2_U3070) );
  AOI22_X1 U23045 ( .A1(n20072), .A2(n20512), .B1(n20071), .B2(n20510), .ZN(
        n20075) );
  AOI22_X1 U23046 ( .A1(n20073), .A2(n20399), .B1(n20097), .B2(n20514), .ZN(
        n20074) );
  OAI211_X1 U23047 ( .C1(n20077), .C2(n20076), .A(n20075), .B(n20074), .ZN(
        P2_U3071) );
  AOI22_X1 U23048 ( .A1(n20470), .A2(n20131), .B1(n20461), .B2(n20104), .ZN(
        n20090) );
  OAI21_X1 U23049 ( .B1(n20144), .B2(n20079), .A(n20266), .ZN(n20088) );
  AND2_X1 U23050 ( .A1(n20080), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20084) );
  INV_X1 U23051 ( .A(n20085), .ZN(n20082) );
  INV_X1 U23052 ( .A(n20104), .ZN(n20081) );
  OAI211_X1 U23053 ( .C1(n20082), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20614), 
        .B(n20081), .ZN(n20083) );
  OAI211_X1 U23054 ( .C1(n20088), .C2(n20084), .A(n20467), .B(n20083), .ZN(
        n20106) );
  INV_X1 U23055 ( .A(n20084), .ZN(n20087) );
  OAI21_X1 U23056 ( .B1(n20085), .B2(n20104), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20086) );
  AOI22_X1 U23057 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20106), .B1(
        n20462), .B2(n20105), .ZN(n20089) );
  OAI211_X1 U23058 ( .C1(n20473), .C2(n20109), .A(n20090), .B(n20089), .ZN(
        P2_U3072) );
  AOI22_X1 U23059 ( .A1(n20097), .A2(n20382), .B1(n20104), .B2(n20474), .ZN(
        n20092) );
  AOI22_X1 U23060 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20106), .B1(
        n20475), .B2(n20105), .ZN(n20091) );
  OAI211_X1 U23061 ( .C1(n20421), .C2(n20143), .A(n20092), .B(n20091), .ZN(
        P2_U3073) );
  AOI22_X1 U23062 ( .A1(n20097), .A2(n20385), .B1(n20104), .B2(n20480), .ZN(
        n20094) );
  AOI22_X1 U23063 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20106), .B1(
        n20481), .B2(n20105), .ZN(n20093) );
  OAI211_X1 U23064 ( .C1(n20426), .C2(n20143), .A(n20094), .B(n20093), .ZN(
        P2_U3074) );
  AOI22_X1 U23065 ( .A1(n20097), .A2(n20388), .B1(n20104), .B2(n20486), .ZN(
        n20096) );
  AOI22_X1 U23066 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20106), .B1(
        n20487), .B2(n20105), .ZN(n20095) );
  OAI211_X1 U23067 ( .C1(n20434), .C2(n20143), .A(n20096), .B(n20095), .ZN(
        P2_U3075) );
  AOI22_X1 U23068 ( .A1(n20097), .A2(n20391), .B1(n20104), .B2(n20492), .ZN(
        n20099) );
  AOI22_X1 U23069 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20106), .B1(
        n20493), .B2(n20105), .ZN(n20098) );
  OAI211_X1 U23070 ( .C1(n20439), .C2(n20143), .A(n20099), .B(n20098), .ZN(
        P2_U3076) );
  AOI22_X1 U23071 ( .A1(n20131), .A2(n20500), .B1(n20104), .B2(n20498), .ZN(
        n20101) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20106), .B1(
        n20499), .B2(n20105), .ZN(n20100) );
  OAI211_X1 U23073 ( .C1(n20503), .C2(n20109), .A(n20101), .B(n20100), .ZN(
        P2_U3077) );
  AOI22_X1 U23074 ( .A1(n20131), .A2(n20506), .B1(n20104), .B2(n20504), .ZN(
        n20103) );
  AOI22_X1 U23075 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20106), .B1(
        n20505), .B2(n20105), .ZN(n20102) );
  OAI211_X1 U23076 ( .C1(n20509), .C2(n20109), .A(n20103), .B(n20102), .ZN(
        P2_U3078) );
  AOI22_X1 U23077 ( .A1(n20131), .A2(n20514), .B1(n20104), .B2(n20510), .ZN(
        n20108) );
  AOI22_X1 U23078 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20106), .B1(
        n20512), .B2(n20105), .ZN(n20107) );
  OAI211_X1 U23079 ( .C1(n20520), .C2(n20109), .A(n20108), .B(n20107), .ZN(
        P2_U3079) );
  INV_X1 U23080 ( .A(n20110), .ZN(n20112) );
  NAND2_X1 U23081 ( .A1(n20112), .A2(n20111), .ZN(n20342) );
  INV_X1 U23082 ( .A(n20342), .ZN(n20117) );
  NAND3_X1 U23083 ( .A1(n20117), .A2(n20618), .A3(n16814), .ZN(n20115) );
  NOR2_X1 U23084 ( .A1(n20113), .A2(n20145), .ZN(n20138) );
  NOR3_X1 U23085 ( .A1(n20114), .A2(n20138), .A3(n20619), .ZN(n20118) );
  AOI21_X1 U23086 ( .B1(n20619), .B2(n20115), .A(n20118), .ZN(n20139) );
  AOI22_X1 U23087 ( .A1(n20139), .A2(n20462), .B1(n20461), .B2(n20138), .ZN(
        n20124) );
  OAI21_X1 U23088 ( .B1(n20131), .B2(n20166), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20121) );
  NAND2_X1 U23089 ( .A1(n20117), .A2(n20618), .ZN(n20120) );
  AOI211_X1 U23090 ( .C1(n20121), .C2(n20120), .A(n20119), .B(n20118), .ZN(
        n20122) );
  AOI22_X1 U23091 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20140), .B1(
        n20166), .B2(n20470), .ZN(n20123) );
  OAI211_X1 U23092 ( .C1(n20473), .C2(n20143), .A(n20124), .B(n20123), .ZN(
        P2_U3080) );
  AOI22_X1 U23093 ( .A1(n20139), .A2(n20475), .B1(n20474), .B2(n20138), .ZN(
        n20126) );
  AOI22_X1 U23094 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20140), .B1(
        n20166), .B2(n20476), .ZN(n20125) );
  OAI211_X1 U23095 ( .C1(n20479), .C2(n20143), .A(n20126), .B(n20125), .ZN(
        P2_U3081) );
  AOI22_X1 U23096 ( .A1(n20139), .A2(n20481), .B1(n20480), .B2(n20138), .ZN(
        n20128) );
  AOI22_X1 U23097 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20140), .B1(
        n20166), .B2(n20482), .ZN(n20127) );
  OAI211_X1 U23098 ( .C1(n20485), .C2(n20143), .A(n20128), .B(n20127), .ZN(
        P2_U3082) );
  AOI22_X1 U23099 ( .A1(n20139), .A2(n20487), .B1(n20486), .B2(n20138), .ZN(
        n20130) );
  AOI22_X1 U23100 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20140), .B1(
        n20166), .B2(n20488), .ZN(n20129) );
  OAI211_X1 U23101 ( .C1(n20491), .C2(n20143), .A(n20130), .B(n20129), .ZN(
        P2_U3083) );
  AOI22_X1 U23102 ( .A1(n20139), .A2(n20493), .B1(n20492), .B2(n20138), .ZN(
        n20133) );
  AOI22_X1 U23103 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20140), .B1(
        n20131), .B2(n20391), .ZN(n20132) );
  OAI211_X1 U23104 ( .C1(n20439), .C2(n20174), .A(n20133), .B(n20132), .ZN(
        P2_U3084) );
  AOI22_X1 U23105 ( .A1(n20139), .A2(n20499), .B1(n20498), .B2(n20138), .ZN(
        n20135) );
  AOI22_X1 U23106 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20140), .B1(
        n20166), .B2(n20500), .ZN(n20134) );
  OAI211_X1 U23107 ( .C1(n20503), .C2(n20143), .A(n20135), .B(n20134), .ZN(
        P2_U3085) );
  AOI22_X1 U23108 ( .A1(n20139), .A2(n20505), .B1(n20504), .B2(n20138), .ZN(
        n20137) );
  AOI22_X1 U23109 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20140), .B1(
        n20166), .B2(n20506), .ZN(n20136) );
  OAI211_X1 U23110 ( .C1(n20509), .C2(n20143), .A(n20137), .B(n20136), .ZN(
        P2_U3086) );
  AOI22_X1 U23111 ( .A1(n20139), .A2(n20512), .B1(n20510), .B2(n20138), .ZN(
        n20142) );
  AOI22_X1 U23112 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20140), .B1(
        n20166), .B2(n20514), .ZN(n20141) );
  OAI211_X1 U23113 ( .C1(n20520), .C2(n20143), .A(n20142), .B(n20141), .ZN(
        P2_U3087) );
  NOR3_X2 U23114 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20627), .A3(
        n20145), .ZN(n20169) );
  AOI22_X1 U23115 ( .A1(n20470), .A2(n20177), .B1(n20461), .B2(n20169), .ZN(
        n20155) );
  OAI21_X1 U23116 ( .B1(n20144), .B2(n20375), .A(n20266), .ZN(n20153) );
  NOR2_X1 U23117 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20145), .ZN(
        n20149) );
  INV_X1 U23118 ( .A(n20150), .ZN(n20147) );
  INV_X1 U23119 ( .A(n20169), .ZN(n20146) );
  OAI211_X1 U23120 ( .C1(n20147), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20614), 
        .B(n20146), .ZN(n20148) );
  OAI211_X1 U23121 ( .C1(n20153), .C2(n20149), .A(n20467), .B(n20148), .ZN(
        n20171) );
  INV_X1 U23122 ( .A(n20149), .ZN(n20152) );
  OAI21_X1 U23123 ( .B1(n20150), .B2(n20169), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20151) );
  AOI22_X1 U23124 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20171), .B1(
        n20462), .B2(n20170), .ZN(n20154) );
  OAI211_X1 U23125 ( .C1(n20473), .C2(n20174), .A(n20155), .B(n20154), .ZN(
        P2_U3088) );
  AOI22_X1 U23126 ( .A1(n20166), .A2(n20382), .B1(n20474), .B2(n20169), .ZN(
        n20157) );
  AOI22_X1 U23127 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20171), .B1(
        n20475), .B2(n20170), .ZN(n20156) );
  OAI211_X1 U23128 ( .C1(n20421), .C2(n20194), .A(n20157), .B(n20156), .ZN(
        P2_U3089) );
  AOI22_X1 U23129 ( .A1(n20177), .A2(n20482), .B1(n20169), .B2(n20480), .ZN(
        n20159) );
  AOI22_X1 U23130 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20171), .B1(
        n20481), .B2(n20170), .ZN(n20158) );
  OAI211_X1 U23131 ( .C1(n20485), .C2(n20174), .A(n20159), .B(n20158), .ZN(
        P2_U3090) );
  AOI22_X1 U23132 ( .A1(n20177), .A2(n20488), .B1(n20169), .B2(n20486), .ZN(
        n20161) );
  AOI22_X1 U23133 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20171), .B1(
        n20487), .B2(n20170), .ZN(n20160) );
  OAI211_X1 U23134 ( .C1(n20491), .C2(n20174), .A(n20161), .B(n20160), .ZN(
        P2_U3091) );
  AOI22_X1 U23135 ( .A1(n20177), .A2(n20494), .B1(n20169), .B2(n20492), .ZN(
        n20163) );
  AOI22_X1 U23136 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20171), .B1(
        n20493), .B2(n20170), .ZN(n20162) );
  OAI211_X1 U23137 ( .C1(n20497), .C2(n20174), .A(n20163), .B(n20162), .ZN(
        P2_U3092) );
  AOI22_X1 U23138 ( .A1(n20440), .A2(n20166), .B1(n20498), .B2(n20169), .ZN(
        n20165) );
  AOI22_X1 U23139 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20171), .B1(
        n20499), .B2(n20170), .ZN(n20164) );
  OAI211_X1 U23140 ( .C1(n20443), .C2(n20194), .A(n20165), .B(n20164), .ZN(
        P2_U3093) );
  AOI22_X1 U23141 ( .A1(n20446), .A2(n20166), .B1(n20504), .B2(n20169), .ZN(
        n20168) );
  AOI22_X1 U23142 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20171), .B1(
        n20505), .B2(n20170), .ZN(n20167) );
  OAI211_X1 U23143 ( .C1(n20449), .C2(n20194), .A(n20168), .B(n20167), .ZN(
        P2_U3094) );
  AOI22_X1 U23144 ( .A1(n20177), .A2(n20514), .B1(n20510), .B2(n20169), .ZN(
        n20173) );
  AOI22_X1 U23145 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20171), .B1(
        n20512), .B2(n20170), .ZN(n20172) );
  OAI211_X1 U23146 ( .C1(n20520), .C2(n20174), .A(n20173), .B(n20172), .ZN(
        P2_U3095) );
  INV_X1 U23147 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n21481) );
  AOI22_X1 U23148 ( .A1(n20190), .A2(n20475), .B1(n20189), .B2(n20474), .ZN(
        n20176) );
  AOI22_X1 U23149 ( .A1(n20218), .A2(n20476), .B1(n20177), .B2(n20382), .ZN(
        n20175) );
  OAI211_X1 U23150 ( .C1(n20180), .C2(n21481), .A(n20176), .B(n20175), .ZN(
        P2_U3097) );
  AOI22_X1 U23151 ( .A1(n20190), .A2(n20481), .B1(n20189), .B2(n20480), .ZN(
        n20179) );
  AOI22_X1 U23152 ( .A1(n20218), .A2(n20482), .B1(n20177), .B2(n20385), .ZN(
        n20178) );
  OAI211_X1 U23153 ( .C1(n20180), .C2(n10624), .A(n20179), .B(n20178), .ZN(
        P2_U3098) );
  AOI22_X1 U23154 ( .A1(n20190), .A2(n20487), .B1(n20189), .B2(n20486), .ZN(
        n20182) );
  AOI22_X1 U23155 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20191), .B1(
        n20218), .B2(n20488), .ZN(n20181) );
  OAI211_X1 U23156 ( .C1(n20491), .C2(n20194), .A(n20182), .B(n20181), .ZN(
        P2_U3099) );
  AOI22_X1 U23157 ( .A1(n20190), .A2(n20493), .B1(n20189), .B2(n20492), .ZN(
        n20184) );
  AOI22_X1 U23158 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20191), .B1(
        n20218), .B2(n20494), .ZN(n20183) );
  OAI211_X1 U23159 ( .C1(n20497), .C2(n20194), .A(n20184), .B(n20183), .ZN(
        P2_U3100) );
  AOI22_X1 U23160 ( .A1(n20190), .A2(n20499), .B1(n20189), .B2(n20498), .ZN(
        n20186) );
  AOI22_X1 U23161 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20191), .B1(
        n20218), .B2(n20500), .ZN(n20185) );
  OAI211_X1 U23162 ( .C1(n20503), .C2(n20194), .A(n20186), .B(n20185), .ZN(
        P2_U3101) );
  AOI22_X1 U23163 ( .A1(n20190), .A2(n20505), .B1(n20189), .B2(n20504), .ZN(
        n20188) );
  AOI22_X1 U23164 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20191), .B1(
        n20218), .B2(n20506), .ZN(n20187) );
  OAI211_X1 U23165 ( .C1(n20509), .C2(n20194), .A(n20188), .B(n20187), .ZN(
        P2_U3102) );
  AOI22_X1 U23166 ( .A1(n20190), .A2(n20512), .B1(n20189), .B2(n20510), .ZN(
        n20193) );
  AOI22_X1 U23167 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20191), .B1(
        n20218), .B2(n20514), .ZN(n20192) );
  OAI211_X1 U23168 ( .C1(n20520), .C2(n20194), .A(n20193), .B(n20192), .ZN(
        P2_U3103) );
  INV_X1 U23169 ( .A(n20228), .ZN(n20231) );
  OAI21_X1 U23170 ( .B1(n20197), .B2(n20231), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20196) );
  OAI21_X1 U23171 ( .B1(n20200), .B2(n20614), .A(n20196), .ZN(n20217) );
  AOI22_X1 U23172 ( .A1(n20217), .A2(n20462), .B1(n20231), .B2(n20461), .ZN(
        n20204) );
  INV_X1 U23173 ( .A(n20197), .ZN(n20198) );
  AOI21_X1 U23174 ( .B1(n20198), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20202) );
  NAND2_X1 U23175 ( .A1(n20199), .A2(n20404), .ZN(n20615) );
  NAND2_X1 U23176 ( .A1(n20615), .A2(n20200), .ZN(n20201) );
  OAI211_X1 U23177 ( .C1(n20231), .C2(n20202), .A(n20201), .B(n20467), .ZN(
        n20219) );
  AOI22_X1 U23178 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20379), .ZN(n20203) );
  OAI211_X1 U23179 ( .C1(n20419), .C2(n20258), .A(n20204), .B(n20203), .ZN(
        P2_U3104) );
  AOI22_X1 U23180 ( .A1(n20217), .A2(n20475), .B1(n20231), .B2(n20474), .ZN(
        n20206) );
  AOI22_X1 U23181 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20382), .ZN(n20205) );
  OAI211_X1 U23182 ( .C1(n20421), .C2(n20258), .A(n20206), .B(n20205), .ZN(
        P2_U3105) );
  AOI22_X1 U23183 ( .A1(n20217), .A2(n20481), .B1(n20231), .B2(n20480), .ZN(
        n20208) );
  AOI22_X1 U23184 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20385), .ZN(n20207) );
  OAI211_X1 U23185 ( .C1(n20426), .C2(n20258), .A(n20208), .B(n20207), .ZN(
        P2_U3106) );
  AOI22_X1 U23186 ( .A1(n20217), .A2(n20487), .B1(n20231), .B2(n20486), .ZN(
        n20210) );
  AOI22_X1 U23187 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20388), .ZN(n20209) );
  OAI211_X1 U23188 ( .C1(n20434), .C2(n20258), .A(n20210), .B(n20209), .ZN(
        P2_U3107) );
  AOI22_X1 U23189 ( .A1(n20217), .A2(n20493), .B1(n20231), .B2(n20492), .ZN(
        n20212) );
  AOI22_X1 U23190 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20391), .ZN(n20211) );
  OAI211_X1 U23191 ( .C1(n20439), .C2(n20258), .A(n20212), .B(n20211), .ZN(
        P2_U3108) );
  AOI22_X1 U23192 ( .A1(n20217), .A2(n20499), .B1(n20231), .B2(n20498), .ZN(
        n20214) );
  AOI22_X1 U23193 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20440), .ZN(n20213) );
  OAI211_X1 U23194 ( .C1(n20443), .C2(n20258), .A(n20214), .B(n20213), .ZN(
        P2_U3109) );
  AOI22_X1 U23195 ( .A1(n20217), .A2(n20505), .B1(n20231), .B2(n20504), .ZN(
        n20216) );
  AOI22_X1 U23196 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20446), .ZN(n20215) );
  OAI211_X1 U23197 ( .C1(n20449), .C2(n20258), .A(n20216), .B(n20215), .ZN(
        P2_U3110) );
  AOI22_X1 U23198 ( .A1(n20217), .A2(n20512), .B1(n20231), .B2(n20510), .ZN(
        n20221) );
  AOI22_X1 U23199 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20399), .ZN(n20220) );
  OAI211_X1 U23200 ( .C1(n20458), .C2(n20258), .A(n20221), .B(n20220), .ZN(
        P2_U3111) );
  INV_X1 U23201 ( .A(n20267), .ZN(n20222) );
  OR2_X1 U23202 ( .A1(n20419), .A2(n20295), .ZN(n20224) );
  NAND2_X1 U23203 ( .A1(n20461), .A2(n20236), .ZN(n20223) );
  AND2_X1 U23204 ( .A1(n20224), .A2(n20223), .ZN(n20235) );
  AOI21_X1 U23205 ( .B1(n20258), .B2(n20295), .A(n20408), .ZN(n20225) );
  NOR2_X1 U23206 ( .A1(n20225), .A2(n20614), .ZN(n20230) );
  OAI21_X1 U23207 ( .B1(n20226), .B2(n20619), .A(n16814), .ZN(n20227) );
  AOI21_X1 U23208 ( .B1(n20230), .B2(n20228), .A(n20227), .ZN(n20229) );
  OAI21_X2 U23209 ( .B1(n20229), .B2(n20236), .A(n20467), .ZN(n20261) );
  OAI21_X1 U23210 ( .B1(n20231), .B2(n20236), .A(n20230), .ZN(n20233) );
  OAI21_X1 U23211 ( .B1(n20226), .B2(n20236), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20232) );
  AOI22_X1 U23212 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20261), .B1(
        n20462), .B2(n20260), .ZN(n20234) );
  OAI211_X1 U23213 ( .C1(n20473), .C2(n20258), .A(n20235), .B(n20234), .ZN(
        P2_U3112) );
  INV_X1 U23214 ( .A(n20236), .ZN(n20257) );
  INV_X1 U23215 ( .A(n20474), .ZN(n20420) );
  OAI22_X1 U23216 ( .A1(n20295), .A2(n20421), .B1(n20257), .B2(n20420), .ZN(
        n20237) );
  INV_X1 U23217 ( .A(n20237), .ZN(n20239) );
  AOI22_X1 U23218 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20261), .B1(
        n20475), .B2(n20260), .ZN(n20238) );
  OAI211_X1 U23219 ( .C1(n20479), .C2(n20258), .A(n20239), .B(n20238), .ZN(
        P2_U3113) );
  INV_X1 U23220 ( .A(n20480), .ZN(n20425) );
  OAI22_X1 U23221 ( .A1(n20295), .A2(n20426), .B1(n20257), .B2(n20425), .ZN(
        n20240) );
  INV_X1 U23222 ( .A(n20240), .ZN(n20242) );
  AOI22_X1 U23223 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20261), .B1(
        n20481), .B2(n20260), .ZN(n20241) );
  OAI211_X1 U23224 ( .C1(n20485), .C2(n20258), .A(n20242), .B(n20241), .ZN(
        P2_U3114) );
  INV_X1 U23225 ( .A(n20486), .ZN(n20430) );
  OAI22_X1 U23226 ( .A1(n20295), .A2(n20434), .B1(n20257), .B2(n20430), .ZN(
        n20243) );
  INV_X1 U23227 ( .A(n20243), .ZN(n20245) );
  AOI22_X1 U23228 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20261), .B1(
        n20487), .B2(n20260), .ZN(n20244) );
  OAI211_X1 U23229 ( .C1(n20491), .C2(n20258), .A(n20245), .B(n20244), .ZN(
        P2_U3115) );
  INV_X1 U23230 ( .A(n20492), .ZN(n20435) );
  OAI22_X1 U23231 ( .A1(n20258), .A2(n20497), .B1(n20257), .B2(n20435), .ZN(
        n20246) );
  INV_X1 U23232 ( .A(n20246), .ZN(n20248) );
  AOI22_X1 U23233 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20261), .B1(
        n20493), .B2(n20260), .ZN(n20247) );
  OAI211_X1 U23234 ( .C1(n20439), .C2(n20295), .A(n20248), .B(n20247), .ZN(
        P2_U3116) );
  INV_X1 U23235 ( .A(n20498), .ZN(n20249) );
  OAI22_X1 U23236 ( .A1(n20295), .A2(n20443), .B1(n20257), .B2(n20249), .ZN(
        n20250) );
  INV_X1 U23237 ( .A(n20250), .ZN(n20252) );
  AOI22_X1 U23238 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20261), .B1(
        n20499), .B2(n20260), .ZN(n20251) );
  OAI211_X1 U23239 ( .C1(n20503), .C2(n20258), .A(n20252), .B(n20251), .ZN(
        P2_U3117) );
  INV_X1 U23240 ( .A(n20504), .ZN(n20253) );
  OAI22_X1 U23241 ( .A1(n20295), .A2(n20449), .B1(n20257), .B2(n20253), .ZN(
        n20254) );
  INV_X1 U23242 ( .A(n20254), .ZN(n20256) );
  AOI22_X1 U23243 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20261), .B1(
        n20505), .B2(n20260), .ZN(n20255) );
  OAI211_X1 U23244 ( .C1(n20509), .C2(n20258), .A(n20256), .B(n20255), .ZN(
        P2_U3118) );
  INV_X1 U23245 ( .A(n20510), .ZN(n20451) );
  OAI22_X1 U23246 ( .A1(n20258), .A2(n20520), .B1(n20257), .B2(n20451), .ZN(
        n20259) );
  INV_X1 U23247 ( .A(n20259), .ZN(n20263) );
  AOI22_X1 U23248 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20261), .B1(
        n20512), .B2(n20260), .ZN(n20262) );
  OAI211_X1 U23249 ( .C1(n20458), .C2(n20295), .A(n20263), .B(n20262), .ZN(
        P2_U3119) );
  OR2_X1 U23250 ( .A1(n20419), .A2(n20308), .ZN(n20265) );
  NAND2_X1 U23251 ( .A1(n20461), .A2(n20290), .ZN(n20264) );
  AND2_X1 U23252 ( .A1(n20265), .A2(n20264), .ZN(n20275) );
  OAI21_X1 U23253 ( .B1(n20466), .B2(n20267), .A(n20266), .ZN(n20273) );
  INV_X1 U23254 ( .A(n20290), .ZN(n20282) );
  OAI211_X1 U23255 ( .C1(n20268), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20614), 
        .B(n20282), .ZN(n20269) );
  OAI211_X1 U23256 ( .C1(n20273), .C2(n20270), .A(n20467), .B(n20269), .ZN(
        n20292) );
  INV_X1 U23257 ( .A(n20270), .ZN(n20272) );
  AOI22_X1 U23258 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20292), .B1(
        n20462), .B2(n20291), .ZN(n20274) );
  OAI211_X1 U23259 ( .C1(n20473), .C2(n20295), .A(n20275), .B(n20274), .ZN(
        P2_U3120) );
  AOI22_X1 U23260 ( .A1(n20311), .A2(n20476), .B1(n20290), .B2(n20474), .ZN(
        n20277) );
  AOI22_X1 U23261 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20292), .B1(
        n20475), .B2(n20291), .ZN(n20276) );
  OAI211_X1 U23262 ( .C1(n20479), .C2(n20295), .A(n20277), .B(n20276), .ZN(
        P2_U3121) );
  AOI22_X1 U23263 ( .A1(n20311), .A2(n20482), .B1(n20290), .B2(n20480), .ZN(
        n20279) );
  AOI22_X1 U23264 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20292), .B1(
        n20481), .B2(n20291), .ZN(n20278) );
  OAI211_X1 U23265 ( .C1(n20485), .C2(n20295), .A(n20279), .B(n20278), .ZN(
        P2_U3122) );
  AOI22_X1 U23266 ( .A1(n20311), .A2(n20488), .B1(n20290), .B2(n20486), .ZN(
        n20281) );
  AOI22_X1 U23267 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20292), .B1(
        n20487), .B2(n20291), .ZN(n20280) );
  OAI211_X1 U23268 ( .C1(n20491), .C2(n20295), .A(n20281), .B(n20280), .ZN(
        P2_U3123) );
  OAI22_X1 U23269 ( .A1(n20295), .A2(n20497), .B1(n20282), .B2(n20435), .ZN(
        n20283) );
  INV_X1 U23270 ( .A(n20283), .ZN(n20285) );
  AOI22_X1 U23271 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20292), .B1(
        n20493), .B2(n20291), .ZN(n20284) );
  OAI211_X1 U23272 ( .C1(n20439), .C2(n20308), .A(n20285), .B(n20284), .ZN(
        P2_U3124) );
  AOI22_X1 U23273 ( .A1(n20311), .A2(n20500), .B1(n20290), .B2(n20498), .ZN(
        n20287) );
  AOI22_X1 U23274 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20292), .B1(
        n20499), .B2(n20291), .ZN(n20286) );
  OAI211_X1 U23275 ( .C1(n20503), .C2(n20295), .A(n20287), .B(n20286), .ZN(
        P2_U3125) );
  AOI22_X1 U23276 ( .A1(n20311), .A2(n20506), .B1(n20290), .B2(n20504), .ZN(
        n20289) );
  AOI22_X1 U23277 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20292), .B1(
        n20505), .B2(n20291), .ZN(n20288) );
  OAI211_X1 U23278 ( .C1(n20509), .C2(n20295), .A(n20289), .B(n20288), .ZN(
        P2_U3126) );
  AOI22_X1 U23279 ( .A1(n20311), .A2(n20514), .B1(n20290), .B2(n20510), .ZN(
        n20294) );
  AOI22_X1 U23280 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20292), .B1(
        n20512), .B2(n20291), .ZN(n20293) );
  OAI211_X1 U23281 ( .C1(n20520), .C2(n20295), .A(n20294), .B(n20293), .ZN(
        P2_U3127) );
  AOI22_X1 U23282 ( .A1(n20310), .A2(n20475), .B1(n20309), .B2(n20474), .ZN(
        n20297) );
  AOI22_X1 U23283 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20312), .B1(
        n20325), .B2(n20476), .ZN(n20296) );
  OAI211_X1 U23284 ( .C1(n20479), .C2(n20308), .A(n20297), .B(n20296), .ZN(
        P2_U3129) );
  AOI22_X1 U23285 ( .A1(n20310), .A2(n20481), .B1(n20309), .B2(n20480), .ZN(
        n20299) );
  AOI22_X1 U23286 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20312), .B1(
        n20325), .B2(n20482), .ZN(n20298) );
  OAI211_X1 U23287 ( .C1(n20485), .C2(n20308), .A(n20299), .B(n20298), .ZN(
        P2_U3130) );
  AOI22_X1 U23288 ( .A1(n20310), .A2(n20487), .B1(n20309), .B2(n20486), .ZN(
        n20301) );
  AOI22_X1 U23289 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20312), .B1(
        n20325), .B2(n20488), .ZN(n20300) );
  OAI211_X1 U23290 ( .C1(n20491), .C2(n20308), .A(n20301), .B(n20300), .ZN(
        P2_U3131) );
  AOI22_X1 U23291 ( .A1(n20310), .A2(n20493), .B1(n20309), .B2(n20492), .ZN(
        n20303) );
  AOI22_X1 U23292 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20312), .B1(
        n20311), .B2(n20391), .ZN(n20302) );
  OAI211_X1 U23293 ( .C1(n20439), .C2(n20333), .A(n20303), .B(n20302), .ZN(
        P2_U3132) );
  AOI22_X1 U23294 ( .A1(n20310), .A2(n20499), .B1(n20309), .B2(n20498), .ZN(
        n20305) );
  AOI22_X1 U23295 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20312), .B1(
        n20325), .B2(n20500), .ZN(n20304) );
  OAI211_X1 U23296 ( .C1(n20503), .C2(n20308), .A(n20305), .B(n20304), .ZN(
        P2_U3133) );
  AOI22_X1 U23297 ( .A1(n20310), .A2(n20505), .B1(n20309), .B2(n20504), .ZN(
        n20307) );
  AOI22_X1 U23298 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20312), .B1(
        n20325), .B2(n20506), .ZN(n20306) );
  OAI211_X1 U23299 ( .C1(n20509), .C2(n20308), .A(n20307), .B(n20306), .ZN(
        P2_U3134) );
  AOI22_X1 U23300 ( .A1(n20310), .A2(n20512), .B1(n20309), .B2(n20510), .ZN(
        n20314) );
  AOI22_X1 U23301 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20312), .B1(
        n20311), .B2(n20399), .ZN(n20313) );
  OAI211_X1 U23302 ( .C1(n20458), .C2(n20333), .A(n20314), .B(n20313), .ZN(
        P2_U3135) );
  AOI22_X1 U23303 ( .A1(n20329), .A2(n20475), .B1(n20328), .B2(n20474), .ZN(
        n20316) );
  AOI22_X1 U23304 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20330), .B1(
        n20340), .B2(n20476), .ZN(n20315) );
  OAI211_X1 U23305 ( .C1(n20479), .C2(n20333), .A(n20316), .B(n20315), .ZN(
        P2_U3137) );
  AOI22_X1 U23306 ( .A1(n20329), .A2(n20481), .B1(n20328), .B2(n20480), .ZN(
        n20318) );
  AOI22_X1 U23307 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20330), .B1(
        n20325), .B2(n20385), .ZN(n20317) );
  OAI211_X1 U23308 ( .C1(n20426), .C2(n20366), .A(n20318), .B(n20317), .ZN(
        P2_U3138) );
  AOI22_X1 U23309 ( .A1(n20329), .A2(n20487), .B1(n20328), .B2(n20486), .ZN(
        n20320) );
  AOI22_X1 U23310 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20330), .B1(
        n20340), .B2(n20488), .ZN(n20319) );
  OAI211_X1 U23311 ( .C1(n20491), .C2(n20333), .A(n20320), .B(n20319), .ZN(
        P2_U3139) );
  AOI22_X1 U23312 ( .A1(n20329), .A2(n20493), .B1(n20328), .B2(n20492), .ZN(
        n20322) );
  AOI22_X1 U23313 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20330), .B1(
        n20340), .B2(n20494), .ZN(n20321) );
  OAI211_X1 U23314 ( .C1(n20497), .C2(n20333), .A(n20322), .B(n20321), .ZN(
        P2_U3140) );
  AOI22_X1 U23315 ( .A1(n20329), .A2(n20499), .B1(n20328), .B2(n20498), .ZN(
        n20324) );
  AOI22_X1 U23316 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20330), .B1(
        n20340), .B2(n20500), .ZN(n20323) );
  OAI211_X1 U23317 ( .C1(n20503), .C2(n20333), .A(n20324), .B(n20323), .ZN(
        P2_U3141) );
  AOI22_X1 U23318 ( .A1(n20329), .A2(n20505), .B1(n20328), .B2(n20504), .ZN(
        n20327) );
  AOI22_X1 U23319 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20330), .B1(
        n20325), .B2(n20446), .ZN(n20326) );
  OAI211_X1 U23320 ( .C1(n20449), .C2(n20366), .A(n20327), .B(n20326), .ZN(
        P2_U3142) );
  AOI22_X1 U23321 ( .A1(n20329), .A2(n20512), .B1(n20328), .B2(n20510), .ZN(
        n20332) );
  AOI22_X1 U23322 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20330), .B1(
        n20340), .B2(n20514), .ZN(n20331) );
  OAI211_X1 U23323 ( .C1(n20520), .C2(n20333), .A(n20332), .B(n20331), .ZN(
        P2_U3143) );
  INV_X1 U23324 ( .A(n20334), .ZN(n20338) );
  NAND2_X1 U23325 ( .A1(n20372), .A2(n20627), .ZN(n20343) );
  OAI21_X1 U23326 ( .B1(n20336), .B2(n20361), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20337) );
  AOI22_X1 U23327 ( .A1(n20362), .A2(n20462), .B1(n20461), .B2(n20361), .ZN(
        n20348) );
  OAI21_X1 U23328 ( .B1(n20400), .B2(n20340), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20341) );
  OAI21_X1 U23329 ( .B1(n20618), .B2(n20342), .A(n20341), .ZN(n20346) );
  OAI211_X1 U23330 ( .C1(n20344), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20614), 
        .B(n20343), .ZN(n20345) );
  NAND3_X1 U23331 ( .A1(n20346), .A2(n20467), .A3(n20345), .ZN(n20363) );
  AOI22_X1 U23332 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20363), .B1(
        n20400), .B2(n20470), .ZN(n20347) );
  OAI211_X1 U23333 ( .C1(n20473), .C2(n20366), .A(n20348), .B(n20347), .ZN(
        P2_U3144) );
  AOI22_X1 U23334 ( .A1(n20362), .A2(n20475), .B1(n20361), .B2(n20474), .ZN(
        n20350) );
  AOI22_X1 U23335 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20363), .B1(
        n20400), .B2(n20476), .ZN(n20349) );
  OAI211_X1 U23336 ( .C1(n20479), .C2(n20366), .A(n20350), .B(n20349), .ZN(
        P2_U3145) );
  AOI22_X1 U23337 ( .A1(n20362), .A2(n20481), .B1(n20361), .B2(n20480), .ZN(
        n20352) );
  AOI22_X1 U23338 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20363), .B1(
        n20400), .B2(n20482), .ZN(n20351) );
  OAI211_X1 U23339 ( .C1(n20485), .C2(n20366), .A(n20352), .B(n20351), .ZN(
        P2_U3146) );
  AOI22_X1 U23340 ( .A1(n20362), .A2(n20487), .B1(n20361), .B2(n20486), .ZN(
        n20354) );
  AOI22_X1 U23341 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20363), .B1(
        n20400), .B2(n20488), .ZN(n20353) );
  OAI211_X1 U23342 ( .C1(n20491), .C2(n20366), .A(n20354), .B(n20353), .ZN(
        P2_U3147) );
  AOI22_X1 U23343 ( .A1(n20362), .A2(n20493), .B1(n20361), .B2(n20492), .ZN(
        n20356) );
  AOI22_X1 U23344 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20363), .B1(
        n20400), .B2(n20494), .ZN(n20355) );
  OAI211_X1 U23345 ( .C1(n20497), .C2(n20366), .A(n20356), .B(n20355), .ZN(
        P2_U3148) );
  AOI22_X1 U23346 ( .A1(n20362), .A2(n20499), .B1(n20361), .B2(n20498), .ZN(
        n20358) );
  AOI22_X1 U23347 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20363), .B1(
        n20400), .B2(n20500), .ZN(n20357) );
  OAI211_X1 U23348 ( .C1(n20503), .C2(n20366), .A(n20358), .B(n20357), .ZN(
        P2_U3149) );
  AOI22_X1 U23349 ( .A1(n20362), .A2(n20505), .B1(n20361), .B2(n20504), .ZN(
        n20360) );
  AOI22_X1 U23350 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20363), .B1(
        n20400), .B2(n20506), .ZN(n20359) );
  OAI211_X1 U23351 ( .C1(n20509), .C2(n20366), .A(n20360), .B(n20359), .ZN(
        P2_U3150) );
  AOI22_X1 U23352 ( .A1(n20362), .A2(n20512), .B1(n20361), .B2(n20510), .ZN(
        n20365) );
  AOI22_X1 U23353 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20363), .B1(
        n20400), .B2(n20514), .ZN(n20364) );
  OAI211_X1 U23354 ( .C1(n20520), .C2(n20366), .A(n20365), .B(n20364), .ZN(
        P2_U3151) );
  INV_X1 U23355 ( .A(n20367), .ZN(n20369) );
  INV_X1 U23356 ( .A(n20375), .ZN(n20368) );
  NAND2_X1 U23357 ( .A1(n20372), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20411) );
  AND2_X1 U23358 ( .A1(n20411), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20370) );
  NAND2_X1 U23359 ( .A1(n20371), .A2(n20370), .ZN(n20377) );
  INV_X1 U23360 ( .A(n20372), .ZN(n20374) );
  OAI21_X1 U23361 ( .B1(n20374), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20619), 
        .ZN(n20373) );
  AND2_X1 U23362 ( .A1(n20377), .A2(n20373), .ZN(n20398) );
  INV_X1 U23363 ( .A(n20411), .ZN(n20414) );
  AOI22_X1 U23364 ( .A1(n20398), .A2(n20462), .B1(n20461), .B2(n20414), .ZN(
        n20381) );
  OAI21_X1 U23365 ( .B1(n20466), .B2(n20375), .A(n20374), .ZN(n20378) );
  NAND2_X1 U23366 ( .A1(n20411), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20376) );
  NAND4_X1 U23367 ( .A1(n20378), .A2(n20467), .A3(n20377), .A4(n20376), .ZN(
        n20401) );
  AOI22_X1 U23368 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20379), .ZN(n20380) );
  OAI211_X1 U23369 ( .C1(n20419), .C2(n20452), .A(n20381), .B(n20380), .ZN(
        P2_U3152) );
  AOI22_X1 U23370 ( .A1(n20398), .A2(n20475), .B1(n20414), .B2(n20474), .ZN(
        n20384) );
  AOI22_X1 U23371 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20382), .ZN(n20383) );
  OAI211_X1 U23372 ( .C1(n20421), .C2(n20452), .A(n20384), .B(n20383), .ZN(
        P2_U3153) );
  AOI22_X1 U23373 ( .A1(n20398), .A2(n20481), .B1(n20414), .B2(n20480), .ZN(
        n20387) );
  AOI22_X1 U23374 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20385), .ZN(n20386) );
  OAI211_X1 U23375 ( .C1(n20426), .C2(n20452), .A(n20387), .B(n20386), .ZN(
        P2_U3154) );
  AOI22_X1 U23376 ( .A1(n20398), .A2(n20487), .B1(n20414), .B2(n20486), .ZN(
        n20390) );
  AOI22_X1 U23377 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20388), .ZN(n20389) );
  OAI211_X1 U23378 ( .C1(n20434), .C2(n20452), .A(n20390), .B(n20389), .ZN(
        P2_U3155) );
  AOI22_X1 U23379 ( .A1(n20398), .A2(n20493), .B1(n20414), .B2(n20492), .ZN(
        n20393) );
  AOI22_X1 U23380 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20391), .ZN(n20392) );
  OAI211_X1 U23381 ( .C1(n20439), .C2(n20452), .A(n20393), .B(n20392), .ZN(
        P2_U3156) );
  AOI22_X1 U23382 ( .A1(n20398), .A2(n20499), .B1(n20414), .B2(n20498), .ZN(
        n20395) );
  AOI22_X1 U23383 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20440), .ZN(n20394) );
  OAI211_X1 U23384 ( .C1(n20443), .C2(n20452), .A(n20395), .B(n20394), .ZN(
        P2_U3157) );
  AOI22_X1 U23385 ( .A1(n20398), .A2(n20505), .B1(n20414), .B2(n20504), .ZN(
        n20397) );
  AOI22_X1 U23386 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20446), .ZN(n20396) );
  OAI211_X1 U23387 ( .C1(n20449), .C2(n20452), .A(n20397), .B(n20396), .ZN(
        P2_U3158) );
  AOI22_X1 U23388 ( .A1(n20398), .A2(n20512), .B1(n20414), .B2(n20510), .ZN(
        n20403) );
  AOI22_X1 U23389 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20399), .ZN(n20402) );
  OAI211_X1 U23390 ( .C1(n20458), .C2(n20452), .A(n20403), .B(n20402), .ZN(
        P2_U3159) );
  NAND3_X1 U23391 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20464) );
  NOR2_X1 U23392 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20464), .ZN(
        n20444) );
  INV_X1 U23393 ( .A(n20444), .ZN(n20450) );
  OAI22_X1 U23394 ( .A1(n20452), .A2(n20473), .B1(n20406), .B2(n20450), .ZN(
        n20407) );
  INV_X1 U23395 ( .A(n20407), .ZN(n20418) );
  AOI21_X1 U23396 ( .B1(n20452), .B2(n20519), .A(n20408), .ZN(n20409) );
  NOR2_X1 U23397 ( .A1(n20409), .A2(n20614), .ZN(n20413) );
  OAI21_X1 U23398 ( .B1(n10890), .B2(n20619), .A(n16814), .ZN(n20410) );
  AOI21_X1 U23399 ( .B1(n20413), .B2(n20411), .A(n20410), .ZN(n20412) );
  OAI21_X2 U23400 ( .B1(n20412), .B2(n20444), .A(n20467), .ZN(n20455) );
  OAI21_X1 U23401 ( .B1(n20444), .B2(n20414), .A(n20413), .ZN(n20416) );
  OAI21_X1 U23402 ( .B1(n10890), .B2(n20444), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20415) );
  AOI22_X1 U23403 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20455), .B1(
        n20462), .B2(n20454), .ZN(n20417) );
  OAI211_X1 U23404 ( .C1(n20419), .C2(n20519), .A(n20418), .B(n20417), .ZN(
        P2_U3160) );
  OAI22_X1 U23405 ( .A1(n20519), .A2(n20421), .B1(n20420), .B2(n20450), .ZN(
        n20422) );
  INV_X1 U23406 ( .A(n20422), .ZN(n20424) );
  AOI22_X1 U23407 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20455), .B1(
        n20475), .B2(n20454), .ZN(n20423) );
  OAI211_X1 U23408 ( .C1(n20479), .C2(n20452), .A(n20424), .B(n20423), .ZN(
        P2_U3161) );
  OAI22_X1 U23409 ( .A1(n20519), .A2(n20426), .B1(n20425), .B2(n20450), .ZN(
        n20427) );
  INV_X1 U23410 ( .A(n20427), .ZN(n20429) );
  AOI22_X1 U23411 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20455), .B1(
        n20481), .B2(n20454), .ZN(n20428) );
  OAI211_X1 U23412 ( .C1(n20485), .C2(n20452), .A(n20429), .B(n20428), .ZN(
        P2_U3162) );
  OAI22_X1 U23413 ( .A1(n20452), .A2(n20491), .B1(n20430), .B2(n20450), .ZN(
        n20431) );
  INV_X1 U23414 ( .A(n20431), .ZN(n20433) );
  AOI22_X1 U23415 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20455), .B1(
        n20487), .B2(n20454), .ZN(n20432) );
  OAI211_X1 U23416 ( .C1(n20434), .C2(n20519), .A(n20433), .B(n20432), .ZN(
        P2_U3163) );
  OAI22_X1 U23417 ( .A1(n20452), .A2(n20497), .B1(n20435), .B2(n20450), .ZN(
        n20436) );
  INV_X1 U23418 ( .A(n20436), .ZN(n20438) );
  AOI22_X1 U23419 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20455), .B1(
        n20493), .B2(n20454), .ZN(n20437) );
  OAI211_X1 U23420 ( .C1(n20439), .C2(n20519), .A(n20438), .B(n20437), .ZN(
        P2_U3164) );
  INV_X1 U23421 ( .A(n20452), .ZN(n20445) );
  AOI22_X1 U23422 ( .A1(n20440), .A2(n20445), .B1(n20498), .B2(n20444), .ZN(
        n20442) );
  AOI22_X1 U23423 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20455), .B1(
        n20499), .B2(n20454), .ZN(n20441) );
  OAI211_X1 U23424 ( .C1(n20443), .C2(n20519), .A(n20442), .B(n20441), .ZN(
        P2_U3165) );
  AOI22_X1 U23425 ( .A1(n20446), .A2(n20445), .B1(n20504), .B2(n20444), .ZN(
        n20448) );
  AOI22_X1 U23426 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20455), .B1(
        n20505), .B2(n20454), .ZN(n20447) );
  OAI211_X1 U23427 ( .C1(n20449), .C2(n20519), .A(n20448), .B(n20447), .ZN(
        P2_U3166) );
  OAI22_X1 U23428 ( .A1(n20452), .A2(n20520), .B1(n20451), .B2(n20450), .ZN(
        n20453) );
  INV_X1 U23429 ( .A(n20453), .ZN(n20457) );
  AOI22_X1 U23430 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20455), .B1(
        n20512), .B2(n20454), .ZN(n20456) );
  OAI211_X1 U23431 ( .C1(n20458), .C2(n20519), .A(n20457), .B(n20456), .ZN(
        P2_U3167) );
  OAI21_X1 U23432 ( .B1(n20459), .B2(n20511), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20460) );
  OAI21_X1 U23433 ( .B1(n20464), .B2(n20614), .A(n20460), .ZN(n20513) );
  AOI22_X1 U23434 ( .A1(n20513), .A2(n20462), .B1(n20461), .B2(n20511), .ZN(
        n20472) );
  AOI21_X1 U23435 ( .B1(n20463), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20469) );
  OAI21_X1 U23436 ( .B1(n20466), .B2(n20465), .A(n20464), .ZN(n20468) );
  OAI211_X1 U23437 ( .C1(n20511), .C2(n20469), .A(n20468), .B(n20467), .ZN(
        n20516) );
  AOI22_X1 U23438 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20470), .ZN(n20471) );
  OAI211_X1 U23439 ( .C1(n20473), .C2(n20519), .A(n20472), .B(n20471), .ZN(
        P2_U3168) );
  AOI22_X1 U23440 ( .A1(n20513), .A2(n20475), .B1(n20511), .B2(n20474), .ZN(
        n20478) );
  AOI22_X1 U23441 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20476), .ZN(n20477) );
  OAI211_X1 U23442 ( .C1(n20479), .C2(n20519), .A(n20478), .B(n20477), .ZN(
        P2_U3169) );
  AOI22_X1 U23443 ( .A1(n20513), .A2(n20481), .B1(n20511), .B2(n20480), .ZN(
        n20484) );
  AOI22_X1 U23444 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20482), .ZN(n20483) );
  OAI211_X1 U23445 ( .C1(n20485), .C2(n20519), .A(n20484), .B(n20483), .ZN(
        P2_U3170) );
  AOI22_X1 U23446 ( .A1(n20513), .A2(n20487), .B1(n20511), .B2(n20486), .ZN(
        n20490) );
  AOI22_X1 U23447 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20488), .ZN(n20489) );
  OAI211_X1 U23448 ( .C1(n20491), .C2(n20519), .A(n20490), .B(n20489), .ZN(
        P2_U3171) );
  AOI22_X1 U23449 ( .A1(n20513), .A2(n20493), .B1(n20511), .B2(n20492), .ZN(
        n20496) );
  AOI22_X1 U23450 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20494), .ZN(n20495) );
  OAI211_X1 U23451 ( .C1(n20497), .C2(n20519), .A(n20496), .B(n20495), .ZN(
        P2_U3172) );
  AOI22_X1 U23452 ( .A1(n20513), .A2(n20499), .B1(n20511), .B2(n20498), .ZN(
        n20502) );
  AOI22_X1 U23453 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20500), .ZN(n20501) );
  OAI211_X1 U23454 ( .C1(n20503), .C2(n20519), .A(n20502), .B(n20501), .ZN(
        P2_U3173) );
  AOI22_X1 U23455 ( .A1(n20513), .A2(n20505), .B1(n20511), .B2(n20504), .ZN(
        n20508) );
  AOI22_X1 U23456 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20506), .ZN(n20507) );
  OAI211_X1 U23457 ( .C1(n20509), .C2(n20519), .A(n20508), .B(n20507), .ZN(
        P2_U3174) );
  AOI22_X1 U23458 ( .A1(n20513), .A2(n20512), .B1(n20511), .B2(n20510), .ZN(
        n20518) );
  AOI22_X1 U23459 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20514), .ZN(n20517) );
  OAI211_X1 U23460 ( .C1(n20520), .C2(n20519), .A(n20518), .B(n20517), .ZN(
        P2_U3175) );
  AND2_X1 U23461 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20521), .ZN(
        P2_U3179) );
  AND2_X1 U23462 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20521), .ZN(
        P2_U3180) );
  AND2_X1 U23463 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20521), .ZN(
        P2_U3181) );
  AND2_X1 U23464 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20521), .ZN(
        P2_U3182) );
  AND2_X1 U23465 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20521), .ZN(
        P2_U3183) );
  AND2_X1 U23466 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20521), .ZN(
        P2_U3184) );
  AND2_X1 U23467 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20521), .ZN(
        P2_U3185) );
  AND2_X1 U23468 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20521), .ZN(
        P2_U3186) );
  AND2_X1 U23469 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20521), .ZN(
        P2_U3187) );
  AND2_X1 U23470 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20521), .ZN(
        P2_U3188) );
  AND2_X1 U23471 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20521), .ZN(
        P2_U3189) );
  AND2_X1 U23472 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20521), .ZN(
        P2_U3190) );
  AND2_X1 U23473 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20521), .ZN(
        P2_U3191) );
  AND2_X1 U23474 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20521), .ZN(
        P2_U3192) );
  AND2_X1 U23475 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20521), .ZN(
        P2_U3193) );
  AND2_X1 U23476 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20521), .ZN(
        P2_U3194) );
  AND2_X1 U23477 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20521), .ZN(
        P2_U3195) );
  AND2_X1 U23478 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20521), .ZN(
        P2_U3196) );
  AND2_X1 U23479 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20521), .ZN(
        P2_U3197) );
  AND2_X1 U23480 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20521), .ZN(
        P2_U3198) );
  AND2_X1 U23481 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20521), .ZN(
        P2_U3199) );
  AND2_X1 U23482 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20521), .ZN(
        P2_U3200) );
  AND2_X1 U23483 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20521), .ZN(P2_U3201) );
  AND2_X1 U23484 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20521), .ZN(P2_U3202) );
  AND2_X1 U23485 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20521), .ZN(P2_U3203) );
  AND2_X1 U23486 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20521), .ZN(P2_U3204) );
  AND2_X1 U23487 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20521), .ZN(P2_U3205) );
  AND2_X1 U23488 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20521), .ZN(P2_U3206) );
  AND2_X1 U23489 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20521), .ZN(P2_U3207) );
  AND2_X1 U23490 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20521), .ZN(P2_U3208) );
  NAND2_X1 U23491 ( .A1(n20532), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20534) );
  NAND3_X1 U23492 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20534), .ZN(n20522) );
  NOR2_X1 U23493 ( .A1(n21362), .A2(n20527), .ZN(n20539) );
  AOI21_X1 U23494 ( .B1(n20540), .B2(n20522), .A(n20539), .ZN(n20523) );
  OAI221_X1 U23495 ( .B1(n20524), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20524), .C2(n21363), .A(n20523), .ZN(P2_U3209) );
  INV_X1 U23496 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20525) );
  AOI21_X1 U23497 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21363), .A(n20540), 
        .ZN(n20531) );
  NOR2_X1 U23498 ( .A1(n20525), .A2(n20531), .ZN(n20528) );
  AOI21_X1 U23499 ( .B1(n20528), .B2(n20527), .A(n20526), .ZN(n20529) );
  OAI211_X1 U23500 ( .C1(n21363), .C2(n20530), .A(n20529), .B(n20534), .ZN(
        P2_U3210) );
  AOI21_X1 U23501 ( .B1(n20533), .B2(n20532), .A(n20531), .ZN(n20538) );
  OAI22_X1 U23502 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20535), .B1(NA), 
        .B2(n20534), .ZN(n20536) );
  OAI211_X1 U23503 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20536), .ZN(n20537) );
  OAI21_X1 U23504 ( .B1(n20539), .B2(n20538), .A(n20537), .ZN(P2_U3211) );
  NAND2_X2 U23505 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20597), .ZN(n20596) );
  INV_X1 U23506 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n21555) );
  OAI222_X1 U23507 ( .A1(n20596), .A2(n20542), .B1(n20541), .B2(n20597), .C1(
        n21555), .C2(n20599), .ZN(P2_U3212) );
  OAI222_X1 U23508 ( .A1(n20596), .A2(n21555), .B1(n20543), .B2(n20597), .C1(
        n20545), .C2(n20599), .ZN(P2_U3213) );
  OAI222_X1 U23509 ( .A1(n20596), .A2(n20545), .B1(n20544), .B2(n20597), .C1(
        n20546), .C2(n20599), .ZN(P2_U3214) );
  INV_X1 U23510 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n20548) );
  OAI222_X1 U23511 ( .A1(n20599), .A2(n20548), .B1(n20547), .B2(n20597), .C1(
        n20546), .C2(n20596), .ZN(P2_U3215) );
  OAI222_X1 U23512 ( .A1(n20599), .A2(n20550), .B1(n20549), .B2(n20597), .C1(
        n20548), .C2(n20596), .ZN(P2_U3216) );
  OAI222_X1 U23513 ( .A1(n20599), .A2(n20552), .B1(n20551), .B2(n20597), .C1(
        n20550), .C2(n20596), .ZN(P2_U3217) );
  OAI222_X1 U23514 ( .A1(n20599), .A2(n20554), .B1(n20553), .B2(n20597), .C1(
        n20552), .C2(n20596), .ZN(P2_U3218) );
  OAI222_X1 U23515 ( .A1(n20599), .A2(n20556), .B1(n20555), .B2(n20597), .C1(
        n20554), .C2(n20596), .ZN(P2_U3219) );
  INV_X1 U23516 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20558) );
  OAI222_X1 U23517 ( .A1(n20599), .A2(n20558), .B1(n20557), .B2(n20597), .C1(
        n20556), .C2(n20596), .ZN(P2_U3220) );
  INV_X1 U23518 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20560) );
  OAI222_X1 U23519 ( .A1(n20599), .A2(n20560), .B1(n20559), .B2(n20597), .C1(
        n20558), .C2(n20596), .ZN(P2_U3221) );
  OAI222_X1 U23520 ( .A1(n20599), .A2(n20562), .B1(n20561), .B2(n20597), .C1(
        n20560), .C2(n20596), .ZN(P2_U3222) );
  INV_X1 U23521 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20564) );
  OAI222_X1 U23522 ( .A1(n20599), .A2(n20564), .B1(n20563), .B2(n20597), .C1(
        n20562), .C2(n20596), .ZN(P2_U3223) );
  INV_X1 U23523 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20566) );
  OAI222_X1 U23524 ( .A1(n20599), .A2(n20566), .B1(n20565), .B2(n20597), .C1(
        n20564), .C2(n20596), .ZN(P2_U3224) );
  OAI222_X1 U23525 ( .A1(n20599), .A2(n20568), .B1(n20567), .B2(n20597), .C1(
        n20566), .C2(n20596), .ZN(P2_U3225) );
  OAI222_X1 U23526 ( .A1(n20599), .A2(n20570), .B1(n20569), .B2(n20597), .C1(
        n20568), .C2(n20596), .ZN(P2_U3226) );
  OAI222_X1 U23527 ( .A1(n20599), .A2(n20572), .B1(n20571), .B2(n20597), .C1(
        n20570), .C2(n20596), .ZN(P2_U3227) );
  OAI222_X1 U23528 ( .A1(n20599), .A2(n20573), .B1(n21463), .B2(n20597), .C1(
        n20572), .C2(n20596), .ZN(P2_U3228) );
  OAI222_X1 U23529 ( .A1(n20599), .A2(n20575), .B1(n20574), .B2(n20597), .C1(
        n20573), .C2(n20596), .ZN(P2_U3229) );
  INV_X1 U23530 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20577) );
  OAI222_X1 U23531 ( .A1(n20599), .A2(n20577), .B1(n20576), .B2(n20597), .C1(
        n20575), .C2(n20596), .ZN(P2_U3230) );
  INV_X1 U23532 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20579) );
  OAI222_X1 U23533 ( .A1(n20599), .A2(n20579), .B1(n20578), .B2(n20597), .C1(
        n20577), .C2(n20596), .ZN(P2_U3231) );
  OAI222_X1 U23534 ( .A1(n20599), .A2(n11798), .B1(n20580), .B2(n20597), .C1(
        n20579), .C2(n20596), .ZN(P2_U3232) );
  OAI222_X1 U23535 ( .A1(n20599), .A2(n20582), .B1(n20581), .B2(n20597), .C1(
        n11798), .C2(n20596), .ZN(P2_U3233) );
  OAI222_X1 U23536 ( .A1(n20599), .A2(n20584), .B1(n20583), .B2(n20597), .C1(
        n20582), .C2(n20596), .ZN(P2_U3234) );
  OAI222_X1 U23537 ( .A1(n20599), .A2(n20586), .B1(n20585), .B2(n20597), .C1(
        n20584), .C2(n20596), .ZN(P2_U3235) );
  OAI222_X1 U23538 ( .A1(n20599), .A2(n20588), .B1(n20587), .B2(n20597), .C1(
        n20586), .C2(n20596), .ZN(P2_U3236) );
  INV_X1 U23539 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20591) );
  OAI222_X1 U23540 ( .A1(n20599), .A2(n20591), .B1(n20589), .B2(n20597), .C1(
        n20588), .C2(n20596), .ZN(P2_U3237) );
  INV_X1 U23541 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20592) );
  OAI222_X1 U23542 ( .A1(n20596), .A2(n20591), .B1(n20590), .B2(n20597), .C1(
        n20592), .C2(n20599), .ZN(P2_U3238) );
  OAI222_X1 U23543 ( .A1(n20599), .A2(n20594), .B1(n20593), .B2(n20597), .C1(
        n20592), .C2(n20596), .ZN(P2_U3239) );
  OAI222_X1 U23544 ( .A1(n20599), .A2(n13357), .B1(n20595), .B2(n20597), .C1(
        n20594), .C2(n20596), .ZN(P2_U3240) );
  OAI222_X1 U23545 ( .A1(n20599), .A2(n14726), .B1(n20598), .B2(n20597), .C1(
        n13357), .C2(n20596), .ZN(P2_U3241) );
  OAI22_X1 U23546 ( .A1(n20638), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20597), .ZN(n20600) );
  INV_X1 U23547 ( .A(n20600), .ZN(P2_U3585) );
  MUX2_X1 U23548 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20638), .Z(P2_U3586) );
  OAI22_X1 U23549 ( .A1(n20638), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20597), .ZN(n20601) );
  INV_X1 U23550 ( .A(n20601), .ZN(P2_U3587) );
  OAI22_X1 U23551 ( .A1(n20638), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20597), .ZN(n20602) );
  INV_X1 U23552 ( .A(n20602), .ZN(P2_U3588) );
  OAI21_X1 U23553 ( .B1(n20606), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20604), 
        .ZN(n20603) );
  INV_X1 U23554 ( .A(n20603), .ZN(P2_U3591) );
  OAI21_X1 U23555 ( .B1(n20606), .B2(n20605), .A(n20604), .ZN(P2_U3592) );
  NAND2_X1 U23556 ( .A1(n20607), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20613) );
  NAND2_X1 U23557 ( .A1(n20609), .A2(n20608), .ZN(n20611) );
  NAND2_X1 U23558 ( .A1(n20611), .A2(n20610), .ZN(n20612) );
  OAI211_X1 U23559 ( .C1(n20615), .C2(n20614), .A(n20613), .B(n20612), .ZN(
        n20616) );
  INV_X1 U23560 ( .A(n20616), .ZN(n20617) );
  AOI22_X1 U23561 ( .A1(n20625), .A2(n20618), .B1(n20617), .B2(n20626), .ZN(
        P2_U3602) );
  OAI22_X1 U23562 ( .A1(n20622), .A2(n20621), .B1(n20620), .B2(n20619), .ZN(
        n20623) );
  AOI21_X1 U23563 ( .B1(n20627), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20623), 
        .ZN(n20624) );
  OAI22_X1 U23564 ( .A1(n20627), .A2(n20626), .B1(n20625), .B2(n20624), .ZN(
        P2_U3605) );
  INV_X1 U23565 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20628) );
  AOI22_X1 U23566 ( .A1(n20597), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20628), 
        .B2(n20638), .ZN(P2_U3608) );
  INV_X1 U23567 ( .A(n20629), .ZN(n20631) );
  AOI22_X1 U23568 ( .A1(n20633), .A2(n20632), .B1(n20631), .B2(n20630), .ZN(
        n20634) );
  NAND2_X1 U23569 ( .A1(n20635), .A2(n20634), .ZN(n20637) );
  MUX2_X1 U23570 ( .A(P2_MORE_REG_SCAN_IN), .B(n20637), .S(n20636), .Z(
        P2_U3609) );
  OAI22_X1 U23571 ( .A1(n20638), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20597), .ZN(n20639) );
  INV_X1 U23572 ( .A(n20639), .ZN(P2_U3611) );
  OAI21_X1 U23573 ( .B1(n20641), .B2(n20640), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20642) );
  OAI21_X1 U23574 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20643), .A(n20642), 
        .ZN(P1_U2803) );
  NOR2_X1 U23575 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20645) );
  OAI21_X1 U23576 ( .B1(n20645), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21407), .ZN(
        n20644) );
  OAI21_X1 U23577 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n13907), .A(n20644), 
        .ZN(P1_U2804) );
  OAI21_X1 U23578 ( .B1(BS16), .B2(n20645), .A(n21385), .ZN(n21383) );
  OAI21_X1 U23579 ( .B1(n21385), .B2(n21397), .A(n21383), .ZN(P1_U2805) );
  OAI21_X1 U23580 ( .B1(n20648), .B2(n20647), .A(n20646), .ZN(P1_U2806) );
  NOR4_X1 U23581 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20652) );
  NOR4_X1 U23582 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20651) );
  NOR4_X1 U23583 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20650) );
  NOR4_X1 U23584 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20649) );
  NAND4_X1 U23585 ( .A1(n20652), .A2(n20651), .A3(n20650), .A4(n20649), .ZN(
        n20658) );
  NOR4_X1 U23586 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20656) );
  AOI211_X1 U23587 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_3__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20655) );
  NOR4_X1 U23588 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20654) );
  NOR4_X1 U23589 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20653) );
  NAND4_X1 U23590 ( .A1(n20656), .A2(n20655), .A3(n20654), .A4(n20653), .ZN(
        n20657) );
  NOR2_X1 U23591 ( .A1(n20658), .A2(n20657), .ZN(n21390) );
  INV_X1 U23592 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20660) );
  NOR3_X1 U23593 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20661) );
  OAI21_X1 U23594 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20661), .A(n21390), .ZN(
        n20659) );
  OAI21_X1 U23595 ( .B1(n21390), .B2(n20660), .A(n20659), .ZN(P1_U2807) );
  INV_X1 U23596 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21384) );
  AOI21_X1 U23597 ( .B1(n21386), .B2(n21384), .A(n20661), .ZN(n20663) );
  INV_X1 U23598 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20662) );
  INV_X1 U23599 ( .A(n21390), .ZN(n21393) );
  AOI22_X1 U23600 ( .A1(n21390), .A2(n20663), .B1(n20662), .B2(n21393), .ZN(
        P1_U2808) );
  OAI22_X1 U23601 ( .A1(n20718), .A2(n20665), .B1(n20702), .B2(n20664), .ZN(
        n20666) );
  AOI211_X1 U23602 ( .C1(n20735), .C2(n20667), .A(n17416), .B(n20666), .ZN(
        n20675) );
  INV_X1 U23603 ( .A(n20668), .ZN(n20670) );
  AOI22_X1 U23604 ( .A1(n20670), .A2(n9887), .B1(n20721), .B2(n20669), .ZN(
        n20674) );
  OAI21_X1 U23605 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20672), .A(n20671), .ZN(
        n20673) );
  NAND3_X1 U23606 ( .A1(n20675), .A2(n20674), .A3(n20673), .ZN(P1_U2831) );
  NAND2_X1 U23607 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20681) );
  OAI21_X1 U23608 ( .B1(n20681), .B2(n20677), .A(n20676), .ZN(n20700) );
  AOI22_X1 U23609 ( .A1(n20735), .A2(n20678), .B1(n20736), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n20679) );
  OAI21_X1 U23610 ( .B1(n20750), .B2(n20680), .A(n20679), .ZN(n20685) );
  NOR3_X1 U23611 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20681), .A3(n20704), .ZN(
        n20682) );
  AOI211_X1 U23612 ( .C1(n20738), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n17416), .B(n20682), .ZN(n20683) );
  INV_X1 U23613 ( .A(n20683), .ZN(n20684) );
  AOI211_X1 U23614 ( .C1(n9887), .C2(n20686), .A(n20685), .B(n20684), .ZN(
        n20687) );
  OAI21_X1 U23615 ( .B1(n20700), .B2(n20688), .A(n20687), .ZN(P1_U2833) );
  AOI22_X1 U23616 ( .A1(n20736), .A2(P1_EBX_REG_6__SCAN_IN), .B1(n20735), .B2(
        n20689), .ZN(n20690) );
  OAI21_X1 U23617 ( .B1(n20750), .B2(n20691), .A(n20690), .ZN(n20696) );
  NOR3_X1 U23618 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20692), .A3(n20704), .ZN(
        n20693) );
  AOI211_X1 U23619 ( .C1(n20738), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17416), .B(n20693), .ZN(n20694) );
  INV_X1 U23620 ( .A(n20694), .ZN(n20695) );
  AOI211_X1 U23621 ( .C1(n9887), .C2(n20697), .A(n20696), .B(n20695), .ZN(
        n20698) );
  OAI21_X1 U23622 ( .B1(n20700), .B2(n20699), .A(n20698), .ZN(P1_U2834) );
  OAI21_X1 U23623 ( .B1(n20718), .B2(n20701), .A(n20716), .ZN(n20706) );
  OAI22_X1 U23624 ( .A1(n20704), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20703), 
        .B2(n20702), .ZN(n20705) );
  AOI211_X1 U23625 ( .C1(n20735), .C2(n20707), .A(n20706), .B(n20705), .ZN(
        n20711) );
  INV_X1 U23626 ( .A(n20708), .ZN(n20722) );
  AOI22_X1 U23627 ( .A1(n20709), .A2(n20723), .B1(n20722), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20710) );
  OAI211_X1 U23628 ( .C1(n20712), .C2(n20750), .A(n20711), .B(n20710), .ZN(
        P1_U2835) );
  INV_X1 U23629 ( .A(n20713), .ZN(n20714) );
  AOI22_X1 U23630 ( .A1(n20715), .A2(n20747), .B1(n20735), .B2(n20714), .ZN(
        n20731) );
  NAND2_X1 U23631 ( .A1(n20736), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n20717) );
  OAI211_X1 U23632 ( .C1(n14539), .C2(n20718), .A(n20717), .B(n20716), .ZN(
        n20719) );
  AOI21_X1 U23633 ( .B1(n20721), .B2(n20720), .A(n20719), .ZN(n20730) );
  AOI22_X1 U23634 ( .A1(n20724), .A2(n20723), .B1(n20722), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20729) );
  NOR2_X1 U23635 ( .A1(n20726), .A2(n20725), .ZN(n20740) );
  NAND3_X1 U23636 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20740), .A3(n20727), 
        .ZN(n20728) );
  NAND4_X1 U23637 ( .A1(n20731), .A2(n20730), .A3(n20729), .A4(n20728), .ZN(
        P1_U2836) );
  INV_X1 U23638 ( .A(n20732), .ZN(n20751) );
  INV_X1 U23639 ( .A(n20733), .ZN(n20734) );
  AOI22_X1 U23640 ( .A1(n20736), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20735), .B2(
        n20734), .ZN(n20749) );
  INV_X1 U23641 ( .A(n20737), .ZN(n20742) );
  AOI22_X1 U23642 ( .A1(n20740), .A2(n20739), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20738), .ZN(n20741) );
  OAI21_X1 U23643 ( .B1(n20742), .B2(n20739), .A(n20741), .ZN(n20746) );
  NOR2_X1 U23644 ( .A1(n20744), .A2(n20743), .ZN(n20745) );
  AOI211_X1 U23645 ( .C1(n20747), .C2(n21063), .A(n20746), .B(n20745), .ZN(
        n20748) );
  OAI211_X1 U23646 ( .C1(n20751), .C2(n20750), .A(n20749), .B(n20748), .ZN(
        P1_U2837) );
  AOI22_X1 U23647 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20766), .B1(n20783), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20752) );
  OAI21_X1 U23648 ( .B1(n20774), .B2(n20753), .A(n20752), .ZN(P1_U2921) );
  INV_X1 U23649 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20755) );
  AOI22_X1 U23650 ( .A1(n20784), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20754) );
  OAI21_X1 U23651 ( .B1(n20755), .B2(n20786), .A(n20754), .ZN(P1_U2922) );
  INV_X1 U23652 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20757) );
  AOI22_X1 U23653 ( .A1(n20784), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20756) );
  OAI21_X1 U23654 ( .B1(n20757), .B2(n20786), .A(n20756), .ZN(P1_U2923) );
  INV_X1 U23655 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20759) );
  AOI22_X1 U23656 ( .A1(n20784), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20758) );
  OAI21_X1 U23657 ( .B1(n20759), .B2(n20786), .A(n20758), .ZN(P1_U2924) );
  INV_X1 U23658 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20761) );
  AOI22_X1 U23659 ( .A1(n20784), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20760) );
  OAI21_X1 U23660 ( .B1(n20761), .B2(n20786), .A(n20760), .ZN(P1_U2925) );
  INV_X1 U23661 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20763) );
  AOI22_X1 U23662 ( .A1(n20784), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20762) );
  OAI21_X1 U23663 ( .B1(n20763), .B2(n20786), .A(n20762), .ZN(P1_U2926) );
  INV_X1 U23664 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20765) );
  AOI22_X1 U23665 ( .A1(n20784), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20764) );
  OAI21_X1 U23666 ( .B1(n20765), .B2(n20786), .A(n20764), .ZN(P1_U2927) );
  AOI222_X1 U23667 ( .A1(n20784), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20766), 
        .B2(P1_EAX_REG_8__SCAN_IN), .C1(P1_DATAO_REG_8__SCAN_IN), .C2(n20783), 
        .ZN(n20767) );
  INV_X1 U23668 ( .A(n20767), .ZN(P1_U2928) );
  AOI22_X1 U23669 ( .A1(n20784), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20768) );
  OAI21_X1 U23670 ( .B1(n20769), .B2(n20786), .A(n20768), .ZN(P1_U2929) );
  AOI22_X1 U23671 ( .A1(n20784), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20770) );
  OAI21_X1 U23672 ( .B1(n12625), .B2(n20786), .A(n20770), .ZN(P1_U2930) );
  INV_X1 U23673 ( .A(P1_LWORD_REG_5__SCAN_IN), .ZN(n21528) );
  OAI222_X1 U23674 ( .A1(n20774), .A2(n21528), .B1(n20786), .B2(n20773), .C1(
        n20772), .C2(n20771), .ZN(P1_U2931) );
  AOI22_X1 U23675 ( .A1(n20784), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20775) );
  OAI21_X1 U23676 ( .B1(n20776), .B2(n20786), .A(n20775), .ZN(P1_U2932) );
  AOI22_X1 U23677 ( .A1(n20784), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20777) );
  OAI21_X1 U23678 ( .B1(n20778), .B2(n20786), .A(n20777), .ZN(P1_U2933) );
  AOI22_X1 U23679 ( .A1(n20784), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20779) );
  OAI21_X1 U23680 ( .B1(n20780), .B2(n20786), .A(n20779), .ZN(P1_U2934) );
  AOI22_X1 U23681 ( .A1(n20784), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20781) );
  OAI21_X1 U23682 ( .B1(n20782), .B2(n20786), .A(n20781), .ZN(P1_U2935) );
  AOI22_X1 U23683 ( .A1(n20784), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20783), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20785) );
  OAI21_X1 U23684 ( .B1(n20787), .B2(n20786), .A(n20785), .ZN(P1_U2936) );
  AOI22_X1 U23685 ( .A1(n20805), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20804), .ZN(n20790) );
  NAND2_X1 U23686 ( .A1(n20807), .A2(n20788), .ZN(n20789) );
  NAND2_X1 U23687 ( .A1(n20790), .A2(n20789), .ZN(P1_U2961) );
  AOI22_X1 U23688 ( .A1(n20805), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20804), .ZN(n20793) );
  NAND2_X1 U23689 ( .A1(n20807), .A2(n20791), .ZN(n20792) );
  NAND2_X1 U23690 ( .A1(n20793), .A2(n20792), .ZN(P1_U2962) );
  AOI22_X1 U23691 ( .A1(n20805), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20804), .ZN(n20796) );
  NAND2_X1 U23692 ( .A1(n20807), .A2(n20794), .ZN(n20795) );
  NAND2_X1 U23693 ( .A1(n20796), .A2(n20795), .ZN(P1_U2963) );
  AOI22_X1 U23694 ( .A1(n20805), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20797), .ZN(n20800) );
  NAND2_X1 U23695 ( .A1(n20807), .A2(n20798), .ZN(n20799) );
  NAND2_X1 U23696 ( .A1(n20800), .A2(n20799), .ZN(P1_U2964) );
  AOI22_X1 U23697 ( .A1(n20805), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20804), .ZN(n20803) );
  NAND2_X1 U23698 ( .A1(n20807), .A2(n20801), .ZN(n20802) );
  NAND2_X1 U23699 ( .A1(n20803), .A2(n20802), .ZN(P1_U2965) );
  AOI22_X1 U23700 ( .A1(n20805), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20804), .ZN(n20809) );
  NAND2_X1 U23701 ( .A1(n20807), .A2(n20806), .ZN(n20808) );
  NAND2_X1 U23702 ( .A1(n20809), .A2(n20808), .ZN(P1_U2966) );
  AND2_X1 U23703 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20810), .ZN(
        P1_U3032) );
  AOI22_X1 U23704 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20849), .B1(DATAI_16_), 
        .B2(n20850), .ZN(n21281) );
  INV_X1 U23705 ( .A(n21155), .ZN(n20813) );
  AOI22_X1 U23706 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20849), .B1(DATAI_24_), 
        .B2(n20850), .ZN(n21311) );
  INV_X1 U23707 ( .A(n21311), .ZN(n21278) );
  NOR2_X2 U23708 ( .A1(n20852), .A2(n11955), .ZN(n21299) );
  NAND2_X1 U23709 ( .A1(n21132), .A2(n21064), .ZN(n20922) );
  OR2_X1 U23710 ( .A1(n21191), .A2(n20922), .ZN(n20818) );
  INV_X1 U23711 ( .A(n20818), .ZN(n20853) );
  AOI22_X1 U23712 ( .A1(n21308), .A2(n21278), .B1(n21299), .B2(n20853), .ZN(
        n20827) );
  INV_X1 U23713 ( .A(n20887), .ZN(n20815) );
  OAI21_X1 U23714 ( .B1(n20815), .B2(n21308), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20816) );
  NAND2_X1 U23715 ( .A1(n20816), .A2(n21265), .ZN(n20825) );
  NOR2_X1 U23716 ( .A1(n20891), .A2(n21273), .ZN(n20822) );
  OR2_X1 U23717 ( .A1(n21066), .A2(n21067), .ZN(n20955) );
  AOI22_X1 U23718 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20955), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20818), .ZN(n20820) );
  INV_X1 U23719 ( .A(n20823), .ZN(n20819) );
  INV_X1 U23720 ( .A(n20822), .ZN(n20824) );
  OR2_X1 U23721 ( .A1(n20823), .A2(n12586), .ZN(n21069) );
  AOI22_X1 U23722 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20857), .B1(
        n21300), .B2(n20856), .ZN(n20826) );
  OAI211_X1 U23723 ( .C1(n21281), .C2(n20887), .A(n20827), .B(n20826), .ZN(
        P1_U3033) );
  AOI22_X1 U23724 ( .A1(DATAI_17_), .A2(n20850), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20849), .ZN(n21317) );
  AOI22_X1 U23725 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20849), .B1(DATAI_25_), 
        .B2(n20850), .ZN(n21102) );
  INV_X1 U23726 ( .A(n21102), .ZN(n21314) );
  NOR2_X2 U23727 ( .A1(n20852), .A2(n20828), .ZN(n21313) );
  AOI22_X1 U23728 ( .A1(n21308), .A2(n21314), .B1(n21313), .B2(n20853), .ZN(
        n20831) );
  AOI22_X1 U23729 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20857), .B1(
        n21312), .B2(n20856), .ZN(n20830) );
  OAI211_X1 U23730 ( .C1(n21317), .C2(n20887), .A(n20831), .B(n20830), .ZN(
        P1_U3034) );
  AOI22_X1 U23731 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20849), .B1(DATAI_18_), 
        .B2(n20850), .ZN(n21416) );
  AOI22_X1 U23732 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20849), .B1(DATAI_26_), 
        .B2(n20850), .ZN(n21418) );
  INV_X1 U23733 ( .A(n21418), .ZN(n21319) );
  NOR2_X2 U23734 ( .A1(n20852), .A2(n20832), .ZN(n21409) );
  AOI22_X1 U23735 ( .A1(n21308), .A2(n21319), .B1(n21409), .B2(n20853), .ZN(
        n20835) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20857), .B1(
        n21318), .B2(n20856), .ZN(n20834) );
  OAI211_X1 U23737 ( .C1(n21416), .C2(n20887), .A(n20835), .B(n20834), .ZN(
        P1_U3035) );
  AOI22_X1 U23738 ( .A1(DATAI_19_), .A2(n20850), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20849), .ZN(n21327) );
  AOI22_X1 U23739 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20849), .B1(DATAI_27_), 
        .B2(n20850), .ZN(n21107) );
  INV_X1 U23740 ( .A(n21107), .ZN(n21324) );
  AOI22_X1 U23741 ( .A1(n21308), .A2(n21324), .B1(n21322), .B2(n20853), .ZN(
        n20838) );
  AOI22_X1 U23742 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20857), .B1(
        n21323), .B2(n20856), .ZN(n20837) );
  OAI211_X1 U23743 ( .C1(n21327), .C2(n20887), .A(n20838), .B(n20837), .ZN(
        P1_U3036) );
  AOI22_X1 U23744 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20849), .B1(DATAI_20_), 
        .B2(n20850), .ZN(n21333) );
  AOI22_X1 U23745 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20849), .B1(DATAI_28_), 
        .B2(n20850), .ZN(n21110) );
  INV_X1 U23746 ( .A(n21110), .ZN(n21330) );
  NOR2_X2 U23747 ( .A1(n20852), .A2(n11957), .ZN(n21328) );
  AOI22_X1 U23748 ( .A1(n21308), .A2(n21330), .B1(n21328), .B2(n20853), .ZN(
        n20841) );
  AOI22_X1 U23749 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20857), .B1(
        n21329), .B2(n20856), .ZN(n20840) );
  OAI211_X1 U23750 ( .C1(n21333), .C2(n20887), .A(n20841), .B(n20840), .ZN(
        P1_U3037) );
  AOI22_X1 U23751 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20849), .B1(DATAI_21_), 
        .B2(n20850), .ZN(n21339) );
  AOI22_X1 U23752 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20849), .B1(DATAI_29_), 
        .B2(n20850), .ZN(n21113) );
  INV_X1 U23753 ( .A(n21113), .ZN(n21336) );
  NOR2_X2 U23754 ( .A1(n20852), .A2(n20842), .ZN(n21334) );
  AOI22_X1 U23755 ( .A1(n21308), .A2(n21336), .B1(n21334), .B2(n20853), .ZN(
        n20845) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20857), .B1(
        n21335), .B2(n20856), .ZN(n20844) );
  OAI211_X1 U23757 ( .C1(n21339), .C2(n20887), .A(n20845), .B(n20844), .ZN(
        P1_U3038) );
  AOI22_X1 U23758 ( .A1(DATAI_22_), .A2(n20850), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20849), .ZN(n21345) );
  AOI22_X1 U23759 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20849), .B1(DATAI_30_), 
        .B2(n20850), .ZN(n21116) );
  INV_X1 U23760 ( .A(n21116), .ZN(n21342) );
  NOR2_X2 U23761 ( .A1(n20852), .A2(n12591), .ZN(n21340) );
  AOI22_X1 U23762 ( .A1(n21308), .A2(n21342), .B1(n21340), .B2(n20853), .ZN(
        n20848) );
  AOI22_X1 U23763 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20857), .B1(
        n21341), .B2(n20856), .ZN(n20847) );
  OAI211_X1 U23764 ( .C1(n21345), .C2(n20887), .A(n20848), .B(n20847), .ZN(
        P1_U3039) );
  AOI22_X1 U23765 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20849), .B1(DATAI_23_), 
        .B2(n20850), .ZN(n21356) );
  AOI22_X1 U23766 ( .A1(DATAI_31_), .A2(n20850), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20849), .ZN(n21123) );
  INV_X1 U23767 ( .A(n21123), .ZN(n21350) );
  NOR2_X2 U23768 ( .A1(n20852), .A2(n20851), .ZN(n21347) );
  AOI22_X1 U23769 ( .A1(n21308), .A2(n21350), .B1(n21347), .B2(n20853), .ZN(
        n20859) );
  AOI22_X1 U23770 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20857), .B1(
        n21349), .B2(n20856), .ZN(n20858) );
  OAI211_X1 U23771 ( .C1(n21356), .C2(n20887), .A(n20859), .B(n20858), .ZN(
        P1_U3040) );
  INV_X1 U23772 ( .A(n20891), .ZN(n20923) );
  INV_X1 U23773 ( .A(n20860), .ZN(n21235) );
  NOR2_X1 U23774 ( .A1(n20922), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20865) );
  INV_X1 U23775 ( .A(n20865), .ZN(n20861) );
  NOR2_X1 U23776 ( .A1(n21234), .A2(n20861), .ZN(n20882) );
  AOI21_X1 U23777 ( .B1(n20923), .B2(n21235), .A(n20882), .ZN(n20863) );
  OAI22_X1 U23778 ( .A1(n20863), .A2(n21302), .B1(n20861), .B2(n12586), .ZN(
        n20883) );
  AOI22_X1 U23779 ( .A1(n21300), .A2(n20883), .B1(n21299), .B2(n20882), .ZN(
        n20869) );
  INV_X1 U23780 ( .A(n20862), .ZN(n21238) );
  OAI21_X1 U23781 ( .B1(n20930), .B2(n21238), .A(n20863), .ZN(n20864) );
  OAI221_X1 U23782 ( .B1(n21265), .B2(n20865), .C1(n21302), .C2(n20864), .A(
        n21306), .ZN(n20884) );
  INV_X1 U23783 ( .A(n14508), .ZN(n20867) );
  INV_X1 U23784 ( .A(n21281), .ZN(n21307) );
  AOI22_X1 U23785 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20884), .B1(
        n20912), .B2(n21307), .ZN(n20868) );
  OAI211_X1 U23786 ( .C1(n21311), .C2(n20887), .A(n20869), .B(n20868), .ZN(
        P1_U3041) );
  AOI22_X1 U23787 ( .A1(n21313), .A2(n20882), .B1(n21312), .B2(n20883), .ZN(
        n20871) );
  INV_X1 U23788 ( .A(n21317), .ZN(n21202) );
  AOI22_X1 U23789 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20884), .B1(
        n20912), .B2(n21202), .ZN(n20870) );
  OAI211_X1 U23790 ( .C1(n21102), .C2(n20887), .A(n20871), .B(n20870), .ZN(
        P1_U3042) );
  AOI22_X1 U23791 ( .A1(n21318), .A2(n20883), .B1(n21409), .B2(n20882), .ZN(
        n20873) );
  INV_X1 U23792 ( .A(n21416), .ZN(n21206) );
  AOI22_X1 U23793 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20884), .B1(
        n20912), .B2(n21206), .ZN(n20872) );
  OAI211_X1 U23794 ( .C1(n21418), .C2(n20887), .A(n20873), .B(n20872), .ZN(
        P1_U3043) );
  AOI22_X1 U23795 ( .A1(n21323), .A2(n20883), .B1(n21322), .B2(n20882), .ZN(
        n20875) );
  INV_X1 U23796 ( .A(n21327), .ZN(n21209) );
  AOI22_X1 U23797 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20884), .B1(
        n20912), .B2(n21209), .ZN(n20874) );
  OAI211_X1 U23798 ( .C1(n21107), .C2(n20887), .A(n20875), .B(n20874), .ZN(
        P1_U3044) );
  AOI22_X1 U23799 ( .A1(n21329), .A2(n20883), .B1(n21328), .B2(n20882), .ZN(
        n20877) );
  INV_X1 U23800 ( .A(n21333), .ZN(n21213) );
  AOI22_X1 U23801 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20884), .B1(
        n20912), .B2(n21213), .ZN(n20876) );
  OAI211_X1 U23802 ( .C1(n21110), .C2(n20887), .A(n20877), .B(n20876), .ZN(
        P1_U3045) );
  AOI22_X1 U23803 ( .A1(n21335), .A2(n20883), .B1(n21334), .B2(n20882), .ZN(
        n20879) );
  INV_X1 U23804 ( .A(n21339), .ZN(n21217) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20884), .B1(
        n20912), .B2(n21217), .ZN(n20878) );
  OAI211_X1 U23806 ( .C1(n21113), .C2(n20887), .A(n20879), .B(n20878), .ZN(
        P1_U3046) );
  AOI22_X1 U23807 ( .A1(n21341), .A2(n20883), .B1(n21340), .B2(n20882), .ZN(
        n20881) );
  INV_X1 U23808 ( .A(n21345), .ZN(n21221) );
  AOI22_X1 U23809 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20884), .B1(
        n20912), .B2(n21221), .ZN(n20880) );
  OAI211_X1 U23810 ( .C1(n21116), .C2(n20887), .A(n20881), .B(n20880), .ZN(
        P1_U3047) );
  AOI22_X1 U23811 ( .A1(n21349), .A2(n20883), .B1(n21347), .B2(n20882), .ZN(
        n20886) );
  INV_X1 U23812 ( .A(n21356), .ZN(n21225) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20884), .B1(
        n20912), .B2(n21225), .ZN(n20885) );
  OAI211_X1 U23814 ( .C1(n21123), .C2(n20887), .A(n20886), .B(n20885), .ZN(
        P1_U3048) );
  INV_X1 U23815 ( .A(n20912), .ZN(n20888) );
  NAND2_X1 U23816 ( .A1(n20888), .A2(n21265), .ZN(n20890) );
  NAND2_X1 U23817 ( .A1(n21265), .A2(n21397), .ZN(n21186) );
  OAI21_X1 U23818 ( .B1(n20890), .B2(n20946), .A(n21186), .ZN(n20895) );
  NOR2_X1 U23819 ( .A1(n20891), .A2(n21065), .ZN(n20892) );
  NOR2_X1 U23820 ( .A1(n21131), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21006) );
  INV_X1 U23821 ( .A(n21069), .ZN(n21126) );
  NOR2_X1 U23822 ( .A1(n21432), .A2(n20922), .ZN(n20925) );
  NAND2_X1 U23823 ( .A1(n21234), .A2(n20925), .ZN(n20893) );
  INV_X1 U23824 ( .A(n20893), .ZN(n20911) );
  AOI22_X1 U23825 ( .A1(n20912), .A2(n21278), .B1(n21299), .B2(n20911), .ZN(
        n20898) );
  INV_X1 U23826 ( .A(n20892), .ZN(n20894) );
  AOI22_X1 U23827 ( .A1(n20895), .A2(n20894), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20893), .ZN(n20896) );
  OAI21_X1 U23828 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n21131), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21012) );
  NAND3_X1 U23829 ( .A1(n21134), .A2(n20896), .A3(n21012), .ZN(n20913) );
  AOI22_X1 U23830 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20913), .B1(
        n20946), .B2(n21307), .ZN(n20897) );
  OAI211_X1 U23831 ( .C1(n20916), .C2(n21201), .A(n20898), .B(n20897), .ZN(
        P1_U3049) );
  INV_X1 U23832 ( .A(n21312), .ZN(n21205) );
  AOI22_X1 U23833 ( .A1(n20912), .A2(n21314), .B1(n21313), .B2(n20911), .ZN(
        n20900) );
  AOI22_X1 U23834 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20913), .B1(
        n20946), .B2(n21202), .ZN(n20899) );
  OAI211_X1 U23835 ( .C1(n20916), .C2(n21205), .A(n20900), .B(n20899), .ZN(
        P1_U3050) );
  INV_X1 U23836 ( .A(n21318), .ZN(n21414) );
  AOI22_X1 U23837 ( .A1(n20946), .A2(n21206), .B1(n21409), .B2(n20911), .ZN(
        n20902) );
  AOI22_X1 U23838 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20913), .B1(
        n20912), .B2(n21319), .ZN(n20901) );
  OAI211_X1 U23839 ( .C1(n20916), .C2(n21414), .A(n20902), .B(n20901), .ZN(
        P1_U3051) );
  INV_X1 U23840 ( .A(n21323), .ZN(n21212) );
  AOI22_X1 U23841 ( .A1(n20912), .A2(n21324), .B1(n21322), .B2(n20911), .ZN(
        n20904) );
  AOI22_X1 U23842 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20913), .B1(
        n20946), .B2(n21209), .ZN(n20903) );
  OAI211_X1 U23843 ( .C1(n20916), .C2(n21212), .A(n20904), .B(n20903), .ZN(
        P1_U3052) );
  INV_X1 U23844 ( .A(n21329), .ZN(n21216) );
  AOI22_X1 U23845 ( .A1(n20946), .A2(n21213), .B1(n21328), .B2(n20911), .ZN(
        n20906) );
  AOI22_X1 U23846 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20913), .B1(
        n20912), .B2(n21330), .ZN(n20905) );
  OAI211_X1 U23847 ( .C1(n20916), .C2(n21216), .A(n20906), .B(n20905), .ZN(
        P1_U3053) );
  AOI22_X1 U23848 ( .A1(n20912), .A2(n21336), .B1(n21334), .B2(n20911), .ZN(
        n20908) );
  AOI22_X1 U23849 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20913), .B1(
        n20946), .B2(n21217), .ZN(n20907) );
  OAI211_X1 U23850 ( .C1(n20916), .C2(n21220), .A(n20908), .B(n20907), .ZN(
        P1_U3054) );
  INV_X1 U23851 ( .A(n21341), .ZN(n21224) );
  AOI22_X1 U23852 ( .A1(n20946), .A2(n21221), .B1(n21340), .B2(n20911), .ZN(
        n20910) );
  AOI22_X1 U23853 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20913), .B1(
        n20912), .B2(n21342), .ZN(n20909) );
  OAI211_X1 U23854 ( .C1(n20916), .C2(n21224), .A(n20910), .B(n20909), .ZN(
        P1_U3055) );
  INV_X1 U23855 ( .A(n21349), .ZN(n21230) );
  AOI22_X1 U23856 ( .A1(n20912), .A2(n21350), .B1(n21347), .B2(n20911), .ZN(
        n20915) );
  AOI22_X1 U23857 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20913), .B1(
        n20946), .B2(n21225), .ZN(n20914) );
  OAI211_X1 U23858 ( .C1(n20916), .C2(n21230), .A(n20915), .B(n20914), .ZN(
        P1_U3056) );
  AOI21_X1 U23859 ( .B1(n20918), .B2(n20917), .A(n21302), .ZN(n20927) );
  INV_X1 U23860 ( .A(n20919), .ZN(n20920) );
  AND2_X1 U23861 ( .A1(n20921), .A2(n20920), .ZN(n21297) );
  NOR2_X1 U23862 ( .A1(n21296), .A2(n20922), .ZN(n20945) );
  AOI21_X1 U23863 ( .B1(n20923), .B2(n21297), .A(n20945), .ZN(n20928) );
  INV_X1 U23864 ( .A(n20928), .ZN(n20924) );
  AOI22_X1 U23865 ( .A1(n20946), .A2(n21278), .B1(n21299), .B2(n20945), .ZN(
        n20932) );
  OAI21_X1 U23866 ( .B1(n21265), .B2(n20925), .A(n21306), .ZN(n20926) );
  AOI21_X1 U23867 ( .B1(n20928), .B2(n20927), .A(n20926), .ZN(n20929) );
  AOI22_X1 U23868 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20947), .B1(
        n20976), .B2(n21307), .ZN(n20931) );
  OAI211_X1 U23869 ( .C1(n20950), .C2(n21201), .A(n20932), .B(n20931), .ZN(
        P1_U3057) );
  AOI22_X1 U23870 ( .A1(n20976), .A2(n21202), .B1(n21313), .B2(n20945), .ZN(
        n20934) );
  AOI22_X1 U23871 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20947), .B1(
        n20946), .B2(n21314), .ZN(n20933) );
  OAI211_X1 U23872 ( .C1(n20950), .C2(n21205), .A(n20934), .B(n20933), .ZN(
        P1_U3058) );
  AOI22_X1 U23873 ( .A1(n20946), .A2(n21319), .B1(n21409), .B2(n20945), .ZN(
        n20936) );
  AOI22_X1 U23874 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20947), .B1(
        n20976), .B2(n21206), .ZN(n20935) );
  OAI211_X1 U23875 ( .C1(n20950), .C2(n21414), .A(n20936), .B(n20935), .ZN(
        P1_U3059) );
  AOI22_X1 U23876 ( .A1(n20946), .A2(n21324), .B1(n21322), .B2(n20945), .ZN(
        n20938) );
  AOI22_X1 U23877 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20947), .B1(
        n20976), .B2(n21209), .ZN(n20937) );
  OAI211_X1 U23878 ( .C1(n20950), .C2(n21212), .A(n20938), .B(n20937), .ZN(
        P1_U3060) );
  AOI22_X1 U23879 ( .A1(n20946), .A2(n21330), .B1(n21328), .B2(n20945), .ZN(
        n20940) );
  AOI22_X1 U23880 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20947), .B1(
        n20976), .B2(n21213), .ZN(n20939) );
  OAI211_X1 U23881 ( .C1(n20950), .C2(n21216), .A(n20940), .B(n20939), .ZN(
        P1_U3061) );
  AOI22_X1 U23882 ( .A1(n20946), .A2(n21336), .B1(n21334), .B2(n20945), .ZN(
        n20942) );
  AOI22_X1 U23883 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20947), .B1(
        n20976), .B2(n21217), .ZN(n20941) );
  OAI211_X1 U23884 ( .C1(n20950), .C2(n21220), .A(n20942), .B(n20941), .ZN(
        P1_U3062) );
  AOI22_X1 U23885 ( .A1(n20946), .A2(n21342), .B1(n21340), .B2(n20945), .ZN(
        n20944) );
  AOI22_X1 U23886 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20947), .B1(
        n20976), .B2(n21221), .ZN(n20943) );
  OAI211_X1 U23887 ( .C1(n20950), .C2(n21224), .A(n20944), .B(n20943), .ZN(
        P1_U3063) );
  AOI22_X1 U23888 ( .A1(n20946), .A2(n21350), .B1(n21347), .B2(n20945), .ZN(
        n20949) );
  AOI22_X1 U23889 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20947), .B1(
        n20976), .B2(n21225), .ZN(n20948) );
  OAI211_X1 U23890 ( .C1(n20950), .C2(n21230), .A(n20949), .B(n20948), .ZN(
        P1_U3064) );
  INV_X1 U23891 ( .A(n21184), .ZN(n20952) );
  INV_X1 U23892 ( .A(n21190), .ZN(n21267) );
  NOR2_X1 U23893 ( .A1(n14078), .A2(n20953), .ZN(n21036) );
  NAND3_X1 U23894 ( .A1(n21036), .A2(n21265), .A3(n21065), .ZN(n20954) );
  AOI22_X1 U23895 ( .A1(n21300), .A2(n20975), .B1(n21299), .B2(n10603), .ZN(
        n20962) );
  INV_X1 U23896 ( .A(n20976), .ZN(n20956) );
  AOI21_X1 U23897 ( .B1(n20956), .B2(n21003), .A(n21397), .ZN(n20957) );
  AOI21_X1 U23898 ( .B1(n21036), .B2(n21065), .A(n20957), .ZN(n20958) );
  NOR2_X1 U23899 ( .A1(n20958), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20960) );
  AOI22_X1 U23900 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20977), .B1(
        n20976), .B2(n21278), .ZN(n20961) );
  OAI211_X1 U23901 ( .C1(n21281), .C2(n21003), .A(n20962), .B(n20961), .ZN(
        P1_U3065) );
  AOI22_X1 U23902 ( .A1(n21313), .A2(n10603), .B1(n21312), .B2(n20975), .ZN(
        n20964) );
  AOI22_X1 U23903 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20977), .B1(
        n20976), .B2(n21314), .ZN(n20963) );
  OAI211_X1 U23904 ( .C1(n21317), .C2(n21003), .A(n20964), .B(n20963), .ZN(
        P1_U3066) );
  AOI22_X1 U23905 ( .A1(n21318), .A2(n20975), .B1(n21409), .B2(n10603), .ZN(
        n20966) );
  AOI22_X1 U23906 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20977), .B1(
        n20976), .B2(n21319), .ZN(n20965) );
  OAI211_X1 U23907 ( .C1(n21416), .C2(n21003), .A(n20966), .B(n20965), .ZN(
        P1_U3067) );
  AOI22_X1 U23908 ( .A1(n21323), .A2(n20975), .B1(n21322), .B2(n10603), .ZN(
        n20968) );
  AOI22_X1 U23909 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20977), .B1(
        n20976), .B2(n21324), .ZN(n20967) );
  OAI211_X1 U23910 ( .C1(n21327), .C2(n21003), .A(n20968), .B(n20967), .ZN(
        P1_U3068) );
  AOI22_X1 U23911 ( .A1(n21329), .A2(n20975), .B1(n21328), .B2(n10603), .ZN(
        n20970) );
  AOI22_X1 U23912 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20977), .B1(
        n20976), .B2(n21330), .ZN(n20969) );
  OAI211_X1 U23913 ( .C1(n21333), .C2(n21003), .A(n20970), .B(n20969), .ZN(
        P1_U3069) );
  AOI22_X1 U23914 ( .A1(n21335), .A2(n20975), .B1(n21334), .B2(n10603), .ZN(
        n20972) );
  AOI22_X1 U23915 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20977), .B1(
        n20976), .B2(n21336), .ZN(n20971) );
  OAI211_X1 U23916 ( .C1(n21339), .C2(n21003), .A(n20972), .B(n20971), .ZN(
        P1_U3070) );
  AOI22_X1 U23917 ( .A1(n21341), .A2(n20975), .B1(n21340), .B2(n10603), .ZN(
        n20974) );
  AOI22_X1 U23918 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20977), .B1(
        n20976), .B2(n21342), .ZN(n20973) );
  OAI211_X1 U23919 ( .C1(n21345), .C2(n21003), .A(n20974), .B(n20973), .ZN(
        P1_U3071) );
  AOI22_X1 U23920 ( .A1(n21349), .A2(n20975), .B1(n21347), .B2(n10603), .ZN(
        n20979) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20977), .B1(
        n20976), .B2(n21350), .ZN(n20978) );
  OAI211_X1 U23922 ( .C1(n21356), .C2(n21003), .A(n20979), .B(n20978), .ZN(
        P1_U3072) );
  NOR2_X1 U23923 ( .A1(n21007), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20983) );
  INV_X1 U23924 ( .A(n20983), .ZN(n20980) );
  NOR2_X1 U23925 ( .A1(n21234), .A2(n20980), .ZN(n20998) );
  AOI21_X1 U23926 ( .B1(n21036), .B2(n21235), .A(n20998), .ZN(n20981) );
  OAI22_X1 U23927 ( .A1(n20981), .A2(n21302), .B1(n20980), .B2(n12586), .ZN(
        n20999) );
  AOI22_X1 U23928 ( .A1(n21300), .A2(n20999), .B1(n21299), .B2(n20998), .ZN(
        n20985) );
  OAI21_X1 U23929 ( .B1(n21039), .B2(n21238), .A(n20981), .ZN(n20982) );
  OAI221_X1 U23930 ( .B1(n21265), .B2(n20983), .C1(n21302), .C2(n20982), .A(
        n21306), .ZN(n21000) );
  AOI22_X1 U23931 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21000), .B1(
        n21030), .B2(n21307), .ZN(n20984) );
  OAI211_X1 U23932 ( .C1(n21311), .C2(n21003), .A(n20985), .B(n20984), .ZN(
        P1_U3073) );
  AOI22_X1 U23933 ( .A1(n21313), .A2(n20998), .B1(n21312), .B2(n20999), .ZN(
        n20987) );
  AOI22_X1 U23934 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21000), .B1(
        n21030), .B2(n21202), .ZN(n20986) );
  OAI211_X1 U23935 ( .C1(n21102), .C2(n21003), .A(n20987), .B(n20986), .ZN(
        P1_U3074) );
  AOI22_X1 U23936 ( .A1(n21318), .A2(n20999), .B1(n21409), .B2(n20998), .ZN(
        n20989) );
  AOI22_X1 U23937 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21000), .B1(
        n21030), .B2(n21206), .ZN(n20988) );
  OAI211_X1 U23938 ( .C1(n21418), .C2(n21003), .A(n20989), .B(n20988), .ZN(
        P1_U3075) );
  AOI22_X1 U23939 ( .A1(n21323), .A2(n20999), .B1(n21322), .B2(n20998), .ZN(
        n20991) );
  AOI22_X1 U23940 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21000), .B1(
        n21030), .B2(n21209), .ZN(n20990) );
  OAI211_X1 U23941 ( .C1(n21107), .C2(n21003), .A(n20991), .B(n20990), .ZN(
        P1_U3076) );
  AOI22_X1 U23942 ( .A1(n21329), .A2(n20999), .B1(n21328), .B2(n20998), .ZN(
        n20993) );
  AOI22_X1 U23943 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21000), .B1(
        n21030), .B2(n21213), .ZN(n20992) );
  OAI211_X1 U23944 ( .C1(n21110), .C2(n21003), .A(n20993), .B(n20992), .ZN(
        P1_U3077) );
  AOI22_X1 U23945 ( .A1(n21335), .A2(n20999), .B1(n21334), .B2(n20998), .ZN(
        n20995) );
  AOI22_X1 U23946 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21000), .B1(
        n21030), .B2(n21217), .ZN(n20994) );
  OAI211_X1 U23947 ( .C1(n21113), .C2(n21003), .A(n20995), .B(n20994), .ZN(
        P1_U3078) );
  AOI22_X1 U23948 ( .A1(n21341), .A2(n20999), .B1(n21340), .B2(n20998), .ZN(
        n20997) );
  AOI22_X1 U23949 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21000), .B1(
        n21030), .B2(n21221), .ZN(n20996) );
  OAI211_X1 U23950 ( .C1(n21116), .C2(n21003), .A(n20997), .B(n20996), .ZN(
        P1_U3079) );
  AOI22_X1 U23951 ( .A1(n21349), .A2(n20999), .B1(n21347), .B2(n20998), .ZN(
        n21002) );
  AOI22_X1 U23952 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21000), .B1(
        n21030), .B2(n21225), .ZN(n21001) );
  OAI211_X1 U23953 ( .C1(n21123), .C2(n21003), .A(n21002), .B(n21001), .ZN(
        P1_U3080) );
  NAND3_X1 U23954 ( .A1(n21014), .A2(n21004), .A3(n21265), .ZN(n21005) );
  NAND2_X1 U23955 ( .A1(n21005), .A2(n21186), .ZN(n21011) );
  AND2_X1 U23956 ( .A1(n21036), .A2(n21273), .ZN(n21008) );
  NOR2_X1 U23957 ( .A1(n21432), .A2(n21007), .ZN(n21041) );
  NAND2_X1 U23958 ( .A1(n21234), .A2(n21041), .ZN(n21009) );
  INV_X1 U23959 ( .A(n21009), .ZN(n21029) );
  AOI22_X1 U23960 ( .A1(n21299), .A2(n21029), .B1(n21030), .B2(n21278), .ZN(
        n21016) );
  INV_X1 U23961 ( .A(n21008), .ZN(n21010) );
  AOI22_X1 U23962 ( .A1(n21011), .A2(n21010), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21009), .ZN(n21013) );
  NAND3_X1 U23963 ( .A1(n21276), .A2(n21013), .A3(n21012), .ZN(n21031) );
  AOI22_X1 U23964 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n21031), .B1(
        n21058), .B2(n21307), .ZN(n21015) );
  OAI211_X1 U23965 ( .C1(n21034), .C2(n21201), .A(n21016), .B(n21015), .ZN(
        P1_U3081) );
  AOI22_X1 U23966 ( .A1(n21313), .A2(n21029), .B1(n21058), .B2(n21202), .ZN(
        n21018) );
  AOI22_X1 U23967 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n21031), .B1(
        n21030), .B2(n21314), .ZN(n21017) );
  OAI211_X1 U23968 ( .C1(n21034), .C2(n21205), .A(n21018), .B(n21017), .ZN(
        P1_U3082) );
  AOI22_X1 U23969 ( .A1(n21409), .A2(n21029), .B1(n21030), .B2(n21319), .ZN(
        n21020) );
  AOI22_X1 U23970 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n21031), .B1(
        n21058), .B2(n21206), .ZN(n21019) );
  OAI211_X1 U23971 ( .C1(n21034), .C2(n21414), .A(n21020), .B(n21019), .ZN(
        P1_U3083) );
  AOI22_X1 U23972 ( .A1(n21322), .A2(n21029), .B1(n21030), .B2(n21324), .ZN(
        n21022) );
  AOI22_X1 U23973 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n21031), .B1(
        n21058), .B2(n21209), .ZN(n21021) );
  OAI211_X1 U23974 ( .C1(n21034), .C2(n21212), .A(n21022), .B(n21021), .ZN(
        P1_U3084) );
  AOI22_X1 U23975 ( .A1(n21328), .A2(n21029), .B1(n21058), .B2(n21213), .ZN(
        n21024) );
  AOI22_X1 U23976 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n21031), .B1(
        n21030), .B2(n21330), .ZN(n21023) );
  OAI211_X1 U23977 ( .C1(n21034), .C2(n21216), .A(n21024), .B(n21023), .ZN(
        P1_U3085) );
  AOI22_X1 U23978 ( .A1(n21334), .A2(n21029), .B1(n21058), .B2(n21217), .ZN(
        n21026) );
  AOI22_X1 U23979 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n21031), .B1(
        n21030), .B2(n21336), .ZN(n21025) );
  OAI211_X1 U23980 ( .C1(n21034), .C2(n21220), .A(n21026), .B(n21025), .ZN(
        P1_U3086) );
  AOI22_X1 U23981 ( .A1(n21340), .A2(n21029), .B1(n21030), .B2(n21342), .ZN(
        n21028) );
  AOI22_X1 U23982 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n21031), .B1(
        n21058), .B2(n21221), .ZN(n21027) );
  OAI211_X1 U23983 ( .C1(n21034), .C2(n21224), .A(n21028), .B(n21027), .ZN(
        P1_U3087) );
  AOI22_X1 U23984 ( .A1(n21347), .A2(n21029), .B1(n21058), .B2(n21225), .ZN(
        n21033) );
  AOI22_X1 U23985 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n21031), .B1(
        n21030), .B2(n21350), .ZN(n21032) );
  OAI211_X1 U23986 ( .C1(n21034), .C2(n21230), .A(n21033), .B(n21032), .ZN(
        P1_U3088) );
  INV_X1 U23987 ( .A(n21035), .ZN(n21056) );
  AOI21_X1 U23988 ( .B1(n21036), .B2(n21297), .A(n21056), .ZN(n21038) );
  INV_X1 U23989 ( .A(n21041), .ZN(n21037) );
  OAI22_X1 U23990 ( .A1(n21038), .A2(n21302), .B1(n21037), .B2(n12586), .ZN(
        n21057) );
  AOI22_X1 U23991 ( .A1(n21300), .A2(n21057), .B1(n21056), .B2(n21299), .ZN(
        n21043) );
  OAI211_X1 U23992 ( .C1(n21039), .C2(n21160), .A(n21265), .B(n21038), .ZN(
        n21040) );
  OAI211_X1 U23993 ( .C1(n21265), .C2(n21041), .A(n21040), .B(n21306), .ZN(
        n21059) );
  AOI22_X1 U23994 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n21059), .B1(
        n21058), .B2(n21278), .ZN(n21042) );
  OAI211_X1 U23995 ( .C1(n21281), .C2(n21070), .A(n21043), .B(n21042), .ZN(
        P1_U3089) );
  AOI22_X1 U23996 ( .A1(n21313), .A2(n21056), .B1(n21312), .B2(n21057), .ZN(
        n21045) );
  AOI22_X1 U23997 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n21059), .B1(
        n21058), .B2(n21314), .ZN(n21044) );
  OAI211_X1 U23998 ( .C1(n21317), .C2(n21070), .A(n21045), .B(n21044), .ZN(
        P1_U3090) );
  AOI22_X1 U23999 ( .A1(n21318), .A2(n21057), .B1(n21056), .B2(n21409), .ZN(
        n21047) );
  AOI22_X1 U24000 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n21059), .B1(
        n21058), .B2(n21319), .ZN(n21046) );
  OAI211_X1 U24001 ( .C1(n21416), .C2(n21070), .A(n21047), .B(n21046), .ZN(
        P1_U3091) );
  AOI22_X1 U24002 ( .A1(n21323), .A2(n21057), .B1(n21056), .B2(n21322), .ZN(
        n21049) );
  AOI22_X1 U24003 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n21059), .B1(
        n21058), .B2(n21324), .ZN(n21048) );
  OAI211_X1 U24004 ( .C1(n21327), .C2(n21070), .A(n21049), .B(n21048), .ZN(
        P1_U3092) );
  AOI22_X1 U24005 ( .A1(n21329), .A2(n21057), .B1(n21056), .B2(n21328), .ZN(
        n21051) );
  AOI22_X1 U24006 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n21059), .B1(
        n21058), .B2(n21330), .ZN(n21050) );
  OAI211_X1 U24007 ( .C1(n21333), .C2(n21070), .A(n21051), .B(n21050), .ZN(
        P1_U3093) );
  AOI22_X1 U24008 ( .A1(n21335), .A2(n21057), .B1(n21056), .B2(n21334), .ZN(
        n21053) );
  AOI22_X1 U24009 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n21059), .B1(
        n21058), .B2(n21336), .ZN(n21052) );
  OAI211_X1 U24010 ( .C1(n21339), .C2(n21070), .A(n21053), .B(n21052), .ZN(
        P1_U3094) );
  AOI22_X1 U24011 ( .A1(n21341), .A2(n21057), .B1(n21056), .B2(n21340), .ZN(
        n21055) );
  AOI22_X1 U24012 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n21059), .B1(
        n21058), .B2(n21342), .ZN(n21054) );
  OAI211_X1 U24013 ( .C1(n21345), .C2(n21070), .A(n21055), .B(n21054), .ZN(
        P1_U3095) );
  AOI22_X1 U24014 ( .A1(n21349), .A2(n21057), .B1(n21056), .B2(n21347), .ZN(
        n21061) );
  AOI22_X1 U24015 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n21059), .B1(
        n21058), .B2(n21350), .ZN(n21060) );
  OAI211_X1 U24016 ( .C1(n21356), .C2(n21070), .A(n21061), .B(n21060), .ZN(
        P1_U3096) );
  INV_X1 U24017 ( .A(n21161), .ZN(n21062) );
  AND2_X1 U24018 ( .A1(n21063), .A2(n14078), .ZN(n21157) );
  NAND2_X1 U24019 ( .A1(n21064), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21156) );
  AOI21_X1 U24020 ( .B1(n21157), .B2(n21065), .A(n10593), .ZN(n21072) );
  INV_X1 U24021 ( .A(n21066), .ZN(n21068) );
  NOR2_X1 U24022 ( .A1(n21068), .A2(n21067), .ZN(n21189) );
  INV_X1 U24023 ( .A(n21189), .ZN(n21193) );
  OAI22_X1 U24024 ( .A1(n21072), .A2(n21302), .B1(n21069), .B2(n21193), .ZN(
        n21089) );
  AOI22_X1 U24025 ( .A1(n21300), .A2(n21089), .B1(n21299), .B2(n10593), .ZN(
        n21076) );
  INV_X1 U24026 ( .A(n21122), .ZN(n21071) );
  OAI21_X1 U24027 ( .B1(n21071), .B2(n21090), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21073) );
  NAND2_X1 U24028 ( .A1(n21073), .A2(n21072), .ZN(n21074) );
  AOI22_X1 U24029 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n21091), .B1(
        n21090), .B2(n21278), .ZN(n21075) );
  OAI211_X1 U24030 ( .C1(n21281), .C2(n21122), .A(n21076), .B(n21075), .ZN(
        P1_U3097) );
  AOI22_X1 U24031 ( .A1(n21313), .A2(n10593), .B1(n21312), .B2(n21089), .ZN(
        n21078) );
  AOI22_X1 U24032 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21091), .B1(
        n21090), .B2(n21314), .ZN(n21077) );
  OAI211_X1 U24033 ( .C1(n21317), .C2(n21122), .A(n21078), .B(n21077), .ZN(
        P1_U3098) );
  AOI22_X1 U24034 ( .A1(n21318), .A2(n21089), .B1(n21409), .B2(n10593), .ZN(
        n21080) );
  AOI22_X1 U24035 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n21091), .B1(
        n21090), .B2(n21319), .ZN(n21079) );
  OAI211_X1 U24036 ( .C1(n21416), .C2(n21122), .A(n21080), .B(n21079), .ZN(
        P1_U3099) );
  AOI22_X1 U24037 ( .A1(n21323), .A2(n21089), .B1(n21322), .B2(n10593), .ZN(
        n21082) );
  AOI22_X1 U24038 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n21091), .B1(
        n21090), .B2(n21324), .ZN(n21081) );
  OAI211_X1 U24039 ( .C1(n21327), .C2(n21122), .A(n21082), .B(n21081), .ZN(
        P1_U3100) );
  AOI22_X1 U24040 ( .A1(n21329), .A2(n21089), .B1(n21328), .B2(n10593), .ZN(
        n21084) );
  AOI22_X1 U24041 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n21091), .B1(
        n21090), .B2(n21330), .ZN(n21083) );
  OAI211_X1 U24042 ( .C1(n21333), .C2(n21122), .A(n21084), .B(n21083), .ZN(
        P1_U3101) );
  AOI22_X1 U24043 ( .A1(n21335), .A2(n21089), .B1(n21334), .B2(n10593), .ZN(
        n21086) );
  AOI22_X1 U24044 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n21091), .B1(
        n21090), .B2(n21336), .ZN(n21085) );
  OAI211_X1 U24045 ( .C1(n21339), .C2(n21122), .A(n21086), .B(n21085), .ZN(
        P1_U3102) );
  AOI22_X1 U24046 ( .A1(n21341), .A2(n21089), .B1(n21340), .B2(n10593), .ZN(
        n21088) );
  AOI22_X1 U24047 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n21091), .B1(
        n21090), .B2(n21342), .ZN(n21087) );
  OAI211_X1 U24048 ( .C1(n21345), .C2(n21122), .A(n21088), .B(n21087), .ZN(
        P1_U3103) );
  AOI22_X1 U24049 ( .A1(n21349), .A2(n21089), .B1(n21347), .B2(n10593), .ZN(
        n21093) );
  AOI22_X1 U24050 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n21091), .B1(
        n21090), .B2(n21350), .ZN(n21092) );
  OAI211_X1 U24051 ( .C1(n21356), .C2(n21122), .A(n21093), .B(n21092), .ZN(
        P1_U3104) );
  NOR2_X1 U24052 ( .A1(n21156), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21096) );
  INV_X1 U24053 ( .A(n21096), .ZN(n21094) );
  NOR2_X1 U24054 ( .A1(n21234), .A2(n21094), .ZN(n21117) );
  AOI21_X1 U24055 ( .B1(n21157), .B2(n21235), .A(n21117), .ZN(n21095) );
  OAI22_X1 U24056 ( .A1(n21095), .A2(n21302), .B1(n21094), .B2(n12586), .ZN(
        n21118) );
  AOI22_X1 U24057 ( .A1(n21300), .A2(n21118), .B1(n21299), .B2(n21117), .ZN(
        n21099) );
  NOR3_X1 U24058 ( .A1(n21161), .A2(n21302), .A3(n21238), .ZN(n21097) );
  AOI22_X1 U24059 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21119), .B1(
        n21150), .B2(n21307), .ZN(n21098) );
  OAI211_X1 U24060 ( .C1(n21311), .C2(n21122), .A(n21099), .B(n21098), .ZN(
        P1_U3105) );
  AOI22_X1 U24061 ( .A1(n21313), .A2(n21117), .B1(n21312), .B2(n21118), .ZN(
        n21101) );
  AOI22_X1 U24062 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21119), .B1(
        n21150), .B2(n21202), .ZN(n21100) );
  OAI211_X1 U24063 ( .C1(n21102), .C2(n21122), .A(n21101), .B(n21100), .ZN(
        P1_U3106) );
  AOI22_X1 U24064 ( .A1(n21318), .A2(n21118), .B1(n21409), .B2(n21117), .ZN(
        n21104) );
  AOI22_X1 U24065 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21119), .B1(
        n21150), .B2(n21206), .ZN(n21103) );
  OAI211_X1 U24066 ( .C1(n21418), .C2(n21122), .A(n21104), .B(n21103), .ZN(
        P1_U3107) );
  AOI22_X1 U24067 ( .A1(n21323), .A2(n21118), .B1(n21322), .B2(n21117), .ZN(
        n21106) );
  AOI22_X1 U24068 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21119), .B1(
        n21150), .B2(n21209), .ZN(n21105) );
  OAI211_X1 U24069 ( .C1(n21107), .C2(n21122), .A(n21106), .B(n21105), .ZN(
        P1_U3108) );
  AOI22_X1 U24070 ( .A1(n21329), .A2(n21118), .B1(n21328), .B2(n21117), .ZN(
        n21109) );
  AOI22_X1 U24071 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21119), .B1(
        n21150), .B2(n21213), .ZN(n21108) );
  OAI211_X1 U24072 ( .C1(n21110), .C2(n21122), .A(n21109), .B(n21108), .ZN(
        P1_U3109) );
  AOI22_X1 U24073 ( .A1(n21335), .A2(n21118), .B1(n21334), .B2(n21117), .ZN(
        n21112) );
  AOI22_X1 U24074 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21119), .B1(
        n21150), .B2(n21217), .ZN(n21111) );
  OAI211_X1 U24075 ( .C1(n21113), .C2(n21122), .A(n21112), .B(n21111), .ZN(
        P1_U3110) );
  AOI22_X1 U24076 ( .A1(n21341), .A2(n21118), .B1(n21340), .B2(n21117), .ZN(
        n21115) );
  AOI22_X1 U24077 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21119), .B1(
        n21150), .B2(n21221), .ZN(n21114) );
  OAI211_X1 U24078 ( .C1(n21116), .C2(n21122), .A(n21115), .B(n21114), .ZN(
        P1_U3111) );
  AOI22_X1 U24079 ( .A1(n21349), .A2(n21118), .B1(n21347), .B2(n21117), .ZN(
        n21121) );
  AOI22_X1 U24080 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21119), .B1(
        n21150), .B2(n21225), .ZN(n21120) );
  OAI211_X1 U24081 ( .C1(n21123), .C2(n21122), .A(n21121), .B(n21120), .ZN(
        P1_U3112) );
  INV_X1 U24082 ( .A(n21150), .ZN(n21124) );
  NAND2_X1 U24083 ( .A1(n21124), .A2(n21265), .ZN(n21125) );
  OAI21_X1 U24084 ( .B1(n21125), .B2(n21180), .A(n21186), .ZN(n21130) );
  AND2_X1 U24085 ( .A1(n21157), .A2(n21273), .ZN(n21127) );
  NOR2_X1 U24086 ( .A1(n21131), .A2(n21132), .ZN(n21266) );
  NOR2_X1 U24087 ( .A1(n21432), .A2(n21156), .ZN(n21163) );
  NAND2_X1 U24088 ( .A1(n21234), .A2(n21163), .ZN(n21128) );
  AOI22_X1 U24089 ( .A1(n21180), .A2(n21307), .B1(n21299), .B2(n21149), .ZN(
        n21136) );
  INV_X1 U24090 ( .A(n21127), .ZN(n21129) );
  AOI22_X1 U24091 ( .A1(n21130), .A2(n21129), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21128), .ZN(n21133) );
  OAI21_X1 U24092 ( .B1(n21132), .B2(n21131), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n21275) );
  NAND3_X1 U24093 ( .A1(n21134), .A2(n21133), .A3(n21275), .ZN(n21151) );
  AOI22_X1 U24094 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21151), .B1(
        n21150), .B2(n21278), .ZN(n21135) );
  OAI211_X1 U24095 ( .C1(n21154), .C2(n21201), .A(n21136), .B(n21135), .ZN(
        P1_U3113) );
  AOI22_X1 U24096 ( .A1(n21180), .A2(n21202), .B1(n21313), .B2(n21149), .ZN(
        n21138) );
  AOI22_X1 U24097 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21151), .B1(
        n21150), .B2(n21314), .ZN(n21137) );
  OAI211_X1 U24098 ( .C1(n21154), .C2(n21205), .A(n21138), .B(n21137), .ZN(
        P1_U3114) );
  AOI22_X1 U24099 ( .A1(n21150), .A2(n21319), .B1(n21409), .B2(n21149), .ZN(
        n21140) );
  AOI22_X1 U24100 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21151), .B1(
        n21180), .B2(n21206), .ZN(n21139) );
  OAI211_X1 U24101 ( .C1(n21154), .C2(n21414), .A(n21140), .B(n21139), .ZN(
        P1_U3115) );
  AOI22_X1 U24102 ( .A1(n21180), .A2(n21209), .B1(n21322), .B2(n21149), .ZN(
        n21142) );
  AOI22_X1 U24103 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21151), .B1(
        n21150), .B2(n21324), .ZN(n21141) );
  OAI211_X1 U24104 ( .C1(n21154), .C2(n21212), .A(n21142), .B(n21141), .ZN(
        P1_U3116) );
  AOI22_X1 U24105 ( .A1(n21150), .A2(n21330), .B1(n21328), .B2(n21149), .ZN(
        n21144) );
  AOI22_X1 U24106 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21151), .B1(
        n21180), .B2(n21213), .ZN(n21143) );
  OAI211_X1 U24107 ( .C1(n21154), .C2(n21216), .A(n21144), .B(n21143), .ZN(
        P1_U3117) );
  AOI22_X1 U24108 ( .A1(n21150), .A2(n21336), .B1(n21334), .B2(n21149), .ZN(
        n21146) );
  AOI22_X1 U24109 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21151), .B1(
        n21180), .B2(n21217), .ZN(n21145) );
  OAI211_X1 U24110 ( .C1(n21154), .C2(n21220), .A(n21146), .B(n21145), .ZN(
        P1_U3118) );
  AOI22_X1 U24111 ( .A1(n21150), .A2(n21342), .B1(n21340), .B2(n21149), .ZN(
        n21148) );
  AOI22_X1 U24112 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21151), .B1(
        n21180), .B2(n21221), .ZN(n21147) );
  OAI211_X1 U24113 ( .C1(n21154), .C2(n21224), .A(n21148), .B(n21147), .ZN(
        P1_U3119) );
  AOI22_X1 U24114 ( .A1(n21150), .A2(n21350), .B1(n21347), .B2(n21149), .ZN(
        n21153) );
  AOI22_X1 U24115 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21151), .B1(
        n21180), .B2(n21225), .ZN(n21152) );
  OAI211_X1 U24116 ( .C1(n21154), .C2(n21230), .A(n21153), .B(n21152), .ZN(
        P1_U3120) );
  NOR2_X1 U24117 ( .A1(n21296), .A2(n21156), .ZN(n21178) );
  AOI21_X1 U24118 ( .B1(n21157), .B2(n21297), .A(n21178), .ZN(n21159) );
  INV_X1 U24119 ( .A(n21163), .ZN(n21158) );
  OAI22_X1 U24120 ( .A1(n21159), .A2(n21302), .B1(n21158), .B2(n12586), .ZN(
        n21179) );
  AOI22_X1 U24121 ( .A1(n21300), .A2(n21179), .B1(n21299), .B2(n21178), .ZN(
        n21165) );
  OAI21_X1 U24122 ( .B1(n21161), .B2(n21160), .A(n21159), .ZN(n21162) );
  OAI221_X1 U24123 ( .B1(n21265), .B2(n21163), .C1(n21302), .C2(n21162), .A(
        n21306), .ZN(n21181) );
  AOI22_X1 U24124 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21278), .ZN(n21164) );
  OAI211_X1 U24125 ( .C1(n21281), .C2(n21198), .A(n21165), .B(n21164), .ZN(
        P1_U3121) );
  AOI22_X1 U24126 ( .A1(n21313), .A2(n21178), .B1(n21312), .B2(n21179), .ZN(
        n21167) );
  AOI22_X1 U24127 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21314), .ZN(n21166) );
  OAI211_X1 U24128 ( .C1(n21317), .C2(n21198), .A(n21167), .B(n21166), .ZN(
        P1_U3122) );
  AOI22_X1 U24129 ( .A1(n21318), .A2(n21179), .B1(n21409), .B2(n21178), .ZN(
        n21169) );
  AOI22_X1 U24130 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21319), .ZN(n21168) );
  OAI211_X1 U24131 ( .C1(n21416), .C2(n21198), .A(n21169), .B(n21168), .ZN(
        P1_U3123) );
  AOI22_X1 U24132 ( .A1(n21323), .A2(n21179), .B1(n21322), .B2(n21178), .ZN(
        n21171) );
  AOI22_X1 U24133 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21324), .ZN(n21170) );
  OAI211_X1 U24134 ( .C1(n21327), .C2(n21198), .A(n21171), .B(n21170), .ZN(
        P1_U3124) );
  AOI22_X1 U24135 ( .A1(n21329), .A2(n21179), .B1(n21328), .B2(n21178), .ZN(
        n21173) );
  AOI22_X1 U24136 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21330), .ZN(n21172) );
  OAI211_X1 U24137 ( .C1(n21333), .C2(n21198), .A(n21173), .B(n21172), .ZN(
        P1_U3125) );
  AOI22_X1 U24138 ( .A1(n21335), .A2(n21179), .B1(n21334), .B2(n21178), .ZN(
        n21175) );
  AOI22_X1 U24139 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21336), .ZN(n21174) );
  OAI211_X1 U24140 ( .C1(n21339), .C2(n21198), .A(n21175), .B(n21174), .ZN(
        P1_U3126) );
  AOI22_X1 U24141 ( .A1(n21341), .A2(n21179), .B1(n21340), .B2(n21178), .ZN(
        n21177) );
  AOI22_X1 U24142 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21342), .ZN(n21176) );
  OAI211_X1 U24143 ( .C1(n21345), .C2(n21198), .A(n21177), .B(n21176), .ZN(
        P1_U3127) );
  AOI22_X1 U24144 ( .A1(n21349), .A2(n21179), .B1(n21347), .B2(n21178), .ZN(
        n21183) );
  AOI22_X1 U24145 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21181), .B1(
        n21180), .B2(n21350), .ZN(n21182) );
  OAI211_X1 U24146 ( .C1(n21356), .C2(n21198), .A(n21183), .B(n21182), .ZN(
        P1_U3128) );
  INV_X1 U24147 ( .A(n21258), .ZN(n21185) );
  NAND3_X1 U24148 ( .A1(n21185), .A2(n21265), .A3(n21198), .ZN(n21187) );
  NAND2_X1 U24149 ( .A1(n21187), .A2(n21186), .ZN(n21195) );
  NOR2_X1 U24150 ( .A1(n21270), .A2(n21273), .ZN(n21192) );
  NAND2_X1 U24151 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21295) );
  AOI22_X1 U24152 ( .A1(n21258), .A2(n21307), .B1(n21299), .B2(n10602), .ZN(
        n21200) );
  INV_X1 U24153 ( .A(n21192), .ZN(n21194) );
  AOI22_X1 U24154 ( .A1(n21195), .A2(n21194), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21193), .ZN(n21196) );
  AOI22_X1 U24155 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21227), .B1(
        n21226), .B2(n21278), .ZN(n21199) );
  OAI211_X1 U24156 ( .C1(n21231), .C2(n21201), .A(n21200), .B(n21199), .ZN(
        P1_U3129) );
  AOI22_X1 U24157 ( .A1(n21258), .A2(n21202), .B1(n21313), .B2(n10602), .ZN(
        n21204) );
  AOI22_X1 U24158 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21227), .B1(
        n21226), .B2(n21314), .ZN(n21203) );
  OAI211_X1 U24159 ( .C1(n21231), .C2(n21205), .A(n21204), .B(n21203), .ZN(
        P1_U3130) );
  AOI22_X1 U24160 ( .A1(n21258), .A2(n21206), .B1(n21409), .B2(n10602), .ZN(
        n21208) );
  AOI22_X1 U24161 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21227), .B1(
        n21226), .B2(n21319), .ZN(n21207) );
  OAI211_X1 U24162 ( .C1(n21231), .C2(n21414), .A(n21208), .B(n21207), .ZN(
        P1_U3131) );
  AOI22_X1 U24163 ( .A1(n21258), .A2(n21209), .B1(n21322), .B2(n10602), .ZN(
        n21211) );
  AOI22_X1 U24164 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21227), .B1(
        n21226), .B2(n21324), .ZN(n21210) );
  OAI211_X1 U24165 ( .C1(n21231), .C2(n21212), .A(n21211), .B(n21210), .ZN(
        P1_U3132) );
  AOI22_X1 U24166 ( .A1(n21258), .A2(n21213), .B1(n21328), .B2(n10602), .ZN(
        n21215) );
  AOI22_X1 U24167 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21227), .B1(
        n21226), .B2(n21330), .ZN(n21214) );
  OAI211_X1 U24168 ( .C1(n21231), .C2(n21216), .A(n21215), .B(n21214), .ZN(
        P1_U3133) );
  AOI22_X1 U24169 ( .A1(n21258), .A2(n21217), .B1(n21334), .B2(n10602), .ZN(
        n21219) );
  AOI22_X1 U24170 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21227), .B1(
        n21226), .B2(n21336), .ZN(n21218) );
  OAI211_X1 U24171 ( .C1(n21231), .C2(n21220), .A(n21219), .B(n21218), .ZN(
        P1_U3134) );
  AOI22_X1 U24172 ( .A1(n21258), .A2(n21221), .B1(n21340), .B2(n10602), .ZN(
        n21223) );
  AOI22_X1 U24173 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21227), .B1(
        n21226), .B2(n21342), .ZN(n21222) );
  OAI211_X1 U24174 ( .C1(n21231), .C2(n21224), .A(n21223), .B(n21222), .ZN(
        P1_U3135) );
  AOI22_X1 U24175 ( .A1(n21258), .A2(n21225), .B1(n21347), .B2(n10602), .ZN(
        n21229) );
  AOI22_X1 U24176 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21227), .B1(
        n21226), .B2(n21350), .ZN(n21228) );
  OAI211_X1 U24177 ( .C1(n21231), .C2(n21230), .A(n21229), .B(n21228), .ZN(
        P1_U3136) );
  INV_X1 U24178 ( .A(n21232), .ZN(n21233) );
  INV_X1 U24179 ( .A(n21270), .ZN(n21298) );
  NOR2_X1 U24180 ( .A1(n21295), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21241) );
  INV_X1 U24181 ( .A(n21241), .ZN(n21236) );
  NOR2_X1 U24182 ( .A1(n21234), .A2(n21236), .ZN(n21256) );
  AOI21_X1 U24183 ( .B1(n21298), .B2(n21235), .A(n21256), .ZN(n21237) );
  OAI22_X1 U24184 ( .A1(n21237), .A2(n21302), .B1(n21236), .B2(n12586), .ZN(
        n21257) );
  AOI22_X1 U24185 ( .A1(n21300), .A2(n21257), .B1(n21299), .B2(n21256), .ZN(
        n21243) );
  INV_X1 U24186 ( .A(n21264), .ZN(n21239) );
  OAI21_X1 U24187 ( .B1(n21239), .B2(n21238), .A(n21237), .ZN(n21240) );
  OAI221_X1 U24188 ( .B1(n21265), .B2(n21241), .C1(n21302), .C2(n21240), .A(
        n21306), .ZN(n21259) );
  AOI22_X1 U24189 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21259), .B1(
        n21258), .B2(n21278), .ZN(n21242) );
  OAI211_X1 U24190 ( .C1(n21281), .C2(n21417), .A(n21243), .B(n21242), .ZN(
        P1_U3137) );
  AOI22_X1 U24191 ( .A1(n21313), .A2(n21256), .B1(n21312), .B2(n21257), .ZN(
        n21245) );
  AOI22_X1 U24192 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21259), .B1(
        n21258), .B2(n21314), .ZN(n21244) );
  OAI211_X1 U24193 ( .C1(n21317), .C2(n21417), .A(n21245), .B(n21244), .ZN(
        P1_U3138) );
  AOI22_X1 U24194 ( .A1(n21318), .A2(n21257), .B1(n21409), .B2(n21256), .ZN(
        n21247) );
  AOI22_X1 U24195 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21259), .B1(
        n21258), .B2(n21319), .ZN(n21246) );
  OAI211_X1 U24196 ( .C1(n21416), .C2(n21417), .A(n21247), .B(n21246), .ZN(
        P1_U3139) );
  AOI22_X1 U24197 ( .A1(n21323), .A2(n21257), .B1(n21322), .B2(n21256), .ZN(
        n21249) );
  AOI22_X1 U24198 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21259), .B1(
        n21258), .B2(n21324), .ZN(n21248) );
  OAI211_X1 U24199 ( .C1(n21327), .C2(n21417), .A(n21249), .B(n21248), .ZN(
        P1_U3140) );
  AOI22_X1 U24200 ( .A1(n21329), .A2(n21257), .B1(n21328), .B2(n21256), .ZN(
        n21251) );
  AOI22_X1 U24201 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21259), .B1(
        n21258), .B2(n21330), .ZN(n21250) );
  OAI211_X1 U24202 ( .C1(n21333), .C2(n21417), .A(n21251), .B(n21250), .ZN(
        P1_U3141) );
  AOI22_X1 U24203 ( .A1(n21335), .A2(n21257), .B1(n21334), .B2(n21256), .ZN(
        n21253) );
  AOI22_X1 U24204 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21259), .B1(
        n21258), .B2(n21336), .ZN(n21252) );
  OAI211_X1 U24205 ( .C1(n21339), .C2(n21417), .A(n21253), .B(n21252), .ZN(
        P1_U3142) );
  AOI22_X1 U24206 ( .A1(n21341), .A2(n21257), .B1(n21340), .B2(n21256), .ZN(
        n21255) );
  AOI22_X1 U24207 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21259), .B1(
        n21258), .B2(n21342), .ZN(n21254) );
  OAI211_X1 U24208 ( .C1(n21345), .C2(n21417), .A(n21255), .B(n21254), .ZN(
        P1_U3143) );
  AOI22_X1 U24209 ( .A1(n21349), .A2(n21257), .B1(n21347), .B2(n21256), .ZN(
        n21261) );
  AOI22_X1 U24210 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21259), .B1(
        n21258), .B2(n21350), .ZN(n21260) );
  OAI211_X1 U24211 ( .C1(n21356), .C2(n21417), .A(n21261), .B(n21260), .ZN(
        P1_U3144) );
  INV_X1 U24212 ( .A(n21262), .ZN(n21263) );
  NAND2_X1 U24213 ( .A1(n21273), .A2(n21265), .ZN(n21269) );
  INV_X1 U24214 ( .A(n21266), .ZN(n21268) );
  OAI22_X1 U24215 ( .A1(n21270), .A2(n21269), .B1(n21268), .B2(n21267), .ZN(
        n21408) );
  INV_X1 U24216 ( .A(n21295), .ZN(n21271) );
  NAND2_X1 U24217 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21271), .ZN(
        n21301) );
  NOR2_X1 U24218 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21301), .ZN(
        n21410) );
  AOI22_X1 U24219 ( .A1(n21300), .A2(n21408), .B1(n21410), .B2(n21299), .ZN(
        n21280) );
  AOI21_X1 U24220 ( .B1(n21415), .B2(n21417), .A(n21397), .ZN(n21272) );
  AOI21_X1 U24221 ( .B1(n21298), .B2(n21273), .A(n21272), .ZN(n21274) );
  NOR2_X1 U24222 ( .A1(n21274), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21277) );
  AOI22_X1 U24223 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21421), .B1(
        n21292), .B2(n21278), .ZN(n21279) );
  OAI211_X1 U24224 ( .C1(n21281), .C2(n21415), .A(n21280), .B(n21279), .ZN(
        P1_U3145) );
  AOI22_X1 U24225 ( .A1(n21313), .A2(n21410), .B1(n21312), .B2(n21408), .ZN(
        n21283) );
  AOI22_X1 U24226 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21421), .B1(
        n21292), .B2(n21314), .ZN(n21282) );
  OAI211_X1 U24227 ( .C1(n21317), .C2(n21415), .A(n21283), .B(n21282), .ZN(
        P1_U3146) );
  AOI22_X1 U24228 ( .A1(n21323), .A2(n21408), .B1(n21322), .B2(n21410), .ZN(
        n21285) );
  AOI22_X1 U24229 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21421), .B1(
        n21292), .B2(n21324), .ZN(n21284) );
  OAI211_X1 U24230 ( .C1(n21327), .C2(n21415), .A(n21285), .B(n21284), .ZN(
        P1_U3148) );
  AOI22_X1 U24231 ( .A1(n21329), .A2(n21408), .B1(n21328), .B2(n21410), .ZN(
        n21287) );
  AOI22_X1 U24232 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21421), .B1(
        n21292), .B2(n21330), .ZN(n21286) );
  OAI211_X1 U24233 ( .C1(n21333), .C2(n21415), .A(n21287), .B(n21286), .ZN(
        P1_U3149) );
  AOI22_X1 U24234 ( .A1(n21335), .A2(n21408), .B1(n21334), .B2(n21410), .ZN(
        n21289) );
  AOI22_X1 U24235 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21421), .B1(
        n21292), .B2(n21336), .ZN(n21288) );
  OAI211_X1 U24236 ( .C1(n21339), .C2(n21415), .A(n21289), .B(n21288), .ZN(
        P1_U3150) );
  AOI22_X1 U24237 ( .A1(n21341), .A2(n21408), .B1(n21340), .B2(n21410), .ZN(
        n21291) );
  AOI22_X1 U24238 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21421), .B1(
        n21292), .B2(n21342), .ZN(n21290) );
  OAI211_X1 U24239 ( .C1(n21345), .C2(n21415), .A(n21291), .B(n21290), .ZN(
        P1_U3151) );
  AOI22_X1 U24240 ( .A1(n21349), .A2(n21408), .B1(n21347), .B2(n21410), .ZN(
        n21294) );
  AOI22_X1 U24241 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21421), .B1(
        n21292), .B2(n21350), .ZN(n21293) );
  OAI211_X1 U24242 ( .C1(n21356), .C2(n21415), .A(n21294), .B(n21293), .ZN(
        P1_U3152) );
  NOR2_X1 U24243 ( .A1(n21296), .A2(n21295), .ZN(n21346) );
  AOI21_X1 U24244 ( .B1(n21298), .B2(n21297), .A(n21346), .ZN(n21304) );
  OAI22_X1 U24245 ( .A1(n21304), .A2(n21302), .B1(n21301), .B2(n12586), .ZN(
        n21348) );
  AOI22_X1 U24246 ( .A1(n21300), .A2(n21348), .B1(n21299), .B2(n21346), .ZN(
        n21310) );
  AOI22_X1 U24247 ( .A1(n21304), .A2(n21303), .B1(n21302), .B2(n21301), .ZN(
        n21305) );
  NAND2_X1 U24248 ( .A1(n21306), .A2(n21305), .ZN(n21352) );
  AOI22_X1 U24249 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21352), .B1(
        n21308), .B2(n21307), .ZN(n21309) );
  OAI211_X1 U24250 ( .C1(n21311), .C2(n21415), .A(n21310), .B(n21309), .ZN(
        P1_U3153) );
  AOI22_X1 U24251 ( .A1(n21313), .A2(n21346), .B1(n21312), .B2(n21348), .ZN(
        n21316) );
  AOI22_X1 U24252 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21314), .ZN(n21315) );
  OAI211_X1 U24253 ( .C1(n21317), .C2(n21355), .A(n21316), .B(n21315), .ZN(
        P1_U3154) );
  AOI22_X1 U24254 ( .A1(n21318), .A2(n21348), .B1(n21409), .B2(n21346), .ZN(
        n21321) );
  AOI22_X1 U24255 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21319), .ZN(n21320) );
  OAI211_X1 U24256 ( .C1(n21416), .C2(n21355), .A(n21321), .B(n21320), .ZN(
        P1_U3155) );
  AOI22_X1 U24257 ( .A1(n21323), .A2(n21348), .B1(n21322), .B2(n21346), .ZN(
        n21326) );
  AOI22_X1 U24258 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21324), .ZN(n21325) );
  OAI211_X1 U24259 ( .C1(n21327), .C2(n21355), .A(n21326), .B(n21325), .ZN(
        P1_U3156) );
  AOI22_X1 U24260 ( .A1(n21329), .A2(n21348), .B1(n21328), .B2(n21346), .ZN(
        n21332) );
  AOI22_X1 U24261 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21330), .ZN(n21331) );
  OAI211_X1 U24262 ( .C1(n21333), .C2(n21355), .A(n21332), .B(n21331), .ZN(
        P1_U3157) );
  AOI22_X1 U24263 ( .A1(n21335), .A2(n21348), .B1(n21334), .B2(n21346), .ZN(
        n21338) );
  AOI22_X1 U24264 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21336), .ZN(n21337) );
  OAI211_X1 U24265 ( .C1(n21339), .C2(n21355), .A(n21338), .B(n21337), .ZN(
        P1_U3158) );
  AOI22_X1 U24266 ( .A1(n21341), .A2(n21348), .B1(n21340), .B2(n21346), .ZN(
        n21344) );
  AOI22_X1 U24267 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21342), .ZN(n21343) );
  OAI211_X1 U24268 ( .C1(n21345), .C2(n21355), .A(n21344), .B(n21343), .ZN(
        P1_U3159) );
  AOI22_X1 U24269 ( .A1(n21349), .A2(n21348), .B1(n21347), .B2(n21346), .ZN(
        n21354) );
  AOI22_X1 U24270 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21352), .B1(
        n21351), .B2(n21350), .ZN(n21353) );
  OAI211_X1 U24271 ( .C1(n21356), .C2(n21355), .A(n21354), .B(n21353), .ZN(
        P1_U3160) );
  NOR2_X1 U24272 ( .A1(n10287), .A2(n21357), .ZN(n21360) );
  INV_X1 U24273 ( .A(n21358), .ZN(n21359) );
  OAI21_X1 U24274 ( .B1(n21360), .B2(n12586), .A(n21359), .ZN(P1_U3163) );
  AND2_X1 U24275 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21361), .ZN(
        P1_U3164) );
  AND2_X1 U24276 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21361), .ZN(
        P1_U3165) );
  AND2_X1 U24277 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21361), .ZN(
        P1_U3166) );
  AND2_X1 U24278 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21361), .ZN(
        P1_U3167) );
  AND2_X1 U24279 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21361), .ZN(
        P1_U3168) );
  AND2_X1 U24280 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21361), .ZN(
        P1_U3169) );
  AND2_X1 U24281 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21361), .ZN(
        P1_U3170) );
  AND2_X1 U24282 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21361), .ZN(
        P1_U3171) );
  AND2_X1 U24283 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21361), .ZN(
        P1_U3172) );
  AND2_X1 U24284 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21361), .ZN(
        P1_U3173) );
  AND2_X1 U24285 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21361), .ZN(
        P1_U3174) );
  AND2_X1 U24286 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21361), .ZN(
        P1_U3175) );
  AND2_X1 U24287 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21361), .ZN(
        P1_U3176) );
  AND2_X1 U24288 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21361), .ZN(
        P1_U3177) );
  AND2_X1 U24289 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21361), .ZN(
        P1_U3178) );
  AND2_X1 U24290 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21361), .ZN(
        P1_U3179) );
  AND2_X1 U24291 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21361), .ZN(
        P1_U3180) );
  AND2_X1 U24292 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21361), .ZN(
        P1_U3181) );
  AND2_X1 U24293 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21361), .ZN(
        P1_U3182) );
  AND2_X1 U24294 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21361), .ZN(
        P1_U3183) );
  AND2_X1 U24295 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21361), .ZN(
        P1_U3184) );
  AND2_X1 U24296 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21361), .ZN(
        P1_U3185) );
  AND2_X1 U24297 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21361), .ZN(P1_U3186) );
  AND2_X1 U24298 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21361), .ZN(P1_U3187) );
  AND2_X1 U24299 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21361), .ZN(P1_U3188) );
  AND2_X1 U24300 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21361), .ZN(P1_U3189) );
  AND2_X1 U24301 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21361), .ZN(P1_U3190) );
  AND2_X1 U24302 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21361), .ZN(P1_U3191) );
  INV_X1 U24303 ( .A(P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21540) );
  NOR2_X1 U24304 ( .A1(n21385), .A2(n21540), .ZN(P1_U3192) );
  AND2_X1 U24305 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21361), .ZN(P1_U3193) );
  OAI22_X1 U24306 ( .A1(n21364), .A2(n21363), .B1(n21362), .B2(
        P1_STATE_REG_0__SCAN_IN), .ZN(n21365) );
  NOR3_X1 U24307 ( .A1(n21366), .A2(n21365), .A3(n21515), .ZN(n21367) );
  OAI22_X1 U24308 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21368), .B1(n21396), 
        .B2(n21367), .ZN(P1_U3194) );
  AOI22_X1 U24309 ( .A1(n21374), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n13907), .ZN(n21369) );
  OAI21_X1 U24310 ( .B1(n13900), .B2(n21376), .A(n21369), .ZN(P1_U3205) );
  AOI22_X1 U24311 ( .A1(n21374), .A2(P1_REIP_REG_17__SCAN_IN), .B1(n21407), 
        .B2(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21370) );
  OAI21_X1 U24312 ( .B1(n21371), .B2(n21376), .A(n21370), .ZN(P1_U3213) );
  AOI22_X1 U24313 ( .A1(n21374), .A2(P1_REIP_REG_22__SCAN_IN), .B1(n21407), 
        .B2(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21372) );
  OAI21_X1 U24314 ( .B1(n21373), .B2(n21376), .A(n21372), .ZN(P1_U3218) );
  AOI22_X1 U24315 ( .A1(n21374), .A2(P1_REIP_REG_26__SCAN_IN), .B1(n21407), 
        .B2(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21375) );
  OAI21_X1 U24316 ( .B1(n21377), .B2(n21376), .A(n21375), .ZN(P1_U3222) );
  OAI22_X1 U24317 ( .A1(n21407), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21396), .ZN(n21378) );
  INV_X1 U24318 ( .A(n21378), .ZN(P1_U3458) );
  OAI22_X1 U24319 ( .A1(n21407), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21396), .ZN(n21379) );
  INV_X1 U24320 ( .A(n21379), .ZN(P1_U3459) );
  OAI22_X1 U24321 ( .A1(n13907), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21396), .ZN(n21380) );
  INV_X1 U24322 ( .A(n21380), .ZN(P1_U3460) );
  OAI22_X1 U24323 ( .A1(n13907), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21396), .ZN(n21381) );
  INV_X1 U24324 ( .A(n21381), .ZN(P1_U3461) );
  OAI21_X1 U24325 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21385), .A(n21383), 
        .ZN(n21382) );
  INV_X1 U24326 ( .A(n21382), .ZN(P1_U3464) );
  OAI21_X1 U24327 ( .B1(n21385), .B2(n21384), .A(n21383), .ZN(P1_U3465) );
  AOI21_X1 U24328 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21387) );
  AOI22_X1 U24329 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21387), .B2(n21386), .ZN(n21389) );
  INV_X1 U24330 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21388) );
  AOI22_X1 U24331 ( .A1(n21390), .A2(n21389), .B1(n21388), .B2(n21393), .ZN(
        P1_U3481) );
  INV_X1 U24332 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21394) );
  NOR2_X1 U24333 ( .A1(n21393), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21391) );
  AOI22_X1 U24334 ( .A1(n21394), .A2(n21393), .B1(n21392), .B2(n21391), .ZN(
        P1_U3482) );
  AOI22_X1 U24335 ( .A1(n21396), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21395), 
        .B2(n13907), .ZN(P1_U3483) );
  AOI21_X1 U24336 ( .B1(n21398), .B2(n21397), .A(n12586), .ZN(n21400) );
  AOI22_X1 U24337 ( .A1(n21401), .A2(n21400), .B1(n21399), .B2(n10287), .ZN(
        n21406) );
  AOI211_X1 U24338 ( .C1(n20784), .C2(n21404), .A(n21403), .B(n21402), .ZN(
        n21405) );
  MUX2_X1 U24339 ( .A(n21406), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21405), 
        .Z(P1_U3485) );
  MUX2_X1 U24340 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21407), .Z(P1_U3486) );
  INV_X1 U24341 ( .A(n21408), .ZN(n21413) );
  INV_X1 U24342 ( .A(n21409), .ZN(n21412) );
  INV_X1 U24343 ( .A(n21410), .ZN(n21411) );
  OAI22_X1 U24344 ( .A1(n21414), .A2(n21413), .B1(n21412), .B2(n21411), .ZN(
        n21420) );
  OAI22_X1 U24345 ( .A1(n21418), .A2(n21417), .B1(n21416), .B2(n21415), .ZN(
        n21419) );
  AOI211_X1 U24346 ( .C1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .C2(n21421), .A(
        n21420), .B(n21419), .ZN(n21574) );
  NAND4_X1 U24347 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(n15125), .A4(n21471), .ZN(n21431) );
  NOR3_X1 U24348 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_LWORD_REG_14__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(
        n21424) );
  NOR4_X1 U24349 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(
        P1_DATAO_REG_8__SCAN_IN), .A3(P2_DATAO_REG_12__SCAN_IN), .A4(n21462), 
        .ZN(n21423) );
  NOR4_X1 U24350 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(
        P2_DATAO_REG_5__SCAN_IN), .A3(n21480), .A4(n21483), .ZN(n21422) );
  NAND4_X1 U24351 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(n21424), .A3(n21423), 
        .A4(n21422), .ZN(n21430) );
  NAND4_X1 U24352 ( .A1(P3_CODEFETCH_REG_SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), 
        .A4(n21538), .ZN(n21429) );
  NOR4_X1 U24353 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n21553), .A3(
        n21509), .A4(n21515), .ZN(n21427) );
  NOR4_X1 U24354 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n21555), .A3(
        n21556), .A4(n21552), .ZN(n21426) );
  INV_X1 U24355 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n21543) );
  NOR3_X1 U24356 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(
        P3_REIP_REG_1__SCAN_IN), .A3(n21543), .ZN(n21425) );
  NAND4_X1 U24357 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21427), .A3(
        n21426), .A4(n21425), .ZN(n21428) );
  NOR4_X1 U24358 ( .A1(n21431), .A2(n21430), .A3(n21429), .A4(n21428), .ZN(
        n21572) );
  OR4_X1 U24359 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(P1_ADDRESS_REG_13__SCAN_IN), 
        .A3(n21432), .A4(n21514), .ZN(n21444) );
  NOR4_X1 U24360 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(
        P2_REIP_REG_26__SCAN_IN), .A3(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A4(
        n21485), .ZN(n21436) );
  NOR4_X1 U24361 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(
        BUF2_REG_29__SCAN_IN), .A3(P3_EAX_REG_21__SCAN_IN), .A4(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n21435) );
  NOR4_X1 U24362 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .A3(P2_DATAO_REG_22__SCAN_IN), .A4(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n21434) );
  NOR4_X1 U24363 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(
        P1_LWORD_REG_5__SCAN_IN), .A3(n18132), .A4(n21512), .ZN(n21433) );
  NAND4_X1 U24364 ( .A1(n21436), .A2(n21435), .A3(n21434), .A4(n21433), .ZN(
        n21443) );
  INV_X1 U24365 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n21452) );
  NAND4_X1 U24366 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_5__7__SCAN_IN), .A3(n21518), .A4(n21452), .ZN(n21442)
         );
  NAND3_X1 U24367 ( .A1(n12593), .A2(n21450), .A3(n21437), .ZN(n21438) );
  NOR3_X1 U24368 ( .A1(n21438), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A3(
        P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n21440) );
  INV_X1 U24369 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n21439) );
  NAND3_X1 U24370 ( .A1(n21440), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A3(
        n21439), .ZN(n21441) );
  NOR4_X1 U24371 ( .A1(n21444), .A2(n21443), .A3(n21442), .A4(n21441), .ZN(
        n21571) );
  AOI22_X1 U24372 ( .A1(n21447), .A2(keyinput57), .B1(keyinput13), .B2(n21446), 
        .ZN(n21445) );
  OAI221_X1 U24373 ( .B1(n21447), .B2(keyinput57), .C1(n21446), .C2(keyinput13), .A(n21445), .ZN(n21460) );
  INV_X1 U24374 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21449) );
  AOI22_X1 U24375 ( .A1(n21450), .A2(keyinput36), .B1(keyinput37), .B2(n21449), 
        .ZN(n21448) );
  OAI221_X1 U24376 ( .B1(n21450), .B2(keyinput36), .C1(n21449), .C2(keyinput37), .A(n21448), .ZN(n21459) );
  AOI22_X1 U24377 ( .A1(n21453), .A2(keyinput61), .B1(n21452), .B2(keyinput0), 
        .ZN(n21451) );
  OAI221_X1 U24378 ( .B1(n21453), .B2(keyinput61), .C1(n21452), .C2(keyinput0), 
        .A(n21451), .ZN(n21458) );
  XOR2_X1 U24379 ( .A(n21454), .B(keyinput17), .Z(n21456) );
  XNOR2_X1 U24380 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B(keyinput34), .ZN(
        n21455) );
  NAND2_X1 U24381 ( .A1(n21456), .A2(n21455), .ZN(n21457) );
  NOR4_X1 U24382 ( .A1(n21460), .A2(n21459), .A3(n21458), .A4(n21457), .ZN(
        n21507) );
  AOI22_X1 U24383 ( .A1(n21463), .A2(keyinput16), .B1(keyinput38), .B2(n21462), 
        .ZN(n21461) );
  OAI221_X1 U24384 ( .B1(n21463), .B2(keyinput16), .C1(n21462), .C2(keyinput38), .A(n21461), .ZN(n21475) );
  AOI22_X1 U24385 ( .A1(n21466), .A2(keyinput3), .B1(keyinput52), .B2(n21465), 
        .ZN(n21464) );
  OAI221_X1 U24386 ( .B1(n21466), .B2(keyinput3), .C1(n21465), .C2(keyinput52), 
        .A(n21464), .ZN(n21474) );
  INV_X1 U24387 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n21469) );
  AOI22_X1 U24388 ( .A1(n21469), .A2(keyinput14), .B1(keyinput23), .B2(n21468), 
        .ZN(n21467) );
  OAI221_X1 U24389 ( .B1(n21469), .B2(keyinput14), .C1(n21468), .C2(keyinput23), .A(n21467), .ZN(n21473) );
  AOI22_X1 U24390 ( .A1(n21471), .A2(keyinput39), .B1(keyinput30), .B2(n15125), 
        .ZN(n21470) );
  OAI221_X1 U24391 ( .B1(n21471), .B2(keyinput39), .C1(n15125), .C2(keyinput30), .A(n21470), .ZN(n21472) );
  NOR4_X1 U24392 ( .A1(n21475), .A2(n21474), .A3(n21473), .A4(n21472), .ZN(
        n21506) );
  INV_X1 U24393 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n21478) );
  AOI22_X1 U24394 ( .A1(n21478), .A2(keyinput54), .B1(keyinput2), .B2(n21477), 
        .ZN(n21476) );
  OAI221_X1 U24395 ( .B1(n21478), .B2(keyinput54), .C1(n21477), .C2(keyinput2), 
        .A(n21476), .ZN(n21489) );
  AOI22_X1 U24396 ( .A1(n21481), .A2(keyinput31), .B1(keyinput6), .B2(n21480), 
        .ZN(n21479) );
  OAI221_X1 U24397 ( .B1(n21481), .B2(keyinput31), .C1(n21480), .C2(keyinput6), 
        .A(n21479), .ZN(n21488) );
  AOI22_X1 U24398 ( .A1(n21483), .A2(keyinput46), .B1(n13463), .B2(keyinput29), 
        .ZN(n21482) );
  OAI221_X1 U24399 ( .B1(n21483), .B2(keyinput46), .C1(n13463), .C2(keyinput29), .A(n21482), .ZN(n21487) );
  AOI22_X1 U24400 ( .A1(n21485), .A2(keyinput28), .B1(n10624), .B2(keyinput50), 
        .ZN(n21484) );
  OAI221_X1 U24401 ( .B1(n21485), .B2(keyinput28), .C1(n10624), .C2(keyinput50), .A(n21484), .ZN(n21486) );
  NOR4_X1 U24402 ( .A1(n21489), .A2(n21488), .A3(n21487), .A4(n21486), .ZN(
        n21505) );
  INV_X1 U24403 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n21492) );
  AOI22_X1 U24404 ( .A1(n21492), .A2(keyinput47), .B1(keyinput22), .B2(n21491), 
        .ZN(n21490) );
  OAI221_X1 U24405 ( .B1(n21492), .B2(keyinput47), .C1(n21491), .C2(keyinput22), .A(n21490), .ZN(n21503) );
  AOI22_X1 U24406 ( .A1(n21495), .A2(keyinput10), .B1(keyinput33), .B2(n21494), 
        .ZN(n21493) );
  OAI221_X1 U24407 ( .B1(n21495), .B2(keyinput10), .C1(n21494), .C2(keyinput33), .A(n21493), .ZN(n21502) );
  XNOR2_X1 U24408 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B(keyinput49), .ZN(
        n21498) );
  XNOR2_X1 U24409 ( .A(P2_REIP_REG_26__SCAN_IN), .B(keyinput59), .ZN(n21497)
         );
  XNOR2_X1 U24410 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B(keyinput27), .ZN(
        n21496) );
  NAND3_X1 U24411 ( .A1(n21498), .A2(n21497), .A3(n21496), .ZN(n21501) );
  XNOR2_X1 U24412 ( .A(n21499), .B(keyinput1), .ZN(n21500) );
  NOR4_X1 U24413 ( .A1(n21503), .A2(n21502), .A3(n21501), .A4(n21500), .ZN(
        n21504) );
  NAND4_X1 U24414 ( .A1(n21507), .A2(n21506), .A3(n21505), .A4(n21504), .ZN(
        n21570) );
  INV_X1 U24415 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21510) );
  AOI22_X1 U24416 ( .A1(n21510), .A2(keyinput25), .B1(keyinput5), .B2(n21509), 
        .ZN(n21508) );
  OAI221_X1 U24417 ( .B1(n21510), .B2(keyinput25), .C1(n21509), .C2(keyinput5), 
        .A(n21508), .ZN(n21522) );
  AOI22_X1 U24418 ( .A1(n21512), .A2(keyinput8), .B1(n18132), .B2(keyinput62), 
        .ZN(n21511) );
  OAI221_X1 U24419 ( .B1(n21512), .B2(keyinput8), .C1(n18132), .C2(keyinput62), 
        .A(n21511), .ZN(n21521) );
  AOI22_X1 U24420 ( .A1(n21515), .A2(keyinput63), .B1(n21514), .B2(keyinput42), 
        .ZN(n21513) );
  OAI221_X1 U24421 ( .B1(n21515), .B2(keyinput63), .C1(n21514), .C2(keyinput42), .A(n21513), .ZN(n21520) );
  INV_X1 U24422 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n21517) );
  AOI22_X1 U24423 ( .A1(n21518), .A2(keyinput40), .B1(keyinput15), .B2(n21517), 
        .ZN(n21516) );
  OAI221_X1 U24424 ( .B1(n21518), .B2(keyinput40), .C1(n21517), .C2(keyinput15), .A(n21516), .ZN(n21519) );
  NOR4_X1 U24425 ( .A1(n21522), .A2(n21521), .A3(n21520), .A4(n21519), .ZN(
        n21568) );
  AOI22_X1 U24426 ( .A1(n13422), .A2(keyinput11), .B1(keyinput51), .B2(n21524), 
        .ZN(n21523) );
  OAI221_X1 U24427 ( .B1(n13422), .B2(keyinput11), .C1(n21524), .C2(keyinput51), .A(n21523), .ZN(n21535) );
  INV_X1 U24428 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n21526) );
  AOI22_X1 U24429 ( .A1(n21527), .A2(keyinput26), .B1(n21526), .B2(keyinput45), 
        .ZN(n21525) );
  OAI221_X1 U24430 ( .B1(n21527), .B2(keyinput26), .C1(n21526), .C2(keyinput45), .A(n21525), .ZN(n21534) );
  XOR2_X1 U24431 ( .A(n21528), .B(keyinput20), .Z(n21532) );
  XNOR2_X1 U24432 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B(keyinput60), .ZN(
        n21531) );
  XNOR2_X1 U24433 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(keyinput43), 
        .ZN(n21530) );
  XNOR2_X1 U24434 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B(keyinput58), .ZN(
        n21529) );
  NAND4_X1 U24435 ( .A1(n21532), .A2(n21531), .A3(n21530), .A4(n21529), .ZN(
        n21533) );
  NOR3_X1 U24436 ( .A1(n21535), .A2(n21534), .A3(n21533), .ZN(n21567) );
  AOI22_X1 U24437 ( .A1(n21538), .A2(keyinput32), .B1(n21537), .B2(keyinput18), 
        .ZN(n21536) );
  OAI221_X1 U24438 ( .B1(n21538), .B2(keyinput32), .C1(n21537), .C2(keyinput18), .A(n21536), .ZN(n21550) );
  AOI22_X1 U24439 ( .A1(n21541), .A2(keyinput21), .B1(keyinput7), .B2(n21540), 
        .ZN(n21539) );
  OAI221_X1 U24440 ( .B1(n21541), .B2(keyinput21), .C1(n21540), .C2(keyinput7), 
        .A(n21539), .ZN(n21549) );
  INV_X1 U24441 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21544) );
  AOI22_X1 U24442 ( .A1(n21544), .A2(keyinput35), .B1(n21543), .B2(keyinput53), 
        .ZN(n21542) );
  OAI221_X1 U24443 ( .B1(n21544), .B2(keyinput35), .C1(n21543), .C2(keyinput53), .A(n21542), .ZN(n21548) );
  XOR2_X1 U24444 ( .A(n18130), .B(keyinput12), .Z(n21546) );
  XNOR2_X1 U24445 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B(keyinput44), .ZN(
        n21545) );
  NAND2_X1 U24446 ( .A1(n21546), .A2(n21545), .ZN(n21547) );
  NOR4_X1 U24447 ( .A1(n21550), .A2(n21549), .A3(n21548), .A4(n21547), .ZN(
        n21566) );
  AOI22_X1 U24448 ( .A1(n21553), .A2(keyinput19), .B1(keyinput56), .B2(n21552), 
        .ZN(n21551) );
  OAI221_X1 U24449 ( .B1(n21553), .B2(keyinput19), .C1(n21552), .C2(keyinput56), .A(n21551), .ZN(n21564) );
  AOI22_X1 U24450 ( .A1(n21556), .A2(keyinput24), .B1(n21555), .B2(keyinput55), 
        .ZN(n21554) );
  OAI221_X1 U24451 ( .B1(n21556), .B2(keyinput24), .C1(n21555), .C2(keyinput55), .A(n21554), .ZN(n21563) );
  XNOR2_X1 U24452 ( .A(n21557), .B(keyinput48), .ZN(n21562) );
  XNOR2_X1 U24453 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B(keyinput4), .ZN(
        n21560) );
  XNOR2_X1 U24454 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B(keyinput41), .ZN(
        n21559) );
  XNOR2_X1 U24455 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput9), 
        .ZN(n21558) );
  NAND3_X1 U24456 ( .A1(n21560), .A2(n21559), .A3(n21558), .ZN(n21561) );
  NOR4_X1 U24457 ( .A1(n21564), .A2(n21563), .A3(n21562), .A4(n21561), .ZN(
        n21565) );
  NAND4_X1 U24458 ( .A1(n21568), .A2(n21567), .A3(n21566), .A4(n21565), .ZN(
        n21569) );
  AOI211_X1 U24459 ( .C1(n21572), .C2(n21571), .A(n21570), .B(n21569), .ZN(
        n21573) );
  XNOR2_X1 U24460 ( .A(n21574), .B(n21573), .ZN(P1_U3147) );
  AND2_X2 U11113 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14087) );
  AND2_X1 U15297 ( .A1(n14481), .A2(n11829), .ZN(n12712) );
  INV_X1 U11052 ( .A(n11255), .ZN(n13361) );
  AND2_X1 U14133 ( .A1(n13133), .A2(n10825), .ZN(n13120) );
  BUF_X2 U14467 ( .A(n11117), .Z(n13778) );
  BUF_X1 U11035 ( .A(n16910), .Z(n17843) );
  AND2_X2 U14121 ( .A1(n10690), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10881) );
  NOR2_X1 U13338 ( .A1(n16695), .A2(n16682), .ZN(n16665) );
  BUF_X2 U11042 ( .A(n11605), .Z(n13434) );
  CLKBUF_X1 U11045 ( .A(n12116), .Z(n12685) );
  CLKBUF_X1 U11064 ( .A(n11876), .Z(n9584) );
  CLKBUF_X1 U11065 ( .A(n9592), .Z(n9581) );
  CLKBUF_X2 U11085 ( .A(n11876), .Z(n9585) );
  CLKBUF_X1 U11093 ( .A(n11953), .Z(n12319) );
  NAND2_X1 U11105 ( .A1(n11853), .A2(n11852), .ZN(n11960) );
  CLKBUF_X1 U11117 ( .A(n11949), .Z(n13853) );
  INV_X1 U11450 ( .A(n14659), .ZN(n17252) );
  CLKBUF_X1 U11707 ( .A(n11970), .Z(n14208) );
  CLKBUF_X1 U11893 ( .A(n14507), .Z(n14508) );
  CLKBUF_X1 U12376 ( .A(n12502), .Z(n19815) );
  CLKBUF_X1 U12563 ( .A(n11255), .Z(n20022) );
  NOR2_X2 U12824 ( .A1(n20267), .A2(n20195), .ZN(n20073) );
endmodule

