

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3419, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207;

  NOR2_X1 U34520 ( .A1(n6340), .A2(n6339), .ZN(n6330) );
  CLKBUF_X2 U3454 ( .A(n3875), .Z(n4700) );
  CLKBUF_X2 U34560 ( .A(n3628), .Z(n4708) );
  CLKBUF_X2 U3457 ( .A(n3954), .Z(n3422) );
  CLKBUF_X2 U3458 ( .A(n3910), .Z(n3949) );
  CLKBUF_X2 U34590 ( .A(n3629), .Z(n4667) );
  BUF_X1 U34600 ( .A(n3836), .Z(n4928) );
  AND4_X1 U34620 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3483)
         );
  AND4_X1 U34630 ( .A1(n3478), .A2(n3477), .A3(n3476), .A4(n3475), .ZN(n3484)
         );
  AND4_X1 U34640 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3485)
         );
  AND4_X1 U34650 ( .A1(n3508), .A2(n3507), .A3(n3506), .A4(n3505), .ZN(n3514)
         );
  AND4_X1 U3466 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3513)
         );
  AND4_X1 U3467 ( .A1(n3604), .A2(n3603), .A3(n3602), .A4(n3601), .ZN(n3605)
         );
  AND2_X1 U34680 ( .A1(n4987), .A2(n4986), .ZN(n3432) );
  AND2_X1 U34700 ( .A1(n3453), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3426) );
  INV_X1 U34720 ( .A(n7205), .ZN(n3419) );
  INV_X2 U34740 ( .A(n7207), .ZN(n3421) );
  AND2_X1 U3475 ( .A1(n3454), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3460)
         );
  BUF_X1 U3476 ( .A(n3655), .Z(n3847) );
  AND4_X1 U3477 ( .A1(n3458), .A2(n3457), .A3(n3456), .A4(n3455), .ZN(n3466)
         );
  XNOR2_X1 U3478 ( .A(n4103), .B(n4090), .ZN(n4248) );
  NAND2_X1 U3479 ( .A1(n3727), .A2(n3812), .ZN(n3813) );
  NAND2_X1 U3480 ( .A1(n4727), .A2(n5946), .ZN(n3821) );
  AND2_X1 U3481 ( .A1(n3690), .A2(n4925), .ZN(n4727) );
  BUF_X1 U3482 ( .A(n5958), .Z(n5907) );
  NAND2_X1 U3483 ( .A1(n5573), .A2(n5572), .ZN(n5571) );
  OR2_X1 U3484 ( .A1(n4742), .A2(n4135), .ZN(n6348) );
  INV_X2 U3485 ( .A(n4116), .ZN(n6418) );
  INV_X1 U3487 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6691) );
  INV_X1 U3488 ( .A(n6950), .ZN(n6923) );
  NAND4_X2 U3489 ( .A1(n3486), .A2(n3485), .A3(n3484), .A4(n3483), .ZN(n3685)
         );
  XNOR2_X1 U3490 ( .A(n5907), .B(n4725), .ZN(n6328) );
  BUF_X1 U3491 ( .A(n4742), .Z(n6410) );
  NAND2_X2 U3492 ( .A1(n4878), .A2(n4877), .ZN(n4212) );
  AND2_X4 U3493 ( .A1(n5829), .A2(n5828), .ZN(n5868) );
  NAND2_X2 U3494 ( .A1(n3918), .A2(n3917), .ZN(n3920) );
  AND2_X2 U3497 ( .A1(n3893), .A2(n3892), .ZN(n3899) );
  NAND2_X1 U3498 ( .A1(n3689), .A2(n4762), .ZN(n3725) );
  INV_X2 U3499 ( .A(n3689), .ZN(n4921) );
  AOI21_X2 U3500 ( .B1(n5571), .B2(n4112), .A(n3442), .ZN(n5660) );
  NAND2_X4 U3502 ( .A1(n3969), .A2(n3968), .ZN(n4906) );
  NAND2_X4 U3504 ( .A1(n4905), .A2(n4006), .ZN(n5261) );
  OR2_X1 U3505 ( .A1(n5913), .A2(n6800), .ZN(n4171) );
  OAI22_X1 U3506 ( .A1(n4176), .A2(n4175), .B1(n6322), .B2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4177) );
  AOI21_X2 U3507 ( .B1(n6348), .B2(n4138), .A(n3443), .ZN(n6340) );
  AND2_X2 U3508 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  NOR2_X1 U3509 ( .A1(n6079), .A2(n6799), .ZN(n4190) );
  CLKBUF_X1 U3510 ( .A(n5571), .Z(n5607) );
  NAND2_X1 U3511 ( .A1(n4361), .A2(n4360), .ZN(n5702) );
  CLKBUF_X1 U3512 ( .A(n4747), .Z(n5831) );
  NAND2_X1 U3513 ( .A1(n4234), .A2(n4233), .ZN(n5092) );
  OAI21_X1 U3514 ( .B1(n4228), .B2(n4062), .A(n4061), .ZN(n4063) );
  OR2_X1 U3515 ( .A1(n4228), .A2(n4420), .ZN(n4234) );
  CLKBUF_X1 U3516 ( .A(n5711), .Z(n5726) );
  NAND2_X1 U3517 ( .A1(n3946), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5525)
         );
  CLKBUF_X1 U3518 ( .A(n5683), .Z(n5808) );
  NAND2_X1 U3520 ( .A1(n4004), .A2(n4003), .ZN(n4954) );
  NAND2_X1 U3521 ( .A1(n4798), .A2(n4205), .ZN(n4815) );
  NOR2_X2 U3522 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4920), .ZN(n5161) );
  NAND2_X2 U3523 ( .A1(n6636), .A2(n5697), .ZN(n6283) );
  NAND2_X1 U3524 ( .A1(n3984), .A2(n3983), .ZN(n5017) );
  INV_X1 U3525 ( .A(n4909), .ZN(n5051) );
  NAND2_X1 U3526 ( .A1(n3737), .A2(n3446), .ZN(n5040) );
  CLKBUF_X1 U3527 ( .A(n3861), .Z(n5019) );
  CLKBUF_X1 U3528 ( .A(n3701), .Z(n5948) );
  OR2_X1 U3529 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3724)
         );
  NAND2_X2 U3530 ( .A1(n3806), .A2(n3434), .ZN(n4178) );
  NAND2_X1 U3531 ( .A1(n3694), .A2(n3693), .ZN(n3833) );
  INV_X2 U3532 ( .A(n3694), .ZN(n3435) );
  INV_X1 U3533 ( .A(n4089), .ZN(n4002) );
  NAND2_X1 U3534 ( .A1(n3518), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4089) );
  BUF_X2 U3535 ( .A(n3831), .Z(n6692) );
  NAND2_X1 U3536 ( .A1(n3659), .A2(n3830), .ZN(n3854) );
  AND2_X1 U3538 ( .A1(n3650), .A2(n5697), .ZN(n3839) );
  OR2_X1 U3539 ( .A1(n3933), .A2(n3932), .ZN(n3971) );
  INV_X2 U3540 ( .A(n3685), .ZN(n4935) );
  INV_X2 U3541 ( .A(n4193), .ZN(n3675) );
  AND4_X1 U3542 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3586)
         );
  AND4_X1 U3543 ( .A1(n3572), .A2(n3571), .A3(n3570), .A4(n3569), .ZN(n3588)
         );
  AND4_X1 U3544 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3607)
         );
  AND4_X1 U3545 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3608)
         );
  AND4_X1 U3546 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3515)
         );
  AND4_X1 U3547 ( .A1(n3464), .A2(n3463), .A3(n3462), .A4(n3461), .ZN(n3465)
         );
  BUF_X2 U3548 ( .A(n3874), .Z(n4706) );
  BUF_X2 U3549 ( .A(n3947), .Z(n4600) );
  BUF_X2 U3550 ( .A(n3955), .Z(n4699) );
  AND2_X2 U3551 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5533), .ZN(n6696) );
  AND2_X2 U3552 ( .A1(n5011), .A2(n4986), .ZN(n3609) );
  NAND2_X1 U3553 ( .A1(n4370), .A2(n4369), .ZN(n3423) );
  AND2_X2 U3554 ( .A1(n3939), .A2(n3940), .ZN(n3919) );
  XNOR2_X2 U3555 ( .A(n3893), .B(n3892), .ZN(n4909) );
  NAND2_X1 U3556 ( .A1(n3873), .A2(n3897), .ZN(n3424) );
  NAND2_X1 U3558 ( .A1(n3873), .A2(n3897), .ZN(n3898) );
  NAND2_X1 U3559 ( .A1(n5525), .A2(n5528), .ZN(n3427) );
  NAND2_X1 U3560 ( .A1(n5775), .A2(n3431), .ZN(n3428) );
  AND2_X1 U3561 ( .A1(n3428), .A2(n3429), .ZN(n5819) );
  OR2_X1 U3562 ( .A1(n3430), .A2(n4122), .ZN(n3429) );
  INV_X1 U3563 ( .A(n5820), .ZN(n3430) );
  AND2_X1 U3564 ( .A1(n5774), .A2(n5820), .ZN(n3431) );
  NAND2_X1 U3565 ( .A1(n6006), .A2(n5920), .ZN(n5919) );
  AOI21_X2 U3567 ( .B1(n4248), .B2(n4304), .A(n4247), .ZN(n5443) );
  OR2_X2 U3568 ( .A1(n4797), .A2(n4204), .ZN(n4798) );
  NAND2_X1 U3569 ( .A1(n4005), .A2(n4954), .ZN(n4040) );
  NOR2_X4 U3570 ( .A1(n5760), .A2(n5759), .ZN(n5829) );
  NAND2_X2 U3571 ( .A1(n4876), .A2(n5435), .ZN(n5437) );
  NAND2_X2 U3572 ( .A1(n4212), .A2(n4211), .ZN(n4876) );
  NOR2_X4 U3573 ( .A1(n5560), .A2(n5561), .ZN(n5591) );
  INV_X1 U3574 ( .A(n3694), .ZN(n3434) );
  AND2_X1 U3575 ( .A1(n4762), .A2(n3438), .ZN(n3727) );
  NOR2_X2 U3576 ( .A1(n6032), .A2(n6019), .ZN(n6004) );
  XNOR2_X2 U3577 ( .A(n3941), .B(n3940), .ZN(n4194) );
  NAND4_X1 U3578 ( .A1(n3486), .A2(n3485), .A3(n3484), .A4(n3483), .ZN(n3437)
         );
  NAND4_X1 U3579 ( .A1(n3486), .A2(n3485), .A3(n3484), .A4(n3483), .ZN(n3438)
         );
  NAND4_X1 U3580 ( .A1(n3486), .A2(n3485), .A3(n3484), .A4(n3483), .ZN(n3439)
         );
  NAND4_X1 U3581 ( .A1(n3486), .A2(n3485), .A3(n3484), .A4(n3483), .ZN(n3440)
         );
  XNOR2_X2 U3582 ( .A(n5702), .B(n4362), .ZN(n5586) );
  CLKBUF_X1 U3583 ( .A(n3927), .Z(n4707) );
  XNOR2_X1 U3584 ( .A(n4040), .B(n4038), .ZN(n4227) );
  CLKBUF_X1 U3585 ( .A(n3859), .Z(n3677) );
  AND2_X1 U3586 ( .A1(n7011), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3864) );
  NOR2_X1 U3587 ( .A1(n5927), .A2(n3706), .ZN(n5942) );
  NAND2_X1 U3588 ( .A1(n4103), .A2(n4102), .ZN(n4140) );
  CLKBUF_X1 U3589 ( .A(n3927), .Z(n4619) );
  OR2_X1 U3590 ( .A1(n3916), .A2(n3915), .ZN(n4009) );
  NAND2_X1 U3591 ( .A1(n4002), .A2(n3847), .ZN(n3843) );
  NAND2_X1 U3592 ( .A1(n4193), .A2(n3657), .ZN(n3655) );
  NAND2_X1 U3593 ( .A1(n4079), .A2(n4078), .ZN(n4103) );
  NOR2_X2 U3594 ( .A1(n5866), .A2(n5883), .ZN(n5881) );
  NAND2_X1 U3595 ( .A1(n4370), .A2(n4369), .ZN(n5708) );
  INV_X1 U3596 ( .A(n5535), .ZN(n4721) );
  CLKBUF_X1 U3597 ( .A(n4213), .Z(n4683) );
  INV_X1 U3598 ( .A(n4420), .ZN(n4304) );
  OR2_X1 U3599 ( .A1(n5874), .A2(n4130), .ZN(n4131) );
  OR2_X1 U3600 ( .A1(n4129), .A2(n4128), .ZN(n4130) );
  NOR2_X1 U3601 ( .A1(n5040), .A2(n5041), .ZN(n5039) );
  NOR2_X1 U3602 ( .A1(n3675), .A2(n3664), .ZN(n3620) );
  XNOR2_X1 U3603 ( .A(n5017), .B(n5015), .ZN(n4908) );
  CLKBUF_X1 U3604 ( .A(n3900), .Z(n3985) );
  AND2_X1 U3605 ( .A1(n3836), .A2(n3440), .ZN(n3831) );
  OR2_X1 U3606 ( .A1(n6694), .A2(n5537), .ZN(n6850) );
  AND2_X1 U3607 ( .A1(n6850), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5971) );
  INV_X1 U3608 ( .A(n4568), .ZN(n5955) );
  NAND2_X1 U3609 ( .A1(n4592), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4636)
         );
  NOR2_X1 U3610 ( .A1(n4390), .A2(n4401), .ZN(n4387) );
  NAND2_X1 U3611 ( .A1(n4387), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4458)
         );
  INV_X1 U3612 ( .A(n4235), .ZN(n4236) );
  NAND2_X1 U3613 ( .A1(n4236), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4242)
         );
  NOR2_X1 U3614 ( .A1(n4223), .A2(n6832), .ZN(n4229) );
  NAND2_X1 U3615 ( .A1(n6330), .A2(n3449), .ZN(n4176) );
  OR2_X1 U3616 ( .A1(n4888), .A2(n4887), .ZN(n6749) );
  NAND2_X1 U3617 ( .A1(n3682), .A2(n3681), .ZN(n4148) );
  OR3_X1 U3618 ( .A1(n4784), .A2(n4900), .A3(n4783), .ZN(n6968) );
  INV_X1 U3619 ( .A(n3556), .ZN(n3566) );
  AND2_X1 U3620 ( .A1(n3517), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4087) );
  NAND2_X1 U3621 ( .A1(n4761), .A2(n4757), .ZN(n6694) );
  OR2_X1 U3622 ( .A1(n4734), .A2(n4162), .ZN(n6081) );
  NAND2_X1 U3623 ( .A1(n4730), .A2(n4729), .ZN(n6636) );
  OR2_X1 U3624 ( .A1(n7017), .A2(n4726), .ZN(n4730) );
  INV_X1 U3625 ( .A(n6287), .ZN(n7062) );
  AND2_X1 U3626 ( .A1(n6287), .A2(n5698), .ZN(n7059) );
  NAND2_X1 U3627 ( .A1(n4902), .A2(n4901), .ZN(n6287) );
  AOI21_X1 U3628 ( .B1(n4900), .B2(n7004), .A(n4899), .ZN(n4901) );
  INV_X1 U3629 ( .A(n5957), .ZN(n4725) );
  AND2_X1 U3630 ( .A1(n3839), .A2(n3838), .ZN(n3840) );
  AOI21_X1 U3631 ( .B1(n3860), .B2(n3625), .A(n3837), .ZN(n3838) );
  INV_X1 U3632 ( .A(n5679), .ZN(n4368) );
  CLKBUF_X1 U3633 ( .A(n3635), .Z(n4666) );
  OR2_X1 U3634 ( .A1(n4050), .A2(n4049), .ZN(n4059) );
  OR2_X1 U3635 ( .A1(n4028), .A2(n4027), .ZN(n4056) );
  CLKBUF_X1 U3636 ( .A(n3921), .Z(n4650) );
  NAND2_X1 U3637 ( .A1(n3890), .A2(n3889), .ZN(n3939) );
  NAND2_X1 U3638 ( .A1(n3888), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3889) );
  MUX2_X1 U3639 ( .A(n3894), .B(n4909), .S(n7020), .Z(n3896) );
  OR2_X1 U3640 ( .A1(n4001), .A2(n4000), .ZN(n4031) );
  AOI21_X1 U3642 ( .B1(n4644), .B2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n3636), 
        .ZN(n3642) );
  AND2_X1 U3643 ( .A1(n3635), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3636) );
  INV_X1 U3644 ( .A(n4087), .ZN(n3537) );
  AND2_X1 U3645 ( .A1(n6067), .A2(n3801), .ZN(n6041) );
  INV_X1 U3646 ( .A(n4128), .ZN(n4124) );
  AND4_X2 U3647 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(n4193)
         );
  AOI21_X1 U3648 ( .B1(n7015), .B2(n4915), .A(n5934), .ZN(n4920) );
  AND2_X2 U3649 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5011) );
  OR2_X1 U3650 ( .A1(n5946), .A2(n3522), .ZN(n3546) );
  NOR2_X1 U3651 ( .A1(n3537), .A2(n3667), .ZN(n3545) );
  INV_X1 U3652 ( .A(n3560), .ZN(n3554) );
  OR2_X1 U3653 ( .A1(n4734), .A2(n3435), .ZN(n4182) );
  AND2_X2 U3654 ( .A1(n4731), .A2(n4161), .ZN(n4734) );
  AND2_X1 U3655 ( .A1(n4502), .A2(n4501), .ZN(n5867) );
  OR2_X1 U3656 ( .A1(n6951), .A2(n5535), .ZN(n4501) );
  AND2_X1 U3657 ( .A1(n5997), .A2(n4721), .ZN(n4662) );
  AND2_X1 U3658 ( .A1(n4822), .A2(n4821), .ZN(n6524) );
  INV_X1 U3659 ( .A(n4902), .ZN(n4858) );
  NOR2_X1 U3660 ( .A1(n4761), .A2(READY_N), .ZN(n4763) );
  AND2_X1 U3661 ( .A1(n6324), .A2(n4721), .ZN(n4722) );
  NOR2_X1 U3662 ( .A1(n4689), .A2(n4688), .ZN(n4690) );
  OR2_X1 U3663 ( .A1(n5987), .A2(n5535), .ZN(n4693) );
  OR2_X1 U3664 ( .A1(n4637), .A2(n6010), .ZN(n4689) );
  INV_X1 U3665 ( .A(n6007), .ZN(n4641) );
  INV_X1 U3666 ( .A(n4590), .ZN(n4591) );
  AND2_X1 U3667 ( .A1(n4597), .A2(n4596), .ZN(n6033) );
  OR2_X1 U3668 ( .A1(n6353), .A2(n5535), .ZN(n4596) );
  AND2_X1 U3669 ( .A1(n4549), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4550)
         );
  INV_X1 U3670 ( .A(n4548), .ZN(n4549) );
  NAND2_X1 U3671 ( .A1(n4550), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4590)
         );
  INV_X1 U3672 ( .A(n6063), .ZN(n4555) );
  AND2_X1 U3673 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n4459), .ZN(n4460)
         );
  INV_X1 U3674 ( .A(n4458), .ZN(n4459) );
  AND2_X1 U3675 ( .A1(n4389), .A2(n4388), .ZN(n5709) );
  NAND2_X1 U3676 ( .A1(n4406), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4390)
         );
  OR2_X1 U3677 ( .A1(n5784), .A2(n5785), .ZN(n5851) );
  NAND2_X1 U3678 ( .A1(n4337), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4363)
         );
  INV_X1 U3679 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4364) );
  NOR2_X1 U3680 ( .A1(n4308), .A2(n4307), .ZN(n4337) );
  NAND2_X1 U3681 ( .A1(n4292), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4308)
         );
  INV_X1 U3682 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4307) );
  AND2_X1 U3683 ( .A1(n4352), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4292)
         );
  AND2_X1 U3684 ( .A1(n4275), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4352)
         );
  AND2_X1 U3685 ( .A1(n5591), .A2(n5590), .ZN(n5678) );
  AND3_X1 U3686 ( .A1(n4263), .A2(n4262), .A3(n4261), .ZN(n5561) );
  NOR2_X1 U3687 ( .A1(n4242), .A2(n4241), .ZN(n4275) );
  INV_X1 U3688 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4241) );
  AOI21_X1 U3689 ( .B1(n4240), .B2(n4304), .A(n4239), .ZN(n5336) );
  NAND2_X1 U3690 ( .A1(n4229), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4235)
         );
  AOI21_X1 U3691 ( .B1(n4227), .B2(n4304), .A(n4226), .ZN(n5029) );
  INV_X1 U3692 ( .A(n4214), .ZN(n4215) );
  NAND2_X1 U3693 ( .A1(n4215), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4223)
         );
  NAND2_X1 U3694 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4214) );
  OAI21_X1 U3695 ( .B1(n5261), .B2(n4062), .A(n3937), .ZN(n3938) );
  CLKBUF_X1 U3696 ( .A(n6041), .Z(n6052) );
  NOR2_X2 U3697 ( .A1(n6065), .A2(n6064), .ZN(n6067) );
  OR2_X1 U3698 ( .A1(n5711), .A2(n5725), .ZN(n5764) );
  NOR2_X2 U3699 ( .A1(n5764), .A2(n5763), .ZN(n5833) );
  CLKBUF_X1 U3700 ( .A(n6416), .Z(n6417) );
  NAND2_X1 U3701 ( .A1(n4121), .A2(n4120), .ZN(n5775) );
  INV_X1 U3702 ( .A(n4140), .ZN(n4116) );
  NAND2_X1 U3703 ( .A1(n6628), .A2(n3751), .ZN(n5593) );
  AND2_X1 U3704 ( .A1(n3741), .A2(n3740), .ZN(n5041) );
  INV_X1 U3705 ( .A(n4194), .ZN(n5299) );
  AND2_X2 U3706 ( .A1(n3452), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4785)
         );
  INV_X1 U3707 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3452) );
  CLKBUF_X1 U3708 ( .A(n4910), .Z(n4911) );
  OR2_X1 U3709 ( .A1(n3705), .A2(n3704), .ZN(n5927) );
  BUF_X1 U3710 ( .A(n4908), .Z(n7083) );
  NAND2_X1 U3711 ( .A1(n3991), .A2(n3990), .ZN(n5015) );
  CLKBUF_X1 U3712 ( .A(n4905), .Z(n5298) );
  INV_X1 U3713 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7103) );
  BUF_X1 U3714 ( .A(n3656), .Z(n4978) );
  CLKBUF_X1 U3715 ( .A(n4193), .Z(n4938) );
  OR2_X1 U3716 ( .A1(n4920), .A2(n7012), .ZN(n4979) );
  NAND2_X1 U3717 ( .A1(n6691), .A2(n7028), .ZN(n5535) );
  AND2_X1 U3718 ( .A1(n3864), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U3719 ( .A1(n5971), .A2(n5543), .ZN(n6884) );
  AND2_X1 U3720 ( .A1(n6850), .A2(n5540), .ZN(n6947) );
  AND2_X1 U3721 ( .A1(n6316), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5554) );
  INV_X1 U3722 ( .A(n6925), .ZN(n6910) );
  INV_X1 U3723 ( .A(n6884), .ZN(n6862) );
  INV_X1 U3724 ( .A(n6943), .ZN(n6907) );
  INV_X1 U3725 ( .A(n6931), .ZN(n6946) );
  NAND2_X1 U3726 ( .A1(n6287), .A2(n3659), .ZN(n5816) );
  NOR2_X1 U3727 ( .A1(n6696), .A2(n6524), .ZN(n6534) );
  NAND2_X1 U3728 ( .A1(n4763), .A2(n4762), .ZN(n4902) );
  XNOR2_X1 U3729 ( .A(n5539), .B(n5974), .ZN(n6316) );
  OR2_X1 U3730 ( .A1(n5538), .A2(n6326), .ZN(n5539) );
  XNOR2_X1 U3731 ( .A(n4142), .B(n3448), .ZN(n5926) );
  NAND2_X1 U3732 ( .A1(n4176), .A2(n4141), .ZN(n4142) );
  INV_X1 U3733 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6832) );
  OR2_X1 U3734 ( .A1(n6669), .A2(n5519), .ZN(n6676) );
  INV_X1 U3735 ( .A(n6676), .ZN(n6665) );
  INV_X1 U3736 ( .A(n6952), .ZN(n6671) );
  OR2_X1 U3737 ( .A1(n6489), .A2(n3721), .ZN(n6466) );
  CLKBUF_X1 U3738 ( .A(n5729), .Z(n5730) );
  OR2_X1 U3739 ( .A1(n5747), .A2(n6749), .ZN(n6794) );
  INV_X1 U3740 ( .A(n6800), .ZN(n6821) );
  CLKBUF_X1 U3741 ( .A(n4909), .Z(n5929) );
  INV_X1 U3742 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7099) );
  CLKBUF_X1 U3743 ( .A(n4788), .Z(n4789) );
  INV_X1 U3744 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6978) );
  INV_X1 U3746 ( .A(n6955), .ZN(n5934) );
  INV_X1 U3747 ( .A(n5447), .ZN(n5510) );
  INV_X1 U3748 ( .A(n5158), .ZN(n5191) );
  NOR2_X1 U3749 ( .A1(n7078), .A2(n4906), .ZN(n7182) );
  INV_X1 U3750 ( .A(n5225), .ZN(n5255) );
  INV_X1 U3751 ( .A(n7120), .ZN(n5462) );
  INV_X1 U3752 ( .A(n7130), .ZN(n5490) );
  INV_X1 U3753 ( .A(n7140), .ZN(n5469) );
  INV_X1 U3754 ( .A(n7150), .ZN(n5476) );
  INV_X1 U3755 ( .A(n7160), .ZN(n5483) );
  INV_X1 U3756 ( .A(n7170), .ZN(n5497) );
  INV_X1 U3757 ( .A(n7180), .ZN(n5515) );
  INV_X1 U3758 ( .A(n7203), .ZN(n5504) );
  NOR2_X1 U3759 ( .A1(n5058), .A2(n4906), .ZN(n5127) );
  NAND2_X1 U3760 ( .A1(n3568), .A2(n3567), .ZN(n7017) );
  INV_X1 U3761 ( .A(n7016), .ZN(n7014) );
  NAND2_X1 U3762 ( .A1(n6328), .A2(n6634), .ZN(n4741) );
  NOR2_X1 U3763 ( .A1(n6636), .A2(n5980), .ZN(n4737) );
  INV_X1 U3764 ( .A(n6328), .ZN(n6293) );
  NOR2_X1 U3765 ( .A1(n4169), .A2(n4168), .ZN(n4170) );
  AND2_X1 U3766 ( .A1(n6428), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4168)
         );
  NAND2_X1 U3767 ( .A1(n5708), .A2(n4422), .ZN(n5696) );
  XOR2_X1 U3768 ( .A(n5960), .B(n5959), .Z(n3441) );
  NOR2_X1 U3769 ( .A1(n4111), .A2(n5609), .ZN(n3442) );
  INV_X1 U3770 ( .A(n4762), .ZN(n3836) );
  AND2_X1 U3771 ( .A1(n3834), .A2(n3833), .ZN(n3851) );
  NOR2_X1 U3772 ( .A1(n4137), .A2(n6350), .ZN(n3443) );
  NOR2_X1 U3773 ( .A1(n5806), .A2(n5626), .ZN(n3444) );
  AND2_X1 U3774 ( .A1(n5197), .A2(n7066), .ZN(n5199) );
  AND4_X1 U3775 ( .A1(n3857), .A2(n3851), .A3(n3856), .A4(n3855), .ZN(n3445)
         );
  INV_X1 U3776 ( .A(n6005), .ZN(n6018) );
  AND2_X2 U3777 ( .A1(n3460), .A2(n4986), .ZN(n3922) );
  AND2_X1 U3778 ( .A1(n4893), .A2(n5669), .ZN(n3446) );
  AND2_X1 U3779 ( .A1(n3632), .A2(n3631), .ZN(n3447) );
  XOR2_X1 U3780 ( .A(n6418), .B(n4152), .Z(n3448) );
  OR2_X1 U3781 ( .A1(n4116), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3449)
         );
  INV_X1 U3782 ( .A(n6427), .ZN(n4739) );
  NAND2_X1 U3783 ( .A1(n4762), .A2(n3657), .ZN(n4062) );
  INV_X1 U3784 ( .A(n4062), .ZN(n4100) );
  OR2_X1 U3785 ( .A1(n5697), .A2(n6691), .ZN(n4213) );
  AND2_X1 U3786 ( .A1(n4441), .A2(n4440), .ZN(n3450) );
  NAND2_X1 U3787 ( .A1(n3904), .A2(n3903), .ZN(n3983) );
  BUF_X1 U3788 ( .A(n3623), .Z(n4143) );
  INV_X1 U3789 ( .A(n4143), .ZN(n3693) );
  INV_X1 U3790 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7020) );
  NAND2_X1 U3791 ( .A1(n6636), .A2(n6288), .ZN(n6629) );
  INV_X1 U3792 ( .A(n6629), .ZN(n4738) );
  INV_X1 U3793 ( .A(n3657), .ZN(n3625) );
  OR2_X1 U3794 ( .A1(n3887), .A2(n3886), .ZN(n3942) );
  INV_X1 U3795 ( .A(n3725), .ZN(n3694) );
  BUF_X1 U3797 ( .A(n4644), .Z(n4601) );
  INV_X1 U3799 ( .A(n4038), .ZN(n4039) );
  AND2_X1 U3800 ( .A1(n3866), .A2(n3865), .ZN(n3870) );
  OR2_X1 U3801 ( .A1(n3867), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3868)
         );
  INV_X1 U3802 ( .A(n3517), .ZN(n3518) );
  INV_X1 U3803 ( .A(n3521), .ZN(n3533) );
  OR2_X1 U3804 ( .A1(n4636), .A2(n6024), .ZN(n4637) );
  OR2_X1 U3805 ( .A1(n4075), .A2(n4074), .ZN(n4092) );
  AND2_X1 U3806 ( .A1(n4077), .A2(n4076), .ZN(n4080) );
  AND2_X1 U3807 ( .A1(n6418), .A2(n6814), .ZN(n4128) );
  OR2_X1 U3808 ( .A1(n4140), .A2(n6788), .ZN(n4110) );
  CLKBUF_X1 U3809 ( .A(n3689), .Z(n3934) );
  OR2_X1 U3810 ( .A1(n4089), .A2(n4062), .ZN(n3556) );
  OR2_X1 U3811 ( .A1(n3561), .A2(n6983), .ZN(n3560) );
  AND2_X1 U3812 ( .A1(n5617), .A2(n4325), .ZN(n4357) );
  AND4_X1 U3813 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3516)
         );
  AND2_X2 U3814 ( .A1(n3426), .A2(n4785), .ZN(n3947) );
  AND2_X1 U3815 ( .A1(n4591), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4592)
         );
  AND2_X1 U3816 ( .A1(n5709), .A2(n5707), .ZN(n4422) );
  AND3_X1 U3817 ( .A1(n4101), .A2(n4100), .A3(n4104), .ZN(n4102) );
  AND2_X1 U3818 ( .A1(n3747), .A2(n3746), .ZN(n6626) );
  OR2_X1 U3819 ( .A1(n4054), .A2(n4053), .ZN(n4055) );
  INV_X1 U3820 ( .A(n4006), .ZN(n4005) );
  NAND2_X1 U3821 ( .A1(n4908), .A2(n7020), .ZN(n4004) );
  AND4_X1 U3822 ( .A1(n3600), .A2(n3599), .A3(n3598), .A4(n3597), .ZN(n3606)
         );
  INV_X1 U3823 ( .A(n3812), .ZN(n4181) );
  NAND2_X1 U3824 ( .A1(n5930), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4686) );
  OR2_X1 U3825 ( .A1(n4904), .A2(n4420), .ZN(n4220) );
  OR2_X1 U3827 ( .A1(n6376), .A2(n5535), .ZN(n4553) );
  NOR2_X1 U3828 ( .A1(n4363), .A2(n4364), .ZN(n4386) );
  INV_X1 U3829 ( .A(n4213), .ZN(n5956) );
  INV_X1 U3830 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6362) );
  AND2_X1 U3831 ( .A1(n3763), .A2(n3762), .ZN(n5805) );
  AND2_X1 U3832 ( .A1(n5625), .A2(n5624), .ZN(n5806) );
  NAND2_X1 U3833 ( .A1(n4016), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6646)
         );
  NAND2_X1 U3834 ( .A1(n3724), .A2(n3723), .ZN(n3728) );
  AND2_X1 U3835 ( .A1(n3648), .A2(n3647), .ZN(n3701) );
  NAND2_X1 U3836 ( .A1(n3701), .A2(n4928), .ZN(n3861) );
  INV_X1 U3837 ( .A(n5261), .ZN(n5263) );
  NAND2_X1 U3838 ( .A1(n5051), .A2(n7020), .ZN(n3969) );
  NAND2_X1 U3839 ( .A1(n3566), .A2(n3669), .ZN(n3567) );
  AND2_X1 U3840 ( .A1(n3859), .A2(n3685), .ZN(n4755) );
  INV_X1 U3841 ( .A(n3436), .ZN(n5552) );
  NOR2_X1 U3842 ( .A1(n4496), .A2(n6400), .ZN(n4497) );
  AND2_X1 U3843 ( .A1(n4386), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4406)
         );
  INV_X1 U3844 ( .A(n6939), .ZN(n6927) );
  AND2_X1 U3845 ( .A1(n6418), .A2(n4152), .ZN(n4155) );
  NAND2_X1 U3846 ( .A1(n4460), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4496)
         );
  OR4_X1 U3847 ( .A1(n6340), .A2(n4116), .A3(n6320), .A4(n6451), .ZN(n6321) );
  OR2_X1 U3848 ( .A1(n6382), .A2(n6360), .ZN(n6364) );
  NAND2_X1 U3849 ( .A1(n5819), .A2(n4123), .ZN(n5874) );
  NOR2_X2 U3850 ( .A1(n5603), .A2(n5604), .ZN(n5625) );
  NAND2_X1 U3851 ( .A1(n3858), .A2(n3445), .ZN(n3892) );
  AND2_X2 U3852 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4986) );
  INV_X1 U3853 ( .A(n5127), .ZN(n5293) );
  NAND2_X1 U3854 ( .A1(n4040), .A2(n4007), .ZN(n4904) );
  OR3_X1 U3855 ( .A1(n5300), .A2(n5263), .A3(n5262), .ZN(n5270) );
  INV_X1 U3856 ( .A(n5456), .ZN(n7084) );
  OR3_X1 U3857 ( .A1(n5300), .A2(n5299), .A3(n5298), .ZN(n7078) );
  INV_X1 U3858 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U3859 ( .A1(n4497), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4548)
         );
  AND2_X1 U3860 ( .A1(n6850), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6939) );
  AND2_X1 U3861 ( .A1(n5971), .A2(n5546), .ZN(n6943) );
  AND2_X1 U3862 ( .A1(n5039), .A2(n5438), .ZN(n6628) );
  INV_X1 U3863 ( .A(n6636), .ZN(n6281) );
  AOI21_X1 U3864 ( .B1(n4176), .B2(n4172), .A(n4155), .ZN(n4157) );
  OR2_X1 U3865 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  NAND2_X1 U3866 ( .A1(n7017), .A2(n7004), .ZN(n4818) );
  NAND2_X1 U3867 ( .A1(n6364), .A2(n6363), .ZN(n6365) );
  OAI21_X1 U3868 ( .B1(n6824), .B2(n4129), .A(n3708), .ZN(n6506) );
  AND2_X1 U3869 ( .A1(n6751), .A2(n3710), .ZN(n5809) );
  OR2_X1 U3870 ( .A1(n5743), .A2(n6748), .ZN(n6796) );
  CLKBUF_X1 U3871 ( .A(n4986), .Z(n5902) );
  NAND2_X1 U3872 ( .A1(n7017), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6955) );
  INV_X1 U3873 ( .A(n7108), .ZN(n7198) );
  OAI211_X1 U3874 ( .C1(n5453), .C2(n5458), .A(n5452), .B(n5451), .ZN(n5508)
         );
  INV_X1 U3875 ( .A(n5299), .ZN(n5262) );
  NOR2_X1 U3876 ( .A1(n5104), .A2(n7077), .ZN(n5394) );
  INV_X1 U3877 ( .A(n4906), .ZN(n7077) );
  INV_X1 U3878 ( .A(n5340), .ZN(n5386) );
  AND2_X1 U3879 ( .A1(n7002), .A2(n7001), .ZN(n7016) );
  OR2_X1 U3880 ( .A1(n4818), .A2(n5949), .ZN(n4761) );
  INV_X1 U3881 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7028) );
  NAND2_X1 U3882 ( .A1(n5971), .A2(n5553), .ZN(n6931) );
  INV_X1 U3883 ( .A(n6947), .ZN(n6077) );
  NAND2_X1 U3884 ( .A1(n6850), .A2(n5554), .ZN(n6950) );
  AOI21_X1 U3885 ( .B1(n4739), .B2(n4738), .A(n4737), .ZN(n4740) );
  INV_X1 U3886 ( .A(n6524), .ZN(n6551) );
  OR2_X1 U3887 ( .A1(n4818), .A2(n7000), .ZN(n4820) );
  OR2_X1 U3888 ( .A1(n4818), .A2(n4802), .ZN(n6952) );
  OR2_X1 U3889 ( .A1(n6319), .A2(n6800), .ZN(n4192) );
  NOR2_X1 U3890 ( .A1(n5809), .A2(n6705), .ZN(n6817) );
  NAND2_X1 U3891 ( .A1(n4148), .A2(n4147), .ZN(n6800) );
  INV_X1 U3892 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5938) );
  INV_X1 U3893 ( .A(n6964), .ZN(n6959) );
  AND2_X1 U3894 ( .A1(n5126), .A2(n5125), .ZN(n5297) );
  OR2_X1 U3895 ( .A1(n7100), .A2(n4906), .ZN(n7108) );
  INV_X1 U3896 ( .A(n5394), .ZN(n5432) );
  OR2_X1 U3897 ( .A1(n5104), .A2(n4906), .ZN(n5158) );
  AND2_X1 U3898 ( .A1(n5165), .A2(n5164), .ZN(n5195) );
  NAND2_X1 U3899 ( .A1(n4955), .A2(n7077), .ZN(n5384) );
  AND2_X1 U3900 ( .A1(n5346), .A2(n5345), .ZN(n5389) );
  NAND2_X1 U3901 ( .A1(n5264), .A2(n4906), .ZN(n5340) );
  AOI22_X1 U3902 ( .A1(n7087), .A2(n7094), .B1(n7086), .B2(n7085), .ZN(n7193)
         );
  INV_X1 U3903 ( .A(n7182), .ZN(n5335) );
  OR2_X1 U3904 ( .A1(n5203), .A2(n4906), .ZN(n5225) );
  AND2_X1 U3905 ( .A1(n5229), .A2(n5228), .ZN(n5260) );
  AND2_X1 U3906 ( .A1(n7116), .A2(n5056), .ZN(n5085) );
  INV_X1 U3907 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7011) );
  NAND2_X1 U3908 ( .A1(n4741), .A2(n4740), .ZN(U2829) );
  INV_X1 U3909 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4152) );
  INV_X1 U3910 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3451) );
  NOR2_X2 U3911 ( .A1(n3451), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4786)
         );
  NOR2_X4 U3912 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4987) );
  AND2_X2 U3913 ( .A1(n4786), .A2(n4987), .ZN(n3874) );
  AND2_X4 U3914 ( .A1(n4785), .A2(n5011), .ZN(n3638) );
  AOI22_X1 U3915 ( .A1(n3874), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3458) );
  INV_X1 U3916 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3453) );
  INV_X1 U3917 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U3918 ( .A1(n3947), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3457) );
  AND2_X2 U3919 ( .A1(n4786), .A2(n5011), .ZN(n3635) );
  NOR2_X4 U3920 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5014) );
  AOI22_X1 U3921 ( .A1(n3635), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4644), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3456) );
  AND2_X2 U3922 ( .A1(n3459), .A2(n4986), .ZN(n3880) );
  AND2_X2 U3923 ( .A1(n5014), .A2(n4987), .ZN(n3910) );
  AOI22_X1 U3924 ( .A1(n3880), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3455) );
  AND2_X2 U3925 ( .A1(n4785), .A2(n4987), .ZN(n3921) );
  AND2_X2 U3926 ( .A1(n5014), .A2(n5011), .ZN(n3927) );
  AOI22_X1 U3927 ( .A1(n3921), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3927), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3464) );
  AND2_X2 U3928 ( .A1(n3460), .A2(n4785), .ZN(n3954) );
  AND2_X2 U3929 ( .A1(n4786), .A2(n3459), .ZN(n3630) );
  AOI22_X1 U3930 ( .A1(n3954), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3463) );
  AND2_X2 U3931 ( .A1(n3460), .A2(n4786), .ZN(n3628) );
  AOI22_X1 U3932 ( .A1(n3628), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3629), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3462) );
  AND2_X2 U3933 ( .A1(n3460), .A2(n5014), .ZN(n3955) );
  AOI22_X1 U3934 ( .A1(n3955), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3609), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3461) );
  NAND2_X2 U3935 ( .A1(n3466), .A2(n3465), .ZN(n3523) );
  BUF_X4 U3936 ( .A(n3523), .Z(n3649) );
  NAND2_X1 U3937 ( .A1(n3955), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3470) );
  NAND2_X1 U3938 ( .A1(n3954), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3469)
         );
  BUF_X2 U3939 ( .A(n3630), .Z(n3875) );
  NAND2_X1 U3940 ( .A1(n3875), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3468) );
  BUF_X4 U3941 ( .A(n3609), .Z(n4698) );
  NAND2_X1 U3942 ( .A1(n4698), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3467)
         );
  AND4_X2 U3943 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(n3486)
         );
  NAND2_X1 U3944 ( .A1(n3874), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3474) );
  NAND2_X1 U3945 ( .A1(n3638), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3473)
         );
  NAND2_X1 U3946 ( .A1(n3947), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3472) );
  NAND2_X1 U3947 ( .A1(n3922), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3471)
         );
  NAND2_X1 U3948 ( .A1(n3880), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3478) );
  NAND2_X1 U3949 ( .A1(n3635), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3477)
         );
  NAND2_X1 U3950 ( .A1(n4644), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3476) );
  NAND2_X1 U3951 ( .A1(n3910), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3475) );
  NAND2_X1 U3952 ( .A1(n3628), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3482) );
  NAND2_X1 U3953 ( .A1(n3921), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U3954 ( .A1(n3927), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3480)
         );
  NAND2_X1 U3955 ( .A1(n3629), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3479) );
  NAND2_X1 U3956 ( .A1(n3649), .A2(n3439), .ZN(n3517) );
  AOI22_X1 U3957 ( .A1(n3638), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3947), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U3958 ( .A1(n3635), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4644), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U3959 ( .A1(n3954), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3927), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U3960 ( .A1(n3880), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3487) );
  NAND4_X1 U3961 ( .A1(n3490), .A2(n3489), .A3(n3488), .A4(n3487), .ZN(n3496)
         );
  AOI22_X1 U3962 ( .A1(n3875), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U3963 ( .A1(n3874), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U3964 ( .A1(n3955), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3609), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U3965 ( .A1(n3628), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3432), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3491) );
  NAND4_X1 U3966 ( .A1(n3494), .A2(n3493), .A3(n3492), .A4(n3491), .ZN(n3495)
         );
  OR2_X4 U3967 ( .A1(n3496), .A2(n3495), .ZN(n4762) );
  NAND2_X1 U3968 ( .A1(n3874), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3500) );
  NAND2_X1 U3969 ( .A1(n3638), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3499)
         );
  NAND2_X1 U3970 ( .A1(n3947), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3498) );
  NAND2_X1 U3971 ( .A1(n3922), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3497)
         );
  NAND2_X1 U3972 ( .A1(n3955), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3504) );
  NAND2_X1 U3973 ( .A1(n3954), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3503)
         );
  NAND2_X1 U3974 ( .A1(n3630), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3502) );
  NAND2_X1 U3975 ( .A1(n3609), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3501)
         );
  NAND2_X1 U3976 ( .A1(n3635), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3508)
         );
  NAND2_X1 U3977 ( .A1(n3880), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3507) );
  NAND2_X1 U3978 ( .A1(n4644), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3506) );
  NAND2_X1 U3979 ( .A1(n3910), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3505) );
  NAND2_X1 U3980 ( .A1(n3628), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U3981 ( .A1(n3921), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3511) );
  NAND2_X1 U3982 ( .A1(n3927), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3510)
         );
  NAND2_X1 U3983 ( .A1(n3629), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3509) );
  NAND4_X4 U3984 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(n3657)
         );
  INV_X1 U3985 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3519) );
  XNOR2_X1 U3986 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3534) );
  NAND2_X1 U3987 ( .A1(n7103), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3521) );
  XNOR2_X1 U3988 ( .A(n3534), .B(n3533), .ZN(n3666) );
  NAND2_X1 U3989 ( .A1(n4002), .A2(n3666), .ZN(n3520) );
  OAI211_X1 U3990 ( .C1(n3537), .C2(n4928), .A(n3657), .B(n3520), .ZN(n3528)
         );
  INV_X1 U3991 ( .A(n3528), .ZN(n3532) );
  OAI21_X1 U3992 ( .B1(n7020), .B2(n3666), .A(n3556), .ZN(n3529) );
  INV_X1 U3993 ( .A(n3529), .ZN(n3531) );
  OAI21_X1 U3994 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7103), .A(n3521), 
        .ZN(n3524) );
  NOR2_X1 U3995 ( .A1(n3537), .A2(n3524), .ZN(n3527) );
  NOR2_X2 U3996 ( .A1(n4762), .A2(n3437), .ZN(n5946) );
  NOR2_X1 U3997 ( .A1(n3625), .A2(n4762), .ZN(n3522) );
  INV_X2 U3998 ( .A(n3523), .ZN(n3656) );
  NAND2_X1 U3999 ( .A1(n3656), .A2(n3657), .ZN(n3623) );
  INV_X1 U4000 ( .A(n3524), .ZN(n3525) );
  AOI21_X1 U4001 ( .B1(n4143), .B2(n3525), .A(n4935), .ZN(n3526) );
  OAI222_X1 U4002 ( .A1(n3529), .A2(n3528), .B1(n3566), .B2(n3527), .C1(n3546), 
        .C2(n3526), .ZN(n3530) );
  OAI21_X1 U4003 ( .B1(n3532), .B2(n3531), .A(n3530), .ZN(n3548) );
  NAND2_X1 U4004 ( .A1(n3534), .A2(n3533), .ZN(n3536) );
  NAND2_X1 U4005 ( .A1(n7099), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3535) );
  NAND2_X1 U4006 ( .A1(n3536), .A2(n3535), .ZN(n3542) );
  XNOR2_X1 U4007 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3541) );
  XNOR2_X1 U4008 ( .A(n3542), .B(n3541), .ZN(n3667) );
  INV_X1 U4009 ( .A(n3667), .ZN(n3540) );
  INV_X1 U4010 ( .A(n3546), .ZN(n3539) );
  INV_X1 U4011 ( .A(n3545), .ZN(n3538) );
  OAI211_X1 U4012 ( .C1(n3540), .C2(n4089), .A(n3539), .B(n3538), .ZN(n3547)
         );
  NAND2_X1 U4013 ( .A1(n3542), .A2(n3541), .ZN(n3544) );
  NAND2_X1 U4014 ( .A1(n6978), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3543) );
  NAND2_X1 U4015 ( .A1(n3544), .A2(n3543), .ZN(n3550) );
  MUX2_X1 U4016 ( .A(n7068), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n3549) );
  XNOR2_X1 U4017 ( .A(n3550), .B(n3549), .ZN(n3665) );
  AOI222_X1 U4018 ( .A1(n3548), .A2(n3547), .B1(n3546), .B2(n3545), .C1(n3665), 
        .C2(n4100), .ZN(n3558) );
  INV_X1 U4019 ( .A(n3665), .ZN(n3555) );
  NAND2_X1 U4020 ( .A1(n3550), .A2(n3549), .ZN(n3552) );
  NAND2_X1 U4021 ( .A1(n7068), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U4022 ( .A1(n3552), .A2(n3551), .ZN(n3561) );
  INV_X1 U4023 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3553) );
  NAND2_X1 U4024 ( .A1(n3554), .A2(n3553), .ZN(n3670) );
  AOI21_X1 U4025 ( .B1(n3555), .B2(n3670), .A(n4002), .ZN(n3557) );
  OAI22_X1 U4026 ( .A1(n3558), .A2(n3557), .B1(n3556), .B2(n3670), .ZN(n3559)
         );
  AOI21_X1 U4027 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7020), .A(n3559), 
        .ZN(n3565) );
  NAND2_X1 U4028 ( .A1(n3560), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3563) );
  NAND2_X1 U4029 ( .A1(n3561), .A2(n6983), .ZN(n3562) );
  NAND2_X1 U4030 ( .A1(n3563), .A2(n3562), .ZN(n3669) );
  NAND2_X1 U4031 ( .A1(n4087), .A2(n3669), .ZN(n3564) );
  NAND2_X1 U4032 ( .A1(n3565), .A2(n3564), .ZN(n3568) );
  NAND2_X1 U4033 ( .A1(n3875), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3572) );
  NAND2_X1 U4034 ( .A1(n3955), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3571) );
  NAND2_X1 U4035 ( .A1(n3628), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3570) );
  NAND2_X1 U4036 ( .A1(n3921), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3569) );
  NAND2_X1 U4037 ( .A1(n3947), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3576) );
  NAND2_X1 U4038 ( .A1(n3638), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3575)
         );
  NAND2_X1 U4040 ( .A1(n4644), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3574) );
  NAND2_X1 U4041 ( .A1(n3880), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3573) );
  NAND2_X1 U4043 ( .A1(n3922), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3580)
         );
  NAND2_X1 U4044 ( .A1(n3874), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3579) );
  NAND2_X1 U4045 ( .A1(n3635), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3578)
         );
  NAND2_X1 U4046 ( .A1(n3910), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3577) );
  NAND2_X1 U4047 ( .A1(n3954), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3584)
         );
  NAND2_X1 U4048 ( .A1(n4698), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3583)
         );
  NAND2_X1 U4049 ( .A1(n3629), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4050 ( .A1(n3927), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3581)
         );
  AND4_X2 U4051 ( .A1(n3584), .A2(n3583), .A3(n3582), .A4(n3581), .ZN(n3585)
         );
  NAND4_X4 U4052 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3654)
         );
  NAND2_X1 U4053 ( .A1(n3649), .A2(n3654), .ZN(n3651) );
  INV_X1 U4054 ( .A(n3651), .ZN(n3621) );
  NAND2_X1 U4055 ( .A1(n3880), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3592) );
  NAND2_X1 U4056 ( .A1(n3635), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3591)
         );
  NAND2_X1 U4057 ( .A1(n4644), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3590) );
  NAND2_X1 U4058 ( .A1(n3910), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4059 ( .A1(n3874), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4060 ( .A1(n3638), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3595)
         );
  NAND2_X1 U4061 ( .A1(n3947), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4062 ( .A1(n3922), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3593)
         );
  NAND2_X1 U4063 ( .A1(n3955), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3600) );
  NAND2_X1 U4064 ( .A1(n3954), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3599)
         );
  NAND2_X1 U4065 ( .A1(n3630), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3598) );
  NAND2_X1 U4066 ( .A1(n3609), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3597)
         );
  NAND2_X1 U4067 ( .A1(n3628), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3604) );
  NAND2_X1 U4068 ( .A1(n3921), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3603) );
  NAND2_X1 U4069 ( .A1(n3927), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3602)
         );
  NAND2_X1 U4070 ( .A1(n3629), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4071 ( .A1(n3628), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4072 ( .A1(n3947), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4073 ( .A1(n3954), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3609), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4074 ( .A1(n3921), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3927), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3610) );
  NAND4_X1 U4075 ( .A1(n3613), .A2(n3612), .A3(n3611), .A4(n3610), .ZN(n3619)
         );
  AOI22_X1 U4076 ( .A1(n3635), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4644), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4077 ( .A1(n3955), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4078 ( .A1(n3874), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3432), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4079 ( .A1(n3880), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3614) );
  NAND4_X1 U4080 ( .A1(n3617), .A2(n3616), .A3(n3615), .A4(n3614), .ZN(n3618)
         );
  OR2_X2 U4081 ( .A1(n3619), .A2(n3618), .ZN(n3664) );
  NAND2_X1 U4082 ( .A1(n3621), .A2(n3620), .ZN(n3626) );
  BUF_X1 U4083 ( .A(n3626), .Z(n3622) );
  INV_X1 U4084 ( .A(n3622), .ZN(n5930) );
  NAND2_X1 U4085 ( .A1(n5930), .A2(n4762), .ZN(n3706) );
  NAND2_X1 U4086 ( .A1(n3623), .A2(n3664), .ZN(n3624) );
  OAI21_X1 U4087 ( .B1(n3664), .B2(n3625), .A(n3624), .ZN(n3627) );
  NAND2_X2 U4088 ( .A1(n3675), .A2(n3654), .ZN(n5699) );
  OAI21_X1 U4089 ( .B1(n3627), .B2(n5699), .A(n3626), .ZN(n3646) );
  AOI22_X1 U4090 ( .A1(n3628), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3432), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4091 ( .A1(n3921), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3927), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4092 ( .A1(n3954), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3630), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4093 ( .A1(n3955), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3633) );
  NAND3_X1 U4094 ( .A1(n3634), .A2(n3447), .A3(n3633), .ZN(n3644) );
  BUF_X1 U4095 ( .A(n3922), .Z(n3637) );
  AOI22_X1 U4096 ( .A1(n3947), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3922), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4097 ( .A1(n3874), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4098 ( .A1(n3880), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3639) );
  NAND4_X1 U4099 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3643)
         );
  OR2_X2 U4100 ( .A1(n3644), .A2(n3643), .ZN(n3689) );
  NAND2_X1 U4101 ( .A1(n3847), .A2(n3689), .ZN(n3645) );
  NAND2_X1 U4102 ( .A1(n3646), .A2(n3645), .ZN(n3683) );
  INV_X1 U4103 ( .A(n3683), .ZN(n3648) );
  NOR2_X1 U4104 ( .A1(n4143), .A2(n3685), .ZN(n3647) );
  INV_X1 U4105 ( .A(n5948), .ZN(n5945) );
  OR2_X1 U4106 ( .A1(n3655), .A2(n3649), .ZN(n3650) );
  OR2_X1 U4107 ( .A1(n3847), .A2(n3651), .ZN(n3853) );
  INV_X2 U4108 ( .A(n3664), .ZN(n4925) );
  AOI21_X1 U4110 ( .B1(n3853), .B2(n4935), .A(n3837), .ZN(n3652) );
  AND2_X1 U4111 ( .A1(n3839), .A2(n3652), .ZN(n4144) );
  INV_X1 U4112 ( .A(n3831), .ZN(n4758) );
  NAND2_X1 U4113 ( .A1(n3847), .A2(n3685), .ZN(n3653) );
  NAND2_X1 U4114 ( .A1(n4758), .A2(n3653), .ZN(n3660) );
  NAND2_X1 U4115 ( .A1(n3655), .A2(n3654), .ZN(n4903) );
  INV_X1 U4116 ( .A(n4903), .ZN(n3659) );
  OAI21_X1 U4117 ( .B1(n4193), .B2(n3657), .A(n3656), .ZN(n3658) );
  INV_X1 U4118 ( .A(n3658), .ZN(n3830) );
  NAND2_X1 U4119 ( .A1(n3660), .A2(n3854), .ZN(n3687) );
  NAND2_X1 U4120 ( .A1(n4144), .A2(n3687), .ZN(n3661) );
  NAND2_X1 U4121 ( .A1(n5945), .A2(n3661), .ZN(n4777) );
  XNOR2_X1 U4122 ( .A(STATE_REG_2__SCAN_IN), .B(STATE_REG_1__SCAN_IN), .ZN(
        n3835) );
  INV_X1 U4123 ( .A(n3835), .ZN(n3663) );
  INV_X1 U4124 ( .A(STATE_REG_0__SCAN_IN), .ZN(n3662) );
  NAND2_X1 U4125 ( .A1(n3663), .A2(n3662), .ZN(n6684) );
  NAND2_X1 U4126 ( .A1(n4762), .A2(n6684), .ZN(n5954) );
  INV_X1 U4127 ( .A(READY_N), .ZN(n7042) );
  NOR3_X1 U4128 ( .A1(n3667), .A2(n3666), .A3(n3665), .ZN(n3668) );
  OR2_X1 U4129 ( .A1(n3669), .A2(n3668), .ZN(n3671) );
  NAND2_X1 U4130 ( .A1(n3671), .A2(n3670), .ZN(n5947) );
  NAND2_X1 U4131 ( .A1(n7042), .A2(n5947), .ZN(n4779) );
  INV_X1 U4132 ( .A(n4779), .ZN(n3672) );
  NAND3_X1 U4133 ( .A1(n5954), .A2(n3664), .A3(n3672), .ZN(n3673) );
  OAI211_X1 U4134 ( .C1(n7017), .C2(n3706), .A(n4777), .B(n3673), .ZN(n3674)
         );
  NAND2_X1 U4135 ( .A1(n3674), .A2(n7004), .ZN(n3682) );
  OR2_X2 U4136 ( .A1(n3837), .A2(n3675), .ZN(n3676) );
  NOR2_X2 U4137 ( .A1(n3676), .A2(n3854), .ZN(n3859) );
  NAND2_X1 U4138 ( .A1(n4928), .A2(n6684), .ZN(n5542) );
  AND2_X1 U4139 ( .A1(n5542), .A2(n7042), .ZN(n3679) );
  AOI21_X1 U4140 ( .B1(n5699), .B2(n3685), .A(n3664), .ZN(n3678) );
  AOI21_X1 U4141 ( .B1(n3677), .B2(n3679), .A(n3678), .ZN(n3680) );
  OR2_X1 U4142 ( .A1(n4818), .A2(n3680), .ZN(n3681) );
  AND2_X1 U4143 ( .A1(n5948), .A2(n4762), .ZN(n6969) );
  NAND2_X1 U4144 ( .A1(n4148), .A2(n6969), .ZN(n5749) );
  OAI21_X2 U4145 ( .B1(n3683), .B2(n4762), .A(n4935), .ZN(n3841) );
  NOR2_X1 U4146 ( .A1(n4143), .A2(n4928), .ZN(n3684) );
  OR2_X1 U4147 ( .A1(n3841), .A2(n3684), .ZN(n3858) );
  NAND2_X1 U4148 ( .A1(n4935), .A2(n4762), .ZN(n5547) );
  NOR2_X1 U4149 ( .A1(n5547), .A2(n3664), .ZN(n4775) );
  NAND2_X4 U4150 ( .A1(n4921), .A2(n3685), .ZN(n3806) );
  OAI21_X1 U4151 ( .B1(n4775), .B2(n4178), .A(n3837), .ZN(n3686) );
  NAND2_X1 U4152 ( .A1(n3664), .A2(n3685), .ZN(n3848) );
  AND4_X1 U4153 ( .A1(n3839), .A2(n3687), .A3(n3686), .A4(n3848), .ZN(n3688)
         );
  NAND2_X1 U4154 ( .A1(n3858), .A2(n3688), .ZN(n3705) );
  NOR2_X1 U4155 ( .A1(n3689), .A2(n3657), .ZN(n3690) );
  INV_X1 U4156 ( .A(n3853), .ZN(n3692) );
  NOR2_X1 U4157 ( .A1(n3934), .A2(n3664), .ZN(n3691) );
  NAND2_X1 U4158 ( .A1(n3692), .A2(n3691), .ZN(n5002) );
  INV_X1 U4159 ( .A(n3833), .ZN(n3695) );
  NAND2_X1 U4160 ( .A1(n3695), .A2(n4935), .ZN(n3696) );
  OAI211_X1 U4161 ( .C1(n3821), .C2(n3675), .A(n5002), .B(n3696), .ZN(n3697)
         );
  OR2_X1 U4162 ( .A1(n3705), .A2(n3697), .ZN(n3698) );
  NAND2_X1 U4163 ( .A1(n4148), .A2(n3698), .ZN(n6702) );
  NAND2_X1 U4164 ( .A1(n5749), .A2(n6702), .ZN(n5743) );
  INV_X1 U4165 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U4166 ( .A1(n5749), .A2(n6745), .ZN(n6719) );
  NAND2_X1 U4167 ( .A1(n5743), .A2(n6719), .ZN(n4889) );
  INV_X1 U4168 ( .A(n4889), .ZN(n6751) );
  INV_X1 U4169 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5043) );
  INV_X1 U4170 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4891) );
  INV_X1 U4171 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4890) );
  NOR3_X1 U4172 ( .A1(n5043), .A2(n4891), .A3(n4890), .ZN(n6734) );
  NAND2_X1 U4173 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6734), .ZN(n5744)
         );
  NAND2_X1 U4174 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6744) );
  INV_X1 U4175 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U4176 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6777) );
  NOR3_X1 U4177 ( .A1(n5661), .A2(n6788), .A3(n6777), .ZN(n5746) );
  INV_X1 U4178 ( .A(n5746), .ZN(n3699) );
  NOR3_X1 U4179 ( .A1(n5744), .A2(n6744), .A3(n3699), .ZN(n3710) );
  INV_X1 U4180 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6814) );
  INV_X1 U4181 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6806) );
  NOR2_X1 U4182 ( .A1(n6814), .A2(n6806), .ZN(n6805) );
  INV_X1 U4183 ( .A(n6805), .ZN(n3700) );
  INV_X1 U4184 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4119) );
  NAND2_X1 U4185 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5750) );
  NOR2_X1 U4186 ( .A1(n4119), .A2(n5750), .ZN(n6700) );
  NAND2_X1 U4187 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6700), .ZN(n6795) );
  NOR2_X1 U4188 ( .A1(n3700), .A2(n6795), .ZN(n3709) );
  NAND2_X1 U4189 ( .A1(n5809), .A2(n3709), .ZN(n6824) );
  NAND2_X1 U4190 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4129) );
  NAND2_X1 U4191 ( .A1(n3821), .A2(n3833), .ZN(n3702) );
  NOR2_X1 U4192 ( .A1(n3677), .A2(n3702), .ZN(n3703) );
  NAND2_X1 U4193 ( .A1(n5019), .A2(n3703), .ZN(n3704) );
  NAND2_X1 U4194 ( .A1(n4148), .A2(n5942), .ZN(n5752) );
  NAND2_X1 U4195 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n3709), .ZN(n6816) );
  INV_X1 U4196 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6741) );
  INV_X1 U4197 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6726) );
  INV_X1 U4198 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6752) );
  OAI21_X1 U4199 ( .B1(n6726), .B2(n6745), .A(n6752), .ZN(n6743) );
  NAND2_X1 U4200 ( .A1(n6734), .A2(n6743), .ZN(n5042) );
  NOR2_X1 U4201 ( .A1(n6741), .A2(n5042), .ZN(n6758) );
  NAND2_X1 U4202 ( .A1(n5746), .A2(n6758), .ZN(n5751) );
  OR2_X1 U4203 ( .A1(n6816), .A2(n5751), .ZN(n6512) );
  INV_X1 U4204 ( .A(n6512), .ZN(n3707) );
  NAND2_X1 U4205 ( .A1(n3707), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3715) );
  OR2_X1 U4206 ( .A1(n5752), .A2(n3715), .ZN(n3708) );
  AND2_X1 U4207 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U4208 ( .A1(n6506), .A2(n4743), .ZN(n4745) );
  AND2_X1 U4209 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3824) );
  OR2_X1 U4210 ( .A1(n4745), .A2(n3824), .ZN(n6486) );
  NAND2_X1 U4211 ( .A1(n3710), .A2(n3709), .ZN(n3711) );
  AND2_X1 U4212 ( .A1(n5743), .A2(n3711), .ZN(n3713) );
  NOR2_X1 U4213 ( .A1(n6702), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3712)
         );
  NOR2_X1 U4214 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7066) );
  AND2_X1 U4215 ( .A1(n7066), .A2(n7011), .ZN(n5596) );
  AND2_X2 U4216 ( .A1(n5596), .A2(n7020), .ZN(n6809) );
  NOR2_X1 U4217 ( .A1(n4148), .A2(n6809), .ZN(n6714) );
  OR2_X1 U4218 ( .A1(n3712), .A2(n6714), .ZN(n4887) );
  OR2_X1 U4219 ( .A1(n3713), .A2(n4887), .ZN(n6511) );
  AND2_X1 U4220 ( .A1(n5743), .A2(n4129), .ZN(n3714) );
  NOR2_X1 U4221 ( .A1(n6511), .A2(n3714), .ZN(n3718) );
  INV_X1 U4222 ( .A(n3715), .ZN(n3716) );
  OR2_X1 U4223 ( .A1(n5752), .A2(n3716), .ZN(n3717) );
  NAND2_X1 U4224 ( .A1(n3718), .A2(n3717), .ZN(n6500) );
  INV_X1 U4225 ( .A(n4743), .ZN(n6495) );
  OR2_X1 U4226 ( .A1(n6500), .A2(n6495), .ZN(n3720) );
  INV_X1 U4227 ( .A(n5752), .ZN(n6748) );
  INV_X1 U4228 ( .A(n6796), .ZN(n6721) );
  NAND2_X1 U4229 ( .A1(n3718), .A2(n6721), .ZN(n3719) );
  NAND2_X1 U4230 ( .A1(n3720), .A2(n3719), .ZN(n4746) );
  NAND2_X1 U4231 ( .A1(n6486), .A2(n4746), .ZN(n6489) );
  AND2_X1 U4232 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3825) );
  AOI21_X1 U4233 ( .B1(n4889), .B2(n5752), .A(n3825), .ZN(n3721) );
  NAND2_X1 U4234 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6446) );
  AND2_X1 U4235 ( .A1(n6796), .A2(n6446), .ZN(n3722) );
  NOR2_X1 U4236 ( .A1(n6466), .A2(n3722), .ZN(n6441) );
  MUX2_X1 U4237 ( .A(n3813), .B(n3812), .S(EBX_REG_1__SCAN_IN), .Z(n3723) );
  INV_X1 U4238 ( .A(EBX_REG_0__SCAN_IN), .ZN(n3726) );
  OAI22_X1 U4239 ( .A1(n3806), .A2(n3726), .B1(n3435), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4769) );
  XNOR2_X1 U4240 ( .A(n3728), .B(n4769), .ZN(n4816) );
  AOI21_X1 U4241 ( .B1(n4816), .B2(n3436), .A(n3728), .ZN(n4881) );
  MUX2_X1 U4242 ( .A(n3813), .B(n3435), .S(EBX_REG_2__SCAN_IN), .Z(n3729) );
  OAI21_X1 U4243 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n4178), .A(n3729), 
        .ZN(n3730) );
  INV_X1 U4244 ( .A(n3730), .ZN(n4880) );
  NAND2_X1 U4245 ( .A1(n4881), .A2(n4880), .ZN(n5670) );
  INV_X1 U4246 ( .A(n5670), .ZN(n3737) );
  MUX2_X1 U4247 ( .A(n3813), .B(n3435), .S(EBX_REG_4__SCAN_IN), .Z(n3731) );
  OAI21_X1 U4248 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n4178), .A(n3731), 
        .ZN(n3732) );
  INV_X1 U4249 ( .A(n3732), .ZN(n4893) );
  NAND2_X1 U4250 ( .A1(n3806), .A2(n4890), .ZN(n3734) );
  INV_X1 U4251 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U4252 ( .A1(n3436), .A2(n6625), .ZN(n3733) );
  NAND3_X1 U4253 ( .A1(n3734), .A2(n3435), .A3(n3733), .ZN(n3736) );
  NAND2_X1 U4254 ( .A1(n4181), .A2(n6625), .ZN(n3735) );
  NAND2_X1 U4255 ( .A1(n3736), .A2(n3735), .ZN(n5669) );
  NAND2_X1 U4256 ( .A1(n3806), .A2(n5043), .ZN(n3739) );
  INV_X1 U4257 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U4258 ( .A1(n3436), .A2(n6848), .ZN(n3738) );
  NAND3_X1 U4259 ( .A1(n3739), .A2(n3435), .A3(n3738), .ZN(n3741) );
  NAND2_X1 U4260 ( .A1(n4181), .A2(n6848), .ZN(n3740) );
  MUX2_X1 U4261 ( .A(n3813), .B(n3435), .S(EBX_REG_6__SCAN_IN), .Z(n3742) );
  OAI21_X1 U4262 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4178), .A(n3742), 
        .ZN(n3743) );
  INV_X1 U4263 ( .A(n3743), .ZN(n5438) );
  INV_X1 U4264 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4097) );
  NAND2_X1 U4265 ( .A1(n3806), .A2(n4097), .ZN(n3745) );
  INV_X1 U4266 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U4267 ( .A1(n3436), .A2(n6632), .ZN(n3744) );
  NAND3_X1 U4268 ( .A1(n3745), .A2(n3435), .A3(n3744), .ZN(n3747) );
  NAND2_X1 U4269 ( .A1(n4181), .A2(n6632), .ZN(n3746) );
  INV_X1 U4270 ( .A(n3813), .ZN(n3786) );
  INV_X1 U4271 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U4272 ( .A1(n3786), .A2(n5637), .ZN(n3750) );
  NAND2_X1 U4273 ( .A1(n3812), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3748)
         );
  OAI211_X1 U4274 ( .C1(n5552), .C2(EBX_REG_8__SCAN_IN), .A(n3806), .B(n3748), 
        .ZN(n3749) );
  NAND2_X1 U4275 ( .A1(n3750), .A2(n3749), .ZN(n5562) );
  NOR2_X1 U4276 ( .A1(n6626), .A2(n5562), .ZN(n3751) );
  NAND2_X1 U4277 ( .A1(n3806), .A2(n6788), .ZN(n3753) );
  INV_X1 U4278 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U4279 ( .A1(n3436), .A2(n5599), .ZN(n3752) );
  NAND3_X1 U4280 ( .A1(n3753), .A2(n3435), .A3(n3752), .ZN(n3755) );
  NAND2_X1 U4281 ( .A1(n4181), .A2(n5599), .ZN(n3754) );
  AND2_X1 U4282 ( .A1(n3755), .A2(n3754), .ZN(n5594) );
  OR2_X2 U4283 ( .A1(n5593), .A2(n5594), .ZN(n5603) );
  MUX2_X1 U4284 ( .A(n3813), .B(n3435), .S(EBX_REG_10__SCAN_IN), .Z(n3756) );
  OAI21_X1 U4285 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n4178), .A(n3756), 
        .ZN(n5604) );
  INV_X1 U4286 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U4287 ( .A1(n3806), .A2(n5799), .ZN(n3758) );
  INV_X1 U4288 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U4289 ( .A1(n3436), .A2(n5628), .ZN(n3757) );
  NAND3_X1 U4290 ( .A1(n3758), .A2(n3435), .A3(n3757), .ZN(n3760) );
  NAND2_X1 U4291 ( .A1(n4181), .A2(n5628), .ZN(n3759) );
  NAND2_X1 U4292 ( .A1(n3760), .A2(n3759), .ZN(n5624) );
  INV_X1 U4293 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U4294 ( .A1(n3786), .A2(n6898), .ZN(n3763) );
  NAND2_X1 U4295 ( .A1(n3435), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3761) );
  OAI211_X1 U4296 ( .C1(n5552), .C2(EBX_REG_12__SCAN_IN), .A(n3806), .B(n3761), 
        .ZN(n3762) );
  NAND2_X1 U4297 ( .A1(n5806), .A2(n5805), .ZN(n5683) );
  MUX2_X1 U4298 ( .A(n3813), .B(n3435), .S(EBX_REG_14__SCAN_IN), .Z(n3764) );
  OAI21_X1 U4299 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n4178), .A(n3764), 
        .ZN(n5684) );
  INV_X1 U4300 ( .A(n5684), .ZN(n3769) );
  NAND2_X1 U4301 ( .A1(n3806), .A2(n4119), .ZN(n3766) );
  INV_X1 U4302 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6908) );
  NAND2_X1 U4303 ( .A1(n3436), .A2(n6908), .ZN(n3765) );
  NAND3_X1 U4304 ( .A1(n3766), .A2(n3435), .A3(n3765), .ZN(n3768) );
  NAND2_X1 U4305 ( .A1(n4181), .A2(n6908), .ZN(n3767) );
  NAND2_X1 U4306 ( .A1(n3768), .A2(n3767), .ZN(n5754) );
  NAND2_X1 U4307 ( .A1(n3769), .A2(n5754), .ZN(n3770) );
  OR2_X2 U4308 ( .A1(n5683), .A2(n3770), .ZN(n5786) );
  NAND2_X1 U4309 ( .A1(n3806), .A2(n6806), .ZN(n3772) );
  INV_X1 U4310 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U4311 ( .A1(n3436), .A2(n5793), .ZN(n3771) );
  NAND3_X1 U4312 ( .A1(n3772), .A2(n3812), .A3(n3771), .ZN(n3774) );
  NAND2_X1 U4313 ( .A1(n4181), .A2(n5793), .ZN(n3773) );
  AND2_X1 U4314 ( .A1(n3774), .A2(n3773), .ZN(n5787) );
  NOR2_X2 U4315 ( .A1(n5786), .A2(n5787), .ZN(n5788) );
  MUX2_X1 U4316 ( .A(n3813), .B(n3812), .S(EBX_REG_16__SCAN_IN), .Z(n3775) );
  OAI21_X1 U4317 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n4178), .A(n3775), 
        .ZN(n5855) );
  INV_X1 U4318 ( .A(n5855), .ZN(n3776) );
  INV_X1 U4320 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3777) );
  NAND2_X1 U4321 ( .A1(n3806), .A2(n3777), .ZN(n3779) );
  INV_X1 U4322 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U4323 ( .A1(n3436), .A2(n5721), .ZN(n3778) );
  NAND3_X1 U4324 ( .A1(n3779), .A2(n3435), .A3(n3778), .ZN(n3781) );
  NAND2_X1 U4325 ( .A1(n4181), .A2(n5721), .ZN(n3780) );
  NAND2_X1 U4326 ( .A1(n3781), .A2(n3780), .ZN(n5713) );
  NAND2_X1 U4327 ( .A1(n5712), .A2(n5713), .ZN(n5711) );
  MUX2_X1 U4328 ( .A(n3813), .B(n3435), .S(EBX_REG_18__SCAN_IN), .Z(n3782) );
  OAI21_X1 U4329 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n4178), .A(n3782), 
        .ZN(n5725) );
  NAND2_X1 U4330 ( .A1(n3435), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3783) );
  NAND2_X1 U4331 ( .A1(n3806), .A2(n3783), .ZN(n3785) );
  INV_X1 U4332 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U4333 ( .A1(n3436), .A2(n5818), .ZN(n3784) );
  AOI22_X1 U4334 ( .A1(n3785), .A2(n3784), .B1(n4181), .B2(n5818), .ZN(n5763)
         );
  INV_X1 U4335 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U4336 ( .A1(n3786), .A2(n5841), .ZN(n3789) );
  NAND2_X1 U4337 ( .A1(n3435), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3787) );
  OAI211_X1 U4338 ( .C1(n5552), .C2(EBX_REG_20__SCAN_IN), .A(n3806), .B(n3787), 
        .ZN(n3788) );
  AND2_X1 U4339 ( .A1(n3789), .A2(n3788), .ZN(n5832) );
  NAND2_X1 U4340 ( .A1(n5833), .A2(n5832), .ZN(n4747) );
  NAND2_X1 U4341 ( .A1(n3435), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3790) );
  NAND2_X1 U4342 ( .A1(n3806), .A2(n3790), .ZN(n3792) );
  INV_X1 U4343 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U4344 ( .A1(n3436), .A2(n5869), .ZN(n3791) );
  AOI22_X1 U4345 ( .A1(n3792), .A2(n3791), .B1(n4181), .B2(n5869), .ZN(n4748)
         );
  OR2_X2 U4346 ( .A1(n4747), .A2(n4748), .ZN(n5885) );
  MUX2_X1 U4347 ( .A(n3813), .B(n3435), .S(EBX_REG_22__SCAN_IN), .Z(n3793) );
  OAI21_X1 U4348 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4178), .A(n3793), 
        .ZN(n5886) );
  OR2_X2 U4349 ( .A1(n5885), .A2(n5886), .ZN(n6065) );
  NAND2_X1 U4350 ( .A1(n3806), .A2(n6362), .ZN(n3794) );
  OAI211_X1 U4351 ( .C1(EBX_REG_23__SCAN_IN), .C2(n5552), .A(n3794), .B(n3435), 
        .ZN(n3797) );
  INV_X1 U4352 ( .A(EBX_REG_23__SCAN_IN), .ZN(n3795) );
  NAND2_X1 U4353 ( .A1(n4181), .A2(n3795), .ZN(n3796) );
  AND2_X1 U4354 ( .A1(n3797), .A2(n3796), .ZN(n6064) );
  MUX2_X1 U4355 ( .A(n3813), .B(n3435), .S(EBX_REG_24__SCAN_IN), .Z(n3800) );
  INV_X1 U4356 ( .A(n4178), .ZN(n4770) );
  INV_X1 U4357 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3798) );
  NAND2_X1 U4358 ( .A1(n4770), .A2(n3798), .ZN(n3799) );
  NAND2_X1 U4359 ( .A1(n3800), .A2(n3799), .ZN(n6054) );
  INV_X1 U4360 ( .A(n6054), .ZN(n3801) );
  INV_X1 U4361 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U4362 ( .A1(n3806), .A2(n6450), .ZN(n3802) );
  OAI211_X1 U4363 ( .C1(EBX_REG_25__SCAN_IN), .C2(n5552), .A(n3802), .B(n3435), 
        .ZN(n3804) );
  INV_X1 U4364 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U4365 ( .A1(n4181), .A2(n6279), .ZN(n3803) );
  NAND2_X1 U4366 ( .A1(n3804), .A2(n3803), .ZN(n6043) );
  NAND2_X1 U4367 ( .A1(n6041), .A2(n6043), .ZN(n6042) );
  MUX2_X1 U4368 ( .A(n3813), .B(n3812), .S(EBX_REG_26__SCAN_IN), .Z(n3805) );
  OAI21_X1 U4369 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n4178), .A(n3805), 
        .ZN(n6022) );
  OR2_X2 U4370 ( .A1(n6042), .A2(n6022), .ZN(n6020) );
  INV_X1 U4371 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U4372 ( .A1(n3806), .A2(n6440), .ZN(n3808) );
  INV_X1 U4373 ( .A(EBX_REG_27__SCAN_IN), .ZN(n3809) );
  NAND2_X1 U4374 ( .A1(n3436), .A2(n3809), .ZN(n3807) );
  NAND3_X1 U4375 ( .A1(n3808), .A2(n3435), .A3(n3807), .ZN(n3811) );
  NAND2_X1 U4376 ( .A1(n4181), .A2(n3809), .ZN(n3810) );
  NAND2_X1 U4377 ( .A1(n3811), .A2(n3810), .ZN(n6008) );
  INV_X1 U4378 ( .A(n6008), .ZN(n3815) );
  MUX2_X1 U4379 ( .A(n3813), .B(n3812), .S(EBX_REG_28__SCAN_IN), .Z(n3814) );
  OAI21_X1 U4380 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n4178), .A(n3814), 
        .ZN(n3817) );
  OAI21_X1 U4381 ( .B1(n6020), .B2(n3815), .A(n3817), .ZN(n3816) );
  INV_X1 U4382 ( .A(n3816), .ZN(n3820) );
  INV_X1 U4383 ( .A(n3817), .ZN(n3818) );
  NAND2_X1 U4384 ( .A1(n3818), .A2(n6008), .ZN(n3819) );
  NOR2_X4 U4385 ( .A1(n6020), .A2(n3819), .ZN(n4731) );
  OR2_X1 U4386 ( .A1(n3820), .A2(n4731), .ZN(n6083) );
  NAND2_X1 U4387 ( .A1(n3677), .A2(n6692), .ZN(n7000) );
  NOR2_X2 U4388 ( .A1(n3821), .A2(n5699), .ZN(n4145) );
  NAND2_X1 U4389 ( .A1(n4145), .A2(n4978), .ZN(n3822) );
  NAND2_X1 U4390 ( .A1(n7000), .A2(n3822), .ZN(n3823) );
  AND2_X2 U4391 ( .A1(n4148), .A2(n3823), .ZN(n6826) );
  INV_X1 U4392 ( .A(n6826), .ZN(n6799) );
  AND2_X1 U4393 ( .A1(n4743), .A2(n3824), .ZN(n6474) );
  NAND2_X1 U4394 ( .A1(n6474), .A2(n3825), .ZN(n6447) );
  NOR2_X1 U4395 ( .A1(n6447), .A2(n6446), .ZN(n3826) );
  AND2_X1 U4396 ( .A1(n6506), .A2(n3826), .ZN(n6438) );
  XNOR2_X1 U4397 ( .A(n6440), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3827)
         );
  AND2_X1 U4398 ( .A1(n6809), .A2(REIP_REG_28__SCAN_IN), .ZN(n5921) );
  AOI21_X1 U4399 ( .B1(n6438), .B2(n3827), .A(n5921), .ZN(n3828) );
  OAI21_X1 U4400 ( .B1(n6083), .B2(n6799), .A(n3828), .ZN(n3829) );
  INV_X1 U4401 ( .A(n3829), .ZN(n4151) );
  NAND2_X1 U4402 ( .A1(n3830), .A2(n5697), .ZN(n3832) );
  NAND2_X1 U4403 ( .A1(n3832), .A2(n3831), .ZN(n3834) );
  NAND2_X1 U4404 ( .A1(n3836), .A2(n3835), .ZN(n3860) );
  NAND3_X1 U4405 ( .A1(n3841), .A2(n3851), .A3(n3840), .ZN(n3842) );
  NAND2_X1 U4406 ( .A1(n3842), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3844) );
  NAND2_X1 U4407 ( .A1(n3844), .A2(n3843), .ZN(n3900) );
  NAND2_X1 U4408 ( .A1(n3900), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3846) );
  NOR2_X1 U4409 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7003) );
  NAND2_X1 U4410 ( .A1(n7003), .A2(n7020), .ZN(n4803) );
  MUX2_X1 U4411 ( .A(n4803), .B(n3864), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3845) );
  NAND2_X1 U4412 ( .A1(n3846), .A2(n3845), .ZN(n3893) );
  INV_X1 U4413 ( .A(n3847), .ZN(n3850) );
  NAND3_X1 U4414 ( .A1(n3848), .A2(n7003), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3849) );
  AOI21_X1 U4415 ( .B1(n6692), .B2(n3850), .A(n3849), .ZN(n3857) );
  NAND3_X1 U4416 ( .A1(n3622), .A2(n4928), .A3(n4758), .ZN(n3852) );
  NAND2_X1 U4417 ( .A1(n3852), .A2(n4921), .ZN(n3856) );
  NAND3_X1 U4418 ( .A1(n3854), .A2(n4762), .A3(n3853), .ZN(n3855) );
  AOI21_X1 U4419 ( .B1(n4755), .B2(n3860), .A(n4145), .ZN(n3862) );
  NAND2_X1 U4420 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  NAND2_X1 U4421 ( .A1(n3863), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3871) );
  INV_X1 U4422 ( .A(n3871), .ZN(n3869) );
  NAND2_X1 U4423 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6972) );
  OAI21_X1 U4424 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6972), .ZN(n5348) );
  OR2_X1 U4425 ( .A1(n4803), .A2(n5348), .ZN(n3866) );
  INV_X1 U4426 ( .A(n3864), .ZN(n3988) );
  NAND2_X1 U4427 ( .A1(n3988), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3865) );
  INV_X1 U4428 ( .A(n3870), .ZN(n3867) );
  NAND2_X1 U4429 ( .A1(n3869), .A2(n3868), .ZN(n3873) );
  NAND2_X1 U4430 ( .A1(n3900), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3872) );
  NAND3_X2 U4431 ( .A1(n3872), .A2(n3871), .A3(n3870), .ZN(n3897) );
  XNOR2_X1 U4432 ( .A(n3899), .B(n3424), .ZN(n4788) );
  NAND2_X1 U4433 ( .A1(n4788), .A2(n7020), .ZN(n3890) );
  AOI22_X1 U4434 ( .A1(n4708), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4435 ( .A1(n3422), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4436 ( .A1(n4706), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4437 ( .A1(n4700), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4438 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3887)
         );
  BUF_X1 U4439 ( .A(n3635), .Z(n4645) );
  AOI22_X1 U4440 ( .A1(n4600), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3885) );
  INV_X1 U4441 ( .A(n3880), .ZN(n3905) );
  AOI22_X1 U4442 ( .A1(n4699), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3884) );
  INV_X1 U4443 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4444 ( .A1(n4601), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4445 ( .A1(n3949), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3882) );
  NAND4_X1 U4446 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3886)
         );
  AND2_X1 U4447 ( .A1(n4978), .A2(n3942), .ZN(n3888) );
  NAND2_X1 U4448 ( .A1(n4935), .A2(n3942), .ZN(n3891) );
  AND2_X1 U4449 ( .A1(n3891), .A2(n3649), .ZN(n3894) );
  NAND2_X1 U4450 ( .A1(n4002), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3895) );
  NAND2_X2 U4451 ( .A1(n3896), .A2(n3895), .ZN(n3940) );
  OAI21_X2 U4452 ( .B1(n3899), .B2(n3898), .A(n3897), .ZN(n3982) );
  NAND2_X1 U4453 ( .A1(n3985), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3904) );
  INV_X1 U4454 ( .A(n6972), .ZN(n3901) );
  AND2_X1 U4455 ( .A1(n3901), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3986)
         );
  INV_X1 U4456 ( .A(n3986), .ZN(n5052) );
  NAND2_X1 U4457 ( .A1(n6972), .A2(n6978), .ZN(n3902) );
  AND2_X1 U4458 ( .A1(n5052), .A2(n3902), .ZN(n5128) );
  INV_X1 U4459 ( .A(n4803), .ZN(n3989) );
  AOI22_X1 U4460 ( .A1(n5128), .A2(n3989), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3988), .ZN(n3903) );
  XNOR2_X1 U4461 ( .A(n3982), .B(n3983), .ZN(n4910) );
  NAND2_X1 U4462 ( .A1(n4910), .A2(n7020), .ZN(n3918) );
  AOI22_X1 U4463 ( .A1(n3422), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4699), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4464 ( .A1(n4708), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4706), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3908) );
  INV_X2 U4465 ( .A(n3905), .ZN(n4697) );
  AOI22_X1 U4466 ( .A1(n3948), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4467 ( .A1(n4707), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4468 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3916)
         );
  AOI22_X1 U4469 ( .A1(n4705), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4470 ( .A1(n4645), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4471 ( .A1(n4700), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4472 ( .A1(n4600), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3911) );
  NAND4_X1 U4473 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3915)
         );
  AOI22_X1 U4474 ( .A1(n4002), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4087), 
        .B2(n4009), .ZN(n3917) );
  OR2_X2 U4475 ( .A1(n3919), .A2(n3920), .ZN(n4905) );
  NAND2_X2 U4476 ( .A1(n3920), .A2(n3919), .ZN(n4006) );
  AOI22_X1 U4477 ( .A1(n3955), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4478 ( .A1(n4706), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3925) );
  CLKBUF_X1 U4479 ( .A(n3922), .Z(n3948) );
  AOI22_X1 U4480 ( .A1(n4600), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4481 ( .A1(n4666), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3923) );
  NAND4_X1 U4482 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(n3933)
         );
  AOI22_X1 U4483 ( .A1(n4700), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4484 ( .A1(n4601), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4485 ( .A1(n4708), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4486 ( .A1(n3422), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U4487 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3932)
         );
  NAND2_X1 U4488 ( .A1(n3971), .A2(n3942), .ZN(n4011) );
  XNOR2_X1 U4489 ( .A(n4011), .B(n4009), .ZN(n3935) );
  NAND2_X1 U4490 ( .A1(n4935), .A2(n3934), .ZN(n3970) );
  OAI21_X1 U4491 ( .B1(n3935), .B2(n4758), .A(n3970), .ZN(n3936) );
  INV_X1 U4492 ( .A(n3936), .ZN(n3937) );
  INV_X1 U4493 ( .A(n3938), .ZN(n6640) );
  INV_X1 U4494 ( .A(n3939), .ZN(n3941) );
  NAND2_X1 U4495 ( .A1(n4194), .A2(n4100), .ZN(n3977) );
  INV_X1 U4496 ( .A(n3942), .ZN(n3943) );
  XNOR2_X1 U4497 ( .A(n3943), .B(n3971), .ZN(n3945) );
  NAND2_X1 U4498 ( .A1(n4925), .A2(n3657), .ZN(n3944) );
  AOI21_X1 U4499 ( .B1(n3945), .B2(n6692), .A(n3944), .ZN(n3975) );
  NAND2_X1 U4500 ( .A1(n3977), .A2(n3975), .ZN(n3946) );
  INV_X1 U4501 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5157) );
  AOI21_X1 U4502 ( .B1(n4935), .B2(n3971), .A(n7020), .ZN(n3963) );
  AOI22_X1 U4503 ( .A1(n4700), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4504 ( .A1(n4708), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4706), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4505 ( .A1(n4600), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4506 ( .A1(n4666), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3950) );
  NAND4_X1 U4507 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3961)
         );
  AOI22_X1 U4508 ( .A1(n4697), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4509 ( .A1(n3422), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4510 ( .A1(n4672), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3432), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4511 ( .A1(n3955), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U4512 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3960)
         );
  NAND2_X1 U4514 ( .A1(n4978), .A2(n4104), .ZN(n3962) );
  OAI211_X1 U4515 ( .C1(n4089), .C2(n5157), .A(n3963), .B(n3962), .ZN(n3967)
         );
  INV_X1 U4516 ( .A(n4104), .ZN(n3964) );
  XNOR2_X1 U4517 ( .A(n3964), .B(n3971), .ZN(n3965) );
  NOR2_X1 U4518 ( .A1(n3649), .A2(n7020), .ZN(n4101) );
  NAND2_X1 U4519 ( .A1(n3965), .A2(n4101), .ZN(n3966) );
  OR2_X1 U4520 ( .A1(n4906), .A2(n4062), .ZN(n3974) );
  OAI21_X1 U4521 ( .B1(n4758), .B2(n3971), .A(n3970), .ZN(n3972) );
  INV_X1 U4522 ( .A(n3972), .ZN(n3973) );
  NAND2_X1 U4523 ( .A1(n3974), .A2(n3973), .ZN(n4766) );
  NAND2_X1 U4524 ( .A1(n4766), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5528)
         );
  NAND2_X1 U4525 ( .A1(n5525), .A2(n5528), .ZN(n3979) );
  AND2_X1 U4526 ( .A1(n3975), .A2(n6726), .ZN(n3976) );
  NAND2_X1 U4527 ( .A1(n3977), .A2(n3976), .ZN(n5526) );
  AND2_X1 U4528 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3978)
         );
  NAND2_X1 U4529 ( .A1(n3979), .A2(n3978), .ZN(n6637) );
  NAND2_X1 U4530 ( .A1(n6640), .A2(n6637), .ZN(n3981) );
  NAND2_X1 U4531 ( .A1(n3427), .A2(n5526), .ZN(n3980) );
  NAND2_X1 U4532 ( .A1(n3980), .A2(n6752), .ZN(n6638) );
  AND2_X1 U4533 ( .A1(n3981), .A2(n6638), .ZN(n4016) );
  INV_X1 U4534 ( .A(n3982), .ZN(n3984) );
  NAND2_X1 U4535 ( .A1(n3985), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3991) );
  NAND2_X1 U4536 ( .A1(n3986), .A2(n7068), .ZN(n4956) );
  NAND2_X1 U4537 ( .A1(n5052), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3987) );
  NAND2_X1 U4538 ( .A1(n4956), .A2(n3987), .ZN(n5347) );
  AOI22_X1 U4539 ( .A1(n5347), .A2(n3989), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3988), .ZN(n3990) );
  AOI22_X1 U4540 ( .A1(n4706), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4541 ( .A1(n4600), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4542 ( .A1(n4645), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4543 ( .A1(n4697), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3992) );
  NAND4_X1 U4544 ( .A1(n3995), .A2(n3994), .A3(n3993), .A4(n3992), .ZN(n4001)
         );
  AOI22_X1 U4545 ( .A1(n3422), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4546 ( .A1(n4705), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4547 ( .A1(n4708), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4548 ( .A1(n4699), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3996) );
  NAND4_X1 U4549 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n4000)
         );
  AOI22_X1 U4550 ( .A1(n4002), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4087), 
        .B2(n4031), .ZN(n4003) );
  INV_X1 U4551 ( .A(n4954), .ZN(n5053) );
  NAND2_X1 U4552 ( .A1(n5053), .A2(n4006), .ZN(n4007) );
  INV_X1 U4553 ( .A(n4904), .ZN(n4008) );
  NAND2_X1 U4554 ( .A1(n4008), .A2(n4100), .ZN(n4015) );
  INV_X1 U4555 ( .A(n4009), .ZN(n4010) );
  NAND2_X1 U4556 ( .A1(n4011), .A2(n4010), .ZN(n4032) );
  INV_X1 U4557 ( .A(n4031), .ZN(n4012) );
  XNOR2_X1 U4558 ( .A(n4032), .B(n4012), .ZN(n4013) );
  NAND2_X1 U4559 ( .A1(n4013), .A2(n6692), .ZN(n4014) );
  AND2_X1 U4560 ( .A1(n4015), .A2(n4014), .ZN(n6648) );
  NAND2_X1 U4561 ( .A1(n6646), .A2(n6648), .ZN(n4018) );
  INV_X1 U4562 ( .A(n4016), .ZN(n4017) );
  NAND2_X1 U4563 ( .A1(n4017), .A2(n4890), .ZN(n6645) );
  NAND2_X1 U4564 ( .A1(n4018), .A2(n6645), .ZN(n4885) );
  INV_X1 U4565 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5296) );
  OR2_X1 U4566 ( .A1(n4089), .A2(n5296), .ZN(n4030) );
  AOI22_X1 U4567 ( .A1(n4706), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4568 ( .A1(n4600), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4569 ( .A1(n4645), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4570 ( .A1(n4697), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4019) );
  NAND4_X1 U4571 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(n4028)
         );
  AOI22_X1 U4572 ( .A1(n3422), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4573 ( .A1(n4705), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4574 ( .A1(n4708), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4575 ( .A1(n4699), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U4576 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4027)
         );
  NAND2_X1 U4577 ( .A1(n4087), .A2(n4056), .ZN(n4029) );
  NAND2_X1 U4578 ( .A1(n4030), .A2(n4029), .ZN(n4038) );
  NAND2_X1 U4579 ( .A1(n4227), .A2(n4100), .ZN(n4035) );
  NAND2_X1 U4580 ( .A1(n4032), .A2(n4031), .ZN(n4058) );
  XNOR2_X1 U4581 ( .A(n4058), .B(n4056), .ZN(n4033) );
  NAND2_X1 U4582 ( .A1(n4033), .A2(n6692), .ZN(n4034) );
  NAND2_X1 U4583 ( .A1(n4035), .A2(n4034), .ZN(n4036) );
  XNOR2_X1 U4584 ( .A(n4036), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4886)
         );
  NAND2_X1 U4585 ( .A1(n4036), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4037)
         );
  OAI21_X1 U4586 ( .B1(n4885), .B2(n4886), .A(n4037), .ZN(n5036) );
  NOR2_X2 U4587 ( .A1(n4040), .A2(n4039), .ZN(n4054) );
  INV_X1 U4588 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5134) );
  OR2_X1 U4589 ( .A1(n4089), .A2(n5134), .ZN(n4052) );
  AOI22_X1 U4590 ( .A1(n4706), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4591 ( .A1(n4708), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4592 ( .A1(n4699), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4593 ( .A1(n4707), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U4594 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4050)
         );
  AOI22_X1 U4595 ( .A1(n3422), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4600), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4596 ( .A1(n4700), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4597 ( .A1(n3637), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U4598 ( .A1(n4672), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U4599 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4049)
         );
  NAND2_X1 U4600 ( .A1(n4087), .A2(n4059), .ZN(n4051) );
  NAND2_X1 U4601 ( .A1(n4052), .A2(n4051), .ZN(n4053) );
  NAND2_X1 U4602 ( .A1(n4054), .A2(n4053), .ZN(n4081) );
  NAND2_X1 U4603 ( .A1(n4081), .A2(n4055), .ZN(n4228) );
  INV_X1 U4604 ( .A(n4056), .ZN(n4057) );
  NOR2_X1 U4605 ( .A1(n4058), .A2(n4057), .ZN(n4060) );
  NAND2_X1 U4606 ( .A1(n4060), .A2(n4059), .ZN(n4091) );
  OAI211_X1 U4607 ( .C1(n4060), .C2(n4059), .A(n4091), .B(n6692), .ZN(n4061)
         );
  XNOR2_X1 U4608 ( .A(n4063), .B(n5043), .ZN(n5038) );
  NAND2_X1 U4609 ( .A1(n5036), .A2(n5038), .ZN(n4065) );
  NAND2_X1 U4610 ( .A1(n4063), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4064)
         );
  NAND2_X1 U4611 ( .A1(n4065), .A2(n4064), .ZN(n6653) );
  INV_X1 U4612 ( .A(n4081), .ZN(n4079) );
  INV_X1 U4613 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5142) );
  OR2_X1 U4614 ( .A1(n4089), .A2(n5142), .ZN(n4077) );
  AOI22_X1 U4615 ( .A1(n4706), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4616 ( .A1(n4600), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U4617 ( .A1(n4645), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U4618 ( .A1(n4697), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4066) );
  NAND4_X1 U4619 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4075)
         );
  AOI22_X1 U4620 ( .A1(n3422), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4621 ( .A1(n4705), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U4622 ( .A1(n4708), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4623 ( .A1(n4699), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4070) );
  NAND4_X1 U4624 ( .A1(n4073), .A2(n4072), .A3(n4071), .A4(n4070), .ZN(n4074)
         );
  NAND2_X1 U4625 ( .A1(n4087), .A2(n4092), .ZN(n4076) );
  INV_X1 U4626 ( .A(n4080), .ZN(n4078) );
  NAND2_X1 U4627 ( .A1(n4081), .A2(n4080), .ZN(n4240) );
  NAND3_X1 U4628 ( .A1(n4103), .A2(n4240), .A3(n4100), .ZN(n4084) );
  XNOR2_X1 U4629 ( .A(n4091), .B(n4092), .ZN(n4082) );
  NAND2_X1 U4630 ( .A1(n4082), .A2(n6692), .ZN(n4083) );
  NAND2_X1 U4631 ( .A1(n4084), .A2(n4083), .ZN(n4085) );
  OR2_X1 U4632 ( .A1(n4085), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6655)
         );
  NAND2_X1 U4633 ( .A1(n6653), .A2(n6655), .ZN(n4086) );
  NAND2_X1 U4634 ( .A1(n4085), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6654)
         );
  NAND2_X1 U4635 ( .A1(n4086), .A2(n6654), .ZN(n6661) );
  INV_X1 U4636 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U4637 ( .A1(n4087), .A2(n4104), .ZN(n4088) );
  OAI21_X1 U4638 ( .B1(n4089), .B2(n5153), .A(n4088), .ZN(n4090) );
  NAND2_X1 U4639 ( .A1(n4248), .A2(n4100), .ZN(n4096) );
  INV_X1 U4640 ( .A(n4091), .ZN(n4093) );
  NAND2_X1 U4641 ( .A1(n4093), .A2(n4092), .ZN(n4106) );
  XNOR2_X1 U4642 ( .A(n4106), .B(n4104), .ZN(n4094) );
  NAND2_X1 U4643 ( .A1(n4094), .A2(n6692), .ZN(n4095) );
  NAND2_X1 U4644 ( .A1(n4096), .A2(n4095), .ZN(n4098) );
  XNOR2_X1 U4645 ( .A(n4098), .B(n4097), .ZN(n6660) );
  NAND2_X1 U4646 ( .A1(n6661), .A2(n6660), .ZN(n6659) );
  NAND2_X1 U4647 ( .A1(n4098), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4099)
         );
  NAND2_X1 U4648 ( .A1(n6659), .A2(n4099), .ZN(n5573) );
  NAND2_X1 U4649 ( .A1(n6692), .A2(n4104), .ZN(n4105) );
  OR2_X1 U4650 ( .A1(n4106), .A2(n4105), .ZN(n4107) );
  NAND2_X1 U4651 ( .A1(n4140), .A2(n4107), .ZN(n4109) );
  INV_X1 U4652 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4108) );
  XNOR2_X1 U4653 ( .A(n4109), .B(n4108), .ZN(n5572) );
  NAND2_X1 U4654 ( .A1(n4109), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5606)
         );
  AND2_X1 U4655 ( .A1(n5606), .A2(n4110), .ZN(n4112) );
  INV_X1 U4656 ( .A(n4110), .ZN(n4111) );
  XNOR2_X1 U4657 ( .A(n4140), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5609)
         );
  INV_X1 U4658 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5803) );
  INV_X1 U4659 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5661) );
  NAND3_X1 U4660 ( .A1(n5803), .A2(n5661), .A3(n5799), .ZN(n4113) );
  OAI21_X1 U4661 ( .B1(n5660), .B2(n4113), .A(n4116), .ZN(n4115) );
  NAND3_X1 U4662 ( .A1(n5660), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4114) );
  NAND2_X1 U4663 ( .A1(n4115), .A2(n4114), .ZN(n4118) );
  NAND2_X1 U4664 ( .A1(n6418), .A2(n5803), .ZN(n4117) );
  NAND2_X1 U4665 ( .A1(n4118), .A2(n4117), .ZN(n5729) );
  XNOR2_X1 U4666 ( .A(n6418), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5731)
         );
  NAND2_X1 U4667 ( .A1(n5729), .A2(n5731), .ZN(n4121) );
  NAND2_X1 U4668 ( .A1(n6418), .A2(n4119), .ZN(n4120) );
  XNOR2_X1 U4669 ( .A(n6418), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5774)
         );
  NAND2_X1 U4670 ( .A1(n5775), .A2(n5774), .ZN(n5773) );
  INV_X1 U4671 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U4672 ( .A1(n6418), .A2(n6699), .ZN(n4122) );
  NAND2_X1 U4673 ( .A1(n5773), .A2(n4122), .ZN(n5821) );
  XNOR2_X1 U4674 ( .A(n6418), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5820)
         );
  NAND2_X1 U4675 ( .A1(n6418), .A2(n6806), .ZN(n4123) );
  INV_X1 U4676 ( .A(n5874), .ZN(n4125) );
  NAND2_X1 U4677 ( .A1(n4125), .A2(n4124), .ZN(n6416) );
  NOR3_X1 U4678 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n4126) );
  NAND2_X1 U4679 ( .A1(n6416), .A2(n4126), .ZN(n4127) );
  NAND2_X1 U4680 ( .A1(n4127), .A2(n4116), .ZN(n4132) );
  NAND2_X1 U4681 ( .A1(n4132), .A2(n4131), .ZN(n4742) );
  INV_X1 U4682 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6487) );
  INV_X1 U4683 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6381) );
  NAND4_X1 U4684 ( .A1(n3798), .A2(n6487), .A3(n6362), .A4(n6381), .ZN(n4133)
         );
  INV_X1 U4685 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6505) );
  INV_X1 U4686 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U4687 ( .A1(n6505), .A2(n6397), .ZN(n6496) );
  NOR2_X1 U4688 ( .A1(n4133), .A2(n6496), .ZN(n4134) );
  NOR2_X1 U4689 ( .A1(n6418), .A2(n4134), .ZN(n4135) );
  NAND2_X1 U4690 ( .A1(n6418), .A2(n6447), .ZN(n6347) );
  NAND2_X1 U4691 ( .A1(n6418), .A2(n6450), .ZN(n4136) );
  AND2_X1 U4692 ( .A1(n6347), .A2(n4136), .ZN(n4138) );
  INV_X1 U4693 ( .A(n4136), .ZN(n4137) );
  XNOR2_X1 U4694 ( .A(n6418), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6350)
         );
  NOR2_X1 U4695 ( .A1(n4116), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6339)
         );
  INV_X1 U4696 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U4697 ( .A1(n6440), .A2(n6451), .ZN(n4153) );
  INV_X1 U4698 ( .A(n4153), .ZN(n4139) );
  OR2_X1 U4699 ( .A1(n4140), .A2(n4139), .ZN(n4141) );
  NAND2_X1 U4700 ( .A1(n4144), .A2(n3693), .ZN(n4802) );
  INV_X1 U4701 ( .A(n4802), .ZN(n6987) );
  AND2_X1 U4702 ( .A1(n4144), .A2(n5946), .ZN(n4985) );
  NOR2_X1 U4703 ( .A1(n6987), .A2(n4985), .ZN(n5940) );
  NAND2_X1 U4704 ( .A1(n3677), .A2(n3436), .ZN(n4773) );
  NAND2_X1 U4705 ( .A1(n4145), .A2(n3649), .ZN(n4146) );
  NAND4_X1 U4706 ( .A1(n5019), .A2(n5940), .A3(n4773), .A4(n4146), .ZN(n4147)
         );
  OAI211_X1 U4709 ( .C1(n4152), .C2(n6441), .A(n4151), .B(n7206), .ZN(U2990)
         );
  NOR2_X1 U4710 ( .A1(n4153), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4154)
         );
  OR2_X1 U4711 ( .A1(n6418), .A2(n4154), .ZN(n4172) );
  XNOR2_X1 U4712 ( .A(n6418), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4156)
         );
  XNOR2_X1 U4713 ( .A(n4157), .B(n4156), .ZN(n5913) );
  OR2_X1 U4714 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4159)
         );
  INV_X1 U4715 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U4716 ( .A1(n3436), .A2(n6082), .ZN(n4158) );
  NAND2_X1 U4717 ( .A1(n4159), .A2(n4158), .ZN(n4732) );
  NAND2_X1 U4718 ( .A1(n4181), .A2(n6082), .ZN(n4160) );
  OAI21_X1 U4719 ( .B1(n4732), .B2(n4181), .A(n4160), .ZN(n4161) );
  NOR2_X1 U4720 ( .A1(n4731), .A2(n4161), .ZN(n4162) );
  AND2_X1 U4721 ( .A1(n6809), .A2(REIP_REG_29__SCAN_IN), .ZN(n5909) );
  INV_X1 U4722 ( .A(n5909), .ZN(n4165) );
  AND2_X1 U4723 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4166) );
  INV_X1 U4724 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4163) );
  NAND3_X1 U4725 ( .A1(n6438), .A2(n4166), .A3(n4163), .ZN(n4164) );
  OAI211_X1 U4726 ( .C1(n6081), .C2(n6799), .A(n4165), .B(n4164), .ZN(n4169)
         );
  NAND2_X1 U4727 ( .A1(n4166), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U4728 ( .A1(n6796), .A2(n6320), .ZN(n4167) );
  NAND2_X1 U4729 ( .A1(n6441), .A2(n4167), .ZN(n6428) );
  NAND2_X1 U4730 ( .A1(n4171), .A2(n4170), .ZN(U2989) );
  NAND4_X1 U4731 ( .A1(n6418), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A4(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n4175) );
  NOR2_X1 U4732 ( .A1(n6418), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4173)
         );
  AND2_X1 U4733 ( .A1(n4173), .A2(n4172), .ZN(n4174) );
  NAND2_X1 U4734 ( .A1(n6340), .A2(n4174), .ZN(n6322) );
  XNOR2_X1 U4735 ( .A(n4177), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6319)
         );
  OR2_X1 U4736 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4180)
         );
  INV_X1 U4737 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U4738 ( .A1(n3436), .A2(n5980), .ZN(n4179) );
  AND2_X1 U4739 ( .A1(n4180), .A2(n4179), .ZN(n4735) );
  NAND2_X1 U4740 ( .A1(n4734), .A2(n4735), .ZN(n4186) );
  NAND2_X1 U4741 ( .A1(n4182), .A2(n4186), .ZN(n4185) );
  INV_X1 U4742 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4787) );
  NOR2_X1 U4743 ( .A1(n5552), .A2(EBX_REG_31__SCAN_IN), .ZN(n4183) );
  AOI21_X1 U4744 ( .B1(n4770), .B2(n4787), .A(n4183), .ZN(n4184) );
  MUX2_X1 U4745 ( .A(n4186), .B(n4185), .S(n4184), .Z(n6079) );
  INV_X1 U4746 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6432) );
  AOI21_X1 U4747 ( .B1(n6796), .B2(n6432), .A(n6428), .ZN(n4188) );
  NAND2_X1 U4748 ( .A1(n6809), .A2(REIP_REG_31__SCAN_IN), .ZN(n6315) );
  INV_X1 U4749 ( .A(n6320), .ZN(n6429) );
  NAND4_X1 U4750 ( .A1(n6438), .A2(n6429), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n4787), .ZN(n4187) );
  OAI211_X1 U4751 ( .C1(n4188), .C2(n4787), .A(n6315), .B(n4187), .ZN(n4189)
         );
  NOR2_X1 U4752 ( .A1(n4190), .A2(n4189), .ZN(n4191) );
  NAND2_X1 U4753 ( .A1(n4192), .A2(n4191), .ZN(U2987) );
  NAND2_X1 U4754 ( .A1(n4938), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4420) );
  NAND2_X1 U4755 ( .A1(n6691), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4568) );
  OAI21_X2 U4756 ( .B1(n5261), .B2(n4420), .A(n4568), .ZN(n4210) );
  NAND2_X1 U4757 ( .A1(n4194), .A2(n4304), .ZN(n4199) );
  INV_X1 U4758 ( .A(n5699), .ZN(n4195) );
  AND2_X1 U4759 ( .A1(n4195), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4221) );
  INV_X1 U4760 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4196) );
  INV_X1 U4761 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5529) );
  OAI22_X1 U4762 ( .A1(n4683), .A2(n4196), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5529), .ZN(n4197) );
  AOI21_X1 U4763 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n4221), .A(n4197), 
        .ZN(n4198) );
  NAND2_X1 U4764 ( .A1(n4199), .A2(n4198), .ZN(n4814) );
  NAND3_X1 U4765 ( .A1(n4906), .A2(n4938), .A3(n5697), .ZN(n4200) );
  NAND2_X1 U4766 ( .A1(n4200), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4797) );
  INV_X1 U4767 ( .A(n4221), .ZN(n4208) );
  NAND2_X1 U4768 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4202)
         );
  NAND2_X1 U4769 ( .A1(n5956), .A2(EAX_REG_0__SCAN_IN), .ZN(n4201) );
  OAI211_X1 U4770 ( .C1(n4208), .C2(n5938), .A(n4202), .B(n4201), .ZN(n4203)
         );
  AOI21_X1 U4771 ( .B1(n5051), .B2(n4304), .A(n4203), .ZN(n4204) );
  INV_X1 U4772 ( .A(n4204), .ZN(n4799) );
  OR2_X1 U4773 ( .A1(n4799), .A2(n5535), .ZN(n4205) );
  AND2_X2 U4774 ( .A1(n4814), .A2(n4815), .ZN(n4209) );
  OR2_X2 U4775 ( .A1(n4210), .A2(n4209), .ZN(n4878) );
  INV_X1 U4776 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5905) );
  OAI21_X1 U4777 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4214), .ZN(n6644) );
  AOI22_X1 U4778 ( .A1(n4721), .A2(n6644), .B1(n5955), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4207) );
  NAND2_X1 U4779 ( .A1(n5956), .A2(EAX_REG_2__SCAN_IN), .ZN(n4206) );
  OAI211_X1 U4780 ( .C1(n4208), .C2(n5905), .A(n4207), .B(n4206), .ZN(n4877)
         );
  NAND2_X1 U4781 ( .A1(n4210), .A2(n4209), .ZN(n4211) );
  INV_X1 U4782 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4217) );
  OAI21_X1 U4783 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4215), .A(n4223), 
        .ZN(n6652) );
  AOI22_X1 U4784 ( .A1(n4721), .A2(n6652), .B1(n5955), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4216) );
  OAI21_X1 U4785 ( .B1(n4683), .B2(n4217), .A(n4216), .ZN(n4218) );
  AOI21_X1 U4786 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n4221), .A(n4218), 
        .ZN(n4219) );
  NAND2_X1 U4787 ( .A1(n4220), .A2(n4219), .ZN(n5435) );
  NAND2_X1 U4788 ( .A1(n4221), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4225) );
  AOI21_X1 U4789 ( .B1(n6832), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4222) );
  AOI21_X1 U4790 ( .B1(n5956), .B2(EAX_REG_4__SCAN_IN), .A(n4222), .ZN(n4224)
         );
  AOI21_X1 U4791 ( .B1(n6832), .B2(n4223), .A(n4229), .ZN(n6836) );
  AOI22_X1 U4792 ( .A1(n4225), .A2(n4224), .B1(n4721), .B2(n6836), .ZN(n4226)
         );
  NOR2_X2 U4793 ( .A1(n5437), .A2(n5029), .ZN(n5028) );
  INV_X1 U4794 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4231) );
  OAI21_X1 U4795 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n4229), .A(n4235), 
        .ZN(n6858) );
  AOI22_X1 U4796 ( .A1(n4721), .A2(n6858), .B1(n5955), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4230) );
  OAI21_X1 U4797 ( .B1(n4683), .B2(n4231), .A(n4230), .ZN(n4232) );
  INV_X1 U4798 ( .A(n4232), .ZN(n4233) );
  NAND2_X1 U4799 ( .A1(n5028), .A2(n5092), .ZN(n5091) );
  INV_X1 U4800 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4238) );
  OAI21_X1 U4801 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n4236), .A(n4242), 
        .ZN(n6869) );
  AOI22_X1 U4802 ( .A1(n4721), .A2(n6869), .B1(n5955), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4237) );
  OAI21_X1 U4803 ( .B1(n4683), .B2(n4238), .A(n4237), .ZN(n4239) );
  OR2_X2 U4804 ( .A1(n5091), .A2(n5336), .ZN(n5444) );
  INV_X1 U4805 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4246) );
  INV_X1 U4806 ( .A(n4242), .ZN(n4244) );
  INV_X1 U4807 ( .A(n4275), .ZN(n4243) );
  OAI21_X1 U4808 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n4244), .A(n4243), 
        .ZN(n6882) );
  AOI22_X1 U4809 ( .A1(n4721), .A2(n6882), .B1(n5955), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4245) );
  OAI21_X1 U4810 ( .B1(n4683), .B2(n4246), .A(n4245), .ZN(n4247) );
  OR2_X2 U4811 ( .A1(n5444), .A2(n5443), .ZN(n5560) );
  NAND2_X1 U4812 ( .A1(n5956), .A2(EAX_REG_8__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U4813 ( .A1(n4700), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U4814 ( .A1(n4706), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U4815 ( .A1(n4708), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U4816 ( .A1(n4666), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4249) );
  NAND4_X1 U4817 ( .A1(n4252), .A2(n4251), .A3(n4250), .A4(n4249), .ZN(n4259)
         );
  AOI22_X1 U4818 ( .A1(n4672), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4600), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U4819 ( .A1(n4697), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U4820 ( .A1(n4699), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U4821 ( .A1(n3422), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4254) );
  NAND4_X1 U4822 ( .A1(n4257), .A2(n4256), .A3(n4255), .A4(n4254), .ZN(n4258)
         );
  NOR2_X1 U4823 ( .A1(n4259), .A2(n4258), .ZN(n4260) );
  OR2_X1 U4824 ( .A1(n4420), .A2(n4260), .ZN(n4262) );
  XNOR2_X1 U4825 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4275), .ZN(n5640) );
  AOI22_X1 U4826 ( .A1(n5955), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4721), 
        .B2(n5640), .ZN(n4261) );
  AOI22_X1 U4827 ( .A1(n4706), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U4828 ( .A1(n4600), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4266) );
  AOI22_X1 U4829 ( .A1(n4645), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4265) );
  AOI22_X1 U4830 ( .A1(n4697), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4264) );
  NAND4_X1 U4831 ( .A1(n4267), .A2(n4266), .A3(n4265), .A4(n4264), .ZN(n4273)
         );
  AOI22_X1 U4832 ( .A1(n3422), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U4833 ( .A1(n4705), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4270) );
  AOI22_X1 U4834 ( .A1(n4708), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4269) );
  AOI22_X1 U4835 ( .A1(n4699), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4268) );
  NAND4_X1 U4836 ( .A1(n4271), .A2(n4270), .A3(n4269), .A4(n4268), .ZN(n4272)
         );
  NOR2_X1 U4837 ( .A1(n4273), .A2(n4272), .ZN(n4274) );
  NOR2_X1 U4838 ( .A1(n4420), .A2(n4274), .ZN(n4362) );
  XNOR2_X1 U4839 ( .A(n4308), .B(n4307), .ZN(n5738) );
  NAND2_X1 U4840 ( .A1(n5738), .A2(n4721), .ZN(n4291) );
  AOI22_X1 U4841 ( .A1(n3422), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4699), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4279) );
  AOI22_X1 U4842 ( .A1(n4700), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4278) );
  AOI22_X1 U4843 ( .A1(n3637), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U4844 ( .A1(n4706), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4276) );
  NAND4_X1 U4845 ( .A1(n4279), .A2(n4278), .A3(n4277), .A4(n4276), .ZN(n4285)
         );
  AOI22_X1 U4846 ( .A1(n4708), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4283) );
  AOI22_X1 U4847 ( .A1(n4697), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4282) );
  AOI22_X1 U4848 ( .A1(n4667), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U4849 ( .A1(n4600), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4280) );
  NAND4_X1 U4850 ( .A1(n4283), .A2(n4282), .A3(n4281), .A4(n4280), .ZN(n4284)
         );
  NOR2_X1 U4851 ( .A1(n4285), .A2(n4284), .ZN(n4288) );
  NAND2_X1 U4852 ( .A1(n5956), .A2(EAX_REG_11__SCAN_IN), .ZN(n4287) );
  NAND2_X1 U4853 ( .A1(n5955), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4286)
         );
  OAI211_X1 U4854 ( .C1(n4420), .C2(n4288), .A(n4287), .B(n4286), .ZN(n4289)
         );
  INV_X1 U4855 ( .A(n4289), .ZN(n4290) );
  NAND2_X1 U4856 ( .A1(n4291), .A2(n4290), .ZN(n5619) );
  XOR2_X1 U4857 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n4292), .Z(n6888) );
  AOI22_X1 U4858 ( .A1(n4700), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U4859 ( .A1(n4672), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U4860 ( .A1(n4666), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4294) );
  AOI22_X1 U4861 ( .A1(n4708), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4293) );
  NAND4_X1 U4862 ( .A1(n4296), .A2(n4295), .A3(n4294), .A4(n4293), .ZN(n4302)
         );
  AOI22_X1 U4863 ( .A1(n4706), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4600), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4300) );
  AOI22_X1 U4864 ( .A1(n3422), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U4865 ( .A1(n4601), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4298) );
  AOI22_X1 U4866 ( .A1(n4699), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4297) );
  NAND4_X1 U4867 ( .A1(n4300), .A2(n4299), .A3(n4298), .A4(n4297), .ZN(n4301)
         );
  OR2_X1 U4868 ( .A1(n4302), .A2(n4301), .ZN(n4303) );
  AOI22_X1 U4869 ( .A1(n4304), .A2(n4303), .B1(n5955), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4306) );
  NAND2_X1 U4870 ( .A1(n5956), .A2(EAX_REG_10__SCAN_IN), .ZN(n4305) );
  OAI211_X1 U4871 ( .C1(n6888), .C2(n5535), .A(n4306), .B(n4305), .ZN(n5618)
         );
  AND2_X1 U4872 ( .A1(n5619), .A2(n5618), .ZN(n5617) );
  XOR2_X1 U4873 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n4337), .Z(n6901) );
  NAND2_X1 U4874 ( .A1(n6901), .A2(n4721), .ZN(n4324) );
  INV_X1 U4875 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4310) );
  OAI21_X1 U4876 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n7028), .A(n6691), 
        .ZN(n4309) );
  OAI21_X1 U4877 ( .B1(n4683), .B2(n4310), .A(n4309), .ZN(n4323) );
  AOI22_X1 U4878 ( .A1(n3422), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4699), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4314) );
  AOI22_X1 U4879 ( .A1(n3638), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4313) );
  AOI22_X1 U4880 ( .A1(n4600), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4312) );
  AOI22_X1 U4881 ( .A1(n4708), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4311) );
  NAND4_X1 U4882 ( .A1(n4314), .A2(n4313), .A3(n4312), .A4(n4311), .ZN(n4320)
         );
  AOI22_X1 U4883 ( .A1(n4666), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4318) );
  AOI22_X1 U4884 ( .A1(n4706), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4317) );
  AOI22_X1 U4885 ( .A1(n4705), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4316) );
  AOI22_X1 U4886 ( .A1(n4700), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4315) );
  NAND4_X1 U4887 ( .A1(n4318), .A2(n4317), .A3(n4316), .A4(n4315), .ZN(n4319)
         );
  NOR2_X1 U4888 ( .A1(n4320), .A2(n4319), .ZN(n4321) );
  NOR2_X1 U4889 ( .A1(n4420), .A2(n4321), .ZN(n4322) );
  AOI21_X1 U4890 ( .B1(n4324), .B2(n4323), .A(n4322), .ZN(n5705) );
  INV_X1 U4891 ( .A(n5705), .ZN(n4325) );
  AND2_X1 U4892 ( .A1(n4362), .A2(n4357), .ZN(n5677) );
  INV_X1 U4893 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U4894 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n3638), .B1(n4706), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4329) );
  AOI22_X1 U4895 ( .A1(n4600), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4328) );
  AOI22_X1 U4896 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n4645), .B1(n4601), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U4897 ( .A1(n4708), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4326) );
  NAND4_X1 U4898 ( .A1(n4329), .A2(n4328), .A3(n4327), .A4(n4326), .ZN(n4335)
         );
  AOI22_X1 U4899 ( .A1(n3422), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4333) );
  AOI22_X1 U4900 ( .A1(n4650), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4332) );
  AOI22_X1 U4901 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n3637), .B1(n3949), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4331) );
  AOI22_X1 U4902 ( .A1(n4699), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4330) );
  NAND4_X1 U4903 ( .A1(n4333), .A2(n4332), .A3(n4331), .A4(n4330), .ZN(n4334)
         );
  NOR2_X1 U4904 ( .A1(n4335), .A2(n4334), .ZN(n4336) );
  OR2_X1 U4905 ( .A1(n4420), .A2(n4336), .ZN(n4339) );
  XNOR2_X1 U4906 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4386), .ZN(n5778)
         );
  AOI22_X1 U4907 ( .A1(n4721), .A2(n5778), .B1(n5955), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4338) );
  OAI211_X1 U4908 ( .C1(n4683), .C2(n4340), .A(n4339), .B(n4338), .ZN(n5681)
         );
  AND2_X1 U4909 ( .A1(n5677), .A2(n5681), .ZN(n4355) );
  AOI22_X1 U4910 ( .A1(n4706), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U4911 ( .A1(n3637), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4343) );
  AOI22_X1 U4912 ( .A1(n4700), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U4913 ( .A1(n4708), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4341) );
  NAND4_X1 U4914 ( .A1(n4344), .A2(n4343), .A3(n4342), .A4(n4341), .ZN(n4350)
         );
  AOI22_X1 U4915 ( .A1(n3422), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4916 ( .A1(n4697), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4347) );
  AOI22_X1 U4917 ( .A1(n4699), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U4918 ( .A1(n4600), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4345) );
  NAND4_X1 U4919 ( .A1(n4348), .A2(n4347), .A3(n4346), .A4(n4345), .ZN(n4349)
         );
  NOR2_X1 U4920 ( .A1(n4350), .A2(n4349), .ZN(n4351) );
  OR2_X1 U4921 ( .A1(n4420), .A2(n4351), .ZN(n4354) );
  XNOR2_X1 U4922 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4352), .ZN(n5613) );
  AOI22_X1 U4923 ( .A1(n4721), .A2(n5613), .B1(n5955), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4353) );
  OAI211_X1 U4924 ( .C1(n4683), .C2(n6540), .A(n4354), .B(n4353), .ZN(n5590)
         );
  AND2_X1 U4925 ( .A1(n4355), .A2(n5590), .ZN(n4356) );
  NAND2_X1 U4926 ( .A1(n5591), .A2(n4356), .ZN(n4370) );
  NOR2_X1 U4927 ( .A1(n5091), .A2(n5336), .ZN(n4361) );
  NAND2_X1 U4928 ( .A1(n4357), .A2(n5590), .ZN(n4358) );
  OR2_X1 U4929 ( .A1(n4358), .A2(n5561), .ZN(n4359) );
  NOR2_X1 U4930 ( .A1(n4359), .A2(n5443), .ZN(n4360) );
  XNOR2_X1 U4931 ( .A(n4363), .B(n4364), .ZN(n6911) );
  NAND2_X1 U4932 ( .A1(n6911), .A2(n4721), .ZN(n4367) );
  OAI22_X1 U4933 ( .A1(n4683), .A2(n6547), .B1(n4568), .B2(n4364), .ZN(n4365)
         );
  INV_X1 U4934 ( .A(n4365), .ZN(n4366) );
  NAND2_X1 U4935 ( .A1(n4367), .A2(n4366), .ZN(n5587) );
  NAND2_X1 U4936 ( .A1(n5586), .A2(n5587), .ZN(n5679) );
  NAND2_X1 U4937 ( .A1(n4368), .A2(n5681), .ZN(n4369) );
  AOI22_X1 U4938 ( .A1(n3422), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U4939 ( .A1(n4708), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U4940 ( .A1(n4645), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4372) );
  AOI22_X1 U4941 ( .A1(n4707), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4371) );
  NAND4_X1 U4942 ( .A1(n4374), .A2(n4373), .A3(n4372), .A4(n4371), .ZN(n4380)
         );
  AOI22_X1 U4943 ( .A1(n4700), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4706), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U4944 ( .A1(n4600), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U4945 ( .A1(n4699), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U4946 ( .A1(n4644), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4375) );
  NAND4_X1 U4947 ( .A1(n4378), .A2(n4377), .A3(n4376), .A4(n4375), .ZN(n4379)
         );
  NOR2_X1 U4948 ( .A1(n4380), .A2(n4379), .ZN(n4385) );
  INV_X1 U4949 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U4950 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4381)
         );
  OAI211_X1 U4951 ( .C1(n4683), .C2(n4382), .A(n5535), .B(n4381), .ZN(n4383)
         );
  INV_X1 U4952 ( .A(n4383), .ZN(n4384) );
  OAI21_X1 U4953 ( .B1(n4686), .B2(n4385), .A(n4384), .ZN(n4389) );
  INV_X1 U4954 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4401) );
  OAI21_X1 U4955 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4387), .A(n4458), 
        .ZN(n6675) );
  OR2_X1 U4956 ( .A1(n5535), .A2(n6675), .ZN(n4388) );
  XNOR2_X1 U4957 ( .A(n4390), .B(n4401), .ZN(n5876) );
  AOI22_X1 U4958 ( .A1(n4706), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4394) );
  AOI22_X1 U4959 ( .A1(n4600), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4393) );
  AOI22_X1 U4960 ( .A1(n4699), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U4961 ( .A1(n4700), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4391) );
  NAND4_X1 U4962 ( .A1(n4394), .A2(n4393), .A3(n4392), .A4(n4391), .ZN(n4400)
         );
  AOI22_X1 U4963 ( .A1(n3422), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4398) );
  AOI22_X1 U4964 ( .A1(n4645), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4397) );
  AOI22_X1 U4965 ( .A1(n4708), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U4966 ( .A1(n3637), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4395) );
  NAND4_X1 U4967 ( .A1(n4398), .A2(n4397), .A3(n4396), .A4(n4395), .ZN(n4399)
         );
  NOR2_X1 U4968 ( .A1(n4400), .A2(n4399), .ZN(n4404) );
  INV_X1 U4969 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4796) );
  OAI22_X1 U4970 ( .A1(n4683), .A2(n4796), .B1(n4568), .B2(n4401), .ZN(n4402)
         );
  INV_X1 U4971 ( .A(n4402), .ZN(n4403) );
  OAI21_X1 U4972 ( .B1(n4686), .B2(n4404), .A(n4403), .ZN(n4405) );
  AOI21_X1 U4973 ( .B1(n5876), .B2(n4721), .A(n4405), .ZN(n5850) );
  XOR2_X1 U4974 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4406), .Z(n5795) );
  INV_X1 U4975 ( .A(n5795), .ZN(n5824) );
  AOI22_X1 U4976 ( .A1(n3422), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U4977 ( .A1(n4708), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U4978 ( .A1(n4697), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4408) );
  AOI22_X1 U4979 ( .A1(n3948), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4407) );
  NAND4_X1 U4980 ( .A1(n4410), .A2(n4409), .A3(n4408), .A4(n4407), .ZN(n4416)
         );
  AOI22_X1 U4981 ( .A1(n4706), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U4982 ( .A1(n4600), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4413) );
  AOI22_X1 U4983 ( .A1(n4699), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4412) );
  AOI22_X1 U4984 ( .A1(n4619), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4411) );
  NAND4_X1 U4985 ( .A1(n4414), .A2(n4413), .A3(n4412), .A4(n4411), .ZN(n4415)
         );
  NOR2_X1 U4986 ( .A1(n4416), .A2(n4415), .ZN(n4419) );
  NAND2_X1 U4987 ( .A1(n5956), .A2(EAX_REG_15__SCAN_IN), .ZN(n4418) );
  NAND2_X1 U4988 ( .A1(n5955), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4417)
         );
  OAI211_X1 U4989 ( .C1(n4420), .C2(n4419), .A(n4418), .B(n4417), .ZN(n4421)
         );
  AOI21_X1 U4990 ( .B1(n5824), .B2(n4721), .A(n4421), .ZN(n5785) );
  NOR2_X1 U4991 ( .A1(n5850), .A2(n5785), .ZN(n5707) );
  INV_X2 U4992 ( .A(n5696), .ZN(n4442) );
  NAND2_X1 U4993 ( .A1(n4686), .A2(n5535), .ZN(n4516) );
  AOI22_X1 U4994 ( .A1(n4708), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4428) );
  NAND2_X1 U4995 ( .A1(n4700), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4424) );
  NAND2_X1 U4996 ( .A1(n4601), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4423) );
  AND3_X1 U4997 ( .A1(n4424), .A2(n4423), .A3(n5535), .ZN(n4427) );
  AOI22_X1 U4998 ( .A1(n4619), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4426) );
  AOI22_X1 U4999 ( .A1(n4666), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4425) );
  NAND4_X1 U5000 ( .A1(n4428), .A2(n4427), .A3(n4426), .A4(n4425), .ZN(n4434)
         );
  AOI22_X1 U5001 ( .A1(n4699), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4706), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U5002 ( .A1(n4672), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4600), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4431) );
  AOI22_X1 U5003 ( .A1(n3948), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U5004 ( .A1(n3422), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4429) );
  NAND4_X1 U5005 ( .A1(n4432), .A2(n4431), .A3(n4430), .A4(n4429), .ZN(n4433)
         );
  OR2_X1 U5006 ( .A1(n4434), .A2(n4433), .ZN(n4435) );
  NAND2_X1 U5007 ( .A1(n4516), .A2(n4435), .ZN(n4439) );
  INV_X1 U5008 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4436) );
  INV_X1 U5009 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6926) );
  OAI22_X1 U5010 ( .A1(n4683), .A2(n4436), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6926), .ZN(n4437) );
  INV_X1 U5011 ( .A(n4437), .ZN(n4438) );
  NAND2_X1 U5012 ( .A1(n4439), .A2(n4438), .ZN(n4441) );
  XNOR2_X1 U5013 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4458), .ZN(n6922)
         );
  NAND2_X1 U5014 ( .A1(n4721), .A2(n6922), .ZN(n4440) );
  NAND2_X2 U5015 ( .A1(n4442), .A2(n3450), .ZN(n5760) );
  AOI22_X1 U5016 ( .A1(n4700), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4446) );
  AOI22_X1 U5017 ( .A1(n4706), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4600), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U5018 ( .A1(n3422), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4444) );
  AOI22_X1 U5019 ( .A1(n4708), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4443) );
  NAND4_X1 U5020 ( .A1(n4446), .A2(n4445), .A3(n4444), .A4(n4443), .ZN(n4452)
         );
  AOI22_X1 U5021 ( .A1(n4672), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4450) );
  AOI22_X1 U5022 ( .A1(n4666), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4644), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4449) );
  AOI22_X1 U5023 ( .A1(n4699), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4448) );
  AOI22_X1 U5024 ( .A1(n4697), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4447) );
  NAND4_X1 U5025 ( .A1(n4450), .A2(n4449), .A3(n4448), .A4(n4447), .ZN(n4451)
         );
  NOR2_X1 U5026 ( .A1(n4452), .A2(n4451), .ZN(n4457) );
  INV_X1 U5027 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U5028 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4453)
         );
  OAI211_X1 U5029 ( .C1(n4683), .C2(n4454), .A(n5535), .B(n4453), .ZN(n4455)
         );
  INV_X1 U5030 ( .A(n4455), .ZN(n4456) );
  OAI21_X1 U5031 ( .B1(n4686), .B2(n4457), .A(n4456), .ZN(n4462) );
  OAI21_X1 U5032 ( .B1(n4460), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n4496), 
        .ZN(n6413) );
  OR2_X1 U5033 ( .A1(n6413), .A2(n5535), .ZN(n4461) );
  NAND2_X1 U5034 ( .A1(n4462), .A2(n4461), .ZN(n5759) );
  AOI22_X1 U5035 ( .A1(n4699), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4468) );
  AOI22_X1 U5036 ( .A1(n4708), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4600), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4467) );
  AOI22_X1 U5037 ( .A1(n4700), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4466) );
  NAND2_X1 U5038 ( .A1(n3949), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U5039 ( .A1(n4707), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4463)
         );
  AND3_X1 U5040 ( .A1(n4464), .A2(n4463), .A3(n5535), .ZN(n4465) );
  NAND4_X1 U5041 ( .A1(n4468), .A2(n4467), .A3(n4466), .A4(n4465), .ZN(n4474)
         );
  AOI22_X1 U5042 ( .A1(n3422), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4706), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U5043 ( .A1(n3637), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4644), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4471) );
  AOI22_X1 U5044 ( .A1(n4697), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4470) );
  AOI22_X1 U5045 ( .A1(n4645), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4469) );
  NAND4_X1 U5046 ( .A1(n4472), .A2(n4471), .A3(n4470), .A4(n4469), .ZN(n4473)
         );
  OR2_X1 U5047 ( .A1(n4474), .A2(n4473), .ZN(n4475) );
  NAND2_X1 U5048 ( .A1(n4516), .A2(n4475), .ZN(n4480) );
  INV_X1 U5049 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4476) );
  INV_X1 U5050 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6400) );
  OAI22_X1 U5051 ( .A1(n4683), .A2(n4476), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6400), .ZN(n4477) );
  INV_X1 U5052 ( .A(n4477), .ZN(n4479) );
  XNOR2_X1 U5053 ( .A(n4496), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6402)
         );
  AND2_X1 U5054 ( .A1(n6402), .A2(n4721), .ZN(n4478) );
  AOI21_X1 U5055 ( .B1(n4480), .B2(n4479), .A(n4478), .ZN(n5828) );
  AOI22_X1 U5056 ( .A1(n3422), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U5057 ( .A1(n4600), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4483) );
  AOI22_X1 U5058 ( .A1(n4697), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4482) );
  AOI22_X1 U5059 ( .A1(n4708), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4481) );
  NAND4_X1 U5060 ( .A1(n4484), .A2(n4483), .A3(n4482), .A4(n4481), .ZN(n4490)
         );
  AOI22_X1 U5061 ( .A1(n4706), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3638), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4488) );
  AOI22_X1 U5062 ( .A1(n4700), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4487) );
  AOI22_X1 U5063 ( .A1(n4666), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4486) );
  AOI22_X1 U5064 ( .A1(n4699), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4485) );
  NAND4_X1 U5065 ( .A1(n4488), .A2(n4487), .A3(n4486), .A4(n4485), .ZN(n4489)
         );
  NOR2_X1 U5066 ( .A1(n4490), .A2(n4489), .ZN(n4495) );
  INV_X1 U5067 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U5068 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4491)
         );
  OAI211_X1 U5069 ( .C1(n4683), .C2(n4492), .A(n5535), .B(n4491), .ZN(n4493)
         );
  INV_X1 U5070 ( .A(n4493), .ZN(n4494) );
  OAI21_X1 U5071 ( .B1(n4686), .B2(n4495), .A(n4494), .ZN(n4502) );
  INV_X1 U5072 ( .A(n4497), .ZN(n4499) );
  INV_X1 U5073 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U5074 ( .A1(n4499), .A2(n4498), .ZN(n4500) );
  NAND2_X1 U5075 ( .A1(n4548), .A2(n4500), .ZN(n6951) );
  NAND2_X2 U5076 ( .A1(n5868), .A2(n5867), .ZN(n5866) );
  NAND2_X1 U5077 ( .A1(n4600), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4504) );
  NAND2_X1 U5078 ( .A1(n4700), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4503) );
  AND3_X1 U5079 ( .A1(n4504), .A2(n4503), .A3(n5535), .ZN(n4508) );
  AOI22_X1 U5080 ( .A1(n4708), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4507) );
  AOI22_X1 U5081 ( .A1(n4667), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U5082 ( .A1(n3638), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4505) );
  NAND4_X1 U5083 ( .A1(n4508), .A2(n4507), .A3(n4506), .A4(n4505), .ZN(n4514)
         );
  AOI22_X1 U5084 ( .A1(n4699), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4706), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4512) );
  AOI22_X1 U5085 ( .A1(n3422), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U5086 ( .A1(n4705), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U5087 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n4601), .B1(n3949), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4509) );
  NAND4_X1 U5088 ( .A1(n4512), .A2(n4511), .A3(n4510), .A4(n4509), .ZN(n4513)
         );
  OR2_X1 U5089 ( .A1(n4514), .A2(n4513), .ZN(n4515) );
  NAND2_X1 U5090 ( .A1(n4516), .A2(n4515), .ZN(n4520) );
  INV_X1 U5091 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4517) );
  INV_X1 U5092 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6384) );
  OAI22_X1 U5093 ( .A1(n4683), .A2(n4517), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6384), .ZN(n4518) );
  INV_X1 U5094 ( .A(n4518), .ZN(n4519) );
  NAND2_X1 U5095 ( .A1(n4520), .A2(n4519), .ZN(n4522) );
  XNOR2_X1 U5096 ( .A(n4548), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6386)
         );
  NAND2_X1 U5097 ( .A1(n6386), .A2(n4721), .ZN(n4521) );
  NAND2_X1 U5098 ( .A1(n4522), .A2(n4521), .ZN(n5883) );
  AOI22_X1 U5099 ( .A1(n4705), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U5100 ( .A1(n3638), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4525) );
  AOI22_X1 U5101 ( .A1(n4708), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4524) );
  AOI22_X1 U5102 ( .A1(n4699), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4523) );
  NAND4_X1 U5103 ( .A1(n4526), .A2(n4525), .A3(n4524), .A4(n4523), .ZN(n4532)
         );
  AOI22_X1 U5104 ( .A1(n3422), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4530) );
  AOI22_X1 U5105 ( .A1(n4706), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4529) );
  AOI22_X1 U5106 ( .A1(n4600), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5107 ( .A1(n4645), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4527) );
  NAND4_X1 U5108 ( .A1(n4530), .A2(n4529), .A3(n4528), .A4(n4527), .ZN(n4531)
         );
  NOR2_X1 U5109 ( .A1(n4532), .A2(n4531), .ZN(n4556) );
  AOI22_X1 U5110 ( .A1(n3422), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4699), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4536) );
  AOI22_X1 U5111 ( .A1(n4708), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5112 ( .A1(n4700), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4534) );
  AOI22_X1 U5113 ( .A1(n4601), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4533) );
  NAND4_X1 U5114 ( .A1(n4536), .A2(n4535), .A3(n4534), .A4(n4533), .ZN(n4542)
         );
  AOI22_X1 U5115 ( .A1(n4600), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4540) );
  AOI22_X1 U5116 ( .A1(n4645), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5117 ( .A1(n4650), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5118 ( .A1(n4706), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4537) );
  NAND4_X1 U5119 ( .A1(n4540), .A2(n4539), .A3(n4538), .A4(n4537), .ZN(n4541)
         );
  NOR2_X1 U5120 ( .A1(n4542), .A2(n4541), .ZN(n4557) );
  XNOR2_X1 U5121 ( .A(n4556), .B(n4557), .ZN(n4547) );
  INV_X1 U5122 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4544) );
  NAND2_X1 U5123 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4543)
         );
  OAI211_X1 U5124 ( .C1(n4683), .C2(n4544), .A(n5535), .B(n4543), .ZN(n4545)
         );
  INV_X1 U5125 ( .A(n4545), .ZN(n4546) );
  OAI21_X1 U5126 ( .B1(n4547), .B2(n4686), .A(n4546), .ZN(n4554) );
  INV_X1 U5127 ( .A(n4550), .ZN(n4551) );
  INV_X1 U5128 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U5129 ( .A1(n4551), .A2(n6070), .ZN(n4552) );
  NAND2_X1 U5130 ( .A1(n4590), .A2(n4552), .ZN(n6376) );
  NAND2_X1 U5131 ( .A1(n4554), .A2(n4553), .ZN(n6063) );
  AND2_X2 U5132 ( .A1(n5881), .A2(n4555), .ZN(n6048) );
  OR2_X1 U5133 ( .A1(n4557), .A2(n4556), .ZN(n4584) );
  AOI22_X1 U5134 ( .A1(n4672), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4600), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4561) );
  AOI22_X1 U5135 ( .A1(n4708), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4706), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5136 ( .A1(n3422), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4559) );
  AOI22_X1 U5137 ( .A1(n4650), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4558) );
  NAND4_X1 U5138 ( .A1(n4561), .A2(n4560), .A3(n4559), .A4(n4558), .ZN(n4567)
         );
  AOI22_X1 U5139 ( .A1(n4699), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5140 ( .A1(n4697), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4644), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4564) );
  AOI22_X1 U5141 ( .A1(n3948), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4563) );
  AOI22_X1 U5142 ( .A1(n4666), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4562) );
  NAND4_X1 U5143 ( .A1(n4565), .A2(n4564), .A3(n4563), .A4(n4562), .ZN(n4566)
         );
  NOR2_X1 U5144 ( .A1(n4567), .A2(n4566), .ZN(n4583) );
  XNOR2_X1 U5145 ( .A(n4584), .B(n4583), .ZN(n4572) );
  INV_X1 U5146 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6056) );
  XNOR2_X1 U5147 ( .A(n4590), .B(n6056), .ZN(n6367) );
  INV_X1 U5148 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4569) );
  OAI22_X1 U5149 ( .A1(n4683), .A2(n4569), .B1(n6056), .B2(n4568), .ZN(n4570)
         );
  AOI21_X1 U5150 ( .B1(n4721), .B2(n6367), .A(n4570), .ZN(n4571) );
  OAI21_X1 U5151 ( .B1(n4572), .B2(n4686), .A(n4571), .ZN(n6047) );
  AOI22_X1 U5152 ( .A1(n3422), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U5153 ( .A1(n4650), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4575) );
  AOI22_X1 U5154 ( .A1(n4666), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5155 ( .A1(n4600), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4573) );
  NAND4_X1 U5156 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(n4582)
         );
  AOI22_X1 U5157 ( .A1(n4708), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4580) );
  AOI22_X1 U5158 ( .A1(n4706), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4579) );
  AOI22_X1 U5159 ( .A1(n4697), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4578) );
  AOI22_X1 U5160 ( .A1(n4699), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4577) );
  NAND4_X1 U5161 ( .A1(n4580), .A2(n4579), .A3(n4578), .A4(n4577), .ZN(n4581)
         );
  NOR2_X1 U5162 ( .A1(n4582), .A2(n4581), .ZN(n4599) );
  OR2_X1 U5163 ( .A1(n4584), .A2(n4583), .ZN(n4598) );
  XNOR2_X1 U5164 ( .A(n4599), .B(n4598), .ZN(n4589) );
  INV_X1 U5165 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4586) );
  NAND2_X1 U5166 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4585)
         );
  OAI211_X1 U5167 ( .C1(n4213), .C2(n4586), .A(n5535), .B(n4585), .ZN(n4587)
         );
  INV_X1 U5168 ( .A(n4587), .ZN(n4588) );
  OAI21_X1 U5169 ( .B1(n4589), .B2(n4686), .A(n4588), .ZN(n4597) );
  INV_X1 U5170 ( .A(n4592), .ZN(n4594) );
  INV_X1 U5171 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4593) );
  NAND2_X1 U5172 ( .A1(n4594), .A2(n4593), .ZN(n4595) );
  NAND2_X1 U5173 ( .A1(n4636), .A2(n4595), .ZN(n6353) );
  NAND2_X2 U5174 ( .A1(n6049), .A2(n6033), .ZN(n6032) );
  NOR2_X1 U5175 ( .A1(n4599), .A2(n4598), .ZN(n4618) );
  AOI22_X1 U5176 ( .A1(n4706), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4605) );
  AOI22_X1 U5177 ( .A1(n4600), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U5178 ( .A1(n4645), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4601), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5179 ( .A1(n4697), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4602) );
  NAND4_X1 U5180 ( .A1(n4605), .A2(n4604), .A3(n4603), .A4(n4602), .ZN(n4611)
         );
  AOI22_X1 U5181 ( .A1(n3422), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4609) );
  AOI22_X1 U5182 ( .A1(n4705), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4608) );
  AOI22_X1 U5183 ( .A1(n4708), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4607) );
  AOI22_X1 U5184 ( .A1(n4699), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4606) );
  NAND4_X1 U5185 ( .A1(n4609), .A2(n4608), .A3(n4607), .A4(n4606), .ZN(n4610)
         );
  OR2_X1 U5186 ( .A1(n4611), .A2(n4610), .ZN(n4617) );
  XNOR2_X1 U5187 ( .A(n4618), .B(n4617), .ZN(n4614) );
  INV_X1 U5188 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U5189 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6024), .A(n5535), .ZN(
        n4612) );
  AOI21_X1 U5190 ( .B1(n5956), .B2(EAX_REG_26__SCAN_IN), .A(n4612), .ZN(n4613)
         );
  OAI21_X1 U5191 ( .B1(n4614), .B2(n4686), .A(n4613), .ZN(n4616) );
  XNOR2_X1 U5192 ( .A(n4636), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6027)
         );
  NAND2_X1 U5193 ( .A1(n6027), .A2(n4721), .ZN(n4615) );
  NAND2_X1 U5194 ( .A1(n4616), .A2(n4615), .ZN(n6019) );
  NAND2_X1 U5195 ( .A1(n4618), .A2(n4617), .ZN(n4642) );
  AOI22_X1 U5196 ( .A1(n3422), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4699), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4623) );
  AOI22_X1 U5197 ( .A1(n4666), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4697), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4622) );
  AOI22_X1 U5198 ( .A1(n4705), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4619), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4621) );
  AOI22_X1 U5199 ( .A1(n4600), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4620) );
  NAND4_X1 U5200 ( .A1(n4623), .A2(n4622), .A3(n4621), .A4(n4620), .ZN(n4630)
         );
  AOI22_X1 U5201 ( .A1(n4708), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5202 ( .A1(n4706), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4627) );
  AOI22_X1 U5203 ( .A1(n4700), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4624), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4626) );
  AOI22_X1 U5204 ( .A1(n4644), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4625) );
  NAND4_X1 U5205 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), .ZN(n4629)
         );
  NOR2_X1 U5206 ( .A1(n4630), .A2(n4629), .ZN(n4643) );
  XNOR2_X1 U5207 ( .A(n4642), .B(n4643), .ZN(n4635) );
  INV_X1 U5208 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U5209 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4631)
         );
  OAI211_X1 U5210 ( .C1(n4213), .C2(n4632), .A(n5535), .B(n4631), .ZN(n4633)
         );
  INV_X1 U5211 ( .A(n4633), .ZN(n4634) );
  OAI21_X1 U5212 ( .B1(n4635), .B2(n4686), .A(n4634), .ZN(n4640) );
  INV_X1 U5213 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U5214 ( .A1(n4637), .A2(n6010), .ZN(n4638) );
  AND2_X1 U5215 ( .A1(n4689), .A2(n4638), .ZN(n6009) );
  NAND2_X1 U5216 ( .A1(n6009), .A2(n4721), .ZN(n4639) );
  NAND2_X1 U5217 ( .A1(n4640), .A2(n4639), .ZN(n6007) );
  AND2_X2 U5218 ( .A1(n6004), .A2(n4641), .ZN(n6006) );
  NOR2_X1 U5219 ( .A1(n4643), .A2(n4642), .ZN(n4680) );
  AOI22_X1 U5220 ( .A1(n4706), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4672), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4649) );
  AOI22_X1 U5221 ( .A1(n4600), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4648) );
  AOI22_X1 U5222 ( .A1(n4645), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4644), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4647) );
  AOI22_X1 U5223 ( .A1(n4697), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4646) );
  NAND4_X1 U5224 ( .A1(n4649), .A2(n4648), .A3(n4647), .A4(n4646), .ZN(n4656)
         );
  AOI22_X1 U5225 ( .A1(n3422), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4654) );
  AOI22_X1 U5226 ( .A1(n4650), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4653) );
  AOI22_X1 U5227 ( .A1(n4708), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4652) );
  AOI22_X1 U5228 ( .A1(n4699), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4651) );
  NAND4_X1 U5229 ( .A1(n4654), .A2(n4653), .A3(n4652), .A4(n4651), .ZN(n4655)
         );
  OR2_X1 U5230 ( .A1(n4656), .A2(n4655), .ZN(n4679) );
  INV_X1 U5231 ( .A(n4679), .ZN(n4657) );
  XNOR2_X1 U5232 ( .A(n4680), .B(n4657), .ZN(n4658) );
  INV_X1 U5233 ( .A(n4686), .ZN(n4717) );
  NAND2_X1 U5234 ( .A1(n4658), .A2(n4717), .ZN(n4664) );
  INV_X1 U5235 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U5236 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4659)
         );
  OAI211_X1 U5237 ( .C1(n4213), .C2(n4660), .A(n5535), .B(n4659), .ZN(n4661)
         );
  INV_X1 U5238 ( .A(n4661), .ZN(n4663) );
  XNOR2_X1 U5239 ( .A(n4689), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5997)
         );
  AOI21_X1 U5240 ( .B1(n4664), .B2(n4663), .A(n4662), .ZN(n5920) );
  AOI22_X1 U5241 ( .A1(n3422), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4700), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4671) );
  AOI22_X1 U5242 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4666), .B1(n4697), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4670) );
  AOI22_X1 U5243 ( .A1(n4699), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4669) );
  AOI22_X1 U5244 ( .A1(n3637), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4668) );
  NAND4_X1 U5245 ( .A1(n4671), .A2(n4670), .A3(n4669), .A4(n4668), .ZN(n4678)
         );
  AOI22_X1 U5246 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4708), .B1(n4672), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U5247 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n4600), .B1(n4706), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4675) );
  AOI22_X1 U5248 ( .A1(n4705), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5249 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n4601), .B1(n3949), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4673) );
  NAND4_X1 U5250 ( .A1(n4676), .A2(n4675), .A3(n4674), .A4(n4673), .ZN(n4677)
         );
  NOR2_X1 U5251 ( .A1(n4678), .A2(n4677), .ZN(n4696) );
  NAND2_X1 U5252 ( .A1(n4680), .A2(n4679), .ZN(n4695) );
  XNOR2_X1 U5253 ( .A(n4696), .B(n4695), .ZN(n4687) );
  INV_X1 U5254 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4682) );
  NAND2_X1 U5255 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4681)
         );
  OAI211_X1 U5256 ( .C1(n4683), .C2(n4682), .A(n5535), .B(n4681), .ZN(n4684)
         );
  INV_X1 U5257 ( .A(n4684), .ZN(n4685) );
  OAI21_X1 U5258 ( .B1(n4687), .B2(n4686), .A(n4685), .ZN(n4694) );
  INV_X1 U5259 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4688) );
  NAND2_X1 U5260 ( .A1(n4690), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5538)
         );
  INV_X1 U5261 ( .A(n4690), .ZN(n4691) );
  INV_X1 U5262 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U5263 ( .A1(n4691), .A2(n5988), .ZN(n4692) );
  NAND2_X1 U5264 ( .A1(n5538), .A2(n4692), .ZN(n5987) );
  NAND2_X1 U5265 ( .A1(n4694), .A2(n4693), .ZN(n5908) );
  NOR2_X2 U5266 ( .A1(n5919), .A2(n5908), .ZN(n5958) );
  NOR2_X1 U5267 ( .A1(n4696), .A2(n4695), .ZN(n4716) );
  AOI22_X1 U5268 ( .A1(n3638), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3948), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5269 ( .A1(n4697), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4644), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4703) );
  AOI22_X1 U5270 ( .A1(n4699), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4698), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4702) );
  AOI22_X1 U5271 ( .A1(n4700), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4701) );
  NAND4_X1 U5272 ( .A1(n4704), .A2(n4703), .A3(n4702), .A4(n4701), .ZN(n4714)
         );
  AOI22_X1 U5273 ( .A1(n3422), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4705), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4712) );
  AOI22_X1 U5274 ( .A1(n4600), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4706), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U5275 ( .A1(n4708), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4707), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4710) );
  AOI22_X1 U5276 ( .A1(n4666), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3949), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4709) );
  NAND4_X1 U5277 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4713)
         );
  NOR2_X1 U5278 ( .A1(n4714), .A2(n4713), .ZN(n4715) );
  XNOR2_X1 U5279 ( .A(n4716), .B(n4715), .ZN(n4718) );
  NAND2_X1 U5280 ( .A1(n4718), .A2(n4717), .ZN(n4724) );
  OAI21_X1 U5281 ( .B1(n7028), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6691), 
        .ZN(n4719) );
  OAI21_X1 U5282 ( .B1(n4213), .B2(n4942), .A(n4719), .ZN(n4720) );
  INV_X1 U5283 ( .A(n4720), .ZN(n4723) );
  XNOR2_X1 U5284 ( .A(n5538), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6324)
         );
  AOI21_X1 U5285 ( .B1(n4724), .B2(n4723), .A(n4722), .ZN(n5957) );
  NAND2_X1 U5286 ( .A1(n5942), .A2(n7004), .ZN(n4726) );
  INV_X1 U5287 ( .A(n5697), .ZN(n6288) );
  NAND4_X1 U5288 ( .A1(n3675), .A2(n6288), .A3(n4978), .A4(n7004), .ZN(n4898)
         );
  INV_X1 U5289 ( .A(n4898), .ZN(n4728) );
  NAND3_X1 U5290 ( .A1(n4728), .A2(n4727), .A3(n3436), .ZN(n4729) );
  INV_X1 U5291 ( .A(n4731), .ZN(n4733) );
  OAI22_X1 U5292 ( .A1(n4734), .A2(n3435), .B1(n4733), .B2(n4732), .ZN(n4736)
         );
  XNOR2_X1 U5293 ( .A(n4736), .B(n4735), .ZN(n6427) );
  XNOR2_X1 U5294 ( .A(n6418), .B(n6505), .ZN(n6409) );
  OR2_X2 U5295 ( .A1(n6410), .A2(n6409), .ZN(n6407) );
  NOR2_X1 U5296 ( .A1(n6418), .A2(n6397), .ZN(n6358) );
  OAI22_X1 U5297 ( .A1(n6407), .A2(n6358), .B1(n4116), .B2(n4743), .ZN(n4744)
         );
  XNOR2_X1 U5298 ( .A(n6418), .B(n6487), .ZN(n6357) );
  XNOR2_X1 U5299 ( .A(n4744), .B(n6357), .ZN(n6395) );
  NOR2_X1 U5300 ( .A1(n6395), .A2(n6800), .ZN(n4753) );
  NOR2_X1 U5301 ( .A1(n4745), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4752)
         );
  NOR2_X1 U5302 ( .A1(n4746), .A2(n6487), .ZN(n4751) );
  NAND2_X1 U5303 ( .A1(n5831), .A2(n4748), .ZN(n4749) );
  NAND2_X1 U5304 ( .A1(n5885), .A2(n4749), .ZN(n6944) );
  NAND2_X1 U5305 ( .A1(n6809), .A2(REIP_REG_21__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U5306 ( .B1(n6944), .B2(n6799), .A(n6392), .ZN(n4750) );
  OR4_X1 U5307 ( .A1(n4753), .A2(n4752), .A3(n4751), .A4(n4750), .ZN(U2997) );
  AND2_X1 U5308 ( .A1(n5947), .A2(n7004), .ZN(n4754) );
  NAND2_X1 U5309 ( .A1(n5948), .A2(n4754), .ZN(n4757) );
  INV_X1 U5310 ( .A(n4757), .ZN(n4756) );
  INV_X1 U5311 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7050) );
  INV_X1 U5312 ( .A(n3425), .ZN(n5949) );
  INV_X1 U5313 ( .A(n5596), .ZN(n6678) );
  OAI211_X1 U5314 ( .C1(n4756), .C2(n7050), .A(n4761), .B(n6678), .ZN(U2788)
         );
  NOR2_X1 U5315 ( .A1(n5596), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4760) );
  NAND3_X1 U5316 ( .A1(n6694), .A2(n4758), .A3(n5547), .ZN(n4759) );
  OAI21_X1 U5317 ( .B1(n6694), .B2(n4760), .A(n4759), .ZN(U3474) );
  INV_X1 U5318 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4765) );
  INV_X2 U5319 ( .A(n4820), .ZN(n4835) );
  OR2_X1 U5320 ( .A1(n4763), .A2(n4835), .ZN(n4833) );
  INV_X1 U5321 ( .A(DATAI_15_), .ZN(n6213) );
  INV_X1 U5322 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4764) );
  OAI222_X1 U5323 ( .A1(n4765), .A2(n4833), .B1(n4902), .B2(n6213), .C1(n4764), 
        .C2(n4820), .ZN(U2954) );
  OAI21_X1 U5324 ( .B1(n4766), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n5528), 
        .ZN(n4808) );
  INV_X1 U5325 ( .A(n6714), .ZN(n4767) );
  NAND2_X1 U5326 ( .A1(n4767), .A2(n5749), .ZN(n4768) );
  NAND2_X1 U5327 ( .A1(n5752), .A2(n6702), .ZN(n6715) );
  AOI22_X1 U5328 ( .A1(n4768), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n6745), 
        .B2(n6715), .ZN(n4772) );
  AOI21_X1 U5329 ( .B1(n4770), .B2(n6745), .A(n4769), .ZN(n5556) );
  AND2_X1 U5330 ( .A1(n6809), .A2(REIP_REG_0__SCAN_IN), .ZN(n4809) );
  AOI21_X1 U5331 ( .B1(n6826), .B2(n5556), .A(n4809), .ZN(n4771) );
  OAI211_X1 U5332 ( .C1(n6800), .C2(n4808), .A(n4772), .B(n4771), .ZN(U3018)
         );
  AOI21_X1 U5333 ( .B1(n4773), .B2(n6684), .A(READY_N), .ZN(n4774) );
  OAI211_X1 U5334 ( .C1(n3677), .C2(n6969), .A(n7017), .B(n4774), .ZN(n4778)
         );
  INV_X1 U5335 ( .A(n4775), .ZN(n4776) );
  NAND3_X1 U5336 ( .A1(n4778), .A2(n4777), .A3(n4776), .ZN(n4784) );
  NAND2_X1 U5337 ( .A1(n7017), .A2(n4985), .ZN(n4781) );
  OR2_X1 U5338 ( .A1(n5019), .A2(n4779), .ZN(n4780) );
  NAND2_X1 U5339 ( .A1(n4781), .A2(n4780), .ZN(n4900) );
  INV_X1 U5340 ( .A(n5942), .ZN(n4782) );
  NOR2_X1 U5341 ( .A1(n7017), .A2(n4782), .ZN(n4783) );
  NAND2_X1 U5342 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n4915) );
  INV_X1 U5343 ( .A(n4915), .ZN(n7007) );
  NAND2_X1 U5344 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7007), .ZN(n7013) );
  INV_X1 U5345 ( .A(n7013), .ZN(n5024) );
  AOI22_X1 U5346 ( .A1(n7004), .A2(n6968), .B1(FLUSH_REG_SCAN_IN), .B2(n5024), 
        .ZN(n6966) );
  NAND2_X1 U5347 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n7020), .ZN(n7012) );
  NAND2_X1 U5348 ( .A1(n6966), .A2(n7012), .ZN(n6964) );
  NOR2_X1 U5349 ( .A1(n4786), .A2(n4785), .ZN(n4791) );
  INV_X1 U5350 ( .A(n4791), .ZN(n4792) );
  AOI22_X1 U5351 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n6726), .B1(
        INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n4787), .ZN(n5899) );
  NOR2_X1 U5352 ( .A1(n7011), .A2(n6745), .ZN(n5933) );
  NAND2_X1 U5353 ( .A1(n4789), .A2(n5927), .ZN(n4790) );
  NAND2_X1 U5354 ( .A1(n6969), .A2(n3519), .ZN(n4999) );
  OAI211_X1 U5355 ( .C1(n4791), .C2(n3622), .A(n4790), .B(n4999), .ZN(n6967)
         );
  AOI222_X1 U5356 ( .A1(n5934), .A2(n4792), .B1(n5899), .B2(n5933), .C1(n6967), 
        .C2(n7003), .ZN(n4794) );
  NAND2_X1 U5357 ( .A1(n6959), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4793) );
  OAI21_X1 U5358 ( .B1(n6959), .B2(n4794), .A(n4793), .ZN(U3460) );
  NAND2_X1 U5359 ( .A1(n4858), .A2(DATAI_0_), .ZN(n4860) );
  INV_X2 U5360 ( .A(n4833), .ZN(n4839) );
  NAND2_X1 U5361 ( .A1(n4839), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4795) );
  OAI211_X1 U5362 ( .C1(n4820), .C2(n4796), .A(n4860), .B(n4795), .ZN(U2924)
         );
  INV_X1 U5363 ( .A(n4797), .ZN(n4800) );
  OAI21_X1 U5364 ( .B1(n4800), .B2(n4799), .A(n4798), .ZN(n5559) );
  NOR2_X1 U5365 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7011), .ZN(n5533) );
  NAND2_X1 U5366 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5533), .ZN(n6689) );
  INV_X1 U5367 ( .A(n6689), .ZN(n4801) );
  NAND2_X1 U5368 ( .A1(n7066), .A2(n4801), .ZN(n6426) );
  INV_X1 U5369 ( .A(n7066), .ZN(n7112) );
  NAND2_X1 U5370 ( .A1(n7112), .A2(n4803), .ZN(n6695) );
  NAND2_X1 U5371 ( .A1(n6695), .A2(n7020), .ZN(n4804) );
  AND2_X2 U5372 ( .A1(n6952), .A2(n4804), .ZN(n6669) );
  NAND2_X1 U5373 ( .A1(n7020), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4806) );
  NAND2_X1 U5374 ( .A1(n7028), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4805) );
  AND2_X1 U5375 ( .A1(n4806), .A2(n4805), .ZN(n5519) );
  INV_X1 U5376 ( .A(n5519), .ZN(n4807) );
  OAI21_X1 U5377 ( .B1(n6669), .B2(n4807), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4812) );
  INV_X1 U5378 ( .A(n4808), .ZN(n4810) );
  AOI21_X1 U5379 ( .B1(n6671), .B2(n4810), .A(n4809), .ZN(n4811) );
  OAI211_X1 U5380 ( .C1(n5559), .C2(n6426), .A(n4812), .B(n4811), .ZN(U2986)
         );
  INV_X1 U5381 ( .A(n4209), .ZN(n4813) );
  OAI21_X1 U5382 ( .B1(n4815), .B2(n4814), .A(n4813), .ZN(n5585) );
  XNOR2_X1 U5383 ( .A(n4816), .B(n3436), .ZN(n6718) );
  AOI22_X1 U5384 ( .A1(n4738), .A2(n6718), .B1(EBX_REG_1__SCAN_IN), .B2(n6281), 
        .ZN(n4817) );
  OAI21_X1 U5385 ( .B1(n5585), .B2(n6283), .A(n4817), .ZN(U2858) );
  INV_X1 U5386 ( .A(n6969), .ZN(n4995) );
  OR2_X1 U5387 ( .A1(n4818), .A2(n4995), .ZN(n4819) );
  NAND2_X1 U5388 ( .A1(n4820), .A2(n4819), .ZN(n4822) );
  INV_X1 U5389 ( .A(n6684), .ZN(n4821) );
  NAND2_X1 U5390 ( .A1(n6524), .A2(n3685), .ZN(n4953) );
  AOI22_X1 U5391 ( .A1(n6696), .A2(UWORD_REG_6__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4823) );
  OAI21_X1 U5392 ( .B1(n4517), .B2(n4953), .A(n4823), .ZN(U2901) );
  AOI22_X1 U5393 ( .A1(n6696), .A2(UWORD_REG_8__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4824) );
  OAI21_X1 U5394 ( .B1(n4569), .B2(n4953), .A(n4824), .ZN(U2899) );
  AOI22_X1 U5395 ( .A1(n6696), .A2(UWORD_REG_5__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4825) );
  OAI21_X1 U5396 ( .B1(n4492), .B2(n4953), .A(n4825), .ZN(U2902) );
  AOI22_X1 U5397 ( .A1(n6696), .A2(UWORD_REG_9__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4826) );
  OAI21_X1 U5398 ( .B1(n4586), .B2(n4953), .A(n4826), .ZN(U2898) );
  AOI22_X1 U5399 ( .A1(n6696), .A2(UWORD_REG_7__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4827) );
  OAI21_X1 U5400 ( .B1(n4544), .B2(n4953), .A(n4827), .ZN(U2900) );
  AOI22_X1 U5401 ( .A1(n4839), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n4835), .ZN(n4828) );
  NAND2_X1 U5402 ( .A1(n4858), .A2(DATAI_5_), .ZN(n4840) );
  NAND2_X1 U5403 ( .A1(n4828), .A2(n4840), .ZN(U2929) );
  AOI22_X1 U5404 ( .A1(n4839), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n4835), .ZN(n4829) );
  NAND2_X1 U5405 ( .A1(n4858), .A2(DATAI_3_), .ZN(n4848) );
  NAND2_X1 U5406 ( .A1(n4829), .A2(n4848), .ZN(U2927) );
  AOI22_X1 U5407 ( .A1(n4839), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n4835), .ZN(n4830) );
  NAND2_X1 U5408 ( .A1(n4858), .A2(DATAI_1_), .ZN(n4866) );
  NAND2_X1 U5409 ( .A1(n4830), .A2(n4866), .ZN(U2925) );
  AOI22_X1 U5410 ( .A1(n4839), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n4835), .ZN(n4831) );
  NAND2_X1 U5411 ( .A1(n4858), .A2(DATAI_2_), .ZN(n4842) );
  NAND2_X1 U5412 ( .A1(n4831), .A2(n4842), .ZN(U2926) );
  AOI22_X1 U5413 ( .A1(n4839), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n4835), .ZN(n4832) );
  INV_X1 U5414 ( .A(DATAI_4_), .ZN(n5433) );
  OR2_X1 U5415 ( .A1(n4902), .A2(n5433), .ZN(n4856) );
  NAND2_X1 U5416 ( .A1(n4832), .A2(n4856), .ZN(U2928) );
  AOI22_X1 U5417 ( .A1(n4839), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n4835), .ZN(n4834) );
  NAND2_X1 U5418 ( .A1(n4858), .A2(DATAI_14_), .ZN(n4874) );
  NAND2_X1 U5419 ( .A1(n4834), .A2(n4874), .ZN(U2953) );
  AOI22_X1 U5420 ( .A1(n4839), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n4835), .ZN(n4836) );
  NAND2_X1 U5421 ( .A1(n4858), .A2(DATAI_8_), .ZN(n4854) );
  NAND2_X1 U5422 ( .A1(n4836), .A2(n4854), .ZN(U2947) );
  AOI22_X1 U5423 ( .A1(n4839), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n4835), .ZN(n4837) );
  NAND2_X1 U5424 ( .A1(n4858), .A2(DATAI_13_), .ZN(n4844) );
  NAND2_X1 U5425 ( .A1(n4837), .A2(n4844), .ZN(U2952) );
  AOI22_X1 U5426 ( .A1(n4839), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n4835), .ZN(n4838) );
  INV_X1 U5427 ( .A(DATAI_11_), .ZN(n5648) );
  OR2_X1 U5428 ( .A1(n4902), .A2(n5648), .ZN(n4868) );
  NAND2_X1 U5429 ( .A1(n4838), .A2(n4868), .ZN(U2950) );
  AOI22_X1 U5430 ( .A1(n4839), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n4835), .ZN(n4841) );
  NAND2_X1 U5431 ( .A1(n4841), .A2(n4840), .ZN(U2944) );
  AOI22_X1 U5432 ( .A1(n4839), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n4835), .ZN(n4843) );
  NAND2_X1 U5433 ( .A1(n4843), .A2(n4842), .ZN(U2941) );
  AOI22_X1 U5434 ( .A1(n4839), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n4835), .ZN(n4845) );
  NAND2_X1 U5435 ( .A1(n4845), .A2(n4844), .ZN(U2937) );
  AOI22_X1 U5436 ( .A1(n4839), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n4835), .ZN(n4846) );
  NAND2_X1 U5437 ( .A1(n4858), .A2(DATAI_9_), .ZN(n4852) );
  NAND2_X1 U5438 ( .A1(n4846), .A2(n4852), .ZN(U2948) );
  AOI22_X1 U5439 ( .A1(n4839), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n4835), .ZN(n4847) );
  NAND2_X1 U5440 ( .A1(n4858), .A2(DATAI_6_), .ZN(n4862) );
  NAND2_X1 U5441 ( .A1(n4847), .A2(n4862), .ZN(U2945) );
  AOI22_X1 U5442 ( .A1(n4839), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n4835), .ZN(n4849) );
  NAND2_X1 U5443 ( .A1(n4849), .A2(n4848), .ZN(U2942) );
  AOI22_X1 U5444 ( .A1(n4839), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n4835), .ZN(n4850) );
  INV_X1 U5445 ( .A(DATAI_10_), .ZN(n5659) );
  OR2_X1 U5446 ( .A1(n4902), .A2(n5659), .ZN(n4872) );
  NAND2_X1 U5447 ( .A1(n4850), .A2(n4872), .ZN(U2949) );
  AOI22_X1 U5448 ( .A1(n4839), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n4835), .ZN(n4851) );
  NAND2_X1 U5449 ( .A1(n4858), .A2(DATAI_7_), .ZN(n4864) );
  NAND2_X1 U5450 ( .A1(n4851), .A2(n4864), .ZN(U2946) );
  AOI22_X1 U5451 ( .A1(n4839), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n4835), .ZN(n4853) );
  NAND2_X1 U5452 ( .A1(n4853), .A2(n4852), .ZN(U2933) );
  AOI22_X1 U5453 ( .A1(n4839), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n4835), .ZN(n4855) );
  NAND2_X1 U5454 ( .A1(n4855), .A2(n4854), .ZN(U2932) );
  AOI22_X1 U5455 ( .A1(n4839), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n4835), .ZN(n4857) );
  NAND2_X1 U5456 ( .A1(n4857), .A2(n4856), .ZN(U2943) );
  AOI22_X1 U5457 ( .A1(n4839), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n4835), .ZN(n4859) );
  NAND2_X1 U5458 ( .A1(n4858), .A2(DATAI_12_), .ZN(n4870) );
  NAND2_X1 U5459 ( .A1(n4859), .A2(n4870), .ZN(U2936) );
  AOI22_X1 U5460 ( .A1(n4839), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n4835), .ZN(n4861) );
  NAND2_X1 U5461 ( .A1(n4861), .A2(n4860), .ZN(U2939) );
  AOI22_X1 U5462 ( .A1(n4839), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n4835), .ZN(n4863) );
  NAND2_X1 U5463 ( .A1(n4863), .A2(n4862), .ZN(U2930) );
  AOI22_X1 U5464 ( .A1(n4839), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n4835), .ZN(n4865) );
  NAND2_X1 U5465 ( .A1(n4865), .A2(n4864), .ZN(U2931) );
  AOI22_X1 U5466 ( .A1(n4839), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n4835), .ZN(n4867) );
  NAND2_X1 U5467 ( .A1(n4867), .A2(n4866), .ZN(U2940) );
  AOI22_X1 U5468 ( .A1(n4839), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n4835), .ZN(n4869) );
  NAND2_X1 U5469 ( .A1(n4869), .A2(n4868), .ZN(U2935) );
  AOI22_X1 U5470 ( .A1(n4839), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n4835), .ZN(n4871) );
  NAND2_X1 U5471 ( .A1(n4871), .A2(n4870), .ZN(U2951) );
  AOI22_X1 U5472 ( .A1(n4839), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n4835), .ZN(n4873) );
  NAND2_X1 U5473 ( .A1(n4873), .A2(n4872), .ZN(U2934) );
  AOI22_X1 U5474 ( .A1(n4839), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n4835), .ZN(n4875) );
  NAND2_X1 U5475 ( .A1(n4875), .A2(n4874), .ZN(U2938) );
  NOR2_X1 U5476 ( .A1(n4878), .A2(n4877), .ZN(n4879) );
  NOR2_X1 U5477 ( .A1(n4876), .A2(n4879), .ZN(n6641) );
  INV_X1 U5478 ( .A(n6641), .ZN(n5658) );
  OR2_X1 U5479 ( .A1(n4881), .A2(n4880), .ZN(n4882) );
  AND2_X1 U5480 ( .A1(n4882), .A2(n5670), .ZN(n6746) );
  AOI22_X1 U5481 ( .A1(n4738), .A2(n6746), .B1(n6281), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4883) );
  OAI21_X1 U5482 ( .B1(n5658), .B2(n6283), .A(n4883), .ZN(U2857) );
  INV_X1 U5483 ( .A(n5556), .ZN(n4884) );
  OAI222_X1 U5484 ( .A1(n4884), .A2(n6629), .B1(n6636), .B2(n3726), .C1(n5559), 
        .C2(n6283), .ZN(U2859) );
  XNOR2_X1 U5485 ( .A(n4885), .B(n4886), .ZN(n5570) );
  AND2_X1 U5486 ( .A1(n5743), .A2(n6744), .ZN(n4888) );
  INV_X1 U5487 ( .A(n6749), .ZN(n6763) );
  OAI21_X1 U5488 ( .B1(n6743), .B2(n5752), .A(n6763), .ZN(n6729) );
  OAI21_X1 U5489 ( .B1(n4889), .B2(n6744), .A(n5752), .ZN(n6757) );
  NAND2_X1 U5490 ( .A1(n6743), .A2(n6757), .ZN(n6735) );
  AOI21_X1 U5491 ( .B1(n4891), .B2(n4890), .A(n6735), .ZN(n4892) );
  NAND2_X1 U5492 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5044) );
  AOI22_X1 U5493 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n6729), .B1(n4892), 
        .B2(n5044), .ZN(n4897) );
  AOI21_X1 U5494 ( .B1(n3737), .B2(n5669), .A(n4893), .ZN(n4895) );
  INV_X1 U5495 ( .A(n5040), .ZN(n4894) );
  NOR2_X1 U5496 ( .A1(n4895), .A2(n4894), .ZN(n6830) );
  INV_X1 U5497 ( .A(n6809), .ZN(n6818) );
  NOR2_X1 U5498 ( .A1(n6818), .A2(n6840), .ZN(n5567) );
  AOI21_X1 U5499 ( .B1(n6826), .B2(n6830), .A(n5567), .ZN(n4896) );
  OAI211_X1 U5500 ( .C1(n5570), .C2(n6800), .A(n4897), .B(n4896), .ZN(U3014)
         );
  NOR2_X1 U5501 ( .A1(n3821), .A2(n4898), .ZN(n4899) );
  INV_X1 U5502 ( .A(DATAI_0_), .ZN(n6177) );
  INV_X1 U5503 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6526) );
  OAI222_X1 U5504 ( .A1(n5559), .A2(n3421), .B1(n5816), .B2(n6177), .C1(n6287), 
        .C2(n6526), .ZN(U2891) );
  INV_X1 U5505 ( .A(DATAI_1_), .ZN(n6089) );
  OAI222_X1 U5506 ( .A1(n5585), .A2(n3421), .B1(n5816), .B2(n6089), .C1(n6287), 
        .C2(n4196), .ZN(U2890) );
  INV_X2 U5507 ( .A(n6426), .ZN(n6670) );
  AND2_X1 U5508 ( .A1(n6670), .A2(DATAI_19_), .ZN(n7146) );
  INV_X1 U5509 ( .A(n7146), .ZN(n5473) );
  NOR2_X1 U5510 ( .A1(n5298), .A2(n4906), .ZN(n4907) );
  NAND3_X1 U5511 ( .A1(n5300), .A2(n5262), .A3(n4907), .ZN(n5426) );
  NOR2_X1 U5512 ( .A1(n7083), .A2(n5929), .ZN(n7105) );
  INV_X1 U5513 ( .A(n4789), .ZN(n5099) );
  OR2_X1 U5514 ( .A1(n4911), .A2(n5099), .ZN(n5456) );
  NOR2_X1 U5515 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7098) );
  INV_X1 U5516 ( .A(n7098), .ZN(n4912) );
  NOR2_X1 U5517 ( .A1(n6972), .A2(n4912), .ZN(n4980) );
  AOI21_X1 U5518 ( .B1(n7105), .B2(n7084), .A(n4980), .ZN(n4919) );
  INV_X1 U5519 ( .A(n4919), .ZN(n4917) );
  INV_X1 U5520 ( .A(n5298), .ZN(n4913) );
  NAND2_X1 U5521 ( .A1(n5300), .A2(n4913), .ZN(n4914) );
  NAND2_X1 U5522 ( .A1(n5262), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5032) );
  OAI21_X1 U5523 ( .B1(n4914), .B2(n5032), .A(n7066), .ZN(n4918) );
  NAND2_X1 U5524 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7098), .ZN(n5450) );
  INV_X1 U5525 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U5526 ( .A1(n6691), .A2(n7011), .ZN(n7015) );
  OAI21_X1 U5527 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n7089), .A(n5161), 
        .ZN(n7073) );
  AOI21_X1 U5528 ( .B1(n7112), .B2(n5450), .A(n7073), .ZN(n4916) );
  OAI21_X1 U5529 ( .B1(n4917), .B2(n4918), .A(n4916), .ZN(n4977) );
  NAND2_X1 U5530 ( .A1(DATAI_3_), .A2(n5161), .ZN(n7150) );
  OAI22_X1 U5531 ( .A1(n4919), .A2(n4918), .B1(n6691), .B2(n5450), .ZN(n4976)
         );
  AOI22_X1 U5532 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n4977), .B1(n5476), 
        .B2(n4976), .ZN(n4924) );
  NOR2_X2 U5533 ( .A1(n4979), .A2(n4921), .ZN(n7145) );
  NOR2_X1 U5534 ( .A1(n5298), .A2(n7077), .ZN(n4922) );
  AND2_X1 U5535 ( .A1(n4922), .A2(n5300), .ZN(n5447) );
  NAND2_X1 U5536 ( .A1(n6670), .A2(DATAI_27_), .ZN(n5479) );
  INV_X1 U5537 ( .A(n5479), .ZN(n7147) );
  AOI22_X1 U5538 ( .A1(n7145), .A2(n4980), .B1(n5447), .B2(n7147), .ZN(n4923)
         );
  OAI211_X1 U5539 ( .C1(n5473), .C2(n5426), .A(n4924), .B(n4923), .ZN(U3047)
         );
  AND2_X1 U5540 ( .A1(n6670), .A2(DATAI_18_), .ZN(n7136) );
  INV_X1 U5541 ( .A(n7136), .ZN(n5466) );
  NAND2_X1 U5542 ( .A1(DATAI_2_), .A2(n5161), .ZN(n7140) );
  AOI22_X1 U5543 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n4977), .B1(n5469), 
        .B2(n4976), .ZN(n4927) );
  NOR2_X2 U5544 ( .A1(n4979), .A2(n4925), .ZN(n7135) );
  NAND2_X1 U5545 ( .A1(n6670), .A2(DATAI_26_), .ZN(n5472) );
  INV_X1 U5546 ( .A(n5472), .ZN(n7137) );
  AOI22_X1 U5547 ( .A1(n7135), .A2(n4980), .B1(n5447), .B2(n7137), .ZN(n4926)
         );
  OAI211_X1 U5548 ( .C1(n5466), .C2(n5426), .A(n4927), .B(n4926), .ZN(U3046)
         );
  AND2_X1 U5549 ( .A1(n6670), .A2(DATAI_17_), .ZN(n7127) );
  INV_X1 U5550 ( .A(n7127), .ZN(n5487) );
  NAND2_X1 U5551 ( .A1(DATAI_1_), .A2(n5161), .ZN(n7130) );
  AOI22_X1 U5552 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4977), .B1(n5490), 
        .B2(n4976), .ZN(n4930) );
  NOR2_X2 U5553 ( .A1(n4979), .A2(n4928), .ZN(n7125) );
  NAND2_X1 U5554 ( .A1(n6670), .A2(DATAI_25_), .ZN(n5493) );
  INV_X1 U5555 ( .A(n5493), .ZN(n7126) );
  AOI22_X1 U5556 ( .A1(n7125), .A2(n4980), .B1(n5447), .B2(n7126), .ZN(n4929)
         );
  OAI211_X1 U5557 ( .C1(n5487), .C2(n5426), .A(n4930), .B(n4929), .ZN(U3045)
         );
  AND2_X1 U5558 ( .A1(n6670), .A2(DATAI_23_), .ZN(n7199) );
  INV_X1 U5559 ( .A(n7199), .ZN(n5501) );
  NAND2_X1 U5560 ( .A1(DATAI_7_), .A2(n5161), .ZN(n7203) );
  AOI22_X1 U5561 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n4977), .B1(n5504), 
        .B2(n4976), .ZN(n4932) );
  NOR2_X2 U5562 ( .A1(n4979), .A2(n6288), .ZN(n7195) );
  NAND2_X1 U5563 ( .A1(n6670), .A2(DATAI_31_), .ZN(n5507) );
  INV_X1 U5564 ( .A(n5507), .ZN(n7196) );
  AOI22_X1 U5565 ( .A1(n7195), .A2(n4980), .B1(n5447), .B2(n7196), .ZN(n4931)
         );
  OAI211_X1 U5566 ( .C1(n5501), .C2(n5426), .A(n4932), .B(n4931), .ZN(U3051)
         );
  AND2_X1 U5567 ( .A1(n6670), .A2(DATAI_21_), .ZN(n7166) );
  INV_X1 U5568 ( .A(n7166), .ZN(n5494) );
  NAND2_X1 U5569 ( .A1(DATAI_5_), .A2(n5161), .ZN(n7170) );
  AOI22_X1 U5570 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n4977), .B1(n5497), 
        .B2(n4976), .ZN(n4934) );
  NOR2_X2 U5571 ( .A1(n4979), .A2(n3625), .ZN(n7165) );
  NAND2_X1 U5572 ( .A1(n6670), .A2(DATAI_29_), .ZN(n5500) );
  INV_X1 U5573 ( .A(n5500), .ZN(n7167) );
  AOI22_X1 U5574 ( .A1(n7165), .A2(n4980), .B1(n5447), .B2(n7167), .ZN(n4933)
         );
  OAI211_X1 U5575 ( .C1(n5494), .C2(n5426), .A(n4934), .B(n4933), .ZN(U3049)
         );
  AND2_X1 U5576 ( .A1(n6670), .A2(DATAI_16_), .ZN(n7110) );
  INV_X1 U5577 ( .A(n7110), .ZN(n5459) );
  NAND2_X1 U5578 ( .A1(DATAI_0_), .A2(n5161), .ZN(n7120) );
  AOI22_X1 U5579 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n4977), .B1(n5462), 
        .B2(n4976), .ZN(n4937) );
  NOR2_X2 U5580 ( .A1(n4979), .A2(n4935), .ZN(n7109) );
  NAND2_X1 U5581 ( .A1(n6670), .A2(DATAI_24_), .ZN(n5465) );
  INV_X1 U5582 ( .A(n5465), .ZN(n7117) );
  AOI22_X1 U5583 ( .A1(n7109), .A2(n4980), .B1(n5447), .B2(n7117), .ZN(n4936)
         );
  OAI211_X1 U5584 ( .C1(n5459), .C2(n5426), .A(n4937), .B(n4936), .ZN(U3044)
         );
  AND2_X1 U5585 ( .A1(n6670), .A2(DATAI_22_), .ZN(n7177) );
  INV_X1 U5586 ( .A(n7177), .ZN(n5509) );
  NAND2_X1 U5587 ( .A1(DATAI_6_), .A2(n5161), .ZN(n7180) );
  AOI22_X1 U5588 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n4977), .B1(n5515), 
        .B2(n4976), .ZN(n4940) );
  NOR2_X2 U5589 ( .A1(n4979), .A2(n4938), .ZN(n7175) );
  NAND2_X1 U5590 ( .A1(n6670), .A2(DATAI_30_), .ZN(n5518) );
  INV_X1 U5591 ( .A(n5518), .ZN(n7176) );
  AOI22_X1 U5592 ( .A1(n7175), .A2(n4980), .B1(n5447), .B2(n7176), .ZN(n4939)
         );
  OAI211_X1 U5593 ( .C1(n5509), .C2(n5426), .A(n4940), .B(n4939), .ZN(U3050)
         );
  INV_X1 U5594 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4942) );
  AOI22_X1 U5595 ( .A1(n6696), .A2(UWORD_REG_14__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4941) );
  OAI21_X1 U5596 ( .B1(n4942), .B2(n4953), .A(n4941), .ZN(U2893) );
  AOI22_X1 U5597 ( .A1(n6696), .A2(UWORD_REG_0__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4943) );
  OAI21_X1 U5598 ( .B1(n4796), .B2(n4953), .A(n4943), .ZN(U2907) );
  AOI22_X1 U5599 ( .A1(n6696), .A2(UWORD_REG_1__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4944) );
  OAI21_X1 U5600 ( .B1(n4382), .B2(n4953), .A(n4944), .ZN(U2906) );
  AOI22_X1 U5601 ( .A1(n6696), .A2(UWORD_REG_2__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4945) );
  OAI21_X1 U5602 ( .B1(n4436), .B2(n4953), .A(n4945), .ZN(U2905) );
  AOI22_X1 U5603 ( .A1(n6696), .A2(UWORD_REG_3__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4946) );
  OAI21_X1 U5604 ( .B1(n4454), .B2(n4953), .A(n4946), .ZN(U2904) );
  AOI22_X1 U5605 ( .A1(n6696), .A2(UWORD_REG_4__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4947) );
  OAI21_X1 U5606 ( .B1(n4476), .B2(n4953), .A(n4947), .ZN(U2903) );
  INV_X1 U5607 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4949) );
  AOI22_X1 U5608 ( .A1(n6696), .A2(UWORD_REG_10__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4948) );
  OAI21_X1 U5609 ( .B1(n4949), .B2(n4953), .A(n4948), .ZN(U2897) );
  AOI22_X1 U5610 ( .A1(n6696), .A2(UWORD_REG_11__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4950) );
  OAI21_X1 U5611 ( .B1(n4632), .B2(n4953), .A(n4950), .ZN(U2896) );
  AOI22_X1 U5612 ( .A1(n6696), .A2(UWORD_REG_12__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4951) );
  OAI21_X1 U5613 ( .B1(n4660), .B2(n4953), .A(n4951), .ZN(U2895) );
  AOI22_X1 U5614 ( .A1(n6696), .A2(UWORD_REG_13__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4952) );
  OAI21_X1 U5615 ( .B1(n4682), .B2(n4953), .A(n4952), .ZN(U2894) );
  NOR2_X1 U5616 ( .A1(n5261), .A2(n4954), .ZN(n5097) );
  NAND2_X1 U5617 ( .A1(n5097), .A2(n5262), .ZN(n4961) );
  INV_X1 U5618 ( .A(n4961), .ZN(n4955) );
  NOR2_X1 U5619 ( .A1(n5261), .A2(n5032), .ZN(n5048) );
  NAND2_X1 U5620 ( .A1(n5048), .A2(n5053), .ZN(n5047) );
  NAND2_X1 U5621 ( .A1(n5047), .A2(n7066), .ZN(n4959) );
  AND2_X1 U5622 ( .A1(n4911), .A2(n4789), .ZN(n5166) );
  INV_X1 U5623 ( .A(n4956), .ZN(n5088) );
  AOI21_X1 U5624 ( .B1(n7105), .B2(n5166), .A(n5088), .ZN(n4960) );
  INV_X1 U5625 ( .A(n4960), .ZN(n4958) );
  INV_X1 U5626 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7068) );
  NAND3_X1 U5627 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7068), .ZN(n5160) );
  AOI21_X1 U5628 ( .B1(n7112), .B2(n5160), .A(n7073), .ZN(n4957) );
  OAI21_X1 U5629 ( .B1(n4959), .B2(n4958), .A(n4957), .ZN(n5087) );
  OAI22_X1 U5630 ( .A1(n4960), .A2(n4959), .B1(n6691), .B2(n5160), .ZN(n5086)
         );
  AOI22_X1 U5631 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5087), .B1(n5469), 
        .B2(n5086), .ZN(n4963) );
  NOR2_X2 U5632 ( .A1(n4961), .A2(n7077), .ZN(n5190) );
  AOI22_X1 U5633 ( .A1(n5190), .A2(n7137), .B1(n5088), .B2(n7135), .ZN(n4962)
         );
  OAI211_X1 U5634 ( .C1(n5466), .C2(n5384), .A(n4963), .B(n4962), .ZN(U3078)
         );
  AOI22_X1 U5635 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5087), .B1(n5476), 
        .B2(n5086), .ZN(n4965) );
  AOI22_X1 U5636 ( .A1(n5190), .A2(n7147), .B1(n5088), .B2(n7145), .ZN(n4964)
         );
  OAI211_X1 U5637 ( .C1(n5473), .C2(n5384), .A(n4965), .B(n4964), .ZN(U3079)
         );
  AOI22_X1 U5638 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5087), .B1(n5497), 
        .B2(n5086), .ZN(n4967) );
  AOI22_X1 U5639 ( .A1(n5190), .A2(n7167), .B1(n5088), .B2(n7165), .ZN(n4966)
         );
  OAI211_X1 U5640 ( .C1(n5494), .C2(n5384), .A(n4967), .B(n4966), .ZN(U3081)
         );
  AOI22_X1 U5641 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5087), .B1(n5515), 
        .B2(n5086), .ZN(n4969) );
  AOI22_X1 U5642 ( .A1(n5190), .A2(n7176), .B1(n5088), .B2(n7175), .ZN(n4968)
         );
  OAI211_X1 U5643 ( .C1(n5509), .C2(n5384), .A(n4969), .B(n4968), .ZN(U3082)
         );
  AOI22_X1 U5644 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5087), .B1(n5504), 
        .B2(n5086), .ZN(n4971) );
  AOI22_X1 U5645 ( .A1(n5190), .A2(n7196), .B1(n5088), .B2(n7195), .ZN(n4970)
         );
  OAI211_X1 U5646 ( .C1(n5501), .C2(n5384), .A(n4971), .B(n4970), .ZN(U3083)
         );
  AOI22_X1 U5647 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5087), .B1(n5462), 
        .B2(n5086), .ZN(n4973) );
  AOI22_X1 U5648 ( .A1(n5190), .A2(n7117), .B1(n5088), .B2(n7109), .ZN(n4972)
         );
  OAI211_X1 U5649 ( .C1(n5459), .C2(n5384), .A(n4973), .B(n4972), .ZN(U3076)
         );
  AOI22_X1 U5650 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5087), .B1(n5490), 
        .B2(n5086), .ZN(n4975) );
  AOI22_X1 U5651 ( .A1(n5190), .A2(n7126), .B1(n5088), .B2(n7125), .ZN(n4974)
         );
  OAI211_X1 U5652 ( .C1(n5487), .C2(n5384), .A(n4975), .B(n4974), .ZN(U3077)
         );
  AND2_X1 U5653 ( .A1(n6670), .A2(DATAI_20_), .ZN(n7157) );
  INV_X1 U5654 ( .A(n7157), .ZN(n5480) );
  NAND2_X1 U5655 ( .A1(DATAI_4_), .A2(n5161), .ZN(n7160) );
  AOI22_X1 U5656 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4977), .B1(n5483), 
        .B2(n4976), .ZN(n4982) );
  NOR2_X2 U5657 ( .A1(n4979), .A2(n4978), .ZN(n7155) );
  NAND2_X1 U5658 ( .A1(n6670), .A2(DATAI_28_), .ZN(n5486) );
  INV_X1 U5659 ( .A(n5486), .ZN(n7156) );
  AOI22_X1 U5660 ( .A1(n7155), .A2(n4980), .B1(n5447), .B2(n7156), .ZN(n4981)
         );
  OAI211_X1 U5661 ( .C1(n5480), .C2(n5426), .A(n4982), .B(n4981), .ZN(U3048)
         );
  XNOR2_X1 U5662 ( .A(n5261), .B(n5032), .ZN(n5027) );
  NAND2_X1 U5663 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4984) );
  INV_X1 U5664 ( .A(n4984), .ZN(n4983) );
  MUX2_X1 U5665 ( .A(n4984), .B(n4983), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4996) );
  OR2_X1 U5666 ( .A1(n5942), .A2(n4985), .ZN(n5005) );
  MUX2_X1 U5667 ( .A(n4987), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5902), 
        .Z(n4988) );
  NOR2_X1 U5668 ( .A1(n4988), .A2(n5011), .ZN(n4989) );
  NAND2_X1 U5669 ( .A1(n5005), .A2(n4989), .ZN(n4994) );
  INV_X1 U5670 ( .A(n5002), .ZN(n4992) );
  NAND2_X1 U5671 ( .A1(n5902), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U5672 ( .A1(n4990), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U5673 ( .A1(n3905), .A2(n4991), .ZN(n6954) );
  NAND2_X1 U5674 ( .A1(n4992), .A2(n6954), .ZN(n4993) );
  OAI211_X1 U5675 ( .C1(n4996), .C2(n4995), .A(n4994), .B(n4993), .ZN(n4997)
         );
  AOI21_X1 U5676 ( .B1(n7083), .B2(n5927), .A(n4997), .ZN(n6958) );
  NAND2_X1 U5677 ( .A1(n6968), .A2(n6958), .ZN(n4998) );
  OAI21_X1 U5678 ( .B1(n6968), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n4998), 
        .ZN(n6982) );
  INV_X1 U5679 ( .A(n6982), .ZN(n5009) );
  NAND2_X1 U5680 ( .A1(n4911), .A2(n5927), .ZN(n5007) );
  XNOR2_X1 U5681 ( .A(n5902), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5004)
         );
  NAND2_X1 U5682 ( .A1(n6969), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5000) );
  MUX2_X1 U5683 ( .A(n5000), .B(n4999), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n5001) );
  OAI21_X1 U5684 ( .B1(n5004), .B2(n5002), .A(n5001), .ZN(n5003) );
  AOI21_X1 U5685 ( .B1(n5005), .B2(n5004), .A(n5003), .ZN(n5006) );
  NAND2_X1 U5686 ( .A1(n5007), .A2(n5006), .ZN(n5900) );
  NAND2_X1 U5687 ( .A1(n6968), .A2(n5900), .ZN(n5008) );
  OAI21_X1 U5688 ( .B1(n6968), .B2(n5905), .A(n5008), .ZN(n6979) );
  NAND3_X1 U5689 ( .A1(n5009), .A2(n7011), .A3(n6979), .ZN(n5013) );
  NOR2_X1 U5690 ( .A1(FLUSH_REG_SCAN_IN), .A2(n7011), .ZN(n5010) );
  NAND2_X1 U5691 ( .A1(n5011), .A2(n5010), .ZN(n5012) );
  NAND2_X1 U5692 ( .A1(n5013), .A2(n5012), .ZN(n6994) );
  INV_X1 U5693 ( .A(n5014), .ZN(n5022) );
  MUX2_X1 U5694 ( .A(n6968), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n5021) );
  INV_X1 U5695 ( .A(n5015), .ZN(n5016) );
  NOR2_X1 U5696 ( .A1(n5017), .A2(n5016), .ZN(n5018) );
  XNOR2_X1 U5697 ( .A(n5018), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6961)
         );
  INV_X1 U5698 ( .A(n5019), .ZN(n6962) );
  NAND2_X1 U5699 ( .A1(n6962), .A2(n7011), .ZN(n5020) );
  OAI22_X1 U5700 ( .A1(n5021), .A2(n3553), .B1(n6961), .B2(n5020), .ZN(n6993)
         );
  AOI21_X1 U5701 ( .B1(n6994), .B2(n5022), .A(n6993), .ZN(n5914) );
  INV_X1 U5702 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5023) );
  NAND2_X1 U5703 ( .A1(n5914), .A2(n5023), .ZN(n5025) );
  AOI21_X1 U5704 ( .B1(n5025), .B2(n5024), .A(n5161), .ZN(n6521) );
  NOR2_X1 U5705 ( .A1(n6521), .A2(n7112), .ZN(n5916) );
  INV_X1 U5706 ( .A(n5916), .ZN(n5026) );
  AOI21_X1 U5707 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n7089), .A(n6521), .ZN(
        n5031) );
  INV_X1 U5708 ( .A(n5031), .ZN(n5918) );
  INV_X1 U5709 ( .A(n4911), .ZN(n5649) );
  INV_X1 U5710 ( .A(n6521), .ZN(n5035) );
  OAI222_X1 U5711 ( .A1(n5027), .A2(n5026), .B1(n5918), .B2(n5649), .C1(n6978), 
        .C2(n5035), .ZN(U3463) );
  CLKBUF_X1 U5712 ( .A(n5028), .Z(n5093) );
  AOI21_X1 U5713 ( .B1(n5029), .B2(n5437), .A(n5093), .ZN(n6837) );
  INV_X1 U5714 ( .A(n6837), .ZN(n5434) );
  AOI22_X1 U5715 ( .A1(n4738), .A2(n6830), .B1(n6281), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n5030) );
  OAI21_X1 U5716 ( .B1(n5434), .B2(n6283), .A(n5030), .ZN(U2855) );
  NAND2_X1 U5717 ( .A1(n5031), .A2(n4789), .ZN(n5034) );
  OAI211_X1 U5718 ( .C1(n5262), .C2(STATEBS16_REG_SCAN_IN), .A(n5916), .B(
        n5032), .ZN(n5033) );
  OAI211_X1 U5719 ( .C1(n5035), .C2(n7099), .A(n5034), .B(n5033), .ZN(U3464)
         );
  CLKBUF_X1 U5720 ( .A(n5036), .Z(n5037) );
  XNOR2_X1 U5721 ( .A(n5037), .B(n5038), .ZN(n5524) );
  CLKBUF_X1 U5722 ( .A(n5039), .Z(n5439) );
  AOI21_X1 U5723 ( .B1(n5041), .B2(n5040), .A(n5439), .ZN(n6846) );
  INV_X1 U5724 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6851) );
  NOR2_X1 U5725 ( .A1(n6818), .A2(n6851), .ZN(n5520) );
  AOI21_X1 U5726 ( .B1(n6796), .B2(n5042), .A(n6749), .ZN(n6742) );
  AOI221_X1 U5727 ( .B1(n5044), .B2(n5043), .C1(n6735), .C2(n5043), .A(n6742), 
        .ZN(n5045) );
  AOI211_X1 U5728 ( .C1(n6826), .C2(n6846), .A(n5520), .B(n5045), .ZN(n5046)
         );
  OAI21_X1 U5729 ( .B1(n6800), .B2(n5524), .A(n5046), .ZN(U3013) );
  INV_X1 U5730 ( .A(n7083), .ZN(n5672) );
  OAI21_X1 U5731 ( .B1(n5048), .B2(n5300), .A(n5047), .ZN(n5049) );
  AOI22_X1 U5732 ( .A1(n5916), .A2(n5049), .B1(n6521), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5050) );
  OAI21_X1 U5733 ( .B1(n5918), .B2(n5672), .A(n5050), .ZN(U3462) );
  INV_X1 U5734 ( .A(n7073), .ZN(n7116) );
  AND2_X1 U5735 ( .A1(n7083), .A2(n5051), .ZN(n7067) );
  NOR2_X1 U5736 ( .A1(n5052), .A2(n7068), .ZN(n5080) );
  AOI21_X1 U5737 ( .B1(n7067), .B2(n5166), .A(n5080), .ZN(n5057) );
  NOR2_X1 U5738 ( .A1(n5261), .A2(n5053), .ZN(n5196) );
  NAND2_X1 U5739 ( .A1(n5196), .A2(n5262), .ZN(n5058) );
  INV_X1 U5740 ( .A(n5058), .ZN(n5054) );
  NOR2_X1 U5741 ( .A1(n7112), .A2(STATEBS16_REG_SCAN_IN), .ZN(n7081) );
  INV_X1 U5742 ( .A(n7081), .ZN(n7101) );
  OAI21_X1 U5743 ( .B1(n5054), .B2(n6426), .A(n7101), .ZN(n5055) );
  NAND3_X1 U5744 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5223) );
  AOI22_X1 U5745 ( .A1(n5057), .A2(n5055), .B1(n7112), .B2(n5223), .ZN(n5056)
         );
  INV_X1 U5746 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5061) );
  OAI22_X1 U5747 ( .A1(n5057), .A2(n7112), .B1(n5223), .B2(n6691), .ZN(n5081)
         );
  AOI22_X1 U5748 ( .A1(n5462), .A2(n5081), .B1(n7109), .B2(n5080), .ZN(n5060)
         );
  NOR2_X2 U5749 ( .A1(n5058), .A2(n7077), .ZN(n5256) );
  AOI22_X1 U5750 ( .A1(n7117), .A2(n5256), .B1(n5127), .B2(n7110), .ZN(n5059)
         );
  OAI211_X1 U5751 ( .C1(n5085), .C2(n5061), .A(n5060), .B(n5059), .ZN(U3140)
         );
  INV_X1 U5752 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5064) );
  AOI22_X1 U5753 ( .A1(n5469), .A2(n5081), .B1(n7135), .B2(n5080), .ZN(n5063)
         );
  AOI22_X1 U5754 ( .A1(n7137), .A2(n5256), .B1(n5127), .B2(n7136), .ZN(n5062)
         );
  OAI211_X1 U5755 ( .C1(n5085), .C2(n5064), .A(n5063), .B(n5062), .ZN(U3142)
         );
  INV_X1 U5756 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5067) );
  AOI22_X1 U5757 ( .A1(n5490), .A2(n5081), .B1(n7125), .B2(n5080), .ZN(n5066)
         );
  AOI22_X1 U5758 ( .A1(n7126), .A2(n5256), .B1(n5127), .B2(n7127), .ZN(n5065)
         );
  OAI211_X1 U5759 ( .C1(n5085), .C2(n5067), .A(n5066), .B(n5065), .ZN(U3141)
         );
  INV_X1 U5760 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5070) );
  AOI22_X1 U5761 ( .A1(n5497), .A2(n5081), .B1(n7165), .B2(n5080), .ZN(n5069)
         );
  AOI22_X1 U5762 ( .A1(n7167), .A2(n5256), .B1(n5127), .B2(n7166), .ZN(n5068)
         );
  OAI211_X1 U5763 ( .C1(n5085), .C2(n5070), .A(n5069), .B(n5068), .ZN(U3145)
         );
  INV_X1 U5764 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5073) );
  AOI22_X1 U5765 ( .A1(n5476), .A2(n5081), .B1(n7145), .B2(n5080), .ZN(n5072)
         );
  AOI22_X1 U5766 ( .A1(n7147), .A2(n5256), .B1(n5127), .B2(n7146), .ZN(n5071)
         );
  OAI211_X1 U5767 ( .C1(n5085), .C2(n5073), .A(n5072), .B(n5071), .ZN(U3143)
         );
  INV_X1 U5768 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5076) );
  AOI22_X1 U5769 ( .A1(n5504), .A2(n5081), .B1(n7195), .B2(n5080), .ZN(n5075)
         );
  AOI22_X1 U5770 ( .A1(n7196), .A2(n5256), .B1(n5127), .B2(n7199), .ZN(n5074)
         );
  OAI211_X1 U5771 ( .C1(n5085), .C2(n5076), .A(n5075), .B(n5074), .ZN(U3147)
         );
  INV_X1 U5772 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5079) );
  AOI22_X1 U5773 ( .A1(n5515), .A2(n5081), .B1(n7175), .B2(n5080), .ZN(n5078)
         );
  AOI22_X1 U5774 ( .A1(n7176), .A2(n5256), .B1(n5127), .B2(n7177), .ZN(n5077)
         );
  OAI211_X1 U5775 ( .C1(n5085), .C2(n5079), .A(n5078), .B(n5077), .ZN(U3146)
         );
  INV_X1 U5776 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5084) );
  AOI22_X1 U5777 ( .A1(n5483), .A2(n5081), .B1(n7155), .B2(n5080), .ZN(n5083)
         );
  AOI22_X1 U5778 ( .A1(n7156), .A2(n5256), .B1(n5127), .B2(n7157), .ZN(n5082)
         );
  OAI211_X1 U5779 ( .C1(n5085), .C2(n5084), .A(n5083), .B(n5082), .ZN(U3144)
         );
  AOI22_X1 U5780 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5087), .B1(n5483), 
        .B2(n5086), .ZN(n5090) );
  AOI22_X1 U5781 ( .A1(n5190), .A2(n7156), .B1(n5088), .B2(n7155), .ZN(n5089)
         );
  OAI211_X1 U5782 ( .C1(n5480), .C2(n5384), .A(n5090), .B(n5089), .ZN(U3080)
         );
  OR2_X1 U5783 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  AND2_X1 U5784 ( .A1(n5091), .A2(n5094), .ZN(n6855) );
  INV_X1 U5785 ( .A(n6855), .ZN(n5096) );
  AOI22_X1 U5786 ( .A1(n4738), .A2(n6846), .B1(n6281), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n5095) );
  OAI21_X1 U5787 ( .B1(n5096), .B2(n6283), .A(n5095), .ZN(U2854) );
  INV_X1 U5788 ( .A(DATAI_5_), .ZN(n6184) );
  OAI222_X1 U5789 ( .A1(n5096), .A2(n3421), .B1(n5816), .B2(n6184), .C1(n6287), 
        .C2(n4231), .ZN(U2886) );
  NAND2_X1 U5790 ( .A1(n5097), .A2(n5299), .ZN(n5104) );
  OR2_X1 U5791 ( .A1(n5104), .A2(n7028), .ZN(n5098) );
  AND2_X1 U5792 ( .A1(n5098), .A2(n7066), .ZN(n5101) );
  AND2_X1 U5793 ( .A1(n4911), .A2(n5099), .ZN(n5400) );
  NAND3_X1 U5794 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7068), .A3(n7099), .ZN(n5390) );
  NOR2_X1 U5795 ( .A1(n7103), .A2(n5390), .ZN(n5121) );
  AOI21_X1 U5796 ( .B1(n7105), .B2(n5400), .A(n5121), .ZN(n5103) );
  AOI22_X1 U5797 ( .A1(n5101), .A2(n5103), .B1(n7112), .B2(n5390), .ZN(n5100)
         );
  NAND2_X1 U5798 ( .A1(n7116), .A2(n5100), .ZN(n5120) );
  INV_X1 U5799 ( .A(n5101), .ZN(n5102) );
  OAI22_X1 U5800 ( .A1(n5103), .A2(n5102), .B1(n6691), .B2(n5390), .ZN(n5119)
         );
  AOI22_X1 U5801 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5120), .B1(n5490), 
        .B2(n5119), .ZN(n5106) );
  AOI22_X1 U5802 ( .A1(n5394), .A2(n7126), .B1(n7125), .B2(n5121), .ZN(n5105)
         );
  OAI211_X1 U5803 ( .C1(n5487), .C2(n5158), .A(n5106), .B(n5105), .ZN(U3061)
         );
  AOI22_X1 U5804 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5120), .B1(n5504), 
        .B2(n5119), .ZN(n5108) );
  AOI22_X1 U5805 ( .A1(n5394), .A2(n7196), .B1(n7195), .B2(n5121), .ZN(n5107)
         );
  OAI211_X1 U5806 ( .C1(n5501), .C2(n5158), .A(n5108), .B(n5107), .ZN(U3067)
         );
  AOI22_X1 U5807 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5120), .B1(n5462), 
        .B2(n5119), .ZN(n5110) );
  AOI22_X1 U5808 ( .A1(n5394), .A2(n7117), .B1(n7109), .B2(n5121), .ZN(n5109)
         );
  OAI211_X1 U5809 ( .C1(n5459), .C2(n5158), .A(n5110), .B(n5109), .ZN(U3060)
         );
  AOI22_X1 U5810 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5120), .B1(n5515), 
        .B2(n5119), .ZN(n5112) );
  AOI22_X1 U5811 ( .A1(n5394), .A2(n7176), .B1(n7175), .B2(n5121), .ZN(n5111)
         );
  OAI211_X1 U5812 ( .C1(n5509), .C2(n5158), .A(n5112), .B(n5111), .ZN(U3066)
         );
  AOI22_X1 U5813 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5120), .B1(n5476), 
        .B2(n5119), .ZN(n5114) );
  AOI22_X1 U5814 ( .A1(n5394), .A2(n7147), .B1(n7145), .B2(n5121), .ZN(n5113)
         );
  OAI211_X1 U5815 ( .C1(n5473), .C2(n5158), .A(n5114), .B(n5113), .ZN(U3063)
         );
  AOI22_X1 U5816 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5120), .B1(n5469), 
        .B2(n5119), .ZN(n5116) );
  AOI22_X1 U5817 ( .A1(n5394), .A2(n7137), .B1(n7135), .B2(n5121), .ZN(n5115)
         );
  OAI211_X1 U5818 ( .C1(n5466), .C2(n5158), .A(n5116), .B(n5115), .ZN(U3062)
         );
  AOI22_X1 U5819 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5120), .B1(n5483), 
        .B2(n5119), .ZN(n5118) );
  AOI22_X1 U5820 ( .A1(n5394), .A2(n7156), .B1(n7155), .B2(n5121), .ZN(n5117)
         );
  OAI211_X1 U5821 ( .C1(n5480), .C2(n5158), .A(n5118), .B(n5117), .ZN(U3064)
         );
  AOI22_X1 U5822 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5120), .B1(n5497), 
        .B2(n5119), .ZN(n5123) );
  AOI22_X1 U5823 ( .A1(n5394), .A2(n7167), .B1(n7165), .B2(n5121), .ZN(n5122)
         );
  OAI211_X1 U5824 ( .C1(n5494), .C2(n5158), .A(n5123), .B(n5122), .ZN(U3065)
         );
  NAND3_X1 U5825 ( .A1(n7099), .A2(n7103), .A3(n7098), .ZN(n5130) );
  INV_X1 U5826 ( .A(n5348), .ZN(n5301) );
  OR2_X1 U5827 ( .A1(n5347), .A2(n5301), .ZN(n5402) );
  AND2_X1 U5828 ( .A1(n5402), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U5829 ( .A1(n5128), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U5830 ( .A1(n5161), .A2(n5401), .ZN(n7091) );
  AOI211_X1 U5831 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5130), .A(n5392), .B(
        n7091), .ZN(n5126) );
  NAND2_X1 U5832 ( .A1(n7083), .A2(n7066), .ZN(n5351) );
  INV_X1 U5833 ( .A(n5351), .ZN(n5397) );
  OR2_X1 U5834 ( .A1(n4911), .A2(n4789), .ZN(n5350) );
  AND2_X1 U5835 ( .A1(n5350), .A2(n7066), .ZN(n5343) );
  NAND3_X1 U5836 ( .A1(n5300), .A2(n5299), .A3(n5261), .ZN(n7100) );
  NOR2_X2 U5837 ( .A1(n7100), .A2(n7077), .ZN(n7197) );
  OAI21_X1 U5838 ( .B1(n5127), .B2(n7197), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5124) );
  OAI21_X1 U5839 ( .B1(n5397), .B2(n5343), .A(n5124), .ZN(n5125) );
  NOR2_X1 U5840 ( .A1(n7083), .A2(n7112), .ZN(n5344) );
  INV_X1 U5841 ( .A(n5344), .ZN(n5457) );
  INV_X1 U5842 ( .A(n5128), .ZN(n5129) );
  NAND2_X1 U5843 ( .A1(n5129), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5454) );
  OAI22_X1 U5844 ( .A1(n5457), .A2(n5350), .B1(n5454), .B2(n5402), .ZN(n5291)
         );
  INV_X1 U5845 ( .A(n5130), .ZN(n5290) );
  AOI22_X1 U5846 ( .A1(n5497), .A2(n5291), .B1(n7165), .B2(n5290), .ZN(n5131)
         );
  OAI21_X1 U5847 ( .B1(n5500), .B2(n5293), .A(n5131), .ZN(n5132) );
  AOI21_X1 U5848 ( .B1(n7166), .B2(n7197), .A(n5132), .ZN(n5133) );
  OAI21_X1 U5849 ( .B1(n5297), .B2(n5134), .A(n5133), .ZN(U3025) );
  INV_X1 U5850 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5138) );
  AOI22_X1 U5851 ( .A1(n5469), .A2(n5291), .B1(n7135), .B2(n5290), .ZN(n5135)
         );
  OAI21_X1 U5852 ( .B1(n5472), .B2(n5293), .A(n5135), .ZN(n5136) );
  AOI21_X1 U5853 ( .B1(n7136), .B2(n7197), .A(n5136), .ZN(n5137) );
  OAI21_X1 U5854 ( .B1(n5297), .B2(n5138), .A(n5137), .ZN(U3022) );
  AOI22_X1 U5855 ( .A1(n5515), .A2(n5291), .B1(n7175), .B2(n5290), .ZN(n5139)
         );
  OAI21_X1 U5856 ( .B1(n5518), .B2(n5293), .A(n5139), .ZN(n5140) );
  AOI21_X1 U5857 ( .B1(n7177), .B2(n7197), .A(n5140), .ZN(n5141) );
  OAI21_X1 U5858 ( .B1(n5297), .B2(n5142), .A(n5141), .ZN(U3026) );
  INV_X1 U5859 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5146) );
  AOI22_X1 U5860 ( .A1(n5476), .A2(n5291), .B1(n7145), .B2(n5290), .ZN(n5143)
         );
  OAI21_X1 U5861 ( .B1(n5479), .B2(n5293), .A(n5143), .ZN(n5144) );
  AOI21_X1 U5862 ( .B1(n7146), .B2(n7197), .A(n5144), .ZN(n5145) );
  OAI21_X1 U5863 ( .B1(n5297), .B2(n5146), .A(n5145), .ZN(U3023) );
  AOI22_X1 U5864 ( .A1(n5490), .A2(n5291), .B1(n7125), .B2(n5290), .ZN(n5147)
         );
  OAI21_X1 U5865 ( .B1(n5493), .B2(n5293), .A(n5147), .ZN(n5148) );
  AOI21_X1 U5866 ( .B1(n7127), .B2(n7197), .A(n5148), .ZN(n5149) );
  OAI21_X1 U5867 ( .B1(n5297), .B2(n3881), .A(n5149), .ZN(U3021) );
  AOI22_X1 U5868 ( .A1(n5504), .A2(n5291), .B1(n7195), .B2(n5290), .ZN(n5150)
         );
  OAI21_X1 U5869 ( .B1(n5507), .B2(n5293), .A(n5150), .ZN(n5151) );
  AOI21_X1 U5870 ( .B1(n7199), .B2(n7197), .A(n5151), .ZN(n5152) );
  OAI21_X1 U5871 ( .B1(n5297), .B2(n5153), .A(n5152), .ZN(U3027) );
  AOI22_X1 U5872 ( .A1(n5462), .A2(n5291), .B1(n7109), .B2(n5290), .ZN(n5154)
         );
  OAI21_X1 U5873 ( .B1(n5465), .B2(n5293), .A(n5154), .ZN(n5155) );
  AOI21_X1 U5874 ( .B1(n7110), .B2(n7197), .A(n5155), .ZN(n5156) );
  OAI21_X1 U5875 ( .B1(n5297), .B2(n5157), .A(n5156), .ZN(U3020) );
  NOR2_X1 U5876 ( .A1(n5166), .A2(n7112), .ZN(n5227) );
  OAI21_X1 U5877 ( .B1(n5190), .B2(n5191), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5159) );
  OAI21_X1 U5878 ( .B1(n5397), .B2(n5227), .A(n5159), .ZN(n5165) );
  NOR2_X1 U5879 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5160), .ZN(n5188)
         );
  OR2_X1 U5880 ( .A1(n5348), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5455)
         );
  NAND2_X1 U5881 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5455), .ZN(n5452) );
  NAND2_X1 U5882 ( .A1(n5161), .A2(n5454), .ZN(n5391) );
  INV_X1 U5883 ( .A(n5391), .ZN(n5162) );
  OAI211_X1 U5884 ( .C1(n7089), .C2(n5188), .A(n5452), .B(n5162), .ZN(n5163)
         );
  INV_X1 U5885 ( .A(n5163), .ZN(n5164) );
  INV_X1 U5886 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5169) );
  INV_X1 U5887 ( .A(n5166), .ZN(n5231) );
  OAI22_X1 U5888 ( .A1(n5457), .A2(n5231), .B1(n5455), .B2(n5401), .ZN(n5189)
         );
  AOI22_X1 U5889 ( .A1(n5504), .A2(n5189), .B1(n7195), .B2(n5188), .ZN(n5168)
         );
  AOI22_X1 U5890 ( .A1(n7196), .A2(n5191), .B1(n5190), .B2(n7199), .ZN(n5167)
         );
  OAI211_X1 U5891 ( .C1(n5195), .C2(n5169), .A(n5168), .B(n5167), .ZN(U3075)
         );
  INV_X1 U5892 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5172) );
  AOI22_X1 U5893 ( .A1(n5515), .A2(n5189), .B1(n7175), .B2(n5188), .ZN(n5171)
         );
  AOI22_X1 U5894 ( .A1(n7176), .A2(n5191), .B1(n5190), .B2(n7177), .ZN(n5170)
         );
  OAI211_X1 U5895 ( .C1(n5195), .C2(n5172), .A(n5171), .B(n5170), .ZN(U3074)
         );
  INV_X1 U5896 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5175) );
  AOI22_X1 U5897 ( .A1(n5483), .A2(n5189), .B1(n7155), .B2(n5188), .ZN(n5174)
         );
  AOI22_X1 U5898 ( .A1(n7156), .A2(n5191), .B1(n5190), .B2(n7157), .ZN(n5173)
         );
  OAI211_X1 U5899 ( .C1(n5195), .C2(n5175), .A(n5174), .B(n5173), .ZN(U3072)
         );
  INV_X1 U5900 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5178) );
  AOI22_X1 U5901 ( .A1(n5490), .A2(n5189), .B1(n7125), .B2(n5188), .ZN(n5177)
         );
  AOI22_X1 U5902 ( .A1(n7126), .A2(n5191), .B1(n5190), .B2(n7127), .ZN(n5176)
         );
  OAI211_X1 U5903 ( .C1(n5195), .C2(n5178), .A(n5177), .B(n5176), .ZN(U3069)
         );
  INV_X1 U5904 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5181) );
  AOI22_X1 U5905 ( .A1(n5476), .A2(n5189), .B1(n7145), .B2(n5188), .ZN(n5180)
         );
  AOI22_X1 U5906 ( .A1(n7147), .A2(n5191), .B1(n5190), .B2(n7146), .ZN(n5179)
         );
  OAI211_X1 U5907 ( .C1(n5195), .C2(n5181), .A(n5180), .B(n5179), .ZN(U3071)
         );
  INV_X1 U5908 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5184) );
  AOI22_X1 U5909 ( .A1(n5497), .A2(n5189), .B1(n7165), .B2(n5188), .ZN(n5183)
         );
  AOI22_X1 U5910 ( .A1(n7167), .A2(n5191), .B1(n5190), .B2(n7166), .ZN(n5182)
         );
  OAI211_X1 U5911 ( .C1(n5195), .C2(n5184), .A(n5183), .B(n5182), .ZN(U3073)
         );
  INV_X1 U5912 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5187) );
  AOI22_X1 U5913 ( .A1(n5462), .A2(n5189), .B1(n7109), .B2(n5188), .ZN(n5186)
         );
  AOI22_X1 U5914 ( .A1(n7117), .A2(n5191), .B1(n5190), .B2(n7110), .ZN(n5185)
         );
  OAI211_X1 U5915 ( .C1(n5195), .C2(n5187), .A(n5186), .B(n5185), .ZN(U3068)
         );
  INV_X1 U5916 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5194) );
  AOI22_X1 U5917 ( .A1(n5469), .A2(n5189), .B1(n7135), .B2(n5188), .ZN(n5193)
         );
  AOI22_X1 U5918 ( .A1(n7137), .A2(n5191), .B1(n5190), .B2(n7136), .ZN(n5192)
         );
  OAI211_X1 U5919 ( .C1(n5195), .C2(n5194), .A(n5193), .B(n5192), .ZN(U3070)
         );
  NAND2_X1 U5920 ( .A1(n5196), .A2(n5299), .ZN(n5203) );
  NOR3_X1 U5921 ( .A1(n6978), .A2(n7068), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5303) );
  INV_X1 U5922 ( .A(n5303), .ZN(n5200) );
  NOR2_X1 U5923 ( .A1(n7103), .A2(n5200), .ZN(n5220) );
  AOI21_X1 U5924 ( .B1(n7067), .B2(n5400), .A(n5220), .ZN(n5202) );
  OR2_X1 U5925 ( .A1(n5203), .A2(n7028), .ZN(n5197) );
  AOI21_X1 U5926 ( .B1(n5202), .B2(n5199), .A(n7073), .ZN(n5198) );
  OAI21_X1 U5927 ( .B1(n7066), .B2(n5303), .A(n5198), .ZN(n5219) );
  INV_X1 U5928 ( .A(n5199), .ZN(n5201) );
  OAI22_X1 U5929 ( .A1(n5202), .A2(n5201), .B1(n6691), .B2(n5200), .ZN(n5218)
         );
  AOI22_X1 U5930 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5219), .B1(n5469), 
        .B2(n5218), .ZN(n5205) );
  NOR2_X2 U5931 ( .A1(n5203), .A2(n7077), .ZN(n5331) );
  AOI22_X1 U5932 ( .A1(n5331), .A2(n7137), .B1(n7135), .B2(n5220), .ZN(n5204)
         );
  OAI211_X1 U5933 ( .C1(n5466), .C2(n5225), .A(n5205), .B(n5204), .ZN(U3126)
         );
  AOI22_X1 U5934 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5219), .B1(n5490), 
        .B2(n5218), .ZN(n5207) );
  AOI22_X1 U5935 ( .A1(n5331), .A2(n7126), .B1(n7125), .B2(n5220), .ZN(n5206)
         );
  OAI211_X1 U5936 ( .C1(n5487), .C2(n5225), .A(n5207), .B(n5206), .ZN(U3125)
         );
  AOI22_X1 U5937 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5219), .B1(n5497), 
        .B2(n5218), .ZN(n5209) );
  AOI22_X1 U5938 ( .A1(n5331), .A2(n7167), .B1(n7165), .B2(n5220), .ZN(n5208)
         );
  OAI211_X1 U5939 ( .C1(n5494), .C2(n5225), .A(n5209), .B(n5208), .ZN(U3129)
         );
  AOI22_X1 U5940 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5219), .B1(n5462), 
        .B2(n5218), .ZN(n5211) );
  AOI22_X1 U5941 ( .A1(n5331), .A2(n7117), .B1(n7109), .B2(n5220), .ZN(n5210)
         );
  OAI211_X1 U5942 ( .C1(n5459), .C2(n5225), .A(n5211), .B(n5210), .ZN(U3124)
         );
  AOI22_X1 U5943 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5219), .B1(n5483), 
        .B2(n5218), .ZN(n5213) );
  AOI22_X1 U5944 ( .A1(n5331), .A2(n7156), .B1(n7155), .B2(n5220), .ZN(n5212)
         );
  OAI211_X1 U5945 ( .C1(n5480), .C2(n5225), .A(n5213), .B(n5212), .ZN(U3128)
         );
  AOI22_X1 U5946 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5219), .B1(n5504), 
        .B2(n5218), .ZN(n5215) );
  AOI22_X1 U5947 ( .A1(n5331), .A2(n7196), .B1(n7195), .B2(n5220), .ZN(n5214)
         );
  OAI211_X1 U5948 ( .C1(n5501), .C2(n5225), .A(n5215), .B(n5214), .ZN(U3131)
         );
  AOI22_X1 U5949 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5219), .B1(n5476), 
        .B2(n5218), .ZN(n5217) );
  AOI22_X1 U5950 ( .A1(n5331), .A2(n7147), .B1(n7145), .B2(n5220), .ZN(n5216)
         );
  OAI211_X1 U5951 ( .C1(n5473), .C2(n5225), .A(n5217), .B(n5216), .ZN(U3127)
         );
  AOI22_X1 U5952 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5219), .B1(n5515), 
        .B2(n5218), .ZN(n5222) );
  AOI22_X1 U5953 ( .A1(n5331), .A2(n7176), .B1(n7175), .B2(n5220), .ZN(n5221)
         );
  OAI211_X1 U5954 ( .C1(n5509), .C2(n5225), .A(n5222), .B(n5221), .ZN(U3130)
         );
  NOR2_X1 U5955 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5223), .ZN(n5253)
         );
  INV_X1 U5956 ( .A(n5253), .ZN(n5224) );
  NAND2_X1 U5957 ( .A1(n5301), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5230) );
  INV_X1 U5958 ( .A(n5230), .ZN(n7085) );
  NOR2_X1 U5959 ( .A1(n7085), .A2(n6691), .ZN(n7090) );
  AOI211_X1 U5960 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5224), .A(n7090), .B(
        n5391), .ZN(n5229) );
  OAI21_X1 U5961 ( .B1(n5256), .B2(n5255), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5226) );
  OAI21_X1 U5962 ( .B1(n5344), .B2(n5227), .A(n5226), .ZN(n5228) );
  INV_X1 U5963 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5234) );
  OAI22_X1 U5964 ( .A1(n5231), .A2(n5351), .B1(n5230), .B2(n5401), .ZN(n5254)
         );
  AOI22_X1 U5965 ( .A1(n5476), .A2(n5254), .B1(n7145), .B2(n5253), .ZN(n5233)
         );
  AOI22_X1 U5966 ( .A1(n7146), .A2(n5256), .B1(n5255), .B2(n7147), .ZN(n5232)
         );
  OAI211_X1 U5967 ( .C1(n5260), .C2(n5234), .A(n5233), .B(n5232), .ZN(U3135)
         );
  INV_X1 U5968 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5237) );
  AOI22_X1 U5969 ( .A1(n5490), .A2(n5254), .B1(n7125), .B2(n5253), .ZN(n5236)
         );
  AOI22_X1 U5970 ( .A1(n7127), .A2(n5256), .B1(n5255), .B2(n7126), .ZN(n5235)
         );
  OAI211_X1 U5971 ( .C1(n5260), .C2(n5237), .A(n5236), .B(n5235), .ZN(U3133)
         );
  INV_X1 U5972 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5240) );
  AOI22_X1 U5973 ( .A1(n5515), .A2(n5254), .B1(n7175), .B2(n5253), .ZN(n5239)
         );
  AOI22_X1 U5974 ( .A1(n7177), .A2(n5256), .B1(n5255), .B2(n7176), .ZN(n5238)
         );
  OAI211_X1 U5975 ( .C1(n5260), .C2(n5240), .A(n5239), .B(n5238), .ZN(U3138)
         );
  INV_X1 U5976 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5243) );
  AOI22_X1 U5977 ( .A1(n5497), .A2(n5254), .B1(n7165), .B2(n5253), .ZN(n5242)
         );
  AOI22_X1 U5978 ( .A1(n7166), .A2(n5256), .B1(n5255), .B2(n7167), .ZN(n5241)
         );
  OAI211_X1 U5979 ( .C1(n5260), .C2(n5243), .A(n5242), .B(n5241), .ZN(U3137)
         );
  INV_X1 U5980 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U5981 ( .A1(n5504), .A2(n5254), .B1(n7195), .B2(n5253), .ZN(n5245)
         );
  AOI22_X1 U5982 ( .A1(n7199), .A2(n5256), .B1(n5255), .B2(n7196), .ZN(n5244)
         );
  OAI211_X1 U5983 ( .C1(n5260), .C2(n5246), .A(n5245), .B(n5244), .ZN(U3139)
         );
  INV_X1 U5984 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5249) );
  AOI22_X1 U5985 ( .A1(n5469), .A2(n5254), .B1(n7135), .B2(n5253), .ZN(n5248)
         );
  AOI22_X1 U5986 ( .A1(n7136), .A2(n5256), .B1(n5255), .B2(n7137), .ZN(n5247)
         );
  OAI211_X1 U5987 ( .C1(n5260), .C2(n5249), .A(n5248), .B(n5247), .ZN(U3134)
         );
  INV_X1 U5988 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5252) );
  AOI22_X1 U5989 ( .A1(n5483), .A2(n5254), .B1(n7155), .B2(n5253), .ZN(n5251)
         );
  AOI22_X1 U5990 ( .A1(n7157), .A2(n5256), .B1(n5255), .B2(n7156), .ZN(n5250)
         );
  OAI211_X1 U5991 ( .C1(n5260), .C2(n5252), .A(n5251), .B(n5250), .ZN(U3136)
         );
  INV_X1 U5992 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5259) );
  AOI22_X1 U5993 ( .A1(n5462), .A2(n5254), .B1(n7109), .B2(n5253), .ZN(n5258)
         );
  AOI22_X1 U5994 ( .A1(n7110), .A2(n5256), .B1(n5255), .B2(n7117), .ZN(n5257)
         );
  OAI211_X1 U5995 ( .C1(n5260), .C2(n5259), .A(n5258), .B(n5257), .ZN(U3132)
         );
  INV_X1 U5996 ( .A(n5270), .ZN(n5264) );
  NOR3_X1 U5997 ( .A1(n7068), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5338) );
  OAI21_X1 U5998 ( .B1(n5270), .B2(n7028), .A(n7066), .ZN(n5268) );
  INV_X1 U5999 ( .A(n5268), .ZN(n5265) );
  INV_X1 U6000 ( .A(n5350), .ZN(n7104) );
  INV_X1 U6001 ( .A(n5338), .ZN(n5267) );
  NOR2_X1 U6002 ( .A1(n7103), .A2(n5267), .ZN(n5287) );
  AOI21_X1 U6003 ( .B1(n7067), .B2(n7104), .A(n5287), .ZN(n5269) );
  NAND2_X1 U6004 ( .A1(n5265), .A2(n5269), .ZN(n5266) );
  OAI211_X1 U6005 ( .C1(n7066), .C2(n5338), .A(n7116), .B(n5266), .ZN(n5286)
         );
  OAI22_X1 U6006 ( .A1(n5269), .A2(n5268), .B1(n6691), .B2(n5267), .ZN(n5285)
         );
  AOI22_X1 U6007 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5286), .B1(n5497), 
        .B2(n5285), .ZN(n5272) );
  AOI22_X1 U6008 ( .A1(n3419), .A2(n7166), .B1(n5287), .B2(n7165), .ZN(n5271)
         );
  OAI211_X1 U6009 ( .C1(n5340), .C2(n5500), .A(n5272), .B(n5271), .ZN(U3097)
         );
  AOI22_X1 U6010 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5286), .B1(n5515), 
        .B2(n5285), .ZN(n5274) );
  AOI22_X1 U6011 ( .A1(n3419), .A2(n7177), .B1(n5287), .B2(n7175), .ZN(n5273)
         );
  OAI211_X1 U6012 ( .C1(n5340), .C2(n5518), .A(n5274), .B(n5273), .ZN(U3098)
         );
  AOI22_X1 U6013 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5286), .B1(n5462), 
        .B2(n5285), .ZN(n5276) );
  AOI22_X1 U6014 ( .A1(n3419), .A2(n7110), .B1(n7109), .B2(n5287), .ZN(n5275)
         );
  OAI211_X1 U6015 ( .C1(n5340), .C2(n5465), .A(n5276), .B(n5275), .ZN(U3092)
         );
  AOI22_X1 U6016 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5286), .B1(n5483), 
        .B2(n5285), .ZN(n5278) );
  AOI22_X1 U6017 ( .A1(n3419), .A2(n7157), .B1(n5287), .B2(n7155), .ZN(n5277)
         );
  OAI211_X1 U6018 ( .C1(n5340), .C2(n5486), .A(n5278), .B(n5277), .ZN(U3096)
         );
  AOI22_X1 U6019 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5286), .B1(n5490), 
        .B2(n5285), .ZN(n5280) );
  AOI22_X1 U6020 ( .A1(n3419), .A2(n7127), .B1(n5287), .B2(n7125), .ZN(n5279)
         );
  OAI211_X1 U6021 ( .C1(n5340), .C2(n5493), .A(n5280), .B(n5279), .ZN(U3093)
         );
  AOI22_X1 U6022 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5286), .B1(n5476), 
        .B2(n5285), .ZN(n5282) );
  AOI22_X1 U6023 ( .A1(n3419), .A2(n7146), .B1(n5287), .B2(n7145), .ZN(n5281)
         );
  OAI211_X1 U6024 ( .C1(n5340), .C2(n5479), .A(n5282), .B(n5281), .ZN(U3095)
         );
  AOI22_X1 U6025 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5286), .B1(n5469), 
        .B2(n5285), .ZN(n5284) );
  AOI22_X1 U6026 ( .A1(n3419), .A2(n7136), .B1(n5287), .B2(n7135), .ZN(n5283)
         );
  OAI211_X1 U6027 ( .C1(n5340), .C2(n5472), .A(n5284), .B(n5283), .ZN(U3094)
         );
  AOI22_X1 U6028 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5286), .B1(n5504), 
        .B2(n5285), .ZN(n5289) );
  AOI22_X1 U6029 ( .A1(n3419), .A2(n7199), .B1(n5287), .B2(n7195), .ZN(n5288)
         );
  OAI211_X1 U6030 ( .C1(n5340), .C2(n5507), .A(n5289), .B(n5288), .ZN(U3099)
         );
  AOI22_X1 U6031 ( .A1(n5483), .A2(n5291), .B1(n7155), .B2(n5290), .ZN(n5292)
         );
  OAI21_X1 U6032 ( .B1(n5486), .B2(n5293), .A(n5292), .ZN(n5294) );
  AOI21_X1 U6033 ( .B1(n7157), .B2(n7197), .A(n5294), .ZN(n5295) );
  OAI21_X1 U6034 ( .B1(n5297), .B2(n5296), .A(n5295), .ZN(U3024) );
  NOR2_X1 U6035 ( .A1(n5401), .A2(n5301), .ZN(n5302) );
  AOI22_X1 U6036 ( .A1(n5397), .A2(n5400), .B1(n5302), .B2(n5347), .ZN(n5329)
         );
  INV_X1 U6037 ( .A(n7145), .ZN(n5474) );
  NAND2_X1 U6038 ( .A1(n7103), .A2(n5303), .ZN(n5328) );
  OAI22_X1 U6039 ( .A1(n7150), .A2(n5329), .B1(n5474), .B2(n5328), .ZN(n5304)
         );
  AOI21_X1 U6040 ( .B1(n7146), .B2(n5331), .A(n5304), .ZN(n5309) );
  AOI21_X1 U6041 ( .B1(n5347), .B2(n5348), .A(n6691), .ZN(n5339) );
  AOI211_X1 U6042 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5328), .A(n5339), .B(
        n5391), .ZN(n5307) );
  NOR2_X1 U6043 ( .A1(n5400), .A2(n7112), .ZN(n5396) );
  OAI21_X1 U6044 ( .B1(n5331), .B2(n7182), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5305) );
  OAI21_X1 U6045 ( .B1(n5344), .B2(n5396), .A(n5305), .ZN(n5306) );
  NAND2_X1 U6046 ( .A1(n5307), .A2(n5306), .ZN(n5332) );
  NAND2_X1 U6047 ( .A1(n5332), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5308)
         );
  OAI211_X1 U6048 ( .C1(n5335), .C2(n5479), .A(n5309), .B(n5308), .ZN(U3119)
         );
  INV_X1 U6049 ( .A(n7125), .ZN(n5488) );
  OAI22_X1 U6050 ( .A1(n7130), .A2(n5329), .B1(n5488), .B2(n5328), .ZN(n5310)
         );
  AOI21_X1 U6051 ( .B1(n7127), .B2(n5331), .A(n5310), .ZN(n5312) );
  NAND2_X1 U6052 ( .A1(n5332), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5311)
         );
  OAI211_X1 U6053 ( .C1(n5335), .C2(n5493), .A(n5312), .B(n5311), .ZN(U3117)
         );
  INV_X1 U6054 ( .A(n7135), .ZN(n5467) );
  OAI22_X1 U6055 ( .A1(n7140), .A2(n5329), .B1(n5467), .B2(n5328), .ZN(n5313)
         );
  AOI21_X1 U6056 ( .B1(n7136), .B2(n5331), .A(n5313), .ZN(n5315) );
  NAND2_X1 U6057 ( .A1(n5332), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5314)
         );
  OAI211_X1 U6058 ( .C1(n5335), .C2(n5472), .A(n5315), .B(n5314), .ZN(U3118)
         );
  INV_X1 U6059 ( .A(n7109), .ZN(n5460) );
  OAI22_X1 U6060 ( .A1(n7120), .A2(n5329), .B1(n5460), .B2(n5328), .ZN(n5316)
         );
  AOI21_X1 U6061 ( .B1(n7110), .B2(n5331), .A(n5316), .ZN(n5318) );
  NAND2_X1 U6062 ( .A1(n5332), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5317)
         );
  OAI211_X1 U6063 ( .C1(n5335), .C2(n5465), .A(n5318), .B(n5317), .ZN(U3116)
         );
  INV_X1 U6064 ( .A(n7195), .ZN(n5502) );
  OAI22_X1 U6065 ( .A1(n7203), .A2(n5329), .B1(n5502), .B2(n5328), .ZN(n5319)
         );
  AOI21_X1 U6066 ( .B1(n7199), .B2(n5331), .A(n5319), .ZN(n5321) );
  NAND2_X1 U6067 ( .A1(n5332), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5320)
         );
  OAI211_X1 U6068 ( .C1(n5335), .C2(n5507), .A(n5321), .B(n5320), .ZN(U3123)
         );
  INV_X1 U6069 ( .A(n7165), .ZN(n5495) );
  OAI22_X1 U6070 ( .A1(n7170), .A2(n5329), .B1(n5495), .B2(n5328), .ZN(n5322)
         );
  AOI21_X1 U6071 ( .B1(n7166), .B2(n5331), .A(n5322), .ZN(n5324) );
  NAND2_X1 U6072 ( .A1(n5332), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5323)
         );
  OAI211_X1 U6073 ( .C1(n5335), .C2(n5500), .A(n5324), .B(n5323), .ZN(U3121)
         );
  INV_X1 U6074 ( .A(n7175), .ZN(n5512) );
  OAI22_X1 U6075 ( .A1(n7180), .A2(n5329), .B1(n5512), .B2(n5328), .ZN(n5325)
         );
  AOI21_X1 U6076 ( .B1(n7177), .B2(n5331), .A(n5325), .ZN(n5327) );
  NAND2_X1 U6077 ( .A1(n5332), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5326)
         );
  OAI211_X1 U6078 ( .C1(n5335), .C2(n5518), .A(n5327), .B(n5326), .ZN(U3122)
         );
  INV_X1 U6079 ( .A(n7155), .ZN(n5481) );
  OAI22_X1 U6080 ( .A1(n7160), .A2(n5329), .B1(n5481), .B2(n5328), .ZN(n5330)
         );
  AOI21_X1 U6081 ( .B1(n7157), .B2(n5331), .A(n5330), .ZN(n5334) );
  NAND2_X1 U6082 ( .A1(n5332), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5333)
         );
  OAI211_X1 U6083 ( .C1(n5335), .C2(n5486), .A(n5334), .B(n5333), .ZN(U3120)
         );
  NAND2_X1 U6084 ( .A1(n5091), .A2(n5336), .ZN(n5337) );
  AND2_X1 U6085 ( .A1(n5444), .A2(n5337), .ZN(n6867) );
  INV_X1 U6086 ( .A(n6867), .ZN(n5441) );
  INV_X1 U6087 ( .A(DATAI_6_), .ZN(n6091) );
  OAI222_X1 U6088 ( .A1(n5441), .A2(n3421), .B1(n5816), .B2(n6091), .C1(n6287), 
        .C2(n4238), .ZN(U2885) );
  NAND2_X1 U6089 ( .A1(n7103), .A2(n5338), .ZN(n5352) );
  AOI211_X1 U6090 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5352), .A(n5339), .B(
        n7091), .ZN(n5346) );
  INV_X1 U6091 ( .A(n5384), .ZN(n5341) );
  OAI21_X1 U6092 ( .B1(n5386), .B2(n5341), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5342) );
  OAI21_X1 U6093 ( .B1(n5344), .B2(n5343), .A(n5342), .ZN(n5345) );
  INV_X1 U6094 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5356) );
  INV_X1 U6095 ( .A(n5454), .ZN(n7086) );
  NAND3_X1 U6096 ( .A1(n7086), .A2(n5348), .A3(n5347), .ZN(n5349) );
  OAI21_X1 U6097 ( .B1(n5351), .B2(n5350), .A(n5349), .ZN(n5382) );
  INV_X1 U6098 ( .A(n5352), .ZN(n5381) );
  AOI22_X1 U6099 ( .A1(n5497), .A2(n5382), .B1(n7165), .B2(n5381), .ZN(n5353)
         );
  OAI21_X1 U6100 ( .B1(n5500), .B2(n5384), .A(n5353), .ZN(n5354) );
  AOI21_X1 U6101 ( .B1(n5386), .B2(n7166), .A(n5354), .ZN(n5355) );
  OAI21_X1 U6102 ( .B1(n5389), .B2(n5356), .A(n5355), .ZN(U3089) );
  INV_X1 U6103 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5360) );
  AOI22_X1 U6104 ( .A1(n5476), .A2(n5382), .B1(n7145), .B2(n5381), .ZN(n5357)
         );
  OAI21_X1 U6105 ( .B1(n5479), .B2(n5384), .A(n5357), .ZN(n5358) );
  AOI21_X1 U6106 ( .B1(n5386), .B2(n7146), .A(n5358), .ZN(n5359) );
  OAI21_X1 U6107 ( .B1(n5389), .B2(n5360), .A(n5359), .ZN(U3087) );
  INV_X1 U6108 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5364) );
  AOI22_X1 U6109 ( .A1(n5490), .A2(n5382), .B1(n7125), .B2(n5381), .ZN(n5361)
         );
  OAI21_X1 U6110 ( .B1(n5493), .B2(n5384), .A(n5361), .ZN(n5362) );
  AOI21_X1 U6111 ( .B1(n5386), .B2(n7127), .A(n5362), .ZN(n5363) );
  OAI21_X1 U6112 ( .B1(n5389), .B2(n5364), .A(n5363), .ZN(U3085) );
  INV_X1 U6113 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5368) );
  AOI22_X1 U6114 ( .A1(n5483), .A2(n5382), .B1(n7155), .B2(n5381), .ZN(n5365)
         );
  OAI21_X1 U6115 ( .B1(n5486), .B2(n5384), .A(n5365), .ZN(n5366) );
  AOI21_X1 U6116 ( .B1(n5386), .B2(n7157), .A(n5366), .ZN(n5367) );
  OAI21_X1 U6117 ( .B1(n5389), .B2(n5368), .A(n5367), .ZN(U3088) );
  INV_X1 U6118 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5372) );
  AOI22_X1 U6119 ( .A1(n5515), .A2(n5382), .B1(n7175), .B2(n5381), .ZN(n5369)
         );
  OAI21_X1 U6120 ( .B1(n5518), .B2(n5384), .A(n5369), .ZN(n5370) );
  AOI21_X1 U6121 ( .B1(n5386), .B2(n7177), .A(n5370), .ZN(n5371) );
  OAI21_X1 U6122 ( .B1(n5389), .B2(n5372), .A(n5371), .ZN(U3090) );
  INV_X1 U6123 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5376) );
  AOI22_X1 U6124 ( .A1(n5469), .A2(n5382), .B1(n7135), .B2(n5381), .ZN(n5373)
         );
  OAI21_X1 U6125 ( .B1(n5472), .B2(n5384), .A(n5373), .ZN(n5374) );
  AOI21_X1 U6126 ( .B1(n5386), .B2(n7136), .A(n5374), .ZN(n5375) );
  OAI21_X1 U6127 ( .B1(n5389), .B2(n5376), .A(n5375), .ZN(U3086) );
  INV_X1 U6128 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5380) );
  AOI22_X1 U6129 ( .A1(n5504), .A2(n5382), .B1(n7195), .B2(n5381), .ZN(n5377)
         );
  OAI21_X1 U6130 ( .B1(n5507), .B2(n5384), .A(n5377), .ZN(n5378) );
  AOI21_X1 U6131 ( .B1(n5386), .B2(n7199), .A(n5378), .ZN(n5379) );
  OAI21_X1 U6132 ( .B1(n5389), .B2(n5380), .A(n5379), .ZN(U3091) );
  INV_X1 U6133 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5388) );
  AOI22_X1 U6134 ( .A1(n5462), .A2(n5382), .B1(n7109), .B2(n5381), .ZN(n5383)
         );
  OAI21_X1 U6135 ( .B1(n5465), .B2(n5384), .A(n5383), .ZN(n5385) );
  AOI21_X1 U6136 ( .B1(n5386), .B2(n7110), .A(n5385), .ZN(n5387) );
  OAI21_X1 U6137 ( .B1(n5389), .B2(n5388), .A(n5387), .ZN(U3084) );
  OR2_X1 U6138 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5390), .ZN(n5427)
         );
  AOI211_X1 U6139 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5427), .A(n5392), .B(
        n5391), .ZN(n5399) );
  INV_X1 U6140 ( .A(n5426), .ZN(n5393) );
  OAI21_X1 U6141 ( .B1(n5394), .B2(n5393), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5395) );
  OAI21_X1 U6142 ( .B1(n5397), .B2(n5396), .A(n5395), .ZN(n5398) );
  NAND2_X1 U6143 ( .A1(n5399), .A2(n5398), .ZN(n5425) );
  NAND2_X1 U6144 ( .A1(n5425), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5406) );
  INV_X1 U6145 ( .A(n5400), .ZN(n5403) );
  OAI22_X1 U6146 ( .A1(n5457), .A2(n5403), .B1(n5402), .B2(n5401), .ZN(n5429)
         );
  OAI22_X1 U6147 ( .A1(n5460), .A2(n5427), .B1(n5465), .B2(n5426), .ZN(n5404)
         );
  AOI21_X1 U6148 ( .B1(n5462), .B2(n5429), .A(n5404), .ZN(n5405) );
  OAI211_X1 U6149 ( .C1(n5432), .C2(n5459), .A(n5406), .B(n5405), .ZN(U3052)
         );
  NAND2_X1 U6150 ( .A1(n5425), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5409) );
  OAI22_X1 U6151 ( .A1(n5481), .A2(n5427), .B1(n5486), .B2(n5426), .ZN(n5407)
         );
  AOI21_X1 U6152 ( .B1(n5483), .B2(n5429), .A(n5407), .ZN(n5408) );
  OAI211_X1 U6153 ( .C1(n5432), .C2(n5480), .A(n5409), .B(n5408), .ZN(U3056)
         );
  NAND2_X1 U6154 ( .A1(n5425), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5412) );
  OAI22_X1 U6155 ( .A1(n5495), .A2(n5427), .B1(n5500), .B2(n5426), .ZN(n5410)
         );
  AOI21_X1 U6156 ( .B1(n5497), .B2(n5429), .A(n5410), .ZN(n5411) );
  OAI211_X1 U6157 ( .C1(n5432), .C2(n5494), .A(n5412), .B(n5411), .ZN(U3057)
         );
  NAND2_X1 U6158 ( .A1(n5425), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5415) );
  OAI22_X1 U6159 ( .A1(n5512), .A2(n5427), .B1(n5518), .B2(n5426), .ZN(n5413)
         );
  AOI21_X1 U6160 ( .B1(n5515), .B2(n5429), .A(n5413), .ZN(n5414) );
  OAI211_X1 U6161 ( .C1(n5432), .C2(n5509), .A(n5415), .B(n5414), .ZN(U3058)
         );
  NAND2_X1 U6162 ( .A1(n5425), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5418) );
  OAI22_X1 U6163 ( .A1(n5502), .A2(n5427), .B1(n5507), .B2(n5426), .ZN(n5416)
         );
  AOI21_X1 U6164 ( .B1(n5504), .B2(n5429), .A(n5416), .ZN(n5417) );
  OAI211_X1 U6165 ( .C1(n5432), .C2(n5501), .A(n5418), .B(n5417), .ZN(U3059)
         );
  NAND2_X1 U6166 ( .A1(n5425), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5421) );
  OAI22_X1 U6167 ( .A1(n5488), .A2(n5427), .B1(n5493), .B2(n5426), .ZN(n5419)
         );
  AOI21_X1 U6168 ( .B1(n5490), .B2(n5429), .A(n5419), .ZN(n5420) );
  OAI211_X1 U6169 ( .C1(n5432), .C2(n5487), .A(n5421), .B(n5420), .ZN(U3053)
         );
  NAND2_X1 U6170 ( .A1(n5425), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5424) );
  OAI22_X1 U6171 ( .A1(n5467), .A2(n5427), .B1(n5472), .B2(n5426), .ZN(n5422)
         );
  AOI21_X1 U6172 ( .B1(n5469), .B2(n5429), .A(n5422), .ZN(n5423) );
  OAI211_X1 U6173 ( .C1(n5432), .C2(n5466), .A(n5424), .B(n5423), .ZN(U3054)
         );
  NAND2_X1 U6174 ( .A1(n5425), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5431) );
  OAI22_X1 U6175 ( .A1(n5474), .A2(n5427), .B1(n5479), .B2(n5426), .ZN(n5428)
         );
  AOI21_X1 U6176 ( .B1(n5476), .B2(n5429), .A(n5428), .ZN(n5430) );
  OAI211_X1 U6177 ( .C1(n5432), .C2(n5473), .A(n5431), .B(n5430), .ZN(U3055)
         );
  INV_X1 U6178 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6532) );
  OAI222_X1 U6179 ( .A1(n5434), .A2(n3421), .B1(n5816), .B2(n5433), .C1(n6287), 
        .C2(n6532), .ZN(U2887) );
  INV_X1 U6180 ( .A(DATAI_2_), .ZN(n6088) );
  INV_X1 U6181 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6529) );
  OAI222_X1 U6182 ( .A1(n5658), .A2(n3421), .B1(n5816), .B2(n6088), .C1(n6287), 
        .C2(n6529), .ZN(U2889) );
  OR2_X1 U6183 ( .A1(n4876), .A2(n5435), .ZN(n5436) );
  NAND2_X1 U6184 ( .A1(n5437), .A2(n5436), .ZN(n6623) );
  INV_X1 U6185 ( .A(DATAI_3_), .ZN(n6232) );
  OAI222_X1 U6186 ( .A1(n6623), .A2(n3421), .B1(n5816), .B2(n6232), .C1(n6287), 
        .C2(n4217), .ZN(U2888) );
  NOR2_X1 U6187 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  OR2_X1 U6188 ( .A1(n6628), .A2(n5440), .ZN(n6860) );
  INV_X1 U6189 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5442) );
  OAI222_X1 U6190 ( .A1(n6860), .A2(n6629), .B1(n5442), .B2(n6636), .C1(n6283), 
        .C2(n5441), .ZN(U2853) );
  NAND2_X1 U6191 ( .A1(n5444), .A2(n5443), .ZN(n5445) );
  AND2_X1 U6192 ( .A1(n5560), .A2(n5445), .ZN(n6877) );
  INV_X1 U6193 ( .A(n6877), .ZN(n5446) );
  INV_X1 U6194 ( .A(DATAI_7_), .ZN(n6186) );
  OAI222_X1 U6195 ( .A1(n5446), .A2(n3421), .B1(n5816), .B2(n6186), .C1(n6287), 
        .C2(n4246), .ZN(U2884) );
  AOI21_X1 U6196 ( .B1(n5510), .B2(n7108), .A(n7081), .ZN(n5448) );
  AOI21_X1 U6197 ( .B1(n5672), .B2(n7084), .A(n5448), .ZN(n5449) );
  NOR2_X1 U6198 ( .A1(n5449), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5453) );
  NOR2_X1 U6199 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5450), .ZN(n5458)
         );
  INV_X1 U6200 ( .A(n7091), .ZN(n5451) );
  NAND2_X1 U6201 ( .A1(n5508), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5464) );
  OAI22_X1 U6202 ( .A1(n5457), .A2(n5456), .B1(n5455), .B2(n5454), .ZN(n5514)
         );
  INV_X1 U6203 ( .A(n5458), .ZN(n5511) );
  OAI22_X1 U6204 ( .A1(n5460), .A2(n5511), .B1(n5510), .B2(n5459), .ZN(n5461)
         );
  AOI21_X1 U6205 ( .B1(n5462), .B2(n5514), .A(n5461), .ZN(n5463) );
  OAI211_X1 U6206 ( .C1(n7108), .C2(n5465), .A(n5464), .B(n5463), .ZN(U3036)
         );
  NAND2_X1 U6207 ( .A1(n5508), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5471) );
  OAI22_X1 U6208 ( .A1(n5467), .A2(n5511), .B1(n5510), .B2(n5466), .ZN(n5468)
         );
  AOI21_X1 U6209 ( .B1(n5469), .B2(n5514), .A(n5468), .ZN(n5470) );
  OAI211_X1 U6210 ( .C1(n7108), .C2(n5472), .A(n5471), .B(n5470), .ZN(U3038)
         );
  NAND2_X1 U6211 ( .A1(n5508), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5478) );
  OAI22_X1 U6212 ( .A1(n5474), .A2(n5511), .B1(n5510), .B2(n5473), .ZN(n5475)
         );
  AOI21_X1 U6213 ( .B1(n5476), .B2(n5514), .A(n5475), .ZN(n5477) );
  OAI211_X1 U6214 ( .C1(n7108), .C2(n5479), .A(n5478), .B(n5477), .ZN(U3039)
         );
  NAND2_X1 U6215 ( .A1(n5508), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5485) );
  OAI22_X1 U6216 ( .A1(n5481), .A2(n5511), .B1(n5510), .B2(n5480), .ZN(n5482)
         );
  AOI21_X1 U6217 ( .B1(n5483), .B2(n5514), .A(n5482), .ZN(n5484) );
  OAI211_X1 U6218 ( .C1(n7108), .C2(n5486), .A(n5485), .B(n5484), .ZN(U3040)
         );
  NAND2_X1 U6219 ( .A1(n5508), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5492) );
  OAI22_X1 U6220 ( .A1(n5488), .A2(n5511), .B1(n5510), .B2(n5487), .ZN(n5489)
         );
  AOI21_X1 U6221 ( .B1(n5490), .B2(n5514), .A(n5489), .ZN(n5491) );
  OAI211_X1 U6222 ( .C1(n7108), .C2(n5493), .A(n5492), .B(n5491), .ZN(U3037)
         );
  NAND2_X1 U6223 ( .A1(n5508), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5499) );
  OAI22_X1 U6224 ( .A1(n5495), .A2(n5511), .B1(n5510), .B2(n5494), .ZN(n5496)
         );
  AOI21_X1 U6225 ( .B1(n5497), .B2(n5514), .A(n5496), .ZN(n5498) );
  OAI211_X1 U6226 ( .C1(n7108), .C2(n5500), .A(n5499), .B(n5498), .ZN(U3041)
         );
  NAND2_X1 U6227 ( .A1(n5508), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5506) );
  OAI22_X1 U6228 ( .A1(n5502), .A2(n5511), .B1(n5510), .B2(n5501), .ZN(n5503)
         );
  AOI21_X1 U6229 ( .B1(n5504), .B2(n5514), .A(n5503), .ZN(n5505) );
  OAI211_X1 U6230 ( .C1(n7108), .C2(n5507), .A(n5506), .B(n5505), .ZN(U3043)
         );
  NAND2_X1 U6231 ( .A1(n5508), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5517) );
  OAI22_X1 U6232 ( .A1(n5512), .A2(n5511), .B1(n5510), .B2(n5509), .ZN(n5513)
         );
  AOI21_X1 U6233 ( .B1(n5515), .B2(n5514), .A(n5513), .ZN(n5516) );
  OAI211_X1 U6234 ( .C1(n7108), .C2(n5518), .A(n5517), .B(n5516), .ZN(U3042)
         );
  AOI21_X1 U6235 ( .B1(n6669), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n5520), 
        .ZN(n5521) );
  OAI21_X1 U6236 ( .B1(n6676), .B2(n6858), .A(n5521), .ZN(n5522) );
  AOI21_X1 U6237 ( .B1(n6855), .B2(n6670), .A(n5522), .ZN(n5523) );
  OAI21_X1 U6238 ( .B1(n5524), .B2(n6952), .A(n5523), .ZN(U2981) );
  NAND2_X1 U6239 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  XOR2_X1 U6240 ( .A(n5528), .B(n5527), .Z(n6723) );
  NAND2_X1 U6241 ( .A1(n6723), .A2(n6671), .ZN(n5532) );
  INV_X1 U6242 ( .A(n6669), .ZN(n6422) );
  NAND2_X1 U6243 ( .A1(n6809), .A2(REIP_REG_1__SCAN_IN), .ZN(n6716) );
  OAI21_X1 U6244 ( .B1(n6422), .B2(n5529), .A(n6716), .ZN(n5530) );
  AOI21_X1 U6245 ( .B1(n6665), .B2(n5529), .A(n5530), .ZN(n5531) );
  OAI211_X1 U6246 ( .C1(n6426), .C2(n5585), .A(n5532), .B(n5531), .ZN(U2985)
         );
  INV_X1 U6247 ( .A(n5533), .ZN(n5534) );
  OR2_X1 U6248 ( .A1(n5535), .A2(n5534), .ZN(n7008) );
  OR3_X1 U6249 ( .A1(n7020), .A2(n7089), .A3(n7015), .ZN(n7023) );
  NAND2_X1 U6250 ( .A1(n7008), .A2(n7023), .ZN(n5536) );
  OR2_X1 U6251 ( .A1(n5536), .A2(n6809), .ZN(n5537) );
  INV_X1 U6252 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6326) );
  INV_X1 U6253 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5974) );
  NOR2_X1 U6254 ( .A1(n6316), .A2(n7011), .ZN(n5540) );
  AOI21_X1 U6255 ( .B1(n5946), .B2(n5971), .A(n6947), .ZN(n6835) );
  NAND2_X1 U6256 ( .A1(n7028), .A2(n7042), .ZN(n5550) );
  INV_X1 U6257 ( .A(n5550), .ZN(n5541) );
  AND3_X1 U6258 ( .A1(n5542), .A2(n3685), .A3(n5541), .ZN(n5543) );
  NAND2_X1 U6259 ( .A1(n6884), .A2(n6850), .ZN(n5964) );
  OR2_X1 U6260 ( .A1(n6684), .A2(n5550), .ZN(n6999) );
  AND2_X1 U6261 ( .A1(n6692), .A2(n6999), .ZN(n5970) );
  INV_X1 U6262 ( .A(n5970), .ZN(n5545) );
  INV_X1 U6263 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6078) );
  NAND3_X1 U6264 ( .A1(n3685), .A2(n5550), .A3(n6078), .ZN(n5544) );
  NAND2_X1 U6265 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  INV_X1 U6266 ( .A(n5547), .ZN(n5548) );
  NAND2_X1 U6267 ( .A1(n5971), .A2(n5548), .ZN(n6831) );
  OAI22_X1 U6268 ( .A1(n6907), .A2(n3726), .B1(n5929), .B2(n6831), .ZN(n5549)
         );
  AOI21_X1 U6269 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5964), .A(n5549), .ZN(n5558)
         );
  NAND2_X1 U6270 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5550), .ZN(n5551) );
  NOR2_X1 U6271 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  NAND2_X1 U6272 ( .A1(n6927), .A2(n6950), .ZN(n5555) );
  AOI22_X1 U6273 ( .A1(n6946), .A2(n5556), .B1(n5555), .B2(
        PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5557) );
  OAI211_X1 U6274 ( .C1(n6835), .C2(n5559), .A(n5558), .B(n5557), .ZN(U2827)
         );
  AOI21_X1 U6275 ( .B1(n5561), .B2(n5560), .A(n5591), .ZN(n5576) );
  INV_X1 U6276 ( .A(n5576), .ZN(n5646) );
  INV_X1 U6277 ( .A(n6628), .ZN(n5563) );
  OAI21_X1 U6278 ( .B1(n5563), .B2(n6626), .A(n5562), .ZN(n5564) );
  NAND2_X1 U6279 ( .A1(n5564), .A2(n5593), .ZN(n5641) );
  INV_X1 U6280 ( .A(n5641), .ZN(n6761) );
  AOI22_X1 U6281 ( .A1(n4738), .A2(n6761), .B1(n6281), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5565) );
  OAI21_X1 U6282 ( .B1(n5646), .B2(n6283), .A(n5565), .ZN(U2851) );
  NAND2_X1 U6283 ( .A1(n6837), .A2(n6670), .ZN(n5569) );
  NOR2_X1 U6284 ( .A1(n6422), .A2(n6832), .ZN(n5566) );
  AOI211_X1 U6285 ( .C1(n6665), .C2(n6836), .A(n5567), .B(n5566), .ZN(n5568)
         );
  OAI211_X1 U6286 ( .C1(n5570), .C2(n6952), .A(n5569), .B(n5568), .ZN(U2982)
         );
  INV_X1 U6287 ( .A(DATAI_8_), .ZN(n6093) );
  INV_X1 U6288 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6538) );
  OAI222_X1 U6289 ( .A1(n5646), .A2(n3421), .B1(n5816), .B2(n6093), .C1(n6287), 
        .C2(n6538), .ZN(U2883) );
  OAI21_X1 U6290 ( .B1(n5573), .B2(n5572), .A(n5607), .ZN(n6762) );
  NAND2_X1 U6291 ( .A1(n6809), .A2(REIP_REG_8__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U6292 ( .A1(n6669), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5574)
         );
  OAI211_X1 U6293 ( .C1(n6676), .C2(n5640), .A(n6759), .B(n5574), .ZN(n5575)
         );
  AOI21_X1 U6294 ( .B1(n5576), .B2(n6670), .A(n5575), .ZN(n5577) );
  OAI21_X1 U6295 ( .B1(n6762), .B2(n6952), .A(n5577), .ZN(U2978) );
  INV_X1 U6296 ( .A(n6831), .ZN(n5581) );
  NOR2_X1 U6297 ( .A1(n6950), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5580)
         );
  INV_X1 U6298 ( .A(n6850), .ZN(n5962) );
  AOI22_X1 U6299 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6943), .B1(n5962), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n5578) );
  OAI21_X1 U6300 ( .B1(n6927), .B2(n5529), .A(n5578), .ZN(n5579) );
  AOI211_X1 U6301 ( .C1(n5581), .C2(n4789), .A(n5580), .B(n5579), .ZN(n5584)
         );
  INV_X1 U6302 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5582) );
  AOI22_X1 U6303 ( .A1(n6946), .A2(n6718), .B1(n6862), .B2(n5582), .ZN(n5583)
         );
  OAI211_X1 U6304 ( .C1(n6835), .C2(n5585), .A(n5584), .B(n5583), .ZN(U2826)
         );
  XOR2_X1 U6305 ( .A(n5587), .B(n5586), .Z(n6913) );
  INV_X1 U6306 ( .A(n6913), .ZN(n5588) );
  INV_X1 U6307 ( .A(DATAI_13_), .ZN(n6222) );
  INV_X1 U6308 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6547) );
  OAI222_X1 U6309 ( .A1(n3421), .A2(n5588), .B1(n5816), .B2(n6222), .C1(n6287), 
        .C2(n6547), .ZN(U2878) );
  INV_X1 U6310 ( .A(n5678), .ZN(n5589) );
  OAI21_X1 U6311 ( .B1(n5591), .B2(n5590), .A(n5589), .ZN(n5647) );
  INV_X1 U6312 ( .A(n5603), .ZN(n5592) );
  AOI21_X1 U6313 ( .B1(n5594), .B2(n5593), .A(n5592), .ZN(n6783) );
  AOI22_X1 U6314 ( .A1(n4738), .A2(n6783), .B1(n6281), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5595) );
  OAI21_X1 U6315 ( .B1(n5647), .B2(n6283), .A(n5595), .ZN(U2850) );
  NOR2_X1 U6316 ( .A1(n6884), .A2(REIP_REG_9__SCAN_IN), .ZN(n6891) );
  NAND4_X1 U6317 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .A4(REIP_REG_4__SCAN_IN), .ZN(n6852) );
  NOR2_X1 U6318 ( .A1(n6852), .A2(n6851), .ZN(n6861) );
  NAND3_X1 U6319 ( .A1(n6861), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .ZN(n5638) );
  INV_X1 U6320 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6561) );
  NOR2_X1 U6321 ( .A1(n5638), .A2(n6561), .ZN(n5639) );
  NAND2_X1 U6322 ( .A1(n6946), .A2(n6783), .ZN(n5597) );
  NAND2_X1 U6323 ( .A1(n6850), .A2(n5596), .ZN(n6925) );
  OAI211_X1 U6324 ( .C1(n6950), .C2(n5613), .A(n5597), .B(n6925), .ZN(n5601)
         );
  OAI21_X1 U6325 ( .B1(n6884), .B2(n5639), .A(n6850), .ZN(n6890) );
  AOI22_X1 U6326 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6939), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6890), .ZN(n5598) );
  OAI21_X1 U6327 ( .B1(n5599), .B2(n6907), .A(n5598), .ZN(n5600) );
  AOI211_X1 U6328 ( .C1(n6891), .C2(n5639), .A(n5601), .B(n5600), .ZN(n5602)
         );
  OAI21_X1 U6329 ( .B1(n6077), .B2(n5647), .A(n5602), .ZN(U2818) );
  XNOR2_X1 U6330 ( .A(n5678), .B(n5618), .ZN(n6887) );
  AOI21_X1 U6331 ( .B1(n5604), .B2(n5603), .A(n5625), .ZN(n6886) );
  AOI22_X1 U6332 ( .A1(n4738), .A2(n6886), .B1(n6281), .B2(EBX_REG_10__SCAN_IN), .ZN(n5605) );
  OAI21_X1 U6333 ( .B1(n6887), .B2(n6283), .A(n5605), .ZN(U2849) );
  NAND2_X1 U6334 ( .A1(n5607), .A2(n5606), .ZN(n5610) );
  NAND2_X1 U6335 ( .A1(n5610), .A2(n5609), .ZN(n5608) );
  OAI21_X1 U6336 ( .B1(n5610), .B2(n5609), .A(n5608), .ZN(n5611) );
  INV_X1 U6337 ( .A(n5611), .ZN(n6785) );
  NAND2_X1 U6338 ( .A1(n6785), .A2(n6671), .ZN(n5616) );
  INV_X1 U6339 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5612) );
  NOR2_X1 U6340 ( .A1(n6818), .A2(n5612), .ZN(n6782) );
  NOR2_X1 U6341 ( .A1(n6676), .A2(n5613), .ZN(n5614) );
  AOI211_X1 U6342 ( .C1(n6669), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6782), 
        .B(n5614), .ZN(n5615) );
  OAI211_X1 U6343 ( .C1(n6426), .C2(n5647), .A(n5616), .B(n5615), .ZN(U2977)
         );
  NAND2_X1 U6344 ( .A1(n5678), .A2(n5617), .ZN(n5704) );
  AND2_X1 U6345 ( .A1(n5678), .A2(n5618), .ZN(n5620) );
  NAND2_X1 U6346 ( .A1(n5704), .A2(n5621), .ZN(n5742) );
  NAND2_X1 U6347 ( .A1(n5639), .A2(REIP_REG_9__SCAN_IN), .ZN(n6883) );
  INV_X1 U6348 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6564) );
  NOR2_X1 U6349 ( .A1(n6883), .A2(n6564), .ZN(n5627) );
  NAND2_X1 U6350 ( .A1(n5627), .A2(REIP_REG_11__SCAN_IN), .ZN(n5838) );
  INV_X1 U6351 ( .A(n5838), .ZN(n5622) );
  NAND2_X1 U6352 ( .A1(n6850), .A2(n5622), .ZN(n5623) );
  NAND2_X1 U6353 ( .A1(n5964), .A2(n5623), .ZN(n6906) );
  INV_X1 U6354 ( .A(n6906), .ZN(n6897) );
  NOR2_X1 U6355 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  NAND2_X1 U6356 ( .A1(n6946), .A2(n3444), .ZN(n5632) );
  NAND2_X1 U6357 ( .A1(n6862), .A2(n5627), .ZN(n5629) );
  OAI22_X1 U6358 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5629), .B1(n5628), .B2(
        n6907), .ZN(n5630) );
  AOI211_X1 U6359 ( .C1(n6939), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5630), 
        .B(n6910), .ZN(n5631) );
  OAI211_X1 U6360 ( .C1(n5738), .C2(n6950), .A(n5632), .B(n5631), .ZN(n5633)
         );
  AOI21_X1 U6361 ( .B1(n6897), .B2(REIP_REG_11__SCAN_IN), .A(n5633), .ZN(n5634) );
  OAI21_X1 U6362 ( .B1(n5742), .B2(n6077), .A(n5634), .ZN(U2816) );
  AOI22_X1 U6363 ( .A1(n4738), .A2(n3444), .B1(n6281), .B2(EBX_REG_11__SCAN_IN), .ZN(n5635) );
  OAI21_X1 U6364 ( .B1(n5742), .B2(n6283), .A(n5635), .ZN(U2848) );
  AOI22_X1 U6365 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6939), .B1(
        REIP_REG_8__SCAN_IN), .B2(n6890), .ZN(n5636) );
  OAI211_X1 U6366 ( .C1(n6907), .C2(n5637), .A(n5636), .B(n6925), .ZN(n5644)
         );
  NOR3_X1 U6367 ( .A1(n6884), .A2(n5639), .A3(n5638), .ZN(n5643) );
  OAI22_X1 U6368 ( .A1(n6931), .A2(n5641), .B1(n6950), .B2(n5640), .ZN(n5642)
         );
  NOR3_X1 U6369 ( .A1(n5644), .A2(n5643), .A3(n5642), .ZN(n5645) );
  OAI21_X1 U6370 ( .B1(n5646), .B2(n6077), .A(n5645), .ZN(U2819) );
  INV_X1 U6371 ( .A(DATAI_9_), .ZN(n6230) );
  INV_X1 U6372 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6540) );
  OAI222_X1 U6373 ( .A1(n5647), .A2(n3421), .B1(n5816), .B2(n6230), .C1(n6287), 
        .C2(n6540), .ZN(U2882) );
  INV_X1 U6374 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6544) );
  OAI222_X1 U6375 ( .A1(n5742), .A2(n3421), .B1(n5816), .B2(n5648), .C1(n6287), 
        .C2(n6544), .ZN(U2880) );
  NOR2_X1 U6376 ( .A1(n6831), .A2(n5649), .ZN(n5656) );
  NAND2_X1 U6377 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n6839) );
  OAI211_X1 U6378 ( .C1(REIP_REG_1__SCAN_IN), .C2(REIP_REG_2__SCAN_IN), .A(
        n6862), .B(n6839), .ZN(n5654) );
  AOI22_X1 U6379 ( .A1(n6939), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5962), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U6380 ( .A1(n6946), .A2(n6746), .ZN(n5652) );
  INV_X1 U6381 ( .A(n6644), .ZN(n5650) );
  NAND2_X1 U6382 ( .A1(n6923), .A2(n5650), .ZN(n5651) );
  NAND4_X1 U6383 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), .ZN(n5655)
         );
  AOI211_X1 U6384 ( .C1(EBX_REG_2__SCAN_IN), .C2(n6943), .A(n5656), .B(n5655), 
        .ZN(n5657) );
  OAI21_X1 U6385 ( .B1(n6835), .B2(n5658), .A(n5657), .ZN(U2825) );
  INV_X1 U6386 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6542) );
  OAI222_X1 U6387 ( .A1(n3421), .A2(n6887), .B1(n5816), .B2(n5659), .C1(n6287), 
        .C2(n6542), .ZN(U2881) );
  INV_X1 U6388 ( .A(n5660), .ZN(n5663) );
  MUX2_X1 U6389 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .B(n5661), .S(n6418), 
        .Z(n5662) );
  NOR2_X1 U6390 ( .A1(n5663), .A2(n5662), .ZN(n5736) );
  AOI21_X1 U6391 ( .B1(n5663), .B2(n5662), .A(n5736), .ZN(n6779) );
  NAND2_X1 U6392 ( .A1(n6779), .A2(n6671), .ZN(n5667) );
  INV_X1 U6393 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U6394 ( .A1(n6809), .A2(REIP_REG_10__SCAN_IN), .ZN(n6774) );
  OAI21_X1 U6395 ( .B1(n6422), .B2(n5664), .A(n6774), .ZN(n5665) );
  AOI21_X1 U6396 ( .B1(n6665), .B2(n6888), .A(n5665), .ZN(n5666) );
  OAI211_X1 U6397 ( .C1(n6887), .C2(n6426), .A(n5667), .B(n5666), .ZN(U2976)
         );
  NOR2_X1 U6398 ( .A1(n5962), .A2(n6839), .ZN(n5668) );
  INV_X1 U6399 ( .A(n5964), .ZN(n6035) );
  AOI21_X1 U6400 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5668), .A(n6035), .ZN(n6834)
         );
  OAI21_X1 U6401 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5668), .A(n6834), .ZN(n5676)
         );
  XNOR2_X1 U6402 ( .A(n5670), .B(n5669), .ZN(n6728) );
  INV_X1 U6403 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5671) );
  OAI22_X1 U6404 ( .A1(n6927), .A2(n5671), .B1(n6652), .B2(n6950), .ZN(n5674)
         );
  OAI22_X1 U6405 ( .A1(n6907), .A2(n6625), .B1(n5672), .B2(n6831), .ZN(n5673)
         );
  AOI211_X1 U6406 ( .C1(n6946), .C2(n6728), .A(n5674), .B(n5673), .ZN(n5675)
         );
  OAI211_X1 U6407 ( .C1(n6835), .C2(n6623), .A(n5676), .B(n5675), .ZN(U2824)
         );
  NAND2_X1 U6408 ( .A1(n5678), .A2(n5677), .ZN(n5680) );
  NAND2_X1 U6409 ( .A1(n5680), .A2(n5679), .ZN(n5682) );
  NAND2_X1 U6410 ( .A1(n5682), .A2(n5681), .ZN(n5784) );
  OAI21_X1 U6411 ( .B1(n5682), .B2(n5681), .A(n5784), .ZN(n5776) );
  INV_X1 U6412 ( .A(n5754), .ZN(n5685) );
  OAI21_X1 U6413 ( .B1(n5808), .B2(n5685), .A(n5684), .ZN(n5686) );
  AND2_X1 U6414 ( .A1(n5686), .A2(n5786), .ZN(n6709) );
  NAND2_X1 U6415 ( .A1(n6939), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5687)
         );
  OAI211_X1 U6416 ( .C1(n6950), .C2(n5778), .A(n5687), .B(n6925), .ZN(n5693)
         );
  NAND3_X1 U6417 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_14__SCAN_IN), .ZN(n5836) );
  OR3_X1 U6418 ( .A1(n5836), .A2(n5838), .A3(n5962), .ZN(n5716) );
  AND2_X1 U6419 ( .A1(n5964), .A2(n5716), .ZN(n5858) );
  AOI22_X1 U6420 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6943), .B1(
        REIP_REG_14__SCAN_IN), .B2(n5858), .ZN(n5691) );
  NAND2_X1 U6421 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n6915) );
  INV_X1 U6422 ( .A(n6915), .ZN(n5689) );
  INV_X1 U6423 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5688) );
  NOR2_X1 U6424 ( .A1(n6884), .A2(n5838), .ZN(n6916) );
  NAND3_X1 U6425 ( .A1(n5689), .A2(n5688), .A3(n6916), .ZN(n5690) );
  NAND2_X1 U6426 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  AOI211_X1 U6427 ( .C1(n6709), .C2(n6946), .A(n5693), .B(n5692), .ZN(n5694)
         );
  OAI21_X1 U6428 ( .B1(n5776), .B2(n6077), .A(n5694), .ZN(U2813) );
  AOI22_X1 U6429 ( .A1(n6709), .A2(n4738), .B1(EBX_REG_14__SCAN_IN), .B2(n6281), .ZN(n5695) );
  OAI21_X1 U6430 ( .B1(n5776), .B2(n6283), .A(n5695), .ZN(U2845) );
  OAI21_X1 U6431 ( .B1(n4442), .B2(n3450), .A(n5760), .ZN(n6921) );
  AND2_X1 U6432 ( .A1(n3625), .A2(n5697), .ZN(n5698) );
  AOI22_X1 U6433 ( .A1(n7059), .A2(DATAI_2_), .B1(n7062), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5701) );
  NOR2_X2 U6434 ( .A1(n7062), .A2(n5699), .ZN(n7063) );
  NAND2_X1 U6435 ( .A1(n7063), .A2(DATAI_18_), .ZN(n5700) );
  OAI211_X1 U6436 ( .C1(n6921), .C2(n3421), .A(n5701), .B(n5700), .ZN(U2873)
         );
  INV_X1 U6437 ( .A(n5702), .ZN(n5703) );
  AOI21_X1 U6438 ( .B1(n5705), .B2(n5704), .A(n5703), .ZN(n6902) );
  INV_X1 U6439 ( .A(n6902), .ZN(n5706) );
  INV_X1 U6440 ( .A(DATAI_12_), .ZN(n6226) );
  OAI222_X1 U6441 ( .A1(n5706), .A2(n3421), .B1(n5816), .B2(n6226), .C1(n6287), 
        .C2(n4310), .ZN(U2879) );
  AND2_X1 U6442 ( .A1(n3423), .A2(n5707), .ZN(n5853) );
  OR2_X1 U6443 ( .A1(n5853), .A2(n5709), .ZN(n5710) );
  AND2_X1 U6444 ( .A1(n5696), .A2(n5710), .ZN(n7053) );
  INV_X1 U6445 ( .A(n7053), .ZN(n5724) );
  OR2_X1 U6446 ( .A1(n5712), .A2(n5713), .ZN(n5714) );
  AND2_X1 U6447 ( .A1(n5726), .A2(n5714), .ZN(n6515) );
  NAND2_X1 U6448 ( .A1(n6939), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5715)
         );
  OAI211_X1 U6449 ( .C1(n6950), .C2(n6675), .A(n5715), .B(n6925), .ZN(n5719)
         );
  NAND2_X1 U6450 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n5859) );
  INV_X1 U6451 ( .A(n6916), .ZN(n6899) );
  NOR3_X1 U6452 ( .A1(n5836), .A2(n5859), .A3(n6899), .ZN(n5762) );
  NOR2_X1 U6453 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5762), .ZN(n5717) );
  NAND3_X1 U6454 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_17__SCAN_IN), .ZN(n5835) );
  OAI21_X1 U6455 ( .B1(n5835), .B2(n5716), .A(n5964), .ZN(n6936) );
  OAI22_X1 U6456 ( .A1(n5717), .A2(n6936), .B1(n5721), .B2(n6907), .ZN(n5718)
         );
  AOI211_X1 U6457 ( .C1(n6515), .C2(n6946), .A(n5719), .B(n5718), .ZN(n5720)
         );
  OAI21_X1 U6458 ( .B1(n5724), .B2(n6077), .A(n5720), .ZN(U2810) );
  NOR2_X1 U6459 ( .A1(n6636), .A2(n5721), .ZN(n5722) );
  AOI21_X1 U6460 ( .B1(n6515), .B2(n4738), .A(n5722), .ZN(n5723) );
  OAI21_X1 U6461 ( .B1(n5724), .B2(n6283), .A(n5723), .ZN(U2842) );
  NAND2_X1 U6462 ( .A1(n5726), .A2(n5725), .ZN(n5727) );
  NAND2_X1 U6463 ( .A1(n5764), .A2(n5727), .ZN(n6930) );
  INV_X1 U6464 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5728) );
  OAI222_X1 U6465 ( .A1(n6930), .A2(n6629), .B1(n5728), .B2(n6636), .C1(n6921), 
        .C2(n6283), .ZN(U2841) );
  INV_X1 U6466 ( .A(DATAI_14_), .ZN(n6216) );
  OAI222_X1 U6467 ( .A1(n5776), .A2(n3421), .B1(n5816), .B2(n6216), .C1(n6287), 
        .C2(n4340), .ZN(U2877) );
  XOR2_X1 U6468 ( .A(n5731), .B(n5730), .Z(n5758) );
  INV_X1 U6469 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5732) );
  NOR2_X1 U6470 ( .A1(n6818), .A2(n5732), .ZN(n5755) );
  AOI21_X1 U6471 ( .B1(n6669), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5755), 
        .ZN(n5733) );
  OAI21_X1 U6472 ( .B1(n6676), .B2(n6911), .A(n5733), .ZN(n5734) );
  AOI21_X1 U6473 ( .B1(n6913), .B2(n6670), .A(n5734), .ZN(n5735) );
  OAI21_X1 U6474 ( .B1(n5758), .B2(n6952), .A(n5735), .ZN(U2973) );
  AOI21_X1 U6475 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n4116), .A(n5736), 
        .ZN(n5800) );
  XNOR2_X1 U6476 ( .A(n6418), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5737)
         );
  XNOR2_X1 U6477 ( .A(n5800), .B(n5737), .ZN(n6791) );
  NAND2_X1 U6478 ( .A1(n6791), .A2(n6671), .ZN(n5741) );
  AND2_X1 U6479 ( .A1(n6809), .A2(REIP_REG_11__SCAN_IN), .ZN(n6790) );
  NOR2_X1 U6480 ( .A1(n6676), .A2(n5738), .ZN(n5739) );
  AOI211_X1 U6481 ( .C1(n6669), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6790), 
        .B(n5739), .ZN(n5740) );
  OAI211_X1 U6482 ( .C1(n6426), .C2(n5742), .A(n5741), .B(n5740), .ZN(U2975)
         );
  INV_X1 U6483 ( .A(n6758), .ZN(n5745) );
  AOI22_X1 U6484 ( .A1(n6748), .A2(n5745), .B1(n5744), .B2(n5743), .ZN(n6764)
         );
  AOI21_X1 U6485 ( .B1(n6764), .B2(n5746), .A(n6721), .ZN(n5747) );
  AOI21_X1 U6486 ( .B1(n6715), .B2(n5750), .A(n6794), .ZN(n5748) );
  OAI21_X1 U6487 ( .B1(n6700), .B2(n5749), .A(n5748), .ZN(n6701) );
  NOR2_X1 U6488 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5750), .ZN(n6703)
         );
  NOR2_X1 U6489 ( .A1(n5752), .A2(n5751), .ZN(n6705) );
  INV_X1 U6490 ( .A(n6817), .ZN(n5753) );
  AOI22_X1 U6491 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6701), .B1(n6703), .B2(n5753), .ZN(n5757) );
  XNOR2_X1 U6492 ( .A(n5808), .B(n5754), .ZN(n6914) );
  AOI21_X1 U6493 ( .B1(n6826), .B2(n6914), .A(n5755), .ZN(n5756) );
  OAI211_X1 U6494 ( .C1(n5758), .C2(n6800), .A(n5757), .B(n5756), .ZN(U3005)
         );
  AND2_X1 U6495 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  OR2_X1 U6496 ( .A1(n5761), .A2(n5829), .ZN(n6411) );
  NAND2_X1 U6497 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5762), .ZN(n5766) );
  OR2_X1 U6498 ( .A1(n5766), .A2(REIP_REG_18__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U6499 ( .A1(n6934), .A2(n6936), .ZN(n5771) );
  AND2_X1 U6500 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  OR2_X1 U6501 ( .A1(n5833), .A2(n5765), .ZN(n6503) );
  OAI22_X1 U6502 ( .A1(n6503), .A2(n6931), .B1(n6907), .B2(n5818), .ZN(n5770)
         );
  INV_X1 U6503 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6937) );
  NOR3_X1 U6504 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6937), .A3(n5766), .ZN(n5767) );
  AOI211_X1 U6505 ( .C1(n6939), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5767), 
        .B(n6910), .ZN(n5768) );
  OAI21_X1 U6506 ( .B1(n6413), .B2(n6950), .A(n5768), .ZN(n5769) );
  AOI211_X1 U6507 ( .C1(REIP_REG_19__SCAN_IN), .C2(n5771), .A(n5770), .B(n5769), .ZN(n5772) );
  OAI21_X1 U6508 ( .B1(n6411), .B2(n6077), .A(n5772), .ZN(U2808) );
  OAI21_X1 U6509 ( .B1(n5775), .B2(n5774), .A(n5773), .ZN(n6710) );
  INV_X1 U6510 ( .A(n6710), .ZN(n5782) );
  INV_X1 U6511 ( .A(n5776), .ZN(n5780) );
  AOI22_X1 U6512 ( .A1(n6669), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6809), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5777) );
  OAI21_X1 U6513 ( .B1(n6676), .B2(n5778), .A(n5777), .ZN(n5779) );
  AOI21_X1 U6514 ( .B1(n5780), .B2(n6670), .A(n5779), .ZN(n5781) );
  OAI21_X1 U6515 ( .B1(n5782), .B2(n6952), .A(n5781), .ZN(U2972) );
  INV_X1 U6516 ( .A(n5851), .ZN(n5783) );
  AOI21_X1 U6517 ( .B1(n5785), .B2(n5784), .A(n5783), .ZN(n5826) );
  INV_X1 U6518 ( .A(n5826), .ZN(n5817) );
  INV_X1 U6519 ( .A(n5786), .ZN(n5790) );
  INV_X1 U6520 ( .A(n5787), .ZN(n5789) );
  INV_X1 U6521 ( .A(n5788), .ZN(n5854) );
  OAI21_X1 U6522 ( .B1(n5790), .B2(n5789), .A(n5854), .ZN(n6798) );
  INV_X1 U6523 ( .A(n6798), .ZN(n5796) );
  AOI22_X1 U6524 ( .A1(n5796), .A2(n4738), .B1(n6281), .B2(EBX_REG_15__SCAN_IN), .ZN(n5791) );
  OAI21_X1 U6525 ( .B1(n5817), .B2(n6283), .A(n5791), .ZN(U2844) );
  NOR2_X1 U6526 ( .A1(n5836), .A2(n6899), .ZN(n5860) );
  INV_X1 U6527 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6797) );
  AOI21_X1 U6528 ( .B1(n6939), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6910), 
        .ZN(n5792) );
  OAI21_X1 U6529 ( .B1(n5793), .B2(n6907), .A(n5792), .ZN(n5794) );
  AOI221_X1 U6530 ( .B1(n5858), .B2(REIP_REG_15__SCAN_IN), .C1(n5860), .C2(
        n6797), .A(n5794), .ZN(n5798) );
  AOI22_X1 U6531 ( .A1(n5796), .A2(n6946), .B1(n6923), .B2(n5795), .ZN(n5797)
         );
  OAI211_X1 U6532 ( .C1(n5817), .C2(n6077), .A(n5798), .B(n5797), .ZN(U2812)
         );
  NAND2_X1 U6533 ( .A1(n6418), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U6534 ( .A1(n4116), .A2(n5799), .ZN(n5801) );
  MUX2_X1 U6535 ( .A(n5802), .B(n5801), .S(n5800), .Z(n5804) );
  XNOR2_X1 U6536 ( .A(n5804), .B(n5803), .ZN(n6668) );
  OR2_X1 U6537 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  AND2_X1 U6538 ( .A1(n5808), .A2(n5807), .ZN(n6896) );
  AOI22_X1 U6539 ( .A1(n6826), .A2(n6896), .B1(n6809), .B2(
        REIP_REG_12__SCAN_IN), .ZN(n5815) );
  NOR2_X1 U6540 ( .A1(n6817), .A2(n5799), .ZN(n5812) );
  AOI221_X1 U6541 ( .B1(n6748), .B2(n5799), .C1(n5809), .C2(n5799), .A(n6794), 
        .ZN(n5810) );
  INV_X1 U6542 ( .A(n5810), .ZN(n5811) );
  MUX2_X1 U6543 ( .A(n5812), .B(n5811), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n5813) );
  INV_X1 U6544 ( .A(n5813), .ZN(n5814) );
  OAI211_X1 U6545 ( .C1(n6668), .C2(n6800), .A(n5815), .B(n5814), .ZN(U3006)
         );
  OAI222_X1 U6546 ( .A1(n5817), .A2(n3421), .B1(n5816), .B2(n6213), .C1(n6287), 
        .C2(n4764), .ZN(U2876) );
  OAI222_X1 U6547 ( .A1(n6503), .A2(n6629), .B1(n5818), .B2(n6636), .C1(n6411), 
        .C2(n6283), .ZN(U2840) );
  OAI21_X1 U6548 ( .B1(n5821), .B2(n5820), .A(n5819), .ZN(n5822) );
  INV_X1 U6549 ( .A(n5822), .ZN(n6801) );
  AOI22_X1 U6550 ( .A1(n6669), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6809), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5823) );
  OAI21_X1 U6551 ( .B1(n6676), .B2(n5824), .A(n5823), .ZN(n5825) );
  AOI21_X1 U6552 ( .B1(n5826), .B2(n6670), .A(n5825), .ZN(n5827) );
  OAI21_X1 U6553 ( .B1(n6801), .B2(n6952), .A(n5827), .ZN(U2971) );
  NOR2_X1 U6554 ( .A1(n5829), .A2(n5828), .ZN(n5830) );
  OR2_X1 U6555 ( .A1(n5868), .A2(n5830), .ZN(n6403) );
  OAI21_X1 U6556 ( .B1(n5833), .B2(n5832), .A(n5831), .ZN(n6492) );
  INV_X1 U6557 ( .A(n6492), .ZN(n5846) );
  INV_X1 U6558 ( .A(n6402), .ZN(n5834) );
  OAI22_X1 U6559 ( .A1(n6927), .A2(n6400), .B1(n5834), .B2(n6950), .ZN(n5844)
         );
  INV_X1 U6560 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6576) );
  NOR4_X1 U6561 ( .A1(n5836), .A2(n6937), .A3(n6576), .A4(n5835), .ZN(n5837)
         );
  AOI21_X1 U6562 ( .B1(n5837), .B2(n6916), .A(REIP_REG_20__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U6563 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5837), .ZN(n5890) );
  NOR2_X1 U6564 ( .A1(n5890), .A2(n5838), .ZN(n5887) );
  INV_X1 U6565 ( .A(n5887), .ZN(n5839) );
  NAND2_X1 U6566 ( .A1(n6862), .A2(n5839), .ZN(n5840) );
  AND2_X1 U6567 ( .A1(n5840), .A2(n6850), .ZN(n5891) );
  OAI22_X1 U6568 ( .A1(n5842), .A2(n5891), .B1(n5841), .B2(n6907), .ZN(n5843)
         );
  AOI211_X1 U6569 ( .C1(n6946), .C2(n5846), .A(n5844), .B(n5843), .ZN(n5845)
         );
  OAI21_X1 U6570 ( .B1(n6403), .B2(n6077), .A(n5845), .ZN(U2807) );
  AOI22_X1 U6571 ( .A1(n5846), .A2(n4738), .B1(n6281), .B2(EBX_REG_20__SCAN_IN), .ZN(n5847) );
  OAI21_X1 U6572 ( .B1(n6403), .B2(n6283), .A(n5847), .ZN(U2839) );
  AOI22_X1 U6573 ( .A1(n7059), .A2(DATAI_4_), .B1(n7062), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U6574 ( .A1(n7063), .A2(DATAI_20_), .ZN(n5848) );
  OAI211_X1 U6575 ( .C1(n6403), .C2(n3421), .A(n5849), .B(n5848), .ZN(U2871)
         );
  AND2_X1 U6576 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  NOR2_X1 U6577 ( .A1(n5853), .A2(n5852), .ZN(n5878) );
  INV_X1 U6578 ( .A(n5878), .ZN(n5872) );
  AOI21_X1 U6579 ( .B1(n5855), .B2(n5854), .A(n5712), .ZN(n6810) );
  AOI22_X1 U6580 ( .A1(n6810), .A2(n4738), .B1(EBX_REG_16__SCAN_IN), .B2(n6281), .ZN(n5856) );
  OAI21_X1 U6581 ( .B1(n5872), .B2(n6283), .A(n5856), .ZN(U2843) );
  NAND2_X1 U6582 ( .A1(n6939), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5857)
         );
  OAI211_X1 U6583 ( .C1(n5876), .C2(n6950), .A(n5857), .B(n6925), .ZN(n5864)
         );
  AOI22_X1 U6584 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6943), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5858), .ZN(n5862) );
  OAI211_X1 U6585 ( .C1(REIP_REG_15__SCAN_IN), .C2(REIP_REG_16__SCAN_IN), .A(
        n5860), .B(n5859), .ZN(n5861) );
  NAND2_X1 U6586 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  AOI211_X1 U6587 ( .C1(n6810), .C2(n6946), .A(n5864), .B(n5863), .ZN(n5865)
         );
  OAI21_X1 U6588 ( .B1(n5872), .B2(n6077), .A(n5865), .ZN(U2811) );
  OAI21_X1 U6589 ( .B1(n5868), .B2(n5867), .A(n5866), .ZN(n6390) );
  OAI222_X1 U6590 ( .A1(n6390), .A2(n6283), .B1(n6636), .B2(n5869), .C1(n6944), 
        .C2(n6629), .ZN(U2838) );
  AOI22_X1 U6591 ( .A1(n7059), .A2(DATAI_0_), .B1(n7062), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U6592 ( .A1(n7063), .A2(DATAI_16_), .ZN(n5870) );
  OAI211_X1 U6593 ( .C1(n5872), .C2(n3421), .A(n5871), .B(n5870), .ZN(U2875)
         );
  MUX2_X1 U6594 ( .A(n6814), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .S(n6418), 
        .Z(n5873) );
  XNOR2_X1 U6595 ( .A(n5874), .B(n5873), .ZN(n6811) );
  INV_X1 U6596 ( .A(n6811), .ZN(n5880) );
  AOI22_X1 U6597 ( .A1(n6669), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6809), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5875) );
  OAI21_X1 U6598 ( .B1(n6676), .B2(n5876), .A(n5875), .ZN(n5877) );
  AOI21_X1 U6599 ( .B1(n5878), .B2(n6670), .A(n5877), .ZN(n5879) );
  OAI21_X1 U6600 ( .B1(n5880), .B2(n6952), .A(n5879), .ZN(U2970) );
  INV_X1 U6601 ( .A(n5881), .ZN(n6062) );
  INV_X1 U6602 ( .A(n6062), .ZN(n5882) );
  AOI21_X1 U6603 ( .B1(n5883), .B2(n5866), .A(n5882), .ZN(n6387) );
  INV_X1 U6604 ( .A(n6387), .ZN(n6284) );
  INV_X1 U6605 ( .A(n6065), .ZN(n5884) );
  AOI21_X1 U6606 ( .B1(n5886), .B2(n5885), .A(n5884), .ZN(n6484) );
  INV_X1 U6607 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U6608 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5887), .ZN(n5961) );
  NOR3_X1 U6609 ( .A1(n6884), .A2(REIP_REG_22__SCAN_IN), .A3(n5961), .ZN(n5888) );
  AOI21_X1 U6610 ( .B1(n6923), .B2(n6386), .A(n5888), .ZN(n5889) );
  OAI21_X1 U6611 ( .B1(n6907), .B2(n6285), .A(n5889), .ZN(n5894) );
  NOR3_X1 U6612 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5890), .A3(n6899), .ZN(n6942) );
  INV_X1 U6613 ( .A(n5891), .ZN(n6938) );
  OAI21_X1 U6614 ( .B1(n6942), .B2(n6938), .A(REIP_REG_22__SCAN_IN), .ZN(n5892) );
  OAI21_X1 U6615 ( .B1(n6927), .B2(n6384), .A(n5892), .ZN(n5893) );
  AOI211_X1 U6616 ( .C1(n6484), .C2(n6946), .A(n5894), .B(n5893), .ZN(n5895)
         );
  OAI21_X1 U6617 ( .B1(n6284), .B2(n6077), .A(n5895), .ZN(U2805) );
  AOI22_X1 U6618 ( .A1(n7059), .A2(DATAI_6_), .B1(n7062), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U6619 ( .A1(n7063), .A2(DATAI_22_), .ZN(n5896) );
  OAI211_X1 U6620 ( .C1(n6284), .C2(n3421), .A(n5897), .B(n5896), .ZN(U2869)
         );
  INV_X1 U6621 ( .A(n5902), .ZN(n5898) );
  AOI21_X1 U6622 ( .B1(n5898), .B2(n5934), .A(n6959), .ZN(n5906) );
  INV_X1 U6623 ( .A(n5899), .ZN(n5903) );
  NOR2_X1 U6624 ( .A1(n6955), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5901)
         );
  AOI222_X1 U6625 ( .A1(n5903), .A2(n5933), .B1(n5902), .B2(n5901), .C1(n5900), 
        .C2(n7003), .ZN(n5904) );
  OAI22_X1 U6626 ( .A1(n5906), .A2(n5905), .B1(n5904), .B2(n6959), .ZN(U3459)
         );
  AOI21_X1 U6627 ( .B1(n5908), .B2(n5919), .A(n5907), .ZN(n6080) );
  AOI21_X1 U6628 ( .B1(n6669), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5909), 
        .ZN(n5910) );
  OAI21_X1 U6629 ( .B1(n6676), .B2(n5987), .A(n5910), .ZN(n5911) );
  AOI21_X1 U6630 ( .B1(n6080), .B2(n6670), .A(n5911), .ZN(n5912) );
  OAI21_X1 U6631 ( .B1(n5913), .B2(n6952), .A(n5912), .ZN(U2957) );
  AND2_X1 U6632 ( .A1(n5914), .A2(n7007), .ZN(n7022) );
  MUX2_X1 U6633 ( .A(n7022), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(n6521), 
        .Z(n5915) );
  AOI21_X1 U6634 ( .B1(n7077), .B2(n5916), .A(n5915), .ZN(n5917) );
  OAI21_X1 U6635 ( .B1(n5918), .B2(n5929), .A(n5917), .ZN(U3465) );
  OAI21_X1 U6636 ( .B1(n6006), .B2(n5920), .A(n5919), .ZN(n6299) );
  INV_X1 U6637 ( .A(n6299), .ZN(n5995) );
  INV_X1 U6638 ( .A(n5997), .ZN(n5923) );
  AOI21_X1 U6639 ( .B1(n6669), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5921), 
        .ZN(n5922) );
  OAI21_X1 U6640 ( .B1(n6676), .B2(n5923), .A(n5922), .ZN(n5924) );
  AOI21_X1 U6641 ( .B1(n5995), .B2(n6670), .A(n5924), .ZN(n5925) );
  OAI21_X1 U6642 ( .B1(n5926), .B2(n6952), .A(n5925), .ZN(U2958) );
  AOI21_X1 U6643 ( .B1(n7003), .B2(n6969), .A(n6959), .ZN(n5939) );
  INV_X1 U6644 ( .A(n5927), .ZN(n5928) );
  OR2_X1 U6645 ( .A1(n5929), .A2(n5928), .ZN(n5932) );
  NAND2_X1 U6646 ( .A1(n5930), .A2(n5938), .ZN(n5931) );
  AND2_X1 U6647 ( .A1(n5932), .A2(n5931), .ZN(n6971) );
  OAI21_X1 U6648 ( .B1(n6971), .B2(STATE2_REG_3__SCAN_IN), .A(n7011), .ZN(
        n5936) );
  INV_X1 U6649 ( .A(n5933), .ZN(n5935) );
  AOI22_X1 U6650 ( .A1(n5936), .A2(n5935), .B1(n5938), .B2(n5934), .ZN(n5937)
         );
  OAI22_X1 U6651 ( .A1(n5939), .A2(n5938), .B1(n5937), .B2(n6959), .ZN(U3461)
         );
  AND2_X1 U6652 ( .A1(n5940), .A2(n5949), .ZN(n5941) );
  OR2_X1 U6653 ( .A1(n7017), .A2(n5941), .ZN(n5944) );
  NAND2_X1 U6654 ( .A1(n7017), .A2(n5942), .ZN(n5943) );
  OAI211_X1 U6655 ( .C1(n5947), .C2(n5945), .A(n5944), .B(n5943), .ZN(n6988)
         );
  OR2_X1 U6656 ( .A1(n7017), .A2(n5946), .ZN(n5952) );
  NAND2_X1 U6657 ( .A1(n5948), .A2(n5947), .ZN(n5950) );
  NAND2_X1 U6658 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  AND2_X1 U6659 ( .A1(n5952), .A2(n5951), .ZN(n6677) );
  NAND2_X1 U6660 ( .A1(n6692), .A2(n6684), .ZN(n5953) );
  OAI211_X1 U6661 ( .C1(n3685), .C2(n5954), .A(n5953), .B(n7042), .ZN(n6690)
         );
  NAND2_X1 U6662 ( .A1(n6677), .A2(n6690), .ZN(n6991) );
  AND2_X1 U6663 ( .A1(n6991), .A2(n7004), .ZN(n6953) );
  MUX2_X1 U6664 ( .A(MORE_REG_SCAN_IN), .B(n6988), .S(n6953), .Z(U3471) );
  AOI22_X1 U6665 ( .A1(n5956), .A2(EAX_REG_31__SCAN_IN), .B1(n5955), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U6666 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  NAND2_X1 U6667 ( .A1(n3441), .A2(n6947), .ZN(n5977) );
  INV_X1 U6668 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6595) );
  INV_X1 U6669 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6599) );
  NOR2_X1 U6670 ( .A1(n6595), .A2(n6599), .ZN(n5969) );
  INV_X1 U6671 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6583) );
  INV_X1 U6672 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6581) );
  NOR2_X1 U6673 ( .A1(n6581), .A2(n5961), .ZN(n6069) );
  NAND2_X1 U6674 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6069), .ZN(n6034) );
  NOR2_X1 U6675 ( .A1(n6583), .A2(n6034), .ZN(n6038) );
  NAND2_X1 U6676 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6038), .ZN(n5966) );
  INV_X1 U6677 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6588) );
  OR3_X1 U6678 ( .A1(n5962), .A2(n5966), .A3(n6588), .ZN(n5963) );
  NAND2_X1 U6679 ( .A1(n5964), .A2(n5963), .ZN(n6026) );
  INV_X1 U6680 ( .A(n6026), .ZN(n6012) );
  NAND2_X1 U6681 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5967) );
  INV_X1 U6682 ( .A(n5967), .ZN(n5965) );
  NOR2_X1 U6683 ( .A1(n6884), .A2(n5965), .ZN(n5996) );
  NOR2_X1 U6684 ( .A1(n6012), .A2(n5996), .ZN(n5986) );
  OAI21_X1 U6685 ( .B1(n5969), .B2(n6884), .A(n5986), .ZN(n5982) );
  NOR2_X1 U6686 ( .A1(n6884), .A2(n5966), .ZN(n6023) );
  NAND2_X1 U6687 ( .A1(n6023), .A2(REIP_REG_26__SCAN_IN), .ZN(n6015) );
  NOR2_X1 U6688 ( .A1(n6015), .A2(n5967), .ZN(n5978) );
  INV_X1 U6689 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5968) );
  NAND3_X1 U6690 ( .A1(n5978), .A2(n5969), .A3(n5968), .ZN(n5973) );
  NAND3_X1 U6691 ( .A1(n5971), .A2(EBX_REG_31__SCAN_IN), .A3(n5970), .ZN(n5972) );
  OAI211_X1 U6692 ( .C1(n5974), .C2(n6927), .A(n5973), .B(n5972), .ZN(n5975)
         );
  AOI21_X1 U6693 ( .B1(REIP_REG_31__SCAN_IN), .B2(n5982), .A(n5975), .ZN(n5976) );
  OAI211_X1 U6694 ( .C1(n6079), .C2(n6931), .A(n5977), .B(n5976), .ZN(U2796)
         );
  NAND2_X1 U6695 ( .A1(n6328), .A2(n6947), .ZN(n5985) );
  INV_X1 U6696 ( .A(n5978), .ZN(n5991) );
  OAI21_X1 U6697 ( .B1(n5991), .B2(n6595), .A(n6599), .ZN(n5983) );
  AOI22_X1 U6698 ( .A1(n6923), .A2(n6324), .B1(n6939), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5979) );
  OAI21_X1 U6699 ( .B1(n6907), .B2(n5980), .A(n5979), .ZN(n5981) );
  AOI21_X1 U6700 ( .B1(n5983), .B2(n5982), .A(n5981), .ZN(n5984) );
  OAI211_X1 U6701 ( .C1(n6427), .C2(n6931), .A(n5985), .B(n5984), .ZN(U2797)
         );
  NAND2_X1 U6702 ( .A1(n6080), .A2(n6947), .ZN(n5994) );
  INV_X1 U6703 ( .A(n5986), .ZN(n6001) );
  OAI22_X1 U6704 ( .A1(n6927), .A2(n5988), .B1(n5987), .B2(n6950), .ZN(n5989)
         );
  AOI21_X1 U6705 ( .B1(n6943), .B2(EBX_REG_29__SCAN_IN), .A(n5989), .ZN(n5990)
         );
  OAI21_X1 U6706 ( .B1(n5991), .B2(REIP_REG_29__SCAN_IN), .A(n5990), .ZN(n5992) );
  AOI21_X1 U6707 ( .B1(REIP_REG_29__SCAN_IN), .B2(n6001), .A(n5992), .ZN(n5993) );
  OAI211_X1 U6708 ( .C1(n6931), .C2(n6081), .A(n5994), .B(n5993), .ZN(U2798)
         );
  NAND2_X1 U6709 ( .A1(n5995), .A2(n6947), .ZN(n6003) );
  INV_X1 U6710 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6084) );
  NAND3_X1 U6711 ( .A1(n6026), .A2(REIP_REG_27__SCAN_IN), .A3(n5996), .ZN(
        n5999) );
  AOI22_X1 U6712 ( .A1(n6923), .A2(n5997), .B1(n6939), .B2(
        PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5998) );
  OAI211_X1 U6713 ( .C1(n6084), .C2(n6907), .A(n5999), .B(n5998), .ZN(n6000)
         );
  AOI21_X1 U6714 ( .B1(n6001), .B2(REIP_REG_28__SCAN_IN), .A(n6000), .ZN(n6002) );
  OAI211_X1 U6715 ( .C1(n6931), .C2(n6083), .A(n6003), .B(n6002), .ZN(U2799)
         );
  AOI21_X1 U6716 ( .B1(n6007), .B2(n6018), .A(n6006), .ZN(n6336) );
  INV_X1 U6717 ( .A(n6336), .ZN(n6302) );
  XNOR2_X1 U6718 ( .A(n6020), .B(n6008), .ZN(n6443) );
  INV_X1 U6719 ( .A(n6009), .ZN(n6334) );
  OAI22_X1 U6720 ( .A1(n6927), .A2(n6010), .B1(n6334), .B2(n6950), .ZN(n6011)
         );
  AOI21_X1 U6721 ( .B1(n6943), .B2(EBX_REG_27__SCAN_IN), .A(n6011), .ZN(n6014)
         );
  NAND2_X1 U6722 ( .A1(n6012), .A2(REIP_REG_27__SCAN_IN), .ZN(n6013) );
  OAI211_X1 U6723 ( .C1(n6015), .C2(REIP_REG_27__SCAN_IN), .A(n6014), .B(n6013), .ZN(n6016) );
  AOI21_X1 U6724 ( .B1(n6443), .B2(n6946), .A(n6016), .ZN(n6017) );
  OAI21_X1 U6725 ( .B1(n6302), .B2(n6077), .A(n6017), .ZN(U2800) );
  AOI21_X1 U6726 ( .B1(n6019), .B2(n6032), .A(n6005), .ZN(n6345) );
  INV_X1 U6727 ( .A(n6345), .ZN(n6305) );
  INV_X1 U6728 ( .A(n6020), .ZN(n6021) );
  AOI21_X1 U6729 ( .B1(n6022), .B2(n6042), .A(n6021), .ZN(n6454) );
  NOR2_X1 U6730 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6023), .ZN(n6025) );
  OAI22_X1 U6731 ( .A1(n6026), .A2(n6025), .B1(n6024), .B2(n6927), .ZN(n6030)
         );
  INV_X1 U6732 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6028) );
  INV_X1 U6733 ( .A(n6027), .ZN(n6343) );
  OAI22_X1 U6734 ( .A1(n6907), .A2(n6028), .B1(n6343), .B2(n6950), .ZN(n6029)
         );
  AOI211_X1 U6735 ( .C1(n6454), .C2(n6946), .A(n6030), .B(n6029), .ZN(n6031)
         );
  OAI21_X1 U6736 ( .B1(n6305), .B2(n6077), .A(n6031), .ZN(U2801) );
  OAI21_X1 U6737 ( .B1(n6049), .B2(n6033), .A(n6032), .ZN(n6351) );
  INV_X1 U6738 ( .A(n6034), .ZN(n6057) );
  AOI21_X1 U6739 ( .B1(n6850), .B2(n6057), .A(n6035), .ZN(n6068) );
  INV_X1 U6740 ( .A(n6353), .ZN(n6036) );
  AOI22_X1 U6741 ( .A1(n6923), .A2(n6036), .B1(n6939), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U6742 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n6037) );
  OAI211_X1 U6743 ( .C1(REIP_REG_25__SCAN_IN), .C2(n6038), .A(n6862), .B(n6037), .ZN(n6039) );
  OAI211_X1 U6744 ( .C1(n6907), .C2(n6279), .A(n6040), .B(n6039), .ZN(n6045)
         );
  OAI21_X1 U6745 ( .B1(n6052), .B2(n6043), .A(n6042), .ZN(n6458) );
  NOR2_X1 U6746 ( .A1(n6458), .A2(n6931), .ZN(n6044) );
  AOI211_X1 U6747 ( .C1(REIP_REG_25__SCAN_IN), .C2(n6068), .A(n6045), .B(n6044), .ZN(n6046) );
  OAI21_X1 U6748 ( .B1(n6351), .B2(n6077), .A(n6046), .ZN(U2802) );
  INV_X1 U6749 ( .A(n6047), .ZN(n6051) );
  INV_X1 U6750 ( .A(n6048), .ZN(n6050) );
  AOI21_X1 U6751 ( .B1(n6051), .B2(n6050), .A(n6049), .ZN(n6369) );
  INV_X1 U6752 ( .A(n6369), .ZN(n6310) );
  INV_X1 U6753 ( .A(n6067), .ZN(n6053) );
  AOI21_X1 U6754 ( .B1(n6054), .B2(n6053), .A(n6052), .ZN(n6471) );
  AOI22_X1 U6755 ( .A1(EBX_REG_24__SCAN_IN), .A2(n6943), .B1(
        REIP_REG_24__SCAN_IN), .B2(n6068), .ZN(n6055) );
  OAI21_X1 U6756 ( .B1(n6056), .B2(n6927), .A(n6055), .ZN(n6060) );
  NAND3_X1 U6757 ( .A1(n6862), .A2(n6057), .A3(n6583), .ZN(n6058) );
  OAI21_X1 U6758 ( .B1(n6950), .B2(n6367), .A(n6058), .ZN(n6059) );
  AOI211_X1 U6759 ( .C1(n6471), .C2(n6946), .A(n6060), .B(n6059), .ZN(n6061)
         );
  OAI21_X1 U6760 ( .B1(n6310), .B2(n6077), .A(n6061), .ZN(U2803) );
  AOI21_X1 U6761 ( .B1(n6063), .B2(n6062), .A(n6048), .ZN(n6378) );
  INV_X1 U6762 ( .A(n6378), .ZN(n6313) );
  AND2_X1 U6763 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  NOR2_X1 U6764 ( .A1(n6067), .A2(n6066), .ZN(n6479) );
  INV_X1 U6765 ( .A(n6068), .ZN(n6074) );
  AOI21_X1 U6766 ( .B1(n6862), .B2(n6069), .A(REIP_REG_23__SCAN_IN), .ZN(n6073) );
  OAI22_X1 U6767 ( .A1(n6927), .A2(n6070), .B1(n6376), .B2(n6950), .ZN(n6071)
         );
  AOI21_X1 U6768 ( .B1(n6943), .B2(EBX_REG_23__SCAN_IN), .A(n6071), .ZN(n6072)
         );
  OAI21_X1 U6769 ( .B1(n6074), .B2(n6073), .A(n6072), .ZN(n6075) );
  AOI21_X1 U6770 ( .B1(n6479), .B2(n6946), .A(n6075), .ZN(n6076) );
  OAI21_X1 U6771 ( .B1(n6313), .B2(n6077), .A(n6076), .ZN(U2804) );
  OAI22_X1 U6772 ( .A1(n6079), .A2(n6629), .B1(n6078), .B2(n6636), .ZN(U2828)
         );
  INV_X1 U6773 ( .A(n6080), .ZN(n6296) );
  OAI222_X1 U6774 ( .A1(n6082), .A2(n6636), .B1(n6629), .B2(n6081), .C1(n6296), 
        .C2(n6283), .ZN(U2830) );
  OAI222_X1 U6775 ( .A1(n6084), .A2(n6636), .B1(n6629), .B2(n6083), .C1(n6299), 
        .C2(n6283), .ZN(U2831) );
  INV_X1 U6776 ( .A(n6283), .ZN(n6634) );
  AOI222_X1 U6777 ( .A1(n6443), .A2(n4738), .B1(n6281), .B2(
        EBX_REG_27__SCAN_IN), .C1(n6634), .C2(n6336), .ZN(n6277) );
  INV_X1 U6778 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6593) );
  OAI22_X1 U6779 ( .A1(n6593), .A2(keyinput_118), .B1(keyinput_117), .B2(
        REIP_REG_29__SCAN_IN), .ZN(n6085) );
  AOI221_X1 U6780 ( .B1(n6593), .B2(keyinput_118), .C1(REIP_REG_29__SCAN_IN), 
        .C2(keyinput_117), .A(n6085), .ZN(n6161) );
  INV_X1 U6781 ( .A(keyinput_112), .ZN(n6154) );
  INV_X1 U6782 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6617) );
  INV_X1 U6783 ( .A(keyinput_111), .ZN(n6152) );
  INV_X1 U6784 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6151) );
  INV_X1 U6785 ( .A(MORE_REG_SCAN_IN), .ZN(n6986) );
  OAI22_X1 U6786 ( .A1(n6986), .A2(keyinput_108), .B1(STATEBS16_REG_SCAN_IN), 
        .B2(keyinput_107), .ZN(n6086) );
  AOI221_X1 U6787 ( .B1(n6986), .B2(keyinput_108), .C1(keyinput_107), .C2(
        STATEBS16_REG_SCAN_IN), .A(n6086), .ZN(n6149) );
  XOR2_X1 U6788 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_96), .Z(n6139) );
  OAI22_X1 U6789 ( .A1(n6089), .A2(keyinput_94), .B1(n6088), .B2(keyinput_93), 
        .ZN(n6087) );
  AOI221_X1 U6790 ( .B1(n6089), .B2(keyinput_94), .C1(keyinput_93), .C2(n6088), 
        .A(n6087), .ZN(n6135) );
  AOI22_X1 U6791 ( .A1(n6091), .A2(keyinput_89), .B1(keyinput_90), .B2(n6184), 
        .ZN(n6090) );
  OAI221_X1 U6792 ( .B1(n6091), .B2(keyinput_89), .C1(n6184), .C2(keyinput_90), 
        .A(n6090), .ZN(n6129) );
  OAI22_X1 U6793 ( .A1(n6093), .A2(keyinput_87), .B1(DATAI_7_), .B2(
        keyinput_88), .ZN(n6092) );
  AOI221_X1 U6794 ( .B1(n6093), .B2(keyinput_87), .C1(keyinput_88), .C2(
        DATAI_7_), .A(n6092), .ZN(n6128) );
  OAI22_X1 U6795 ( .A1(DATAI_11_), .A2(keyinput_84), .B1(DATAI_10_), .B2(
        keyinput_85), .ZN(n6094) );
  AOI221_X1 U6796 ( .B1(DATAI_11_), .B2(keyinput_84), .C1(keyinput_85), .C2(
        DATAI_10_), .A(n6094), .ZN(n6123) );
  INV_X1 U6797 ( .A(keyinput_83), .ZN(n6121) );
  INV_X1 U6798 ( .A(DATAI_16_), .ZN(n6214) );
  OAI22_X1 U6799 ( .A1(n6214), .A2(keyinput_79), .B1(n6213), .B2(keyinput_80), 
        .ZN(n6095) );
  AOI221_X1 U6800 ( .B1(n6214), .B2(keyinput_79), .C1(keyinput_80), .C2(n6213), 
        .A(n6095), .ZN(n6118) );
  INV_X1 U6801 ( .A(DATAI_20_), .ZN(n6208) );
  OAI22_X1 U6802 ( .A1(n6208), .A2(keyinput_75), .B1(DATAI_19_), .B2(
        keyinput_76), .ZN(n6096) );
  AOI221_X1 U6803 ( .B1(n6208), .B2(keyinput_75), .C1(keyinput_76), .C2(
        DATAI_19_), .A(n6096), .ZN(n6113) );
  OAI22_X1 U6804 ( .A1(DATAI_23_), .A2(keyinput_72), .B1(DATAI_22_), .B2(
        keyinput_73), .ZN(n6097) );
  AOI221_X1 U6805 ( .B1(DATAI_23_), .B2(keyinput_72), .C1(keyinput_73), .C2(
        DATAI_22_), .A(n6097), .ZN(n6110) );
  INV_X1 U6806 ( .A(DATAI_24_), .ZN(n6203) );
  INV_X1 U6807 ( .A(keyinput_71), .ZN(n6108) );
  INV_X1 U6808 ( .A(keyinput_70), .ZN(n6106) );
  INV_X1 U6809 ( .A(DATAI_25_), .ZN(n6200) );
  OAI22_X1 U6810 ( .A1(DATAI_27_), .A2(keyinput_68), .B1(DATAI_28_), .B2(
        keyinput_67), .ZN(n6098) );
  AOI221_X1 U6811 ( .B1(DATAI_27_), .B2(keyinput_68), .C1(keyinput_67), .C2(
        DATAI_28_), .A(n6098), .ZN(n6103) );
  INV_X1 U6812 ( .A(DATAI_29_), .ZN(n6194) );
  INV_X1 U6813 ( .A(keyinput_66), .ZN(n6101) );
  AOI22_X1 U6814 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(DATAI_31_), .B2(
        keyinput_64), .ZN(n6099) );
  OAI221_X1 U6815 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n6099), .ZN(n6100) );
  OAI221_X1 U6816 ( .B1(DATAI_29_), .B2(keyinput_66), .C1(n6194), .C2(n6101), 
        .A(n6100), .ZN(n6102) );
  AOI22_X1 U6817 ( .A1(n6103), .A2(n6102), .B1(keyinput_69), .B2(DATAI_26_), 
        .ZN(n6104) );
  OAI21_X1 U6818 ( .B1(keyinput_69), .B2(DATAI_26_), .A(n6104), .ZN(n6105) );
  OAI221_X1 U6819 ( .B1(DATAI_25_), .B2(n6106), .C1(n6200), .C2(keyinput_70), 
        .A(n6105), .ZN(n6107) );
  OAI221_X1 U6820 ( .B1(DATAI_24_), .B2(keyinput_71), .C1(n6203), .C2(n6108), 
        .A(n6107), .ZN(n6109) );
  AOI22_X1 U6821 ( .A1(n6110), .A2(n6109), .B1(keyinput_74), .B2(DATAI_21_), 
        .ZN(n6111) );
  OAI21_X1 U6822 ( .B1(keyinput_74), .B2(DATAI_21_), .A(n6111), .ZN(n6112) );
  AOI22_X1 U6823 ( .A1(keyinput_77), .A2(DATAI_18_), .B1(n6113), .B2(n6112), 
        .ZN(n6116) );
  AOI22_X1 U6824 ( .A1(DATAI_17_), .A2(keyinput_78), .B1(DATAI_14_), .B2(
        keyinput_81), .ZN(n6114) );
  OAI221_X1 U6825 ( .B1(DATAI_17_), .B2(keyinput_78), .C1(DATAI_14_), .C2(
        keyinput_81), .A(n6114), .ZN(n6115) );
  AOI221_X1 U6826 ( .B1(DATAI_18_), .B2(n6116), .C1(keyinput_77), .C2(n6116), 
        .A(n6115), .ZN(n6117) );
  AOI22_X1 U6827 ( .A1(n6118), .A2(n6117), .B1(keyinput_82), .B2(DATAI_13_), 
        .ZN(n6119) );
  OAI21_X1 U6828 ( .B1(keyinput_82), .B2(DATAI_13_), .A(n6119), .ZN(n6120) );
  OAI221_X1 U6829 ( .B1(DATAI_12_), .B2(n6121), .C1(n6226), .C2(keyinput_83), 
        .A(n6120), .ZN(n6122) );
  AOI22_X1 U6830 ( .A1(keyinput_86), .A2(n6230), .B1(n6123), .B2(n6122), .ZN(
        n6124) );
  OAI21_X1 U6831 ( .B1(n6230), .B2(keyinput_86), .A(n6124), .ZN(n6127) );
  OAI22_X1 U6832 ( .A1(DATAI_3_), .A2(keyinput_92), .B1(DATAI_4_), .B2(
        keyinput_91), .ZN(n6125) );
  AOI221_X1 U6833 ( .B1(DATAI_3_), .B2(keyinput_92), .C1(keyinput_91), .C2(
        DATAI_4_), .A(n6125), .ZN(n6126) );
  OAI221_X1 U6834 ( .B1(n6129), .B2(n6128), .C1(n6129), .C2(n6127), .A(n6126), 
        .ZN(n6134) );
  AOI22_X1 U6835 ( .A1(keyinput_97), .A2(NA_N), .B1(n6177), .B2(keyinput_95), 
        .ZN(n6130) );
  OAI221_X1 U6836 ( .B1(keyinput_97), .B2(NA_N), .C1(n6177), .C2(keyinput_95), 
        .A(n6130), .ZN(n6133) );
  INV_X1 U6837 ( .A(BS16_N), .ZN(n6519) );
  AOI22_X1 U6838 ( .A1(READY_N), .A2(keyinput_99), .B1(n6519), .B2(keyinput_98), .ZN(n6131) );
  OAI221_X1 U6839 ( .B1(READY_N), .B2(keyinput_99), .C1(n6519), .C2(
        keyinput_98), .A(n6131), .ZN(n6132) );
  AOI211_X1 U6840 ( .C1(n6135), .C2(n6134), .A(n6133), .B(n6132), .ZN(n6138)
         );
  INV_X1 U6841 ( .A(HOLD), .ZN(n7033) );
  AOI22_X1 U6842 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_101), .B1(n7033), 
        .B2(keyinput_100), .ZN(n6136) );
  OAI221_X1 U6843 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_101), .C1(n7033), .C2(keyinput_100), .A(n6136), .ZN(n6137) );
  AOI21_X1 U6844 ( .B1(n6139), .B2(n6138), .A(n6137), .ZN(n6145) );
  INV_X1 U6845 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6679) );
  AOI22_X1 U6846 ( .A1(keyinput_102), .A2(ADS_N_REG_SCAN_IN), .B1(n6679), .B2(
        keyinput_103), .ZN(n6140) );
  OAI221_X1 U6847 ( .B1(keyinput_102), .B2(ADS_N_REG_SCAN_IN), .C1(n6679), 
        .C2(keyinput_103), .A(n6140), .ZN(n6144) );
  INV_X1 U6848 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7035) );
  OAI22_X1 U6849 ( .A1(n7035), .A2(keyinput_106), .B1(D_C_N_REG_SCAN_IN), .B2(
        keyinput_105), .ZN(n6141) );
  AOI221_X1 U6850 ( .B1(n7035), .B2(keyinput_106), .C1(keyinput_105), .C2(
        D_C_N_REG_SCAN_IN), .A(n6141), .ZN(n6143) );
  XNOR2_X1 U6851 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_104), .ZN(n6142) );
  OAI211_X1 U6852 ( .C1(n6145), .C2(n6144), .A(n6143), .B(n6142), .ZN(n6148)
         );
  AOI22_X1 U6853 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_109), .B1(
        W_R_N_REG_SCAN_IN), .B2(keyinput_110), .ZN(n6146) );
  OAI221_X1 U6854 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_109), .C1(
        W_R_N_REG_SCAN_IN), .C2(keyinput_110), .A(n6146), .ZN(n6147) );
  AOI21_X1 U6855 ( .B1(n6149), .B2(n6148), .A(n6147), .ZN(n6150) );
  AOI221_X1 U6856 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(n6152), .C1(n6151), 
        .C2(keyinput_111), .A(n6150), .ZN(n6153) );
  AOI221_X1 U6857 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6154), .C1(n6617), 
        .C2(keyinput_112), .A(n6153), .ZN(n6159) );
  AOI22_X1 U6858 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_114), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_113), .ZN(n6155) );
  OAI221_X1 U6859 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_114), .C1(
        BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_113), .A(n6155), .ZN(n6158)
         );
  OAI22_X1 U6860 ( .A1(n6599), .A2(keyinput_116), .B1(REIP_REG_31__SCAN_IN), 
        .B2(keyinput_115), .ZN(n6156) );
  AOI221_X1 U6861 ( .B1(n6599), .B2(keyinput_116), .C1(keyinput_115), .C2(
        REIP_REG_31__SCAN_IN), .A(n6156), .ZN(n6157) );
  OAI21_X1 U6862 ( .B1(n6159), .B2(n6158), .A(n6157), .ZN(n6160) );
  AOI22_X1 U6863 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput_119), .B1(n6161), 
        .B2(n6160), .ZN(n6164) );
  AOI22_X1 U6864 ( .A1(REIP_REG_23__SCAN_IN), .A2(keyinput_123), .B1(n6588), 
        .B2(keyinput_120), .ZN(n6162) );
  OAI221_X1 U6865 ( .B1(REIP_REG_23__SCAN_IN), .B2(keyinput_123), .C1(n6588), 
        .C2(keyinput_120), .A(n6162), .ZN(n6163) );
  AOI221_X1 U6866 ( .B1(REIP_REG_27__SCAN_IN), .B2(n6164), .C1(keyinput_119), 
        .C2(n6164), .A(n6163), .ZN(n6171) );
  INV_X1 U6867 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6586) );
  OAI22_X1 U6868 ( .A1(n6583), .A2(keyinput_122), .B1(n6586), .B2(keyinput_121), .ZN(n6165) );
  AOI221_X1 U6869 ( .B1(n6583), .B2(keyinput_122), .C1(keyinput_121), .C2(
        n6586), .A(n6165), .ZN(n6170) );
  INV_X1 U6870 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6579) );
  AOI22_X1 U6871 ( .A1(n6579), .A2(keyinput_125), .B1(n6581), .B2(keyinput_124), .ZN(n6166) );
  OAI221_X1 U6872 ( .B1(n6579), .B2(keyinput_125), .C1(n6581), .C2(
        keyinput_124), .A(n6166), .ZN(n6169) );
  AOI22_X1 U6873 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput_127), .B1(
        REIP_REG_20__SCAN_IN), .B2(keyinput_126), .ZN(n6167) );
  OAI221_X1 U6874 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_127), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput_126), .A(n6167), .ZN(n6168) );
  AOI211_X1 U6875 ( .C1(n6171), .C2(n6170), .A(n6169), .B(n6168), .ZN(n6275)
         );
  INV_X1 U6876 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6262) );
  AOI22_X1 U6877 ( .A1(n6593), .A2(keyinput_54), .B1(n6595), .B2(keyinput_53), 
        .ZN(n6172) );
  OAI221_X1 U6878 ( .B1(n6593), .B2(keyinput_54), .C1(n6595), .C2(keyinput_53), 
        .A(n6172), .ZN(n6260) );
  OAI22_X1 U6879 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_49), .B1(
        keyinput_50), .B2(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6173) );
  AOI221_X1 U6880 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_49), .C1(
        BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_50), .A(n6173), .ZN(n6258) );
  INV_X1 U6881 ( .A(keyinput_48), .ZN(n6254) );
  INV_X1 U6882 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6683) );
  OAI22_X1 U6883 ( .A1(n6683), .A2(keyinput_46), .B1(n5023), .B2(keyinput_45), 
        .ZN(n6174) );
  AOI221_X1 U6884 ( .B1(n6683), .B2(keyinput_46), .C1(keyinput_45), .C2(n5023), 
        .A(n6174), .ZN(n6251) );
  OAI22_X1 U6885 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_39), .B1(
        keyinput_38), .B2(ADS_N_REG_SCAN_IN), .ZN(n6175) );
  AOI221_X1 U6886 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_39), .C1(
        ADS_N_REG_SCAN_IN), .C2(keyinput_38), .A(n6175), .ZN(n6243) );
  INV_X1 U6887 ( .A(NA_N), .ZN(n7040) );
  AOI22_X1 U6888 ( .A1(n7040), .A2(keyinput_33), .B1(keyinput_31), .B2(n6177), 
        .ZN(n6176) );
  OAI221_X1 U6889 ( .B1(n7040), .B2(keyinput_33), .C1(n6177), .C2(keyinput_31), 
        .A(n6176), .ZN(n6180) );
  AOI22_X1 U6890 ( .A1(n6519), .A2(keyinput_34), .B1(n7042), .B2(keyinput_35), 
        .ZN(n6178) );
  OAI221_X1 U6891 ( .B1(n6519), .B2(keyinput_34), .C1(n7042), .C2(keyinput_35), 
        .A(n6178), .ZN(n6179) );
  AOI211_X1 U6892 ( .C1(keyinput_32), .C2(MEMORYFETCH_REG_SCAN_IN), .A(n6180), 
        .B(n6179), .ZN(n6181) );
  OAI21_X1 U6893 ( .B1(keyinput_32), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n6181), 
        .ZN(n6241) );
  OAI22_X1 U6894 ( .A1(DATAI_1_), .A2(keyinput_30), .B1(DATAI_2_), .B2(
        keyinput_29), .ZN(n6182) );
  AOI221_X1 U6895 ( .B1(DATAI_1_), .B2(keyinput_30), .C1(keyinput_29), .C2(
        DATAI_2_), .A(n6182), .ZN(n6240) );
  AOI22_X1 U6896 ( .A1(DATAI_6_), .A2(keyinput_25), .B1(n6184), .B2(
        keyinput_26), .ZN(n6183) );
  OAI221_X1 U6897 ( .B1(DATAI_6_), .B2(keyinput_25), .C1(n6184), .C2(
        keyinput_26), .A(n6183), .ZN(n6236) );
  OAI22_X1 U6898 ( .A1(n6186), .A2(keyinput_24), .B1(keyinput_23), .B2(
        DATAI_8_), .ZN(n6185) );
  AOI221_X1 U6899 ( .B1(n6186), .B2(keyinput_24), .C1(DATAI_8_), .C2(
        keyinput_23), .A(n6185), .ZN(n6235) );
  OAI22_X1 U6900 ( .A1(DATAI_11_), .A2(keyinput_20), .B1(DATAI_10_), .B2(
        keyinput_21), .ZN(n6187) );
  AOI221_X1 U6901 ( .B1(DATAI_11_), .B2(keyinput_20), .C1(keyinput_21), .C2(
        DATAI_10_), .A(n6187), .ZN(n6228) );
  INV_X1 U6902 ( .A(keyinput_19), .ZN(n6225) );
  INV_X1 U6903 ( .A(keyinput_18), .ZN(n6223) );
  OAI22_X1 U6904 ( .A1(DATAI_23_), .A2(keyinput_8), .B1(DATAI_22_), .B2(
        keyinput_9), .ZN(n6188) );
  AOI221_X1 U6905 ( .B1(DATAI_23_), .B2(keyinput_8), .C1(keyinput_9), .C2(
        DATAI_22_), .A(n6188), .ZN(n6206) );
  INV_X1 U6906 ( .A(keyinput_7), .ZN(n6204) );
  INV_X1 U6907 ( .A(keyinput_6), .ZN(n6201) );
  INV_X1 U6908 ( .A(DATAI_27_), .ZN(n6191) );
  INV_X1 U6909 ( .A(DATAI_28_), .ZN(n6190) );
  OAI22_X1 U6910 ( .A1(n6191), .A2(keyinput_4), .B1(n6190), .B2(keyinput_3), 
        .ZN(n6189) );
  AOI221_X1 U6911 ( .B1(n6191), .B2(keyinput_4), .C1(keyinput_3), .C2(n6190), 
        .A(n6189), .ZN(n6197) );
  INV_X1 U6912 ( .A(keyinput_2), .ZN(n6195) );
  AOI22_X1 U6913 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(DATAI_31_), .B2(
        keyinput_0), .ZN(n6192) );
  OAI221_X1 U6914 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n6192), .ZN(n6193) );
  OAI221_X1 U6915 ( .B1(DATAI_29_), .B2(n6195), .C1(n6194), .C2(keyinput_2), 
        .A(n6193), .ZN(n6196) );
  AOI22_X1 U6916 ( .A1(n6197), .A2(n6196), .B1(keyinput_5), .B2(DATAI_26_), 
        .ZN(n6198) );
  OAI21_X1 U6917 ( .B1(keyinput_5), .B2(DATAI_26_), .A(n6198), .ZN(n6199) );
  OAI221_X1 U6918 ( .B1(DATAI_25_), .B2(n6201), .C1(n6200), .C2(keyinput_6), 
        .A(n6199), .ZN(n6202) );
  OAI221_X1 U6919 ( .B1(DATAI_24_), .B2(n6204), .C1(n6203), .C2(keyinput_7), 
        .A(n6202), .ZN(n6205) );
  AOI22_X1 U6920 ( .A1(DATAI_21_), .A2(keyinput_10), .B1(n6206), .B2(n6205), 
        .ZN(n6211) );
  INV_X1 U6921 ( .A(DATAI_19_), .ZN(n6209) );
  AOI22_X1 U6922 ( .A1(n6209), .A2(keyinput_12), .B1(keyinput_11), .B2(n6208), 
        .ZN(n6207) );
  OAI221_X1 U6923 ( .B1(n6209), .B2(keyinput_12), .C1(n6208), .C2(keyinput_11), 
        .A(n6207), .ZN(n6210) );
  AOI221_X1 U6924 ( .B1(DATAI_21_), .B2(n6211), .C1(keyinput_10), .C2(n6211), 
        .A(n6210), .ZN(n6220) );
  XOR2_X1 U6925 ( .A(DATAI_18_), .B(keyinput_13), .Z(n6219) );
  OAI22_X1 U6926 ( .A1(n6214), .A2(keyinput_15), .B1(n6213), .B2(keyinput_16), 
        .ZN(n6212) );
  AOI221_X1 U6927 ( .B1(n6214), .B2(keyinput_15), .C1(keyinput_16), .C2(n6213), 
        .A(n6212), .ZN(n6218) );
  OAI22_X1 U6928 ( .A1(n6216), .A2(keyinput_17), .B1(DATAI_17_), .B2(
        keyinput_14), .ZN(n6215) );
  AOI221_X1 U6929 ( .B1(n6216), .B2(keyinput_17), .C1(keyinput_14), .C2(
        DATAI_17_), .A(n6215), .ZN(n6217) );
  OAI211_X1 U6930 ( .C1(n6220), .C2(n6219), .A(n6218), .B(n6217), .ZN(n6221)
         );
  OAI221_X1 U6931 ( .B1(DATAI_13_), .B2(n6223), .C1(n6222), .C2(keyinput_18), 
        .A(n6221), .ZN(n6224) );
  OAI221_X1 U6932 ( .B1(DATAI_12_), .B2(keyinput_19), .C1(n6226), .C2(n6225), 
        .A(n6224), .ZN(n6227) );
  AOI22_X1 U6933 ( .A1(keyinput_22), .A2(n6230), .B1(n6228), .B2(n6227), .ZN(
        n6229) );
  OAI21_X1 U6934 ( .B1(n6230), .B2(keyinput_22), .A(n6229), .ZN(n6234) );
  OAI22_X1 U6935 ( .A1(n6232), .A2(keyinput_28), .B1(DATAI_4_), .B2(
        keyinput_27), .ZN(n6231) );
  AOI221_X1 U6936 ( .B1(n6232), .B2(keyinput_28), .C1(keyinput_27), .C2(
        DATAI_4_), .A(n6231), .ZN(n6233) );
  OAI221_X1 U6937 ( .B1(n6236), .B2(n6235), .C1(n6236), .C2(n6234), .A(n6233), 
        .ZN(n6239) );
  OAI22_X1 U6938 ( .A1(HOLD), .A2(keyinput_36), .B1(keyinput_37), .B2(
        READREQUEST_REG_SCAN_IN), .ZN(n6237) );
  AOI221_X1 U6939 ( .B1(HOLD), .B2(keyinput_36), .C1(READREQUEST_REG_SCAN_IN), 
        .C2(keyinput_37), .A(n6237), .ZN(n6238) );
  OAI221_X1 U6940 ( .B1(n6241), .B2(n6240), .C1(n6241), .C2(n6239), .A(n6238), 
        .ZN(n6242) );
  AOI22_X1 U6941 ( .A1(n6243), .A2(n6242), .B1(keyinput_42), .B2(n7035), .ZN(
        n6244) );
  OAI21_X1 U6942 ( .B1(keyinput_42), .B2(n7035), .A(n6244), .ZN(n6249) );
  AOI22_X1 U6943 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_41), .B1(
        M_IO_N_REG_SCAN_IN), .B2(keyinput_40), .ZN(n6245) );
  OAI221_X1 U6944 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_41), .C1(
        M_IO_N_REG_SCAN_IN), .C2(keyinput_40), .A(n6245), .ZN(n6248) );
  OAI22_X1 U6945 ( .A1(n7028), .A2(keyinput_43), .B1(MORE_REG_SCAN_IN), .B2(
        keyinput_44), .ZN(n6246) );
  AOI221_X1 U6946 ( .B1(n7028), .B2(keyinput_43), .C1(keyinput_44), .C2(
        MORE_REG_SCAN_IN), .A(n6246), .ZN(n6247) );
  OAI21_X1 U6947 ( .B1(n6249), .B2(n6248), .A(n6247), .ZN(n6250) );
  AOI22_X1 U6948 ( .A1(n6251), .A2(n6250), .B1(keyinput_47), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n6252) );
  OAI21_X1 U6949 ( .B1(keyinput_47), .B2(BYTEENABLE_REG_0__SCAN_IN), .A(n6252), 
        .ZN(n6253) );
  OAI221_X1 U6950 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_48), .C1(
        n6617), .C2(n6254), .A(n6253), .ZN(n6257) );
  AOI22_X1 U6951 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_51), .B1(n6599), 
        .B2(keyinput_52), .ZN(n6255) );
  OAI221_X1 U6952 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_51), .C1(n6599), 
        .C2(keyinput_52), .A(n6255), .ZN(n6256) );
  AOI21_X1 U6953 ( .B1(n6258), .B2(n6257), .A(n6256), .ZN(n6259) );
  OAI22_X1 U6954 ( .A1(keyinput_55), .A2(n6262), .B1(n6260), .B2(n6259), .ZN(
        n6261) );
  AOI21_X1 U6955 ( .B1(keyinput_55), .B2(n6262), .A(n6261), .ZN(n6267) );
  AOI22_X1 U6956 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_57), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_58), .ZN(n6263) );
  OAI221_X1 U6957 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_57), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_58), .A(n6263), .ZN(n6266) );
  AOI22_X1 U6958 ( .A1(REIP_REG_26__SCAN_IN), .A2(keyinput_56), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_59), .ZN(n6264) );
  OAI221_X1 U6959 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_56), .C1(
        REIP_REG_23__SCAN_IN), .C2(keyinput_59), .A(n6264), .ZN(n6265) );
  NOR3_X1 U6960 ( .A1(n6267), .A2(n6266), .A3(n6265), .ZN(n6274) );
  OAI22_X1 U6961 ( .A1(n6581), .A2(keyinput_60), .B1(REIP_REG_20__SCAN_IN), 
        .B2(keyinput_62), .ZN(n6273) );
  AOI22_X1 U6962 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput_62), .B1(n6579), 
        .B2(keyinput_61), .ZN(n6269) );
  AOI22_X1 U6963 ( .A1(n6581), .A2(keyinput_60), .B1(keyinput_63), .B2(n6576), 
        .ZN(n6268) );
  OAI211_X1 U6964 ( .C1(n6579), .C2(keyinput_61), .A(n6269), .B(n6268), .ZN(
        n6270) );
  INV_X1 U6965 ( .A(n6270), .ZN(n6271) );
  OAI21_X1 U6966 ( .B1(keyinput_63), .B2(n6576), .A(n6271), .ZN(n6272) );
  NOR4_X1 U6967 ( .A1(n6275), .A2(n6274), .A3(n6273), .A4(n6272), .ZN(n6276)
         );
  XNOR2_X1 U6968 ( .A(n6277), .B(n6276), .ZN(U2832) );
  AOI22_X1 U6969 ( .A1(n6454), .A2(n4738), .B1(n6281), .B2(EBX_REG_26__SCAN_IN), .ZN(n6278) );
  OAI21_X1 U6970 ( .B1(n6305), .B2(n6283), .A(n6278), .ZN(U2833) );
  OAI222_X1 U6971 ( .A1(n6458), .A2(n6629), .B1(n6279), .B2(n6636), .C1(n6351), 
        .C2(n6283), .ZN(U2834) );
  AOI22_X1 U6972 ( .A1(n6471), .A2(n4738), .B1(EBX_REG_24__SCAN_IN), .B2(n6281), .ZN(n6280) );
  OAI21_X1 U6973 ( .B1(n6310), .B2(n6283), .A(n6280), .ZN(U2835) );
  AOI22_X1 U6974 ( .A1(n6479), .A2(n4738), .B1(n6281), .B2(EBX_REG_23__SCAN_IN), .ZN(n6282) );
  OAI21_X1 U6975 ( .B1(n6313), .B2(n6283), .A(n6282), .ZN(U2836) );
  INV_X1 U6976 ( .A(n6484), .ZN(n6286) );
  OAI222_X1 U6977 ( .A1(n6286), .A2(n6629), .B1(n6285), .B2(n6636), .C1(n6284), 
        .C2(n6283), .ZN(U2837) );
  NAND3_X1 U6978 ( .A1(n3441), .A2(n6288), .A3(n6287), .ZN(n6290) );
  AOI22_X1 U6979 ( .A1(n7063), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7062), .ZN(n6289) );
  NAND2_X1 U6980 ( .A1(n6290), .A2(n6289), .ZN(U2860) );
  AOI22_X1 U6981 ( .A1(n7059), .A2(DATAI_14_), .B1(n7062), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U6982 ( .A1(n7063), .A2(DATAI_30_), .ZN(n6291) );
  OAI211_X1 U6983 ( .C1(n6293), .C2(n3421), .A(n6292), .B(n6291), .ZN(U2861)
         );
  AOI22_X1 U6984 ( .A1(n7059), .A2(DATAI_13_), .B1(n7062), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U6985 ( .A1(n7063), .A2(DATAI_29_), .ZN(n6294) );
  OAI211_X1 U6986 ( .C1(n6296), .C2(n3421), .A(n6295), .B(n6294), .ZN(U2862)
         );
  AOI22_X1 U6987 ( .A1(n7059), .A2(DATAI_12_), .B1(n7062), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U6988 ( .A1(n7063), .A2(DATAI_28_), .ZN(n6297) );
  OAI211_X1 U6989 ( .C1(n6299), .C2(n3421), .A(n6298), .B(n6297), .ZN(U2863)
         );
  AOI22_X1 U6990 ( .A1(n7059), .A2(DATAI_11_), .B1(n7062), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U6991 ( .A1(n7063), .A2(DATAI_27_), .ZN(n6300) );
  OAI211_X1 U6992 ( .C1(n6302), .C2(n3421), .A(n6301), .B(n6300), .ZN(U2864)
         );
  AOI22_X1 U6993 ( .A1(n7059), .A2(DATAI_10_), .B1(n7062), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U6994 ( .A1(n7063), .A2(DATAI_26_), .ZN(n6303) );
  OAI211_X1 U6995 ( .C1(n6305), .C2(n3421), .A(n6304), .B(n6303), .ZN(U2865)
         );
  AOI22_X1 U6996 ( .A1(n7059), .A2(DATAI_9_), .B1(n7062), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U6997 ( .A1(n7063), .A2(DATAI_25_), .ZN(n6306) );
  OAI211_X1 U6998 ( .C1(n6351), .C2(n3421), .A(n6307), .B(n6306), .ZN(U2866)
         );
  AOI22_X1 U6999 ( .A1(n7059), .A2(DATAI_8_), .B1(n7062), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7000 ( .A1(n7063), .A2(DATAI_24_), .ZN(n6308) );
  OAI211_X1 U7001 ( .C1(n6310), .C2(n3421), .A(n6309), .B(n6308), .ZN(U2867)
         );
  AOI22_X1 U7002 ( .A1(n7059), .A2(DATAI_7_), .B1(n7062), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7003 ( .A1(n7063), .A2(DATAI_23_), .ZN(n6311) );
  OAI211_X1 U7004 ( .C1(n6313), .C2(n3421), .A(n6312), .B(n6311), .ZN(U2868)
         );
  NAND2_X1 U7005 ( .A1(n6669), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6314)
         );
  OAI211_X1 U7006 ( .C1(n6676), .C2(n6316), .A(n6315), .B(n6314), .ZN(n6317)
         );
  OAI21_X1 U7007 ( .B1(n6319), .B2(n6952), .A(n6318), .ZN(U2955) );
  NAND2_X1 U7008 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  XNOR2_X1 U7009 ( .A(n6323), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6436)
         );
  NAND2_X1 U7010 ( .A1(n6665), .A2(n6324), .ZN(n6325) );
  NAND2_X1 U7011 ( .A1(n6809), .A2(REIP_REG_30__SCAN_IN), .ZN(n6430) );
  OAI211_X1 U7012 ( .C1(n6326), .C2(n6422), .A(n6325), .B(n6430), .ZN(n6327)
         );
  AOI21_X1 U7013 ( .B1(n6328), .B2(n6670), .A(n6327), .ZN(n6329) );
  OAI21_X1 U7014 ( .B1(n6436), .B2(n6952), .A(n6329), .ZN(U2956) );
  NOR2_X1 U7015 ( .A1(n6418), .A2(n6451), .ZN(n6338) );
  NOR2_X1 U7016 ( .A1(n6330), .A2(n6338), .ZN(n6332) );
  XNOR2_X1 U7017 ( .A(n6418), .B(n6440), .ZN(n6331) );
  XNOR2_X1 U7018 ( .A(n6332), .B(n6331), .ZN(n6445) );
  AND2_X1 U7019 ( .A1(n6809), .A2(REIP_REG_27__SCAN_IN), .ZN(n6437) );
  AOI21_X1 U7020 ( .B1(n6669), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6437), 
        .ZN(n6333) );
  OAI21_X1 U7021 ( .B1(n6676), .B2(n6334), .A(n6333), .ZN(n6335) );
  AOI21_X1 U7022 ( .B1(n6336), .B2(n6670), .A(n6335), .ZN(n6337) );
  OAI21_X1 U7023 ( .B1(n6445), .B2(n6952), .A(n6337), .ZN(U2959) );
  NOR2_X1 U7024 ( .A1(n6339), .A2(n6338), .ZN(n6341) );
  XOR2_X1 U7025 ( .A(n6341), .B(n6340), .Z(n6457) );
  AND2_X1 U7026 ( .A1(n6809), .A2(REIP_REG_26__SCAN_IN), .ZN(n6453) );
  AOI21_X1 U7027 ( .B1(n6669), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6453), 
        .ZN(n6342) );
  OAI21_X1 U7028 ( .B1(n6676), .B2(n6343), .A(n6342), .ZN(n6344) );
  AOI21_X1 U7029 ( .B1(n6345), .B2(n6670), .A(n6344), .ZN(n6346) );
  OAI21_X1 U7030 ( .B1(n6952), .B2(n6457), .A(n6346), .ZN(U2960) );
  NAND2_X1 U7031 ( .A1(n6348), .A2(n6347), .ZN(n6349) );
  XOR2_X1 U7032 ( .A(n6350), .B(n6349), .Z(n6465) );
  INV_X1 U7033 ( .A(n6351), .ZN(n6355) );
  AND2_X1 U7034 ( .A1(n6809), .A2(REIP_REG_25__SCAN_IN), .ZN(n6461) );
  AOI21_X1 U7035 ( .B1(n6669), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n6461), 
        .ZN(n6352) );
  OAI21_X1 U7036 ( .B1(n6676), .B2(n6353), .A(n6352), .ZN(n6354) );
  AOI21_X1 U7037 ( .B1(n6355), .B2(n6670), .A(n6354), .ZN(n6356) );
  OAI21_X1 U7038 ( .B1(n6952), .B2(n6465), .A(n6356), .ZN(U2961) );
  OR3_X2 U7039 ( .A1(n6407), .A2(n6358), .A3(n6357), .ZN(n6361) );
  OAI21_X1 U7040 ( .B1(n6495), .B2(n6487), .A(n6418), .ZN(n6359) );
  NAND2_X1 U7041 ( .A1(n6361), .A2(n6359), .ZN(n6382) );
  NAND3_X1 U7042 ( .A1(n6418), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U7043 ( .A1(n4116), .A2(n6381), .ZN(n6380) );
  NOR2_X2 U7044 ( .A1(n6361), .A2(n6380), .ZN(n6371) );
  NAND2_X1 U7045 ( .A1(n6371), .A2(n6362), .ZN(n6363) );
  XNOR2_X1 U7046 ( .A(n6365), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6473)
         );
  AND2_X1 U7047 ( .A1(n6809), .A2(REIP_REG_24__SCAN_IN), .ZN(n6470) );
  AOI21_X1 U7048 ( .B1(n6669), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6470), 
        .ZN(n6366) );
  OAI21_X1 U7049 ( .B1(n6676), .B2(n6367), .A(n6366), .ZN(n6368) );
  AOI21_X1 U7050 ( .B1(n6369), .B2(n6670), .A(n6368), .ZN(n6370) );
  OAI21_X1 U7051 ( .B1(n6473), .B2(n6952), .A(n6370), .ZN(U2962) );
  INV_X1 U7052 ( .A(n6371), .ZN(n6373) );
  NAND3_X1 U7053 ( .A1(n6410), .A2(n6474), .A3(n6418), .ZN(n6372) );
  NAND2_X1 U7054 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  XNOR2_X1 U7055 ( .A(n6374), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6482)
         );
  AND2_X1 U7056 ( .A1(n6809), .A2(REIP_REG_23__SCAN_IN), .ZN(n6478) );
  AOI21_X1 U7057 ( .B1(n6669), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6478), 
        .ZN(n6375) );
  OAI21_X1 U7058 ( .B1(n6676), .B2(n6376), .A(n6375), .ZN(n6377) );
  AOI21_X1 U7059 ( .B1(n6378), .B2(n6670), .A(n6377), .ZN(n6379) );
  OAI21_X1 U7060 ( .B1(n6482), .B2(n6952), .A(n6379), .ZN(U2963) );
  OAI21_X1 U7061 ( .B1(n4116), .B2(n6381), .A(n6380), .ZN(n6383) );
  XOR2_X1 U7062 ( .A(n6383), .B(n6382), .Z(n6491) );
  NOR2_X1 U7063 ( .A1(n6818), .A2(n6581), .ZN(n6483) );
  NOR2_X1 U7064 ( .A1(n6422), .A2(n6384), .ZN(n6385) );
  AOI211_X1 U7065 ( .C1(n6665), .C2(n6386), .A(n6483), .B(n6385), .ZN(n6389)
         );
  NAND2_X1 U7066 ( .A1(n6387), .A2(n6670), .ZN(n6388) );
  OAI211_X1 U7067 ( .C1(n6491), .C2(n6952), .A(n6389), .B(n6388), .ZN(U2964)
         );
  INV_X1 U7068 ( .A(n6390), .ZN(n7061) );
  NAND2_X1 U7069 ( .A1(n6669), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6391)
         );
  OAI211_X1 U7070 ( .C1(n6676), .C2(n6951), .A(n6392), .B(n6391), .ZN(n6393)
         );
  AOI21_X1 U7071 ( .B1(n7061), .B2(n6670), .A(n6393), .ZN(n6394) );
  OAI21_X1 U7072 ( .B1(n6395), .B2(n6952), .A(n6394), .ZN(U2965) );
  NAND2_X1 U7073 ( .A1(n6407), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6396) );
  MUX2_X1 U7074 ( .A(n6407), .B(n6396), .S(n6418), .Z(n6398) );
  XNOR2_X1 U7075 ( .A(n6398), .B(n6397), .ZN(n6499) );
  INV_X1 U7076 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6399) );
  NOR2_X1 U7077 ( .A1(n6818), .A2(n6399), .ZN(n6494) );
  NOR2_X1 U7078 ( .A1(n6422), .A2(n6400), .ZN(n6401) );
  AOI211_X1 U7079 ( .C1(n6665), .C2(n6402), .A(n6494), .B(n6401), .ZN(n6406)
         );
  INV_X1 U7080 ( .A(n6403), .ZN(n6404) );
  NAND2_X1 U7081 ( .A1(n6404), .A2(n6670), .ZN(n6405) );
  OAI211_X1 U7082 ( .C1(n6499), .C2(n6952), .A(n6406), .B(n6405), .ZN(U2966)
         );
  INV_X1 U7083 ( .A(n6407), .ZN(n6408) );
  AOI21_X1 U7084 ( .B1(n6410), .B2(n6409), .A(n6408), .ZN(n6508) );
  INV_X1 U7085 ( .A(n6411), .ZN(n7056) );
  NAND2_X1 U7086 ( .A1(n6809), .A2(REIP_REG_19__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U7087 ( .A1(n6669), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6412)
         );
  OAI211_X1 U7088 ( .C1(n6676), .C2(n6413), .A(n6502), .B(n6412), .ZN(n6414)
         );
  AOI21_X1 U7089 ( .B1(n7056), .B2(n6670), .A(n6414), .ZN(n6415) );
  OAI21_X1 U7090 ( .B1(n6508), .B2(n6952), .A(n6415), .ZN(U2967) );
  NOR2_X1 U7091 ( .A1(n6417), .A2(n3777), .ZN(n6420) );
  OAI21_X1 U7092 ( .B1(n6814), .B2(n6418), .A(n6417), .ZN(n6509) );
  NOR2_X1 U7093 ( .A1(n6509), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6419)
         );
  MUX2_X1 U7094 ( .A(n6420), .B(n6419), .S(n4116), .Z(n6421) );
  XOR2_X1 U7095 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n6421), .Z(n6822) );
  NAND2_X1 U7096 ( .A1(n6822), .A2(n6671), .ZN(n6425) );
  OAI22_X1 U7097 ( .A1(n6422), .A2(n6926), .B1(n6818), .B2(n6937), .ZN(n6423)
         );
  AOI21_X1 U7098 ( .B1(n6665), .B2(n6922), .A(n6423), .ZN(n6424) );
  OAI211_X1 U7099 ( .C1(n6426), .C2(n6921), .A(n6425), .B(n6424), .ZN(U2968)
         );
  INV_X1 U7100 ( .A(n6428), .ZN(n6433) );
  NAND3_X1 U7101 ( .A1(n6438), .A2(n6429), .A3(n6432), .ZN(n6431) );
  OAI211_X1 U7102 ( .C1(n6433), .C2(n6432), .A(n6431), .B(n6430), .ZN(n6434)
         );
  AOI21_X1 U7103 ( .B1(n4739), .B2(n6826), .A(n6434), .ZN(n6435) );
  OAI21_X1 U7104 ( .B1(n6436), .B2(n6800), .A(n6435), .ZN(U2988) );
  AOI21_X1 U7105 ( .B1(n6438), .B2(n6440), .A(n6437), .ZN(n6439) );
  OAI21_X1 U7106 ( .B1(n6441), .B2(n6440), .A(n6439), .ZN(n6442) );
  AOI21_X1 U7107 ( .B1(n6826), .B2(n6443), .A(n6442), .ZN(n6444) );
  OAI21_X1 U7108 ( .B1(n6445), .B2(n6800), .A(n6444), .ZN(U2991) );
  INV_X1 U7109 ( .A(n6446), .ZN(n6449) );
  INV_X1 U7110 ( .A(n6447), .ZN(n6448) );
  NAND2_X1 U7111 ( .A1(n6506), .A2(n6448), .ZN(n6459) );
  AOI211_X1 U7112 ( .C1(n6451), .C2(n6450), .A(n6449), .B(n6459), .ZN(n6452)
         );
  AOI211_X1 U7113 ( .C1(n6454), .C2(n6826), .A(n6453), .B(n6452), .ZN(n6456)
         );
  NAND2_X1 U7114 ( .A1(n6466), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6455) );
  OAI211_X1 U7115 ( .C1(n6457), .C2(n6800), .A(n6456), .B(n6455), .ZN(U2992)
         );
  INV_X1 U7116 ( .A(n6458), .ZN(n6462) );
  NOR2_X1 U7117 ( .A1(n6459), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6460)
         );
  AOI211_X1 U7118 ( .C1(n6462), .C2(n6826), .A(n6461), .B(n6460), .ZN(n6464)
         );
  NAND2_X1 U7119 ( .A1(n6466), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6463) );
  OAI211_X1 U7120 ( .C1(n6465), .C2(n6800), .A(n6464), .B(n6463), .ZN(U2993)
         );
  NAND3_X1 U7121 ( .A1(n6506), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n6474), .ZN(n6468) );
  INV_X1 U7122 ( .A(n6466), .ZN(n6467) );
  AOI21_X1 U7123 ( .B1(n3798), .B2(n6468), .A(n6467), .ZN(n6469) );
  AOI211_X1 U7124 ( .C1(n6826), .C2(n6471), .A(n6470), .B(n6469), .ZN(n6472)
         );
  OAI21_X1 U7125 ( .B1(n6473), .B2(n6800), .A(n6472), .ZN(U2994) );
  INV_X1 U7126 ( .A(n6506), .ZN(n6476) );
  INV_X1 U7127 ( .A(n6474), .ZN(n6475) );
  NOR3_X1 U7128 ( .A1(n6476), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n6475), 
        .ZN(n6477) );
  AOI211_X1 U7129 ( .C1(n6826), .C2(n6479), .A(n6478), .B(n6477), .ZN(n6481)
         );
  NAND2_X1 U7130 ( .A1(n6489), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6480) );
  OAI211_X1 U7131 ( .C1(n6482), .C2(n6800), .A(n6481), .B(n6480), .ZN(U2995)
         );
  AOI21_X1 U7132 ( .B1(n6484), .B2(n6826), .A(n6483), .ZN(n6485) );
  OAI21_X1 U7133 ( .B1(n6487), .B2(n6486), .A(n6485), .ZN(n6488) );
  AOI21_X1 U7134 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6489), .A(n6488), 
        .ZN(n6490) );
  OAI21_X1 U7135 ( .B1(n6491), .B2(n6800), .A(n6490), .ZN(U2996) );
  NOR2_X1 U7136 ( .A1(n6492), .A2(n6799), .ZN(n6493) );
  AOI211_X1 U7137 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n6500), .A(n6494), .B(n6493), .ZN(n6498) );
  NAND3_X1 U7138 ( .A1(n6506), .A2(n6496), .A3(n6495), .ZN(n6497) );
  OAI211_X1 U7139 ( .C1(n6499), .C2(n6800), .A(n6498), .B(n6497), .ZN(U2998)
         );
  NAND2_X1 U7140 ( .A1(n6500), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6501) );
  OAI211_X1 U7141 ( .C1(n6503), .C2(n6799), .A(n6502), .B(n6501), .ZN(n6504)
         );
  AOI21_X1 U7142 ( .B1(n6506), .B2(n6505), .A(n6504), .ZN(n6507) );
  OAI21_X1 U7143 ( .B1(n6508), .B2(n6800), .A(n6507), .ZN(U2999) );
  NOR2_X1 U7144 ( .A1(n6817), .A2(n6795), .ZN(n6808) );
  NAND2_X1 U7145 ( .A1(n6808), .A2(n6805), .ZN(n6518) );
  MUX2_X1 U7146 ( .A(n3777), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .S(n6418), 
        .Z(n6510) );
  XOR2_X1 U7147 ( .A(n6510), .B(n6509), .Z(n6672) );
  NAND2_X1 U7148 ( .A1(n6672), .A2(n6821), .ZN(n6517) );
  AOI21_X1 U7149 ( .B1(n6748), .B2(n6512), .A(n6511), .ZN(n6823) );
  NAND2_X1 U7150 ( .A1(n6809), .A2(REIP_REG_17__SCAN_IN), .ZN(n6513) );
  OAI21_X1 U7151 ( .B1(n3777), .B2(n6823), .A(n6513), .ZN(n6514) );
  AOI21_X1 U7152 ( .B1(n6515), .B2(n6826), .A(n6514), .ZN(n6516) );
  OAI211_X1 U7153 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n6518), .A(n6517), .B(n6516), .ZN(U3001) );
  INV_X1 U7154 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6614) );
  INV_X1 U7155 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7034) );
  NOR2_X1 U7156 ( .A1(n7034), .A2(STATE_REG_0__SCAN_IN), .ZN(n7051) );
  INV_X1 U7157 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7032) );
  AOI21_X1 U7158 ( .B1(n7032), .B2(STATE_REG_1__SCAN_IN), .A(n3662), .ZN(n6523) );
  NOR2_X1 U7159 ( .A1(n7051), .A2(n6523), .ZN(n7031) );
  INV_X1 U7160 ( .A(n7031), .ZN(n6520) );
  NAND2_X1 U7161 ( .A1(n7032), .A2(n3662), .ZN(n6682) );
  AOI21_X1 U7162 ( .B1(n6519), .B2(n6682), .A(n6520), .ZN(n7027) );
  AOI21_X1 U7163 ( .B1(n6614), .B2(n6520), .A(n7027), .ZN(U3451) );
  AND2_X1 U7164 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6520), .ZN(U3180) );
  AND2_X1 U7165 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6520), .ZN(U3179) );
  AND2_X1 U7166 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6520), .ZN(U3178) );
  AND2_X1 U7167 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6520), .ZN(U3177) );
  AND2_X1 U7168 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6520), .ZN(U3176) );
  AND2_X1 U7169 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6520), .ZN(U3175) );
  AND2_X1 U7170 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6520), .ZN(U3174) );
  AND2_X1 U7171 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6520), .ZN(U3173) );
  AND2_X1 U7172 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6520), .ZN(U3172) );
  AND2_X1 U7173 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6520), .ZN(U3171) );
  AND2_X1 U7174 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6520), .ZN(U3170) );
  AND2_X1 U7175 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6520), .ZN(U3169) );
  AND2_X1 U7176 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6520), .ZN(U3168) );
  AND2_X1 U7177 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6520), .ZN(U3167) );
  AND2_X1 U7178 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6520), .ZN(U3166) );
  AND2_X1 U7179 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6520), .ZN(U3165) );
  AND2_X1 U7180 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6520), .ZN(U3164) );
  AND2_X1 U7181 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6520), .ZN(U3163) );
  AND2_X1 U7182 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6520), .ZN(U3162) );
  AND2_X1 U7183 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6520), .ZN(U3161) );
  AND2_X1 U7184 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6520), .ZN(U3160) );
  AND2_X1 U7185 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6520), .ZN(U3159) );
  AND2_X1 U7186 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6520), .ZN(U3158) );
  AND2_X1 U7187 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6520), .ZN(U3157) );
  AND2_X1 U7188 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6520), .ZN(U3156) );
  AND2_X1 U7189 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6520), .ZN(U3155) );
  AND2_X1 U7190 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6520), .ZN(U3154) );
  AND2_X1 U7191 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6520), .ZN(U3153) );
  AND2_X1 U7192 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6520), .ZN(U3152) );
  AND2_X1 U7193 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6520), .ZN(U3151) );
  AND2_X1 U7194 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6521), .ZN(U3019)
         );
  AND2_X1 U7195 ( .A1(n6534), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7196 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6522) );
  AOI21_X1 U7197 ( .B1(n6523), .B2(n6522), .A(n7051), .ZN(U2789) );
  AOI22_X1 U7198 ( .A1(n6696), .A2(LWORD_REG_0__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6525) );
  OAI21_X1 U7199 ( .B1(n6526), .B2(n6551), .A(n6525), .ZN(U2923) );
  AOI22_X1 U7200 ( .A1(n6696), .A2(LWORD_REG_1__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6527) );
  OAI21_X1 U7201 ( .B1(n4196), .B2(n6551), .A(n6527), .ZN(U2922) );
  AOI22_X1 U7202 ( .A1(n6696), .A2(LWORD_REG_2__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6528) );
  OAI21_X1 U7203 ( .B1(n6529), .B2(n6551), .A(n6528), .ZN(U2921) );
  AOI22_X1 U7204 ( .A1(n6696), .A2(LWORD_REG_3__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6530) );
  OAI21_X1 U7205 ( .B1(n4217), .B2(n6551), .A(n6530), .ZN(U2920) );
  AOI22_X1 U7206 ( .A1(n6696), .A2(LWORD_REG_4__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6531) );
  OAI21_X1 U7207 ( .B1(n6532), .B2(n6551), .A(n6531), .ZN(U2919) );
  AOI22_X1 U7208 ( .A1(n6696), .A2(LWORD_REG_5__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6533) );
  OAI21_X1 U7209 ( .B1(n4231), .B2(n6551), .A(n6533), .ZN(U2918) );
  AOI22_X1 U7210 ( .A1(n6696), .A2(LWORD_REG_6__SCAN_IN), .B1(n6534), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6535) );
  OAI21_X1 U7211 ( .B1(n4238), .B2(n6551), .A(n6535), .ZN(U2917) );
  AOI22_X1 U7212 ( .A1(n6696), .A2(LWORD_REG_7__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6536) );
  OAI21_X1 U7213 ( .B1(n4246), .B2(n6551), .A(n6536), .ZN(U2916) );
  AOI22_X1 U7214 ( .A1(n6696), .A2(LWORD_REG_8__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6537) );
  OAI21_X1 U7215 ( .B1(n6538), .B2(n6551), .A(n6537), .ZN(U2915) );
  AOI22_X1 U7216 ( .A1(n6696), .A2(LWORD_REG_9__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6539) );
  OAI21_X1 U7217 ( .B1(n6540), .B2(n6551), .A(n6539), .ZN(U2914) );
  AOI22_X1 U7218 ( .A1(n6696), .A2(LWORD_REG_10__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6541) );
  OAI21_X1 U7219 ( .B1(n6542), .B2(n6551), .A(n6541), .ZN(U2913) );
  AOI22_X1 U7220 ( .A1(n6696), .A2(LWORD_REG_11__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6543) );
  OAI21_X1 U7221 ( .B1(n6544), .B2(n6551), .A(n6543), .ZN(U2912) );
  AOI22_X1 U7222 ( .A1(n6696), .A2(LWORD_REG_12__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6545) );
  OAI21_X1 U7223 ( .B1(n4310), .B2(n6551), .A(n6545), .ZN(U2911) );
  AOI22_X1 U7224 ( .A1(n6696), .A2(LWORD_REG_13__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6546) );
  OAI21_X1 U7225 ( .B1(n6547), .B2(n6551), .A(n6546), .ZN(U2910) );
  AOI22_X1 U7226 ( .A1(n6696), .A2(LWORD_REG_14__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6548) );
  OAI21_X1 U7227 ( .B1(n4340), .B2(n6551), .A(n6548), .ZN(U2909) );
  AOI22_X1 U7228 ( .A1(n6696), .A2(LWORD_REG_15__SCAN_IN), .B1(n6549), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6550) );
  OAI21_X1 U7229 ( .B1(n4764), .B2(n6551), .A(n6550), .ZN(U2908) );
  INV_X2 U7230 ( .A(n7051), .ZN(n7048) );
  NOR2_X1 U7231 ( .A1(n7032), .A2(n7048), .ZN(n6589) );
  INV_X1 U7232 ( .A(n6589), .ZN(n6598) );
  NAND2_X1 U7233 ( .A1(n7032), .A2(n7051), .ZN(n6591) );
  INV_X1 U7234 ( .A(n6591), .ZN(n6596) );
  AOI22_X1 U7235 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n7048), .ZN(n6552) );
  OAI21_X1 U7236 ( .B1(n5582), .B2(n6598), .A(n6552), .ZN(U3184) );
  INV_X1 U7237 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6554) );
  AOI22_X1 U7238 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n7048), .ZN(n6553) );
  OAI21_X1 U7239 ( .B1(n6554), .B2(n6598), .A(n6553), .ZN(U3185) );
  INV_X1 U7240 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U7241 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n7048), .ZN(n6555) );
  OAI21_X1 U7242 ( .B1(n6838), .B2(n6598), .A(n6555), .ZN(U3186) );
  INV_X1 U7243 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6840) );
  AOI22_X1 U7244 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n7048), .ZN(n6556) );
  OAI21_X1 U7245 ( .B1(n6840), .B2(n6598), .A(n6556), .ZN(U3187) );
  AOI22_X1 U7246 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n7048), .ZN(n6557) );
  OAI21_X1 U7247 ( .B1(n6851), .B2(n6598), .A(n6557), .ZN(U3188) );
  INV_X1 U7248 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6870) );
  AOI22_X1 U7249 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n7048), .ZN(n6558) );
  OAI21_X1 U7250 ( .B1(n6870), .B2(n6598), .A(n6558), .ZN(U3189) );
  AOI22_X1 U7251 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n7048), .ZN(n6559) );
  OAI21_X1 U7252 ( .B1(n6561), .B2(n6591), .A(n6559), .ZN(U3190) );
  AOI22_X1 U7253 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n7048), .ZN(n6560) );
  OAI21_X1 U7254 ( .B1(n6561), .B2(n6598), .A(n6560), .ZN(U3191) );
  AOI22_X1 U7255 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n7048), .ZN(n6562) );
  OAI21_X1 U7256 ( .B1(n6564), .B2(n6591), .A(n6562), .ZN(U3192) );
  AOI22_X1 U7257 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n7048), .ZN(n6563) );
  OAI21_X1 U7258 ( .B1(n6564), .B2(n6598), .A(n6563), .ZN(U3193) );
  INV_X1 U7259 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6566) );
  AOI22_X1 U7260 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n7048), .ZN(n6565) );
  OAI21_X1 U7261 ( .B1(n6566), .B2(n6591), .A(n6565), .ZN(U3194) );
  AOI22_X1 U7262 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n7048), .ZN(n6567) );
  OAI21_X1 U7263 ( .B1(n5732), .B2(n6591), .A(n6567), .ZN(U3195) );
  AOI22_X1 U7264 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n7048), .ZN(n6568) );
  OAI21_X1 U7265 ( .B1(n5732), .B2(n6598), .A(n6568), .ZN(U3196) );
  AOI22_X1 U7266 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n7048), .ZN(n6569) );
  OAI21_X1 U7267 ( .B1(n6797), .B2(n6591), .A(n6569), .ZN(U3197) );
  AOI22_X1 U7268 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n7048), .ZN(n6570) );
  OAI21_X1 U7269 ( .B1(n6797), .B2(n6598), .A(n6570), .ZN(U3198) );
  INV_X1 U7270 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6573) );
  AOI22_X1 U7271 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n7048), .ZN(n6571) );
  OAI21_X1 U7272 ( .B1(n6573), .B2(n6591), .A(n6571), .ZN(U3199) );
  AOI22_X1 U7273 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n7048), .ZN(n6572) );
  OAI21_X1 U7274 ( .B1(n6573), .B2(n6598), .A(n6572), .ZN(U3200) );
  AOI22_X1 U7275 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n7048), .ZN(n6574) );
  OAI21_X1 U7276 ( .B1(n6576), .B2(n6591), .A(n6574), .ZN(U3201) );
  AOI22_X1 U7277 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n7048), .ZN(n6575) );
  OAI21_X1 U7278 ( .B1(n6576), .B2(n6598), .A(n6575), .ZN(U3202) );
  AOI22_X1 U7279 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n7048), .ZN(n6577) );
  OAI21_X1 U7280 ( .B1(n6579), .B2(n6591), .A(n6577), .ZN(U3203) );
  AOI22_X1 U7281 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n7048), .ZN(n6578) );
  OAI21_X1 U7282 ( .B1(n6579), .B2(n6598), .A(n6578), .ZN(U3204) );
  AOI22_X1 U7283 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n7048), .ZN(n6580) );
  OAI21_X1 U7284 ( .B1(n6581), .B2(n6598), .A(n6580), .ZN(U3205) );
  AOI22_X1 U7285 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n7048), .ZN(n6582) );
  OAI21_X1 U7286 ( .B1(n6583), .B2(n6591), .A(n6582), .ZN(U3206) );
  AOI22_X1 U7287 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n7048), .ZN(n6584) );
  OAI21_X1 U7288 ( .B1(n6586), .B2(n6591), .A(n6584), .ZN(U3207) );
  AOI22_X1 U7289 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n7048), .ZN(n6585) );
  OAI21_X1 U7290 ( .B1(n6586), .B2(n6598), .A(n6585), .ZN(U3208) );
  AOI22_X1 U7291 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n7048), .ZN(n6587) );
  OAI21_X1 U7292 ( .B1(n6588), .B2(n6598), .A(n6587), .ZN(U3209) );
  AOI22_X1 U7293 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6589), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n7048), .ZN(n6590) );
  OAI21_X1 U7294 ( .B1(n6593), .B2(n6591), .A(n6590), .ZN(U3210) );
  AOI22_X1 U7295 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n7048), .ZN(n6592) );
  OAI21_X1 U7296 ( .B1(n6593), .B2(n6598), .A(n6592), .ZN(U3211) );
  AOI22_X1 U7297 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n7048), .ZN(n6594) );
  OAI21_X1 U7298 ( .B1(n6595), .B2(n6598), .A(n6594), .ZN(U3212) );
  AOI22_X1 U7299 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6596), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n7048), .ZN(n6597) );
  OAI21_X1 U7300 ( .B1(n6599), .B2(n6598), .A(n6597), .ZN(U3213) );
  MUX2_X1 U7301 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n7048), .Z(U3445) );
  NOR4_X1 U7302 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6609) );
  NOR4_X1 U7303 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6608) );
  INV_X1 U7304 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7030) );
  NOR4_X1 U7305 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6600) );
  OAI21_X1 U7306 ( .B1(n6614), .B2(n7030), .A(n6600), .ZN(n6606) );
  NOR4_X1 U7307 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6604) );
  NOR4_X1 U7308 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6603) );
  NOR4_X1 U7309 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6602) );
  NOR4_X1 U7310 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6601) );
  NAND4_X1 U7311 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n6605)
         );
  NOR4_X1 U7312 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(
        DATAWIDTH_REG_30__SCAN_IN), .A3(n6606), .A4(n6605), .ZN(n6607) );
  NAND3_X1 U7313 ( .A1(n6609), .A2(n6608), .A3(n6607), .ZN(n6616) );
  INV_X1 U7314 ( .A(n6616), .ZN(n6621) );
  INV_X1 U7315 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6610) );
  NOR2_X1 U7316 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6616), .ZN(n6619) );
  NAND2_X1 U7317 ( .A1(n6619), .A2(n7030), .ZN(n6615) );
  INV_X1 U7318 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6611) );
  NAND4_X1 U7319 ( .A1(n6621), .A2(n6611), .A3(n6614), .A4(n7030), .ZN(n6618)
         );
  OAI211_X1 U7320 ( .C1(n6621), .C2(n6610), .A(n6615), .B(n6618), .ZN(U2795)
         );
  MUX2_X1 U7321 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n7048), .Z(U3446) );
  NAND2_X1 U7322 ( .A1(n6619), .A2(n6611), .ZN(n6620) );
  NOR2_X1 U7323 ( .A1(n6616), .A2(n5582), .ZN(n6612) );
  AOI22_X1 U7324 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(n6616), .B1(
        REIP_REG_0__SCAN_IN), .B2(n6612), .ZN(n6613) );
  OAI221_X1 U7325 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6615), .C1(n6614), 
        .C2(n6620), .A(n6613), .ZN(U3468) );
  MUX2_X1 U7326 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n7048), .Z(U3447) );
  AOI22_X1 U7327 ( .A1(n6619), .A2(n6618), .B1(n6617), .B2(n6616), .ZN(U2794)
         );
  MUX2_X1 U7328 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n7048), .Z(U3448) );
  OAI21_X1 U7329 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(n6621), .A(n6620), .ZN(
        n6622) );
  INV_X1 U7330 ( .A(n6622), .ZN(U3469) );
  INV_X1 U7331 ( .A(n6623), .ZN(n6649) );
  AOI22_X1 U7332 ( .A1(n6649), .A2(n6634), .B1(n4738), .B2(n6728), .ZN(n6624)
         );
  OAI21_X1 U7333 ( .B1(n6636), .B2(n6625), .A(n6624), .ZN(U2856) );
  INV_X1 U7334 ( .A(n6626), .ZN(n6627) );
  XNOR2_X1 U7335 ( .A(n6628), .B(n6627), .ZN(n6874) );
  NOR2_X1 U7336 ( .A1(n6629), .A2(n6874), .ZN(n6630) );
  AOI21_X1 U7337 ( .B1(n6877), .B2(n6634), .A(n6630), .ZN(n6631) );
  OAI21_X1 U7338 ( .B1(n6636), .B2(n6632), .A(n6631), .ZN(U2852) );
  AOI22_X1 U7339 ( .A1(n6902), .A2(n6634), .B1(n4738), .B2(n6896), .ZN(n6633)
         );
  OAI21_X1 U7340 ( .B1(n6636), .B2(n6898), .A(n6633), .ZN(U2847) );
  AOI22_X1 U7341 ( .A1(n6913), .A2(n6634), .B1(n4738), .B2(n6914), .ZN(n6635)
         );
  OAI21_X1 U7342 ( .B1(n6636), .B2(n6908), .A(n6635), .ZN(U2846) );
  AOI22_X1 U7343 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6669), .B1(n6809), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U7344 ( .A1(n6637), .A2(n6638), .ZN(n6639) );
  XOR2_X1 U7345 ( .A(n6640), .B(n6639), .Z(n6750) );
  AOI22_X1 U7346 ( .A1(n6750), .A2(n6671), .B1(n6670), .B2(n6641), .ZN(n6642)
         );
  OAI211_X1 U7347 ( .C1(n6676), .C2(n6644), .A(n6643), .B(n6642), .ZN(U2984)
         );
  AOI22_X1 U7348 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6669), .B1(n6809), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U7349 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  XOR2_X1 U7350 ( .A(n6648), .B(n6647), .Z(n6730) );
  AOI22_X1 U7351 ( .A1(n6730), .A2(n6671), .B1(n6670), .B2(n6649), .ZN(n6650)
         );
  OAI211_X1 U7352 ( .C1(n6676), .C2(n6652), .A(n6651), .B(n6650), .ZN(U2983)
         );
  AOI22_X1 U7353 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6669), .B1(n6809), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U7354 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  XNOR2_X1 U7355 ( .A(n6653), .B(n6656), .ZN(n6738) );
  AOI22_X1 U7356 ( .A1(n6738), .A2(n6671), .B1(n6670), .B2(n6867), .ZN(n6657)
         );
  OAI211_X1 U7357 ( .C1(n6676), .C2(n6869), .A(n6658), .B(n6657), .ZN(U2980)
         );
  AOI22_X1 U7358 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6669), .B1(n6809), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6664) );
  OAI21_X1 U7359 ( .B1(n6661), .B2(n6660), .A(n6659), .ZN(n6662) );
  INV_X1 U7360 ( .A(n6662), .ZN(n6770) );
  AOI22_X1 U7361 ( .A1(n6770), .A2(n6671), .B1(n6670), .B2(n6877), .ZN(n6663)
         );
  OAI211_X1 U7362 ( .C1(n6676), .C2(n6882), .A(n6664), .B(n6663), .ZN(U2979)
         );
  AOI22_X1 U7363 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6669), .B1(n6809), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n6667) );
  AOI22_X1 U7364 ( .A1(n6902), .A2(n6670), .B1(n6901), .B2(n6665), .ZN(n6666)
         );
  OAI211_X1 U7365 ( .C1(n6668), .C2(n6952), .A(n6667), .B(n6666), .ZN(U2974)
         );
  AOI22_X1 U7366 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6669), .B1(n6809), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n6674) );
  AOI22_X1 U7367 ( .A1(n6672), .A2(n6671), .B1(n6670), .B2(n7053), .ZN(n6673)
         );
  OAI211_X1 U7368 ( .C1(n6676), .C2(n6675), .A(n6674), .B(n6673), .ZN(U2969)
         );
  AND2_X1 U7369 ( .A1(n6677), .A2(n7004), .ZN(n6680) );
  OAI22_X1 U7370 ( .A1(n6680), .A2(n6679), .B1(n7020), .B2(n6678), .ZN(U2790)
         );
  NOR2_X1 U7371 ( .A1(n7051), .A2(D_C_N_REG_SCAN_IN), .ZN(n6681) );
  AOI22_X1 U7372 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7051), .B1(n6682), .B2(
        n6681), .ZN(U2791) );
  AOI22_X1 U7373 ( .A1(n7051), .A2(READREQUEST_REG_SCAN_IN), .B1(n6683), .B2(
        n7048), .ZN(U3470) );
  NAND2_X1 U7374 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n7038) );
  INV_X1 U7375 ( .A(n7038), .ZN(n6686) );
  NOR2_X1 U7376 ( .A1(n3662), .A2(n7035), .ZN(n7041) );
  AOI21_X1 U7377 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n7041), .ZN(n6685)
         );
  NAND2_X1 U7378 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n7046) );
  OAI211_X1 U7379 ( .C1(n6686), .C2(n6685), .A(n6684), .B(n7046), .ZN(U3182)
         );
  NOR2_X1 U7380 ( .A1(READY_N), .A2(n7020), .ZN(n6687) );
  OAI211_X1 U7381 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6687), .A(n7013), .B(
        n7015), .ZN(n6688) );
  NAND2_X1 U7382 ( .A1(n6689), .A2(n6688), .ZN(U3150) );
  AOI211_X1 U7383 ( .C1(n6692), .C2(n7028), .A(n6691), .B(n6690), .ZN(n6693)
         );
  OAI21_X1 U7384 ( .B1(n6693), .B2(n7020), .A(n7015), .ZN(n6698) );
  AOI211_X1 U7385 ( .C1(n6696), .C2(n7042), .A(n6695), .B(n6694), .ZN(n6697)
         );
  MUX2_X1 U7386 ( .A(n6698), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6697), .Z(
        U3472) );
  NAND2_X1 U7387 ( .A1(n6700), .A2(n6699), .ZN(n6713) );
  INV_X1 U7388 ( .A(n6701), .ZN(n6707) );
  INV_X1 U7389 ( .A(n6702), .ZN(n6704) );
  OAI21_X1 U7390 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6706) );
  NAND2_X1 U7391 ( .A1(n6707), .A2(n6706), .ZN(n6708) );
  AOI222_X1 U7392 ( .A1(n6710), .A2(n6821), .B1(n6826), .B2(n6709), .C1(n6708), 
        .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U7393 ( .A1(n6809), .A2(REIP_REG_14__SCAN_IN), .ZN(n6711) );
  OAI211_X1 U7394 ( .C1(n6817), .C2(n6713), .A(n6712), .B(n6711), .ZN(U3004)
         );
  AOI21_X1 U7395 ( .B1(n6745), .B2(n6715), .A(n6714), .ZN(n6727) );
  INV_X1 U7396 ( .A(n6716), .ZN(n6717) );
  AOI21_X1 U7397 ( .B1(n6826), .B2(n6718), .A(n6717), .ZN(n6725) );
  INV_X1 U7398 ( .A(n6719), .ZN(n6720) );
  NOR3_X1 U7399 ( .A1(n6721), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6720), 
        .ZN(n6722) );
  AOI21_X1 U7400 ( .B1(n6821), .B2(n6723), .A(n6722), .ZN(n6724) );
  OAI211_X1 U7401 ( .C1(n6727), .C2(n6726), .A(n6725), .B(n6724), .ZN(U3017)
         );
  AOI22_X1 U7402 ( .A1(n6826), .A2(n6728), .B1(n6809), .B2(REIP_REG_3__SCAN_IN), .ZN(n6732) );
  AOI22_X1 U7403 ( .A1(n6730), .A2(n6821), .B1(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n6729), .ZN(n6731) );
  OAI211_X1 U7404 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6735), .A(n6732), 
        .B(n6731), .ZN(U3015) );
  INV_X1 U7405 ( .A(n6860), .ZN(n6733) );
  AOI22_X1 U7406 ( .A1(n6826), .A2(n6733), .B1(n6809), .B2(REIP_REG_6__SCAN_IN), .ZN(n6740) );
  INV_X1 U7407 ( .A(n6734), .ZN(n6736) );
  NOR3_X1 U7408 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6736), .A3(n6735), 
        .ZN(n6737) );
  AOI21_X1 U7409 ( .B1(n6738), .B2(n6821), .A(n6737), .ZN(n6739) );
  OAI211_X1 U7410 ( .C1(n6742), .C2(n6741), .A(n6740), .B(n6739), .ZN(U3012)
         );
  OAI21_X1 U7411 ( .B1(n6745), .B2(n6744), .A(n6743), .ZN(n6747) );
  AOI22_X1 U7412 ( .A1(n6748), .A2(n6747), .B1(n6826), .B2(n6746), .ZN(n6756)
         );
  AOI22_X1 U7413 ( .A1(n6750), .A2(n6821), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6749), .ZN(n6755) );
  NAND2_X1 U7414 ( .A1(n6809), .A2(REIP_REG_2__SCAN_IN), .ZN(n6754) );
  NAND3_X1 U7415 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6752), .A3(n6751), 
        .ZN(n6753) );
  NAND4_X1 U7416 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(U3016)
         );
  NAND2_X1 U7417 ( .A1(n6758), .A2(n6757), .ZN(n6776) );
  OAI21_X1 U7418 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6777), .ZN(n6768) );
  INV_X1 U7419 ( .A(n6759), .ZN(n6760) );
  AOI21_X1 U7420 ( .B1(n6826), .B2(n6761), .A(n6760), .ZN(n6767) );
  INV_X1 U7421 ( .A(n6762), .ZN(n6765) );
  NAND2_X1 U7422 ( .A1(n6764), .A2(n6763), .ZN(n6773) );
  AOI22_X1 U7423 ( .A1(n6765), .A2(n6821), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6773), .ZN(n6766) );
  OAI211_X1 U7424 ( .C1(n6776), .C2(n6768), .A(n6767), .B(n6766), .ZN(U3010)
         );
  INV_X1 U7425 ( .A(n6874), .ZN(n6769) );
  AOI22_X1 U7426 ( .A1(n6826), .A2(n6769), .B1(n6809), .B2(REIP_REG_7__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U7427 ( .A1(n6770), .A2(n6821), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6773), .ZN(n6771) );
  OAI211_X1 U7428 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6776), .A(n6772), 
        .B(n6771), .ZN(U3011) );
  AOI21_X1 U7429 ( .B1(n6796), .B2(n6777), .A(n6773), .ZN(n6789) );
  INV_X1 U7430 ( .A(n6774), .ZN(n6775) );
  AOI21_X1 U7431 ( .B1(n6826), .B2(n6886), .A(n6775), .ZN(n6781) );
  NOR2_X1 U7432 ( .A1(n6777), .A2(n6776), .ZN(n6784) );
  AOI22_X1 U7433 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n6788), .B2(n5661), .ZN(n6778) );
  AOI22_X1 U7434 ( .A1(n6779), .A2(n6821), .B1(n6784), .B2(n6778), .ZN(n6780)
         );
  OAI211_X1 U7435 ( .C1(n6789), .C2(n5661), .A(n6781), .B(n6780), .ZN(U3008)
         );
  AOI21_X1 U7436 ( .B1(n6826), .B2(n6783), .A(n6782), .ZN(n6787) );
  AOI22_X1 U7437 ( .A1(n6785), .A2(n6821), .B1(n6784), .B2(n6788), .ZN(n6786)
         );
  OAI211_X1 U7438 ( .C1(n6789), .C2(n6788), .A(n6787), .B(n6786), .ZN(U3009)
         );
  AOI21_X1 U7439 ( .B1(n6826), .B2(n3444), .A(n6790), .ZN(n6793) );
  AOI22_X1 U7440 ( .A1(n6791), .A2(n6821), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6794), .ZN(n6792) );
  OAI211_X1 U7441 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6817), .A(n6793), .B(n6792), .ZN(U3007) );
  AOI21_X1 U7442 ( .B1(n6796), .B2(n6795), .A(n6794), .ZN(n6815) );
  NOR2_X1 U7443 ( .A1(n6818), .A2(n6797), .ZN(n6803) );
  OAI22_X1 U7444 ( .A1(n6801), .A2(n6800), .B1(n6799), .B2(n6798), .ZN(n6802)
         );
  AOI211_X1 U7445 ( .C1(n6808), .C2(n6806), .A(n6803), .B(n6802), .ZN(n6804)
         );
  OAI21_X1 U7446 ( .B1(n6815), .B2(n6806), .A(n6804), .ZN(U3003) );
  AOI21_X1 U7447 ( .B1(n6814), .B2(n6806), .A(n6805), .ZN(n6807) );
  AOI22_X1 U7448 ( .A1(n6809), .A2(REIP_REG_16__SCAN_IN), .B1(n6808), .B2(
        n6807), .ZN(n6813) );
  AOI22_X1 U7449 ( .A1(n6811), .A2(n6821), .B1(n6826), .B2(n6810), .ZN(n6812)
         );
  OAI211_X1 U7450 ( .C1(n6815), .C2(n6814), .A(n6813), .B(n6812), .ZN(U3002)
         );
  NOR3_X1 U7451 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6817), .A3(n6816), 
        .ZN(n6820) );
  NOR2_X1 U7452 ( .A1(n6818), .A2(n6937), .ZN(n6819) );
  AOI211_X1 U7453 ( .C1(n6822), .C2(n6821), .A(n6820), .B(n6819), .ZN(n6829)
         );
  INV_X1 U7454 ( .A(n6930), .ZN(n6827) );
  OAI21_X1 U7455 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6824), .A(n6823), 
        .ZN(n6825) );
  AOI22_X1 U7456 ( .A1(n6827), .A2(n6826), .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6825), .ZN(n6828) );
  NAND2_X1 U7457 ( .A1(n6829), .A2(n6828), .ZN(U3000) );
  AOI22_X1 U7458 ( .A1(n6946), .A2(n6830), .B1(n6943), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n6845) );
  OAI22_X1 U7459 ( .A1(n6832), .A2(n6927), .B1(n6961), .B2(n6831), .ZN(n6833)
         );
  AOI211_X1 U7460 ( .C1(REIP_REG_4__SCAN_IN), .C2(n6834), .A(n6910), .B(n6833), 
        .ZN(n6844) );
  INV_X1 U7461 ( .A(n6835), .ZN(n6854) );
  AOI22_X1 U7462 ( .A1(n6837), .A2(n6854), .B1(n6836), .B2(n6923), .ZN(n6843)
         );
  NOR2_X1 U7463 ( .A1(n6839), .A2(n6838), .ZN(n6841) );
  NAND3_X1 U7464 ( .A1(n6862), .A2(n6841), .A3(n6840), .ZN(n6842) );
  NAND4_X1 U7465 ( .A1(n6845), .A2(n6844), .A3(n6843), .A4(n6842), .ZN(U2823)
         );
  INV_X1 U7466 ( .A(n6846), .ZN(n6847) );
  OAI22_X1 U7467 ( .A1(n6907), .A2(n6848), .B1(n6847), .B2(n6931), .ZN(n6849)
         );
  AOI211_X1 U7468 ( .C1(n6939), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6910), 
        .B(n6849), .ZN(n6857) );
  OAI21_X1 U7469 ( .B1(n6884), .B2(n6861), .A(n6850), .ZN(n6878) );
  OAI21_X1 U7470 ( .B1(n6884), .B2(n6852), .A(n6851), .ZN(n6853) );
  AOI22_X1 U7471 ( .A1(n6855), .A2(n6854), .B1(n6878), .B2(n6853), .ZN(n6856)
         );
  OAI211_X1 U7472 ( .C1(n6858), .C2(n6950), .A(n6857), .B(n6856), .ZN(U2822)
         );
  INV_X1 U7473 ( .A(n6878), .ZN(n6865) );
  AOI21_X1 U7474 ( .B1(n6939), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6910), 
        .ZN(n6859) );
  OAI21_X1 U7475 ( .B1(n6931), .B2(n6860), .A(n6859), .ZN(n6863) );
  NAND2_X1 U7476 ( .A1(n6862), .A2(n6861), .ZN(n6871) );
  NOR2_X1 U7477 ( .A1(n6871), .A2(REIP_REG_6__SCAN_IN), .ZN(n6879) );
  AOI211_X1 U7478 ( .C1(n6943), .C2(EBX_REG_6__SCAN_IN), .A(n6863), .B(n6879), 
        .ZN(n6864) );
  OAI21_X1 U7479 ( .B1(n6865), .B2(n6870), .A(n6864), .ZN(n6866) );
  AOI21_X1 U7480 ( .B1(n6947), .B2(n6867), .A(n6866), .ZN(n6868) );
  OAI21_X1 U7481 ( .B1(n6869), .B2(n6950), .A(n6868), .ZN(U2821) );
  NOR3_X1 U7482 ( .A1(n6871), .A2(n6870), .A3(REIP_REG_7__SCAN_IN), .ZN(n6876)
         );
  NAND2_X1 U7483 ( .A1(n6943), .A2(EBX_REG_7__SCAN_IN), .ZN(n6873) );
  AOI21_X1 U7484 ( .B1(n6939), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6910), 
        .ZN(n6872) );
  OAI211_X1 U7485 ( .C1(n6874), .C2(n6931), .A(n6873), .B(n6872), .ZN(n6875)
         );
  AOI211_X1 U7486 ( .C1(n6877), .C2(n6947), .A(n6876), .B(n6875), .ZN(n6881)
         );
  OAI21_X1 U7487 ( .B1(n6879), .B2(n6878), .A(REIP_REG_7__SCAN_IN), .ZN(n6880)
         );
  OAI211_X1 U7488 ( .C1(n6950), .C2(n6882), .A(n6881), .B(n6880), .ZN(U2820)
         );
  NOR3_X1 U7489 ( .A1(n6884), .A2(REIP_REG_10__SCAN_IN), .A3(n6883), .ZN(n6885) );
  AOI211_X1 U7490 ( .C1(n6939), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6910), 
        .B(n6885), .ZN(n6895) );
  AOI22_X1 U7491 ( .A1(n6946), .A2(n6886), .B1(n6943), .B2(EBX_REG_10__SCAN_IN), .ZN(n6894) );
  INV_X1 U7492 ( .A(n6887), .ZN(n6889) );
  AOI22_X1 U7493 ( .A1(n6889), .A2(n6947), .B1(n6923), .B2(n6888), .ZN(n6893)
         );
  OAI21_X1 U7494 ( .B1(n6891), .B2(n6890), .A(REIP_REG_10__SCAN_IN), .ZN(n6892) );
  NAND4_X1 U7495 ( .A1(n6895), .A2(n6894), .A3(n6893), .A4(n6892), .ZN(U2817)
         );
  AOI22_X1 U7496 ( .A1(n6897), .A2(REIP_REG_12__SCAN_IN), .B1(n6946), .B2(
        n6896), .ZN(n6905) );
  OAI22_X1 U7497 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6899), .B1(n6898), .B2(
        n6907), .ZN(n6900) );
  AOI211_X1 U7498 ( .C1(n6939), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6910), 
        .B(n6900), .ZN(n6904) );
  AOI22_X1 U7499 ( .A1(n6902), .A2(n6947), .B1(n6901), .B2(n6923), .ZN(n6903)
         );
  NAND3_X1 U7500 ( .A1(n6905), .A2(n6904), .A3(n6903), .ZN(U2815) );
  OAI22_X1 U7501 ( .A1(n6908), .A2(n6907), .B1(n5732), .B2(n6906), .ZN(n6909)
         );
  AOI211_X1 U7502 ( .C1(n6939), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6910), 
        .B(n6909), .ZN(n6920) );
  INV_X1 U7503 ( .A(n6911), .ZN(n6912) );
  AOI22_X1 U7504 ( .A1(n6913), .A2(n6947), .B1(n6923), .B2(n6912), .ZN(n6919)
         );
  NAND2_X1 U7505 ( .A1(n6946), .A2(n6914), .ZN(n6918) );
  OAI211_X1 U7506 ( .C1(REIP_REG_12__SCAN_IN), .C2(REIP_REG_13__SCAN_IN), .A(
        n6916), .B(n6915), .ZN(n6917) );
  NAND4_X1 U7507 ( .A1(n6920), .A2(n6919), .A3(n6918), .A4(n6917), .ZN(U2814)
         );
  INV_X1 U7508 ( .A(n6921), .ZN(n6933) );
  NAND2_X1 U7509 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  OAI211_X1 U7510 ( .C1(n6927), .C2(n6926), .A(n6925), .B(n6924), .ZN(n6928)
         );
  AOI21_X1 U7511 ( .B1(n6943), .B2(EBX_REG_18__SCAN_IN), .A(n6928), .ZN(n6929)
         );
  OAI21_X1 U7512 ( .B1(n6931), .B2(n6930), .A(n6929), .ZN(n6932) );
  AOI21_X1 U7513 ( .B1(n6933), .B2(n6947), .A(n6932), .ZN(n6935) );
  OAI211_X1 U7514 ( .C1(n6937), .C2(n6936), .A(n6935), .B(n6934), .ZN(U2809)
         );
  AOI22_X1 U7515 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6939), .B1(
        REIP_REG_21__SCAN_IN), .B2(n6938), .ZN(n6940) );
  INV_X1 U7516 ( .A(n6940), .ZN(n6941) );
  AOI211_X1 U7517 ( .C1(n6943), .C2(EBX_REG_21__SCAN_IN), .A(n6942), .B(n6941), 
        .ZN(n6949) );
  INV_X1 U7518 ( .A(n6944), .ZN(n6945) );
  AOI22_X1 U7519 ( .A1(n7061), .A2(n6947), .B1(n6946), .B2(n6945), .ZN(n6948)
         );
  OAI211_X1 U7520 ( .C1(n6951), .C2(n6950), .A(n6949), .B(n6948), .ZN(U2806)
         );
  OAI21_X1 U7521 ( .B1(n6953), .B2(n5023), .A(n6952), .ZN(U2793) );
  INV_X1 U7522 ( .A(n7003), .ZN(n6957) );
  INV_X1 U7523 ( .A(n6954), .ZN(n6956) );
  OAI22_X1 U7524 ( .A1(n6958), .A2(n6957), .B1(n6956), .B2(n6955), .ZN(n6960)
         );
  MUX2_X1 U7525 ( .A(n6960), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6959), 
        .Z(U3456) );
  INV_X1 U7526 ( .A(n6961), .ZN(n6963) );
  NAND4_X1 U7527 ( .A1(n6963), .A2(n6962), .A3(n7089), .A4(n7011), .ZN(n6965)
         );
  OAI22_X1 U7528 ( .A1(n6966), .A2(n6965), .B1(n3553), .B2(n6964), .ZN(U3455)
         );
  NAND2_X1 U7529 ( .A1(n6968), .A2(n6967), .ZN(n6976) );
  NAND2_X1 U7530 ( .A1(n6969), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6970) );
  NAND2_X1 U7531 ( .A1(n6971), .A2(n6970), .ZN(n6973) );
  OAI21_X1 U7532 ( .B1(n6973), .B2(n7103), .A(n7099), .ZN(n6975) );
  NOR2_X1 U7533 ( .A1(n6973), .A2(n6972), .ZN(n6974) );
  AOI21_X1 U7534 ( .B1(n6976), .B2(n6975), .A(n6974), .ZN(n6977) );
  OAI21_X1 U7535 ( .B1(n6979), .B2(n6978), .A(n6977), .ZN(n6981) );
  NAND2_X1 U7536 ( .A1(n6979), .A2(n6978), .ZN(n6980) );
  AOI22_X1 U7537 ( .A1(n6981), .A2(n6980), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6982), .ZN(n6985) );
  NOR2_X1 U7538 ( .A1(n6982), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6984)
         );
  OAI21_X1 U7539 ( .B1(n6985), .B2(n6984), .A(n6983), .ZN(n6996) );
  AND2_X1 U7540 ( .A1(n5023), .A2(n6986), .ZN(n6990) );
  NOR2_X1 U7541 ( .A1(n6988), .A2(n6987), .ZN(n6989) );
  OAI21_X1 U7542 ( .B1(n6991), .B2(n6990), .A(n6989), .ZN(n6992) );
  NOR3_X1 U7543 ( .A1(n6994), .A2(n6993), .A3(n6992), .ZN(n6995) );
  AND2_X1 U7544 ( .A1(n6996), .A2(n6995), .ZN(n7026) );
  NAND2_X1 U7545 ( .A1(n7026), .A2(n7004), .ZN(n6998) );
  NAND2_X1 U7546 ( .A1(READY_N), .A2(n6696), .ZN(n6997) );
  NAND2_X1 U7547 ( .A1(n6998), .A2(n6997), .ZN(n7002) );
  OR2_X1 U7548 ( .A1(n7000), .A2(n6999), .ZN(n7001) );
  AOI221_X1 U7549 ( .B1(n7014), .B2(n7042), .C1(n7014), .C2(
        STATE2_REG_2__SCAN_IN), .A(n7020), .ZN(n7019) );
  INV_X1 U7550 ( .A(n7019), .ZN(n7010) );
  NAND3_X1 U7551 ( .A1(n7003), .A2(STATE2_REG_0__SCAN_IN), .A3(n7042), .ZN(
        n7005) );
  INV_X1 U7552 ( .A(n7004), .ZN(n7025) );
  NAND3_X1 U7553 ( .A1(n7005), .A2(n7025), .A3(n7014), .ZN(n7006) );
  OAI21_X1 U7554 ( .B1(n7007), .B2(n7014), .A(n7006), .ZN(n7009) );
  OAI211_X1 U7555 ( .C1(n7011), .C2(n7010), .A(n7009), .B(n7008), .ZN(U3149)
         );
  OAI211_X1 U7556 ( .C1(n7014), .C2(n7089), .A(n7013), .B(n7012), .ZN(U3453)
         );
  NOR2_X1 U7557 ( .A1(n7089), .A2(n7015), .ZN(n7018) );
  AOI21_X1 U7558 ( .B1(n7018), .B2(n7017), .A(n7016), .ZN(n7021) );
  AOI221_X1 U7559 ( .B1(n7022), .B2(STATE2_REG_0__SCAN_IN), .C1(n7021), .C2(
        n7020), .A(n7019), .ZN(n7024) );
  OAI211_X1 U7560 ( .C1(n7026), .C2(n7025), .A(n7024), .B(n7023), .ZN(U3148)
         );
  INV_X1 U7561 ( .A(n7027), .ZN(n7029) );
  OAI21_X1 U7562 ( .B1(n7031), .B2(n7028), .A(n7029), .ZN(U2792) );
  OAI21_X1 U7563 ( .B1(n7031), .B2(n7030), .A(n7029), .ZN(U3452) );
  NOR2_X1 U7564 ( .A1(n7032), .A2(n7034), .ZN(n7039) );
  NOR2_X1 U7565 ( .A1(n7034), .A2(n7033), .ZN(n7036) );
  AOI221_X1 U7566 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7040), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7045) );
  AOI221_X1 U7567 ( .B1(n7036), .B2(n7048), .C1(n7035), .C2(n7048), .A(n7045), 
        .ZN(n7037) );
  OAI221_X1 U7568 ( .B1(n7039), .B2(n7038), .C1(n7039), .C2(n7046), .A(n7037), 
        .ZN(U3181) );
  AOI21_X1 U7569 ( .B1(n7041), .B2(n7040), .A(STATE_REG_2__SCAN_IN), .ZN(n7047) );
  AOI221_X1 U7570 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7042), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7043) );
  AOI221_X1 U7571 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7043), .C2(HOLD), .A(n3662), .ZN(n7044) );
  OAI22_X1 U7572 ( .A1(n7047), .A2(n7046), .B1(n7045), .B2(n7044), .ZN(U3183)
         );
  INV_X1 U7573 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7049) );
  AOI22_X1 U7574 ( .A1(n7051), .A2(n7050), .B1(n7049), .B2(n7048), .ZN(U3473)
         );
  AOI22_X1 U7576 ( .A1(n7053), .A2(n7207), .B1(n7059), .B2(DATAI_1_), .ZN(
        n7055) );
  AOI22_X1 U7577 ( .A1(n7063), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n7062), .ZN(n7054) );
  NAND2_X1 U7578 ( .A1(n7055), .A2(n7054), .ZN(U2874) );
  AOI22_X1 U7579 ( .A1(n7056), .A2(n7207), .B1(n7059), .B2(DATAI_3_), .ZN(
        n7058) );
  AOI22_X1 U7580 ( .A1(n7063), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n7062), .ZN(n7057) );
  NAND2_X1 U7581 ( .A1(n7058), .A2(n7057), .ZN(U2872) );
  AOI22_X1 U7582 ( .A1(n7061), .A2(n7207), .B1(n7059), .B2(DATAI_5_), .ZN(
        n7065) );
  AOI22_X1 U7583 ( .A1(n7063), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n7062), .ZN(n7064) );
  NAND2_X1 U7584 ( .A1(n7065), .A2(n7064), .ZN(U2870) );
  AOI21_X1 U7585 ( .B1(n7078), .B2(n7066), .A(n7081), .ZN(n7076) );
  INV_X1 U7586 ( .A(n7076), .ZN(n7070) );
  NAND2_X1 U7587 ( .A1(n7067), .A2(n7084), .ZN(n7069) );
  NOR3_X1 U7588 ( .A1(n7068), .A2(n7099), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n7072) );
  NAND2_X1 U7589 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7072), .ZN(n7071) );
  NAND2_X1 U7590 ( .A1(n7069), .A2(n7071), .ZN(n7075) );
  AOI22_X1 U7591 ( .A1(n7070), .A2(n7075), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7072), .ZN(n7186) );
  INV_X1 U7592 ( .A(n7071), .ZN(n7181) );
  AOI22_X1 U7593 ( .A1(n7182), .A2(n7110), .B1(n7109), .B2(n7181), .ZN(n7080)
         );
  INV_X1 U7594 ( .A(n7072), .ZN(n7088) );
  AOI21_X1 U7595 ( .B1(n7112), .B2(n7088), .A(n7073), .ZN(n7074) );
  OAI21_X1 U7596 ( .B1(n7076), .B2(n7075), .A(n7074), .ZN(n7183) );
  NOR2_X2 U7597 ( .A1(n7078), .A2(n7077), .ZN(n7189) );
  AOI22_X1 U7598 ( .A1(n7183), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n7117), 
        .B2(n7189), .ZN(n7079) );
  OAI211_X1 U7599 ( .C1(n7186), .C2(n7120), .A(n7080), .B(n7079), .ZN(U3108)
         );
  NOR3_X1 U7600 ( .A1(n3419), .A2(n7189), .A3(n7112), .ZN(n7082) );
  NOR2_X1 U7601 ( .A1(n7082), .A2(n7081), .ZN(n7095) );
  INV_X1 U7602 ( .A(n7095), .ZN(n7087) );
  AND2_X1 U7603 ( .A1(n7084), .A2(n7083), .ZN(n7094) );
  NOR2_X1 U7604 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7088), .ZN(n7187)
         );
  AOI22_X1 U7605 ( .A1(n3419), .A2(n7117), .B1(n7109), .B2(n7187), .ZN(n7097)
         );
  INV_X1 U7606 ( .A(n7187), .ZN(n7092) );
  AOI211_X1 U7607 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n7092), .A(n7091), .B(
        n7090), .ZN(n7093) );
  OAI21_X1 U7608 ( .B1(n7095), .B2(n7094), .A(n7093), .ZN(n7190) );
  AOI22_X1 U7609 ( .A1(n7190), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n7110), 
        .B2(n7189), .ZN(n7096) );
  OAI211_X1 U7610 ( .C1(n7193), .C2(n7120), .A(n7097), .B(n7096), .ZN(U3100)
         );
  NAND2_X1 U7611 ( .A1(n7099), .A2(n7098), .ZN(n7111) );
  INV_X1 U7612 ( .A(n7111), .ZN(n7107) );
  INV_X1 U7613 ( .A(n7100), .ZN(n7102) );
  OAI21_X1 U7614 ( .B1(n7102), .B2(n7112), .A(n7101), .ZN(n7114) );
  NOR2_X1 U7615 ( .A1(n7103), .A2(n7111), .ZN(n7194) );
  AOI21_X1 U7616 ( .B1(n7105), .B2(n7104), .A(n7194), .ZN(n7113) );
  INV_X1 U7617 ( .A(n7113), .ZN(n7106) );
  AOI22_X1 U7618 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7107), .B1(n7114), .B2(
        n7106), .ZN(n7204) );
  AOI22_X1 U7619 ( .A1(n7198), .A2(n7110), .B1(n7109), .B2(n7194), .ZN(n7119)
         );
  AOI22_X1 U7620 ( .A1(n7114), .A2(n7113), .B1(n7112), .B2(n7111), .ZN(n7115)
         );
  NAND2_X1 U7621 ( .A1(n7116), .A2(n7115), .ZN(n7200) );
  AOI22_X1 U7622 ( .A1(n7200), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n7117), 
        .B2(n7197), .ZN(n7118) );
  OAI211_X1 U7623 ( .C1(n7204), .C2(n7120), .A(n7119), .B(n7118), .ZN(U3028)
         );
  AOI22_X1 U7624 ( .A1(n7189), .A2(n7126), .B1(n7125), .B2(n7181), .ZN(n7122)
         );
  AOI22_X1 U7625 ( .A1(n7183), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n7127), 
        .B2(n7182), .ZN(n7121) );
  OAI211_X1 U7626 ( .C1(n7186), .C2(n7130), .A(n7122), .B(n7121), .ZN(U3109)
         );
  AOI22_X1 U7627 ( .A1(n3419), .A2(n7126), .B1(n7125), .B2(n7187), .ZN(n7124)
         );
  AOI22_X1 U7628 ( .A1(n7190), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n7127), 
        .B2(n7189), .ZN(n7123) );
  OAI211_X1 U7629 ( .C1(n7193), .C2(n7130), .A(n7124), .B(n7123), .ZN(U3101)
         );
  AOI22_X1 U7630 ( .A1(n7197), .A2(n7126), .B1(n7125), .B2(n7194), .ZN(n7129)
         );
  AOI22_X1 U7631 ( .A1(n7200), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n7127), 
        .B2(n7198), .ZN(n7128) );
  OAI211_X1 U7632 ( .C1(n7204), .C2(n7130), .A(n7129), .B(n7128), .ZN(U3029)
         );
  AOI22_X1 U7633 ( .A1(n7189), .A2(n7137), .B1(n7135), .B2(n7181), .ZN(n7132)
         );
  AOI22_X1 U7634 ( .A1(n7183), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n7136), 
        .B2(n7182), .ZN(n7131) );
  OAI211_X1 U7635 ( .C1(n7186), .C2(n7140), .A(n7132), .B(n7131), .ZN(U3110)
         );
  AOI22_X1 U7636 ( .A1(n3419), .A2(n7137), .B1(n7135), .B2(n7187), .ZN(n7134)
         );
  AOI22_X1 U7637 ( .A1(n7190), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n7136), 
        .B2(n7189), .ZN(n7133) );
  OAI211_X1 U7638 ( .C1(n7193), .C2(n7140), .A(n7134), .B(n7133), .ZN(U3102)
         );
  AOI22_X1 U7639 ( .A1(n7198), .A2(n7136), .B1(n7135), .B2(n7194), .ZN(n7139)
         );
  AOI22_X1 U7640 ( .A1(n7200), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n7137), 
        .B2(n7197), .ZN(n7138) );
  OAI211_X1 U7641 ( .C1(n7204), .C2(n7140), .A(n7139), .B(n7138), .ZN(U3030)
         );
  AOI22_X1 U7642 ( .A1(n7189), .A2(n7147), .B1(n7145), .B2(n7181), .ZN(n7142)
         );
  AOI22_X1 U7643 ( .A1(n7183), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n7146), 
        .B2(n7182), .ZN(n7141) );
  OAI211_X1 U7644 ( .C1(n7186), .C2(n7150), .A(n7142), .B(n7141), .ZN(U3111)
         );
  AOI22_X1 U7645 ( .A1(n3419), .A2(n7147), .B1(n7145), .B2(n7187), .ZN(n7144)
         );
  AOI22_X1 U7646 ( .A1(n7190), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n7146), 
        .B2(n7189), .ZN(n7143) );
  OAI211_X1 U7647 ( .C1(n7193), .C2(n7150), .A(n7144), .B(n7143), .ZN(U3103)
         );
  AOI22_X1 U7648 ( .A1(n7198), .A2(n7146), .B1(n7145), .B2(n7194), .ZN(n7149)
         );
  AOI22_X1 U7649 ( .A1(n7200), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n7147), 
        .B2(n7197), .ZN(n7148) );
  OAI211_X1 U7650 ( .C1(n7204), .C2(n7150), .A(n7149), .B(n7148), .ZN(U3031)
         );
  AOI22_X1 U7651 ( .A1(n7189), .A2(n7156), .B1(n7155), .B2(n7181), .ZN(n7152)
         );
  AOI22_X1 U7652 ( .A1(n7183), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n7157), 
        .B2(n7182), .ZN(n7151) );
  OAI211_X1 U7653 ( .C1(n7186), .C2(n7160), .A(n7152), .B(n7151), .ZN(U3112)
         );
  AOI22_X1 U7654 ( .A1(n3419), .A2(n7156), .B1(n7155), .B2(n7187), .ZN(n7154)
         );
  AOI22_X1 U7655 ( .A1(n7190), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n7157), 
        .B2(n7189), .ZN(n7153) );
  OAI211_X1 U7656 ( .C1(n7193), .C2(n7160), .A(n7154), .B(n7153), .ZN(U3104)
         );
  AOI22_X1 U7657 ( .A1(n7197), .A2(n7156), .B1(n7155), .B2(n7194), .ZN(n7159)
         );
  AOI22_X1 U7658 ( .A1(n7200), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n7157), 
        .B2(n7198), .ZN(n7158) );
  OAI211_X1 U7659 ( .C1(n7204), .C2(n7160), .A(n7159), .B(n7158), .ZN(U3032)
         );
  AOI22_X1 U7660 ( .A1(n7182), .A2(n7166), .B1(n7165), .B2(n7181), .ZN(n7162)
         );
  AOI22_X1 U7661 ( .A1(n7183), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n7167), 
        .B2(n7189), .ZN(n7161) );
  OAI211_X1 U7662 ( .C1(n7186), .C2(n7170), .A(n7162), .B(n7161), .ZN(U3113)
         );
  AOI22_X1 U7663 ( .A1(n3419), .A2(n7167), .B1(n7165), .B2(n7187), .ZN(n7164)
         );
  AOI22_X1 U7664 ( .A1(n7190), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n7166), 
        .B2(n7189), .ZN(n7163) );
  OAI211_X1 U7665 ( .C1(n7193), .C2(n7170), .A(n7164), .B(n7163), .ZN(U3105)
         );
  AOI22_X1 U7666 ( .A1(n7198), .A2(n7166), .B1(n7165), .B2(n7194), .ZN(n7169)
         );
  AOI22_X1 U7667 ( .A1(n7200), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n7167), 
        .B2(n7197), .ZN(n7168) );
  OAI211_X1 U7668 ( .C1(n7204), .C2(n7170), .A(n7169), .B(n7168), .ZN(U3033)
         );
  AOI22_X1 U7669 ( .A1(n7189), .A2(n7176), .B1(n7175), .B2(n7181), .ZN(n7172)
         );
  AOI22_X1 U7670 ( .A1(n7183), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n7177), 
        .B2(n7182), .ZN(n7171) );
  OAI211_X1 U7671 ( .C1(n7186), .C2(n7180), .A(n7172), .B(n7171), .ZN(U3114)
         );
  AOI22_X1 U7672 ( .A1(n3419), .A2(n7176), .B1(n7175), .B2(n7187), .ZN(n7174)
         );
  AOI22_X1 U7673 ( .A1(n7190), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n7177), 
        .B2(n7189), .ZN(n7173) );
  OAI211_X1 U7674 ( .C1(n7193), .C2(n7180), .A(n7174), .B(n7173), .ZN(U3106)
         );
  AOI22_X1 U7675 ( .A1(n7197), .A2(n7176), .B1(n7175), .B2(n7194), .ZN(n7179)
         );
  AOI22_X1 U7676 ( .A1(n7200), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n7177), 
        .B2(n7198), .ZN(n7178) );
  OAI211_X1 U7677 ( .C1(n7204), .C2(n7180), .A(n7179), .B(n7178), .ZN(U3034)
         );
  AOI22_X1 U7678 ( .A1(n7182), .A2(n7199), .B1(n7195), .B2(n7181), .ZN(n7185)
         );
  AOI22_X1 U7679 ( .A1(n7183), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n7196), 
        .B2(n7189), .ZN(n7184) );
  OAI211_X1 U7680 ( .C1(n7186), .C2(n7203), .A(n7185), .B(n7184), .ZN(U3115)
         );
  AOI22_X1 U7681 ( .A1(n3419), .A2(n7196), .B1(n7195), .B2(n7187), .ZN(n7192)
         );
  AOI22_X1 U7682 ( .A1(n7190), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n7199), 
        .B2(n7189), .ZN(n7191) );
  OAI211_X1 U7683 ( .C1(n7193), .C2(n7203), .A(n7192), .B(n7191), .ZN(U3107)
         );
  AOI22_X1 U7684 ( .A1(n7197), .A2(n7196), .B1(n7195), .B2(n7194), .ZN(n7202)
         );
  AOI22_X1 U7685 ( .A1(n7200), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n7199), 
        .B2(n7198), .ZN(n7201) );
  OAI211_X1 U7686 ( .C1(n7204), .C2(n7203), .A(n7202), .B(n7201), .ZN(U3035)
         );
  AND2_X1 U3641 ( .A1(n3453), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3459)
         );
  NAND2_X1 U4109 ( .A1(n4925), .A2(n3689), .ZN(n3837) );
  BUF_X1 U34610 ( .A(n3654), .Z(n5697) );
  CLKBUF_X1 U34550 ( .A(n3638), .Z(n4672) );
  AND2_X4 U3566 ( .A1(n3426), .A2(n5014), .ZN(n4644) );
  AND4_X1 U4042 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3587)
         );
  OR2_X1 U4513 ( .A1(n3961), .A2(n3960), .ZN(n4104) );
  XNOR2_X1 U3503 ( .A(n3967), .B(n3966), .ZN(n3968) );
  CLKBUF_X1 U34530 ( .A(n4698), .Z(n4624) );
  CLKBUF_X1 U34690 ( .A(n3921), .Z(n4705) );
  AND2_X1 U34710 ( .A1(n4987), .A2(n4986), .ZN(n3629) );
  CLKBUF_X2 U34730 ( .A(n3725), .Z(n3812) );
  CLKBUF_X1 U3486 ( .A(n4755), .Z(n3425) );
  CLKBUF_X1 U3495 ( .A(n6004), .Z(n6005) );
  AND2_X1 U3496 ( .A1(n5788), .A2(n3776), .ZN(n5712) );
  CLKBUF_X1 U3501 ( .A(n3727), .Z(n3436) );
  CLKBUF_X1 U3519 ( .A(n6534), .Z(n6549) );
  CLKBUF_X1 U3537 ( .A(n4904), .Z(n5300) );
  AOI21_X1 U3557 ( .B1(n3441), .B2(n6670), .A(n6317), .ZN(n6318) );
  OR2_X1 U3745 ( .A1(n5270), .A2(n4906), .ZN(n7205) );
  OR2_X1 U3796 ( .A1(n5926), .A2(n6800), .ZN(n7206) );
  AND2_X1 U3798 ( .A1(n6287), .A2(n4903), .ZN(n7207) );
endmodule

