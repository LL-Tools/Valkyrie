

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4380, n4381, n4383, n4384, n4385, n4386, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10481;

  NAND2_X1 U4885 ( .A1(n8811), .A2(n6562), .ZN(n8820) );
  NAND2_X1 U4886 ( .A1(n5454), .A2(n5453), .ZN(n10138) );
  BUF_X1 U4887 ( .A(n6588), .Z(n6598) );
  NAND2_X1 U4888 ( .A1(n5408), .A2(n5407), .ZN(n5424) );
  CLKBUF_X2 U4889 ( .A(n6659), .Z(n4396) );
  INV_X1 U4890 ( .A(n6875), .ZN(n6663) );
  INV_X2 U4891 ( .A(n6847), .ZN(n6690) );
  CLKBUF_X2 U4892 ( .A(n5831), .Z(n6043) );
  NAND2_X1 U4893 ( .A1(n5478), .A2(n5660), .ZN(n9857) );
  CLKBUF_X2 U4894 ( .A(n8454), .Z(n4394) );
  INV_X1 U4895 ( .A(n8445), .ZN(n5777) );
  CLKBUF_X2 U4896 ( .A(n5952), .Z(n5984) );
  NAND2_X1 U4897 ( .A1(n4973), .A2(n10216), .ZN(n5083) );
  NOR2_X1 U4898 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5065) );
  CLKBUF_X1 U4899 ( .A(n9545), .Z(n4380) );
  OAI21_X1 U4900 ( .B1(n6882), .B2(n6887), .A(n9898), .ZN(n9545) );
  INV_X1 U4901 ( .A(n10481), .ZN(n4381) );
  INV_X2 U4902 ( .A(n4381), .ZN(P1_U3084) );
  INV_X1 U4903 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n10481) );
  AND3_X1 U4904 ( .A1(n5663), .A2(n4758), .A3(n4681), .ZN(n4660) );
  NAND2_X1 U4905 ( .A1(n6487), .A2(n6486), .ZN(n6588) );
  NAND2_X1 U4906 ( .A1(n7313), .A2(n10326), .ZN(n10309) );
  INV_X1 U4907 ( .A(n6588), .ZN(n6603) );
  NAND2_X1 U4908 ( .A1(n9148), .A2(n6201), .ZN(n9130) );
  INV_X1 U4909 ( .A(n5799), .ZN(n6021) );
  AND2_X1 U4910 ( .A1(n7679), .A2(n6308), .ZN(n7745) );
  NAND2_X1 U4911 ( .A1(n8699), .A2(n9765), .ZN(n8470) );
  OAI21_X1 U4912 ( .B1(n8820), .B2(n4457), .A(n4955), .ZN(n4954) );
  NOR2_X1 U4913 ( .A1(n4418), .A2(n9394), .ZN(n9133) );
  AND2_X1 U4914 ( .A1(n5952), .A2(n5747), .ZN(n5015) );
  INV_X2 U4915 ( .A(n6875), .ZN(n6868) );
  INV_X1 U4916 ( .A(n9673), .ZN(n7461) );
  NOR2_X1 U4917 ( .A1(n7797), .A2(n10174), .ZN(n7796) );
  NAND2_X2 U4918 ( .A1(n4560), .A2(n5699), .ZN(n7358) );
  AND2_X1 U4919 ( .A1(n5614), .A2(n5613), .ZN(n9519) );
  AND4_X1 U4920 ( .A1(n5140), .A2(n5139), .A3(n5138), .A4(n5137), .ZN(n7445)
         );
  OAI21_X1 U4922 ( .B1(n5326), .B2(P1_IR_REG_0__SCAN_IN), .A(n4526), .ZN(n7366) );
  INV_X1 U4923 ( .A(n7649), .ZN(n9671) );
  NAND2_X1 U4924 ( .A1(n5778), .A2(n5777), .ZN(n4383) );
  OR2_X1 U4925 ( .A1(n8681), .A2(n8702), .ZN(n4384) );
  OR2_X1 U4926 ( .A1(n9863), .A2(n8682), .ZN(n5005) );
  AND4_X2 U4927 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n5793)
         );
  AND2_X2 U4928 ( .A1(n6452), .A2(n4472), .ZN(n4824) );
  AND2_X2 U4929 ( .A1(n5220), .A2(n5219), .ZN(n5281) );
  OAI21_X2 U4930 ( .B1(n7610), .B2(n4459), .A(n4947), .ZN(n8870) );
  NOR2_X1 U4931 ( .A1(n9676), .A2(n7366), .ZN(n7361) );
  XNOR2_X2 U4932 ( .A(n5424), .B(n5055), .ZN(n7184) );
  NAND2_X2 U4933 ( .A1(n4995), .A2(n4992), .ZN(n9785) );
  NOR4_X2 U4934 ( .A1(n6452), .A2(n8316), .A3(n8371), .A4(n6451), .ZN(n6454)
         );
  INV_X1 U4935 ( .A(n4383), .ZN(n4385) );
  INV_X2 U4936 ( .A(n4383), .ZN(n4386) );
  BUF_X4 U4938 ( .A(n5218), .Z(n8464) );
  NAND2_X1 U4939 ( .A1(n6487), .A2(n6486), .ZN(n4388) );
  NAND2_X1 U4940 ( .A1(n6487), .A2(n6486), .ZN(n4389) );
  XNOR2_X2 U4941 ( .A(n6161), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6168) );
  OAI211_X4 U4942 ( .C1(n5813), .C2(n4727), .A(n5814), .B(n4726), .ZN(n8931)
         );
  OR2_X1 U4943 ( .A1(n9130), .A2(n9137), .ZN(n4815) );
  NAND2_X1 U4944 ( .A1(n7458), .A2(n7459), .ZN(n4509) );
  NAND2_X1 U4945 ( .A1(n5512), .A2(n5511), .ZN(n10118) );
  NAND2_X1 U4946 ( .A1(n4515), .A2(n4444), .ZN(n7393) );
  AND2_X1 U4947 ( .A1(n4504), .A2(n4503), .ZN(n4502) );
  INV_X1 U4948 ( .A(n9455), .ZN(n9357) );
  NAND2_X1 U4949 ( .A1(n4532), .A2(n5262), .ZN(n10174) );
  NAND2_X1 U4950 ( .A1(n5222), .A2(n5221), .ZN(n7640) );
  CLKBUF_X2 U4951 ( .A(n6658), .Z(n4395) );
  AND4_X1 U4952 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n7876)
         );
  INV_X1 U4953 ( .A(n7688), .ZN(n6497) );
  INV_X2 U4954 ( .A(n5631), .ZN(n5718) );
  INV_X1 U4955 ( .A(n7176), .ZN(n10286) );
  CLKBUF_X2 U4956 ( .A(n5174), .Z(n5631) );
  INV_X2 U4957 ( .A(n5716), .ZN(n8456) );
  INV_X1 U4958 ( .A(n7720), .ZN(n10365) );
  INV_X4 U4959 ( .A(n5154), .ZN(n5179) );
  INV_X1 U4960 ( .A(n6488), .ZN(n10326) );
  INV_X4 U4962 ( .A(n5840), .ZN(n6056) );
  CLKBUF_X2 U4963 ( .A(n8454), .Z(n4393) );
  INV_X1 U4964 ( .A(n6986), .ZN(n8454) );
  INV_X1 U4965 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5744) );
  INV_X1 U4966 ( .A(n6870), .ZN(n9517) );
  NAND2_X1 U4967 ( .A1(n4512), .A2(n6857), .ZN(n9638) );
  OR2_X1 U4968 ( .A1(n4820), .A2(n10405), .ZN(n4520) );
  AND2_X1 U4969 ( .A1(n4521), .A2(n9384), .ZN(n4820) );
  NAND2_X1 U4970 ( .A1(n6836), .A2(n6835), .ZN(n9526) );
  NAND2_X1 U4971 ( .A1(n9525), .A2(n9528), .ZN(n6837) );
  OAI21_X1 U4972 ( .B1(n9130), .B2(n4811), .A(n4808), .ZN(n6223) );
  AND2_X1 U4973 ( .A1(n4643), .A2(n4565), .ZN(n9799) );
  OR2_X1 U4974 ( .A1(n4981), .A2(n4982), .ZN(n4980) );
  AOI21_X1 U4975 ( .B1(n4833), .B2(n9180), .A(n4460), .ZN(n4831) );
  NAND2_X1 U4976 ( .A1(n5522), .A2(n5521), .ZN(n9885) );
  NAND2_X1 U4977 ( .A1(n9890), .A2(n9889), .ZN(n5522) );
  NAND2_X1 U4978 ( .A1(n8597), .A2(n8594), .ZN(n9851) );
  NAND2_X1 U4979 ( .A1(n9220), .A2(n9222), .ZN(n9221) );
  NAND2_X1 U4980 ( .A1(n5588), .A2(n5587), .ZN(n10099) );
  NAND2_X1 U4981 ( .A1(n9970), .A2(n5444), .ZN(n4971) );
  NAND2_X1 U4982 ( .A1(n6088), .A2(n6418), .ZN(n9137) );
  NAND2_X1 U4983 ( .A1(n9989), .A2(n5423), .ZN(n9970) );
  INV_X1 U4984 ( .A(n6587), .ZN(n4943) );
  INV_X1 U4985 ( .A(n9519), .ZN(n9829) );
  NAND2_X1 U4986 ( .A1(n4693), .A2(n4692), .ZN(n4697) );
  AND2_X1 U4987 ( .A1(n9778), .A2(n5645), .ZN(n6890) );
  OR2_X1 U4988 ( .A1(n5644), .A2(n8047), .ZN(n9778) );
  NAND2_X1 U4989 ( .A1(n5550), .A2(n5549), .ZN(n10109) );
  OR2_X1 U4990 ( .A1(n9934), .A2(n10124), .ZN(n9917) );
  AND2_X1 U4991 ( .A1(n5708), .A2(n4694), .ZN(n4692) );
  XNOR2_X1 U4992 ( .A(n5579), .B(n5577), .ZN(n8395) );
  AND2_X1 U4993 ( .A1(n5596), .A2(n5595), .ZN(n9853) );
  NAND2_X1 U4994 ( .A1(n6049), .A2(n6048), .ZN(n9415) );
  NAND2_X1 U4995 ( .A1(n6040), .A2(n6039), .ZN(n9420) );
  AOI21_X1 U4996 ( .B1(n4824), .B2(n4483), .A(n4425), .ZN(n4482) );
  NAND2_X1 U4997 ( .A1(n4589), .A2(n4594), .ZN(n5561) );
  NAND2_X1 U4998 ( .A1(n9238), .A2(n6371), .ZN(n9292) );
  NAND2_X1 U4999 ( .A1(n5494), .A2(n5493), .ZN(n10124) );
  NOR2_X1 U5000 ( .A1(n5031), .A2(n10164), .ZN(n10050) );
  NAND2_X1 U5001 ( .A1(n5481), .A2(n5480), .ZN(n10133) );
  NAND2_X1 U5002 ( .A1(n5510), .A2(n5509), .ZN(n5528) );
  OR2_X1 U5003 ( .A1(n10159), .A2(n9656), .ZN(n8619) );
  NAND2_X1 U5004 ( .A1(n5415), .A2(n5414), .ZN(n10149) );
  NAND2_X1 U5005 ( .A1(n5989), .A2(n5988), .ZN(n9445) );
  NAND2_X2 U5006 ( .A1(n6000), .A2(n5999), .ZN(n9442) );
  NAND2_X1 U5007 ( .A1(n5967), .A2(n5966), .ZN(n9455) );
  NAND2_X1 U5008 ( .A1(n5435), .A2(n5434), .ZN(n10144) );
  NAND2_X1 U5009 ( .A1(n5566), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U5010 ( .A1(n5393), .A2(n5392), .ZN(n10154) );
  XNOR2_X1 U5011 ( .A(n5465), .B(n5464), .ZN(n7351) );
  AND2_X1 U5012 ( .A1(n8618), .A2(n8320), .ZN(n8627) );
  XNOR2_X1 U5013 ( .A(n5359), .B(n5377), .ZN(n7145) );
  NAND2_X1 U5014 ( .A1(n5955), .A2(n5954), .ZN(n9460) );
  XNOR2_X1 U5015 ( .A(n5388), .B(n5402), .ZN(n7152) );
  NAND2_X2 U5016 ( .A1(n7657), .A2(n9359), .ZN(n10335) );
  NAND2_X1 U5017 ( .A1(n7507), .A2(n4426), .ZN(n7591) );
  XNOR2_X1 U5018 ( .A(n5356), .B(n5355), .ZN(n7125) );
  NAND2_X1 U5019 ( .A1(n5305), .A2(n5304), .ZN(n8411) );
  NAND2_X1 U5020 ( .A1(n5916), .A2(n5915), .ZN(n9470) );
  NAND2_X1 U5021 ( .A1(n5406), .A2(n5405), .ZN(n5408) );
  NAND2_X1 U5022 ( .A1(n7444), .A2(n8477), .ZN(n7507) );
  NAND2_X1 U5023 ( .A1(n5381), .A2(n5373), .ZN(n5356) );
  NAND2_X1 U5024 ( .A1(n4615), .A2(n5922), .ZN(n8229) );
  AND2_X1 U5025 ( .A1(n5898), .A2(n5897), .ZN(n7828) );
  AND2_X1 U5026 ( .A1(n4979), .A2(n7634), .ZN(n4409) );
  NAND2_X1 U5027 ( .A1(n4841), .A2(n5876), .ZN(n10397) );
  NAND2_X1 U5028 ( .A1(n5416), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U5029 ( .A1(n5243), .A2(n5242), .ZN(n10179) );
  INV_X2 U5030 ( .A(n9940), .ZN(n10062) );
  INV_X1 U5031 ( .A(n5418), .ZN(n5416) );
  NOR2_X1 U5032 ( .A1(n6882), .A2(n6872), .ZN(n9650) );
  NAND2_X1 U5033 ( .A1(n5891), .A2(n5890), .ZN(n7622) );
  INV_X1 U5034 ( .A(n6679), .ZN(n7553) );
  AND2_X1 U5035 ( .A1(n8568), .A2(n8563), .ZN(n8474) );
  NAND2_X1 U5036 ( .A1(n6287), .A2(n6288), .ZN(n7681) );
  AND2_X1 U5037 ( .A1(n7758), .A2(n7632), .ZN(n8578) );
  NAND2_X1 U5038 ( .A1(n8929), .A2(n6497), .ZN(n6287) );
  OR2_X1 U5039 ( .A1(n7257), .A2(n7176), .ZN(n7452) );
  NAND2_X1 U5040 ( .A1(n4612), .A2(n5232), .ZN(n4611) );
  INV_X1 U5041 ( .A(n7445), .ZN(n9675) );
  NAND2_X1 U5042 ( .A1(n5857), .A2(n5856), .ZN(n7738) );
  NAND2_X1 U5043 ( .A1(n5092), .A2(n5091), .ZN(n9676) );
  NAND2_X1 U5044 ( .A1(n5763), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6009) );
  AND4_X1 U5045 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n7730)
         );
  INV_X1 U5046 ( .A(n8930), .ZN(n5808) );
  NAND4_X1 U5047 ( .A1(n5183), .A2(n5182), .A3(n5181), .A4(n5180), .ZN(n9673)
         );
  INV_X1 U5048 ( .A(n7315), .ZN(n6293) );
  NAND2_X1 U5049 ( .A1(n5306), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5331) );
  INV_X1 U5050 ( .A(n7366), .ZN(n7179) );
  AOI21_X1 U5051 ( .B1(n5090), .B2(P1_REG0_REG_0__SCAN_IN), .A(n5089), .ZN(
        n5091) );
  AND3_X2 U5052 ( .A1(n5134), .A2(n5133), .A3(n4648), .ZN(n7424) );
  NAND3_X1 U5053 ( .A1(n6485), .A2(n6484), .A3(n7768), .ZN(n6486) );
  OAI211_X1 U5054 ( .C1(n7008), .C2(n5166), .A(n5152), .B(n5151), .ZN(n7176)
         );
  AOI21_X1 U5055 ( .B1(n8976), .B2(n8975), .A(n8974), .ZN(n8991) );
  NAND2_X1 U5056 ( .A1(n4848), .A2(n4846), .ZN(n8726) );
  BUF_X2 U5057 ( .A(n5179), .Z(n8457) );
  OR2_X1 U5058 ( .A1(n5432), .A2(n7018), .ZN(n5112) );
  INV_X1 U5059 ( .A(n9154), .ZN(n6278) );
  INV_X2 U5060 ( .A(n5326), .ZN(n5479) );
  NAND2_X1 U5061 ( .A1(n6160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6161) );
  NAND2_X2 U5062 ( .A1(n6160), .A2(n6020), .ZN(n9154) );
  CLKBUF_X1 U5063 ( .A(n5841), .Z(n6248) );
  XNOR2_X1 U5064 ( .A(n6165), .B(n5744), .ZN(n7768) );
  NAND2_X1 U5065 ( .A1(n6019), .A2(n6127), .ZN(n6160) );
  NAND2_X1 U5066 ( .A1(n5672), .A2(n4551), .ZN(n8433) );
  NAND2_X1 U5067 ( .A1(n4910), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U5068 ( .A1(n5799), .A2(n8454), .ZN(n5841) );
  NAND2_X1 U5069 ( .A1(n6018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6019) );
  NAND2_X2 U5070 ( .A1(n4394), .A2(P1_U3084), .ZN(n10232) );
  NAND2_X1 U5071 ( .A1(n5244), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U5073 ( .A1(n5080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4972) );
  OR2_X1 U5074 ( .A1(n5674), .A2(n5673), .ZN(n4551) );
  MUX2_X1 U5075 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5770), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5773) );
  MUX2_X1 U5076 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5477), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5478) );
  NAND2_X1 U5077 ( .A1(n5235), .A2(n8198), .ZN(n5295) );
  NOR2_X1 U5078 ( .A1(n4537), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U5079 ( .A1(n4936), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6017) );
  NOR2_X1 U5080 ( .A1(n5475), .A2(n4908), .ZN(n4912) );
  XNOR2_X1 U5081 ( .A(n5150), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6984) );
  AND2_X1 U5082 ( .A1(n4511), .A2(n4510), .ZN(n5672) );
  NAND2_X1 U5083 ( .A1(n5774), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5776) );
  INV_X1 U5084 ( .A(n5184), .ZN(n4390) );
  AND3_X2 U5085 ( .A1(n5474), .A2(n5473), .A3(n5472), .ZN(n5668) );
  AND2_X1 U5086 ( .A1(n5738), .A2(n5737), .ZN(n5933) );
  AND3_X1 U5087 ( .A1(n4919), .A2(n4918), .A3(n4917), .ZN(n5740) );
  CLKBUF_X1 U5088 ( .A(n5785), .Z(n5838) );
  INV_X1 U5089 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5673) );
  NOR2_X1 U5090 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5066) );
  INV_X1 U5091 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5678) );
  NOR2_X1 U5092 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5738) );
  NOR2_X1 U5093 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5737) );
  INV_X2 U5094 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5110) );
  INV_X2 U5095 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10240) );
  NOR2_X1 U5096 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5785) );
  NOR2_X1 U5097 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5069) );
  NOR2_X1 U5098 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5070) );
  INV_X1 U5099 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5167) );
  NAND3_X1 U5100 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5206) );
  INV_X4 U5101 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5102 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5279) );
  INV_X1 U5103 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5278) );
  INV_X1 U5104 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9751) );
  NOR2_X1 U5105 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5741) );
  INV_X1 U5106 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6131) );
  INV_X1 U5107 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6144) );
  NOR2_X1 U5108 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5736) );
  NOR2_X1 U5109 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4917) );
  NOR2_X1 U5110 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4918) );
  NOR2_X1 U5111 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4919) );
  INV_X1 U5112 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U5113 ( .A1(n5660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U5114 ( .A1(n5793), .A2(n7720), .ZN(n7746) );
  NAND2_X1 U5115 ( .A1(n5101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5103) );
  AND2_X1 U5116 ( .A1(n5778), .A2(n8445), .ZN(n5818) );
  XNOR2_X1 U5117 ( .A(n5103), .B(n5102), .ZN(n5720) );
  AOI21_X1 U5118 ( .B1(n6317), .B2(n6316), .A(n6315), .ZN(n6334) );
  OAI22_X2 U5119 ( .A1(n8838), .A2(n8837), .B1(n6577), .B2(n6576), .ZN(n8771)
         );
  NOR2_X2 U5120 ( .A1(n4397), .A2(n9455), .ZN(n9355) );
  NAND2_X2 U5121 ( .A1(n7393), .A2(n6687), .ZN(n7458) );
  AND2_X1 U5122 ( .A1(n6413), .A2(n4583), .ZN(n4547) );
  INV_X1 U5123 ( .A(n5668), .ZN(n5475) );
  NOR2_X1 U5124 ( .A1(n5471), .A2(n5470), .ZN(n4658) );
  OAI21_X2 U5125 ( .B1(n5408), .B2(n4605), .A(n4603), .ZN(n5450) );
  XNOR2_X1 U5126 ( .A(n5662), .B(n5661), .ZN(n5699) );
  AOI21_X1 U5127 ( .B1(n6830), .B2(n9676), .A(n6641), .ZN(n7119) );
  NOR2_X2 U5128 ( .A1(n6279), .A2(n6278), .ZN(n6496) );
  NAND2_X4 U5129 ( .A1(n6173), .A2(n6229), .ZN(n6279) );
  XNOR2_X1 U5130 ( .A(n5131), .B(n5130), .ZN(n6991) );
  NOR2_X1 U5131 ( .A1(n7358), .A2(n6640), .ZN(n6658) );
  OAI21_X2 U5132 ( .B1(n4509), .B2(n4506), .A(n4502), .ZN(n7943) );
  INV_X1 U5133 ( .A(n6830), .ZN(n6659) );
  BUF_X4 U5134 ( .A(n5090), .Z(n7002) );
  NAND2_X1 U5135 ( .A1(n4750), .A2(n4749), .ZN(n8635) );
  NAND2_X1 U5136 ( .A1(n7789), .A2(n8702), .ZN(n4750) );
  NAND2_X1 U5137 ( .A1(n8611), .A2(n8714), .ZN(n4749) );
  NAND2_X1 U5138 ( .A1(n5467), .A2(n8069), .ZN(n5487) );
  NOR2_X1 U5139 ( .A1(n5338), .A2(n4881), .ZN(n4880) );
  INV_X1 U5140 ( .A(n5317), .ZN(n4881) );
  OR2_X1 U5141 ( .A1(n10099), .A2(n9853), .ZN(n9804) );
  OR2_X1 U5142 ( .A1(n10154), .A2(n10016), .ZN(n8640) );
  OR2_X1 U5143 ( .A1(n10077), .A2(n8469), .ZN(n8704) );
  NAND2_X1 U5144 ( .A1(n4872), .A2(n4871), .ZN(n6244) );
  AOI21_X1 U5145 ( .B1(n4874), .B2(n4876), .A(n4474), .ZN(n4871) );
  NAND2_X1 U5146 ( .A1(n5639), .A2(n4874), .ZN(n4872) );
  NAND2_X1 U5147 ( .A1(n5799), .A2(n6986), .ZN(n5840) );
  INV_X1 U5148 ( .A(n7290), .ZN(n4723) );
  NAND2_X1 U5149 ( .A1(n6222), .A2(n4809), .ZN(n9387) );
  NAND2_X1 U5150 ( .A1(n9813), .A2(n5039), .ZN(n9775) );
  NOR2_X1 U5151 ( .A1(n5040), .A2(n10077), .ZN(n5039) );
  NAND2_X1 U5152 ( .A1(n10154), .A2(n10016), .ZN(n9975) );
  OAI21_X1 U5153 ( .B1(n8635), .B2(n8614), .A(n4747), .ZN(n8616) );
  NOR2_X1 U5154 ( .A1(n4748), .A2(n5011), .ZN(n4747) );
  NOR2_X1 U5155 ( .A1(n4853), .A2(n6399), .ZN(n4852) );
  INV_X1 U5156 ( .A(n9242), .ZN(n4853) );
  AND2_X1 U5157 ( .A1(n4591), .A2(n4598), .ZN(n4590) );
  NOR2_X1 U5158 ( .A1(n4423), .A2(n4599), .ZN(n4598) );
  NAND2_X1 U5159 ( .A1(n4594), .A2(n4592), .ZN(n4591) );
  INV_X1 U5160 ( .A(n5560), .ZN(n4599) );
  NOR2_X1 U5161 ( .A1(n4602), .A2(n4451), .ZN(n4601) );
  INV_X1 U5162 ( .A(n4866), .ZN(n4602) );
  INV_X1 U5163 ( .A(n4604), .ZN(n4603) );
  OAI21_X1 U5164 ( .B1(n5407), .B2(n4605), .A(n5425), .ZN(n4604) );
  INV_X1 U5165 ( .A(n4489), .ZN(n5259) );
  AOI21_X1 U5166 ( .B1(n4831), .B2(n4832), .A(n6458), .ZN(n4829) );
  AND2_X1 U5167 ( .A1(n9199), .A2(n6395), .ZN(n4805) );
  OR2_X1 U5168 ( .A1(n9432), .A2(n9247), .ZN(n6398) );
  INV_X1 U5169 ( .A(n5990), .ZN(n5763) );
  NAND2_X1 U5170 ( .A1(n4796), .A2(n6347), .ZN(n4798) );
  NAND2_X1 U5171 ( .A1(n6188), .A2(n4803), .ZN(n4796) );
  NAND2_X1 U5172 ( .A1(n6339), .A2(n6337), .ZN(n5930) );
  AOI21_X1 U5173 ( .B1(n6328), .B2(n4793), .A(n6330), .ZN(n4792) );
  INV_X1 U5174 ( .A(n6324), .ZN(n6328) );
  NAND2_X1 U5175 ( .A1(n7692), .A2(n6186), .ZN(n5021) );
  NAND2_X1 U5176 ( .A1(n6716), .A2(n6717), .ZN(n4508) );
  NAND2_X1 U5177 ( .A1(n9611), .A2(n9613), .ZN(n6833) );
  INV_X1 U5178 ( .A(n5666), .ZN(n5663) );
  OR2_X1 U5179 ( .A1(n10089), .A2(n9641), .ZN(n8694) );
  OR2_X1 U5180 ( .A1(n5616), .A2(n9818), .ZN(n4646) );
  NAND2_X1 U5181 ( .A1(n9519), .A2(n4568), .ZN(n8689) );
  AND2_X1 U5182 ( .A1(n9883), .A2(n9894), .ZN(n8544) );
  OR2_X1 U5183 ( .A1(n10149), .A2(n9653), .ZN(n8650) );
  AND2_X1 U5184 ( .A1(n5707), .A2(n4695), .ZN(n4694) );
  INV_X1 U5185 ( .A(n8627), .ZN(n4696) );
  NAND2_X1 U5186 ( .A1(n10159), .A2(n9656), .ZN(n8532) );
  INV_X1 U5187 ( .A(n5254), .ZN(n4977) );
  OR2_X1 U5188 ( .A1(n8399), .A2(n8270), .ZN(n8636) );
  AND2_X1 U5189 ( .A1(n5252), .A2(n7573), .ZN(n5253) );
  INV_X1 U5190 ( .A(n8521), .ZN(n4688) );
  INV_X1 U5191 ( .A(n8604), .ZN(n4687) );
  NOR2_X1 U5192 ( .A1(n4690), .A2(n8578), .ZN(n4689) );
  AND2_X1 U5193 ( .A1(n4392), .A2(n9857), .ZN(n6871) );
  OAI21_X1 U5194 ( .B1(n6244), .B2(n6243), .A(n6246), .ZN(n6264) );
  AND2_X1 U5195 ( .A1(n5640), .A2(n5625), .ZN(n5638) );
  NAND2_X1 U5196 ( .A1(n5620), .A2(n5619), .ZN(n5639) );
  NAND2_X1 U5197 ( .A1(n5280), .A2(n4914), .ZN(n4913) );
  NAND2_X1 U5198 ( .A1(n5487), .A2(n5469), .ZN(n5488) );
  AND2_X1 U5199 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  OR2_X1 U5200 ( .A1(n5476), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U5201 ( .A1(n5295), .A2(n5237), .ZN(n5255) );
  NAND2_X1 U5202 ( .A1(n4611), .A2(n5234), .ZN(n5256) );
  NAND4_X2 U5203 ( .A1(n4533), .A2(n10240), .A3(n5110), .A4(n5167), .ZN(n5190)
         );
  NOR2_X2 U5204 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4533) );
  INV_X1 U5205 ( .A(n7611), .ZN(n4952) );
  NAND2_X1 U5206 ( .A1(n7782), .A2(n4951), .ZN(n4950) );
  INV_X1 U5207 ( .A(n5061), .ZN(n4951) );
  OR3_X1 U5208 ( .A1(n8410), .A2(n9512), .A3(n8435), .ZN(n6903) );
  NAND2_X1 U5209 ( .A1(n4926), .A2(n4925), .ZN(n4924) );
  INV_X1 U5210 ( .A(n8791), .ZN(n4925) );
  INV_X1 U5211 ( .A(n8792), .ZN(n4926) );
  AND2_X1 U5212 ( .A1(n6173), .A2(n9154), .ZN(n6626) );
  OAI21_X1 U5213 ( .B1(n8991), .B2(n8990), .A(n8989), .ZN(n9005) );
  AND2_X1 U5214 ( .A1(n4718), .A2(n4466), .ZN(n4715) );
  INV_X1 U5215 ( .A(n4725), .ZN(n9080) );
  OR2_X1 U5216 ( .A1(n9400), .A2(n9165), .ZN(n6080) );
  NAND2_X1 U5217 ( .A1(n4822), .A2(n4449), .ZN(n4826) );
  NAND2_X1 U5218 ( .A1(n8371), .A2(n8367), .ZN(n4822) );
  OR2_X1 U5219 ( .A1(n9470), .A2(n8785), .ZN(n8309) );
  INV_X2 U5220 ( .A(n5841), .ZN(n6022) );
  OR2_X1 U5221 ( .A1(n6205), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5750) );
  OR2_X1 U5222 ( .A1(n9389), .A2(n8915), .ZN(n6097) );
  NAND2_X1 U5223 ( .A1(n6223), .A2(n6424), .ZN(n6241) );
  NAND2_X1 U5224 ( .A1(n6143), .A2(n6142), .ZN(n6625) );
  AND2_X1 U5225 ( .A1(n6903), .A2(n6148), .ZN(n10339) );
  AND2_X1 U5226 ( .A1(n5785), .A2(n5736), .ZN(n5739) );
  INV_X1 U5227 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6138) );
  NOR2_X1 U5228 ( .A1(n5872), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5874) );
  INV_X1 U5229 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4727) );
  XNOR2_X1 U5230 ( .A(n6700), .B(n6847), .ZN(n6702) );
  NAND2_X1 U5231 ( .A1(n6640), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n4556) );
  NAND2_X1 U5232 ( .A1(n9676), .A2(n4395), .ZN(n6644) );
  NAND2_X1 U5233 ( .A1(n5455), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5498) );
  AND2_X1 U5234 ( .A1(n9756), .A2(n9664), .ZN(n8720) );
  NAND2_X1 U5235 ( .A1(n4754), .A2(n8702), .ZN(n4753) );
  INV_X1 U5236 ( .A(n8715), .ZN(n4754) );
  INV_X1 U5237 ( .A(n5716), .ZN(n7001) );
  INV_X1 U5238 ( .A(n5156), .ZN(n5716) );
  INV_X1 U5239 ( .A(n5611), .ZN(n5090) );
  NAND2_X1 U5240 ( .A1(n8468), .A2(n8467), .ZN(n10077) );
  AND2_X1 U5241 ( .A1(n5001), .A2(n5000), .ZN(n9806) );
  INV_X1 U5242 ( .A(n8673), .ZN(n4563) );
  NAND2_X1 U5243 ( .A1(n4570), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U5244 ( .A1(n4663), .A2(n4662), .ZN(n9997) );
  AND2_X1 U5245 ( .A1(n5400), .A2(n5372), .ZN(n4662) );
  AND2_X1 U5246 ( .A1(n8640), .A2(n9975), .ZN(n9994) );
  INV_X1 U5247 ( .A(n5166), .ZN(n5218) );
  OAI21_X1 U5248 ( .B1(n5136), .B2(n8474), .A(n5135), .ZN(n7409) );
  INV_X1 U5249 ( .A(n10014), .ZN(n10041) );
  INV_X1 U5250 ( .A(n10045), .ZN(n4705) );
  MUX2_X1 U5251 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5079), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n4973) );
  XNOR2_X1 U5252 ( .A(n5639), .B(n5638), .ZN(n9504) );
  XNOR2_X1 U5253 ( .A(n5671), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U5254 ( .A1(n5672), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U5255 ( .A1(n5280), .A2(n4909), .ZN(n4908) );
  INV_X1 U5256 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4909) );
  XNOR2_X1 U5257 ( .A(n5256), .B(n5255), .ZN(n6999) );
  XNOR2_X1 U5258 ( .A(n5162), .B(SI_3_), .ZN(n5161) );
  NAND2_X1 U5259 ( .A1(n10240), .A2(n5110), .ZN(n5170) );
  INV_X1 U5260 ( .A(n9641), .ZN(n9807) );
  INV_X1 U5261 ( .A(n9656), .ZN(n10042) );
  NAND2_X1 U5262 ( .A1(n6307), .A2(n4583), .ZN(n4582) );
  NAND2_X1 U5263 ( .A1(n6442), .A2(n6435), .ZN(n4581) );
  INV_X1 U5264 ( .A(n6339), .ZN(n6332) );
  INV_X1 U5265 ( .A(n9292), .ZN(n4855) );
  NOR2_X1 U5266 ( .A1(n6369), .A2(n6370), .ZN(n4854) );
  NAND2_X1 U5267 ( .A1(n6406), .A2(n6407), .ZN(n4879) );
  OR2_X1 U5268 ( .A1(n8693), .A2(n8692), .ZN(n4762) );
  NAND2_X1 U5269 ( .A1(n8690), .A2(n8691), .ZN(n4765) );
  OR2_X1 U5270 ( .A1(n6429), .A2(n4893), .ZN(n4892) );
  AND2_X1 U5271 ( .A1(n6430), .A2(n4583), .ZN(n4893) );
  NAND2_X1 U5272 ( .A1(n8229), .A2(n7831), .ZN(n6339) );
  OR2_X1 U5273 ( .A1(n9756), .A2(n9664), .ZN(n8708) );
  NAND2_X1 U5274 ( .A1(n5530), .A2(n5529), .ZN(n5541) );
  INV_X1 U5275 ( .A(n5055), .ZN(n4605) );
  NAND2_X1 U5276 ( .A1(n5409), .A2(n8057), .ZN(n5425) );
  AOI21_X1 U5277 ( .B1(n5019), .B2(n6426), .A(n5018), .ZN(n5017) );
  INV_X1 U5278 ( .A(n5020), .ZN(n5019) );
  AOI21_X1 U5279 ( .B1(n4813), .B2(n9137), .A(n6425), .ZN(n4812) );
  OR2_X1 U5280 ( .A1(n6050), .A2(n5768), .ZN(n6058) );
  OR2_X1 U5281 ( .A1(n9425), .A2(n8774), .ZN(n6404) );
  NAND2_X1 U5282 ( .A1(n5766), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6050) );
  INV_X1 U5283 ( .A(n6041), .ZN(n5766) );
  OR2_X1 U5284 ( .A1(n6034), .A2(n8839), .ZN(n6041) );
  AND2_X1 U5285 ( .A1(n6404), .A2(n6401), .ZN(n9241) );
  NAND2_X1 U5286 ( .A1(n9343), .A2(n4484), .ZN(n4487) );
  NOR2_X1 U5287 ( .A1(n4837), .A2(n4485), .ZN(n4484) );
  NAND2_X1 U5288 ( .A1(n4408), .A2(n6005), .ZN(n4837) );
  INV_X1 U5289 ( .A(n5997), .ZN(n4485) );
  INV_X1 U5290 ( .A(n9442), .ZN(n4777) );
  AND2_X1 U5291 ( .A1(n9292), .A2(n9293), .ZN(n4840) );
  OR2_X1 U5292 ( .A1(n9442), .A2(n9313), .ZN(n9238) );
  NOR2_X1 U5293 ( .A1(n9445), .A2(n9450), .ZN(n4778) );
  OR2_X1 U5294 ( .A1(n5977), .A2(n5762), .ZN(n5990) );
  INV_X1 U5295 ( .A(n4827), .ZN(n4483) );
  NOR2_X1 U5296 ( .A1(n5948), .A2(n4826), .ZN(n4823) );
  NAND2_X1 U5297 ( .A1(n5760), .A2(n5759), .ZN(n5956) );
  INV_X1 U5298 ( .A(n5942), .ZN(n5760) );
  NAND2_X1 U5299 ( .A1(n4615), .A2(n4613), .ZN(n6337) );
  NOR2_X1 U5300 ( .A1(n4614), .A2(n7831), .ZN(n4613) );
  INV_X1 U5301 ( .A(n5922), .ZN(n4614) );
  OR2_X1 U5302 ( .A1(n10397), .A2(n7832), .ZN(n6322) );
  INV_X1 U5303 ( .A(n7679), .ZN(n6441) );
  INV_X1 U5304 ( .A(n5778), .ZN(n5022) );
  INV_X1 U5305 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6126) );
  AND2_X1 U5306 ( .A1(n8163), .A2(n5983), .ZN(n4938) );
  NOR2_X1 U5307 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5983) );
  NAND2_X1 U5308 ( .A1(n7840), .A2(n6715), .ZN(n4507) );
  INV_X1 U5309 ( .A(n6904), .ZN(n6640) );
  NAND2_X1 U5310 ( .A1(n4859), .A2(n4419), .ZN(n4858) );
  NAND2_X1 U5311 ( .A1(n4860), .A2(n6820), .ZN(n4859) );
  OR2_X1 U5312 ( .A1(n4861), .A2(n6802), .ZN(n4860) );
  NAND2_X1 U5313 ( .A1(n9538), .A2(n4442), .ZN(n4857) );
  AND2_X1 U5314 ( .A1(n9603), .A2(n6797), .ZN(n4514) );
  NAND2_X1 U5315 ( .A1(n9595), .A2(n6844), .ZN(n4887) );
  OR2_X1 U5316 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  INV_X1 U5317 ( .A(n6919), .ZN(n4670) );
  AND2_X1 U5318 ( .A1(n6876), .A2(n9786), .ZN(n9764) );
  INV_X1 U5319 ( .A(n9764), .ZN(n8699) );
  NAND2_X1 U5320 ( .A1(n10085), .A2(n9768), .ZN(n9765) );
  NOR2_X1 U5321 ( .A1(n8505), .A2(n4990), .ZN(n4989) );
  INV_X1 U5322 ( .A(n9930), .ZN(n4987) );
  OR2_X1 U5323 ( .A1(n10124), .A2(n9543), .ZN(n8671) );
  OR2_X1 U5324 ( .A1(n10144), .A2(n5044), .ZN(n5043) );
  OR2_X1 U5325 ( .A1(n10149), .A2(n10154), .ZN(n5044) );
  OR2_X1 U5326 ( .A1(n10164), .A2(n10015), .ZN(n8531) );
  OR2_X1 U5327 ( .A1(n8411), .A2(n7948), .ZN(n8527) );
  OR2_X1 U5328 ( .A1(n10170), .A2(n7909), .ZN(n8638) );
  NAND2_X1 U5329 ( .A1(n7134), .A2(n7424), .ZN(n8568) );
  NAND2_X1 U5330 ( .A1(n7258), .A2(n7173), .ZN(n8563) );
  NAND2_X1 U5331 ( .A1(n4588), .A2(n4587), .ZN(n5618) );
  AOI21_X1 U5332 ( .B1(n4590), .B2(n4593), .A(n4903), .ZN(n4587) );
  AND2_X1 U5333 ( .A1(n5619), .A2(n5604), .ZN(n5617) );
  NOR2_X1 U5334 ( .A1(n5542), .A2(n4597), .ZN(n4596) );
  INV_X1 U5335 ( .A(n5526), .ZN(n4597) );
  NAND2_X1 U5336 ( .A1(n4865), .A2(n4863), .ZN(n5508) );
  AOI21_X1 U5337 ( .B1(n4866), .B2(n4868), .A(n4864), .ZN(n4863) );
  INV_X1 U5338 ( .A(n5487), .ZN(n4864) );
  AND2_X1 U5339 ( .A1(n5509), .A2(n5492), .ZN(n5507) );
  INV_X1 U5340 ( .A(n5446), .ZN(n4870) );
  INV_X1 U5341 ( .A(SI_15_), .ZN(n5384) );
  AND2_X1 U5342 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  NAND2_X1 U5343 ( .A1(n5274), .A2(n5273), .ZN(n5300) );
  INV_X1 U5344 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U5345 ( .A1(n5217), .A2(n5216), .ZN(n4612) );
  NAND2_X1 U5346 ( .A1(n5165), .A2(n5164), .ZN(n5185) );
  NAND2_X1 U5347 ( .A1(n5757), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U5348 ( .A1(n4934), .A2(n4935), .ZN(n4933) );
  NAND2_X1 U5349 ( .A1(n4933), .A2(n4398), .ZN(n8804) );
  NAND2_X1 U5350 ( .A1(n7026), .A2(n6056), .ZN(n4615) );
  NOR2_X1 U5351 ( .A1(n4965), .A2(n8819), .ZN(n4957) );
  NAND2_X1 U5352 ( .A1(n4967), .A2(n4961), .ZN(n4960) );
  NOR2_X1 U5353 ( .A1(n4966), .A2(n4964), .ZN(n4961) );
  NAND2_X1 U5354 ( .A1(n4965), .A2(n4970), .ZN(n4959) );
  AND2_X1 U5355 ( .A1(n8757), .A2(n4963), .ZN(n4962) );
  AOI21_X1 U5356 ( .B1(n8879), .B2(n4964), .A(n4966), .ZN(n4963) );
  NOR2_X1 U5357 ( .A1(n4434), .A2(n4942), .ZN(n4941) );
  INV_X1 U5358 ( .A(n4944), .ZN(n4942) );
  AND2_X1 U5359 ( .A1(n8810), .A2(n6558), .ZN(n6559) );
  INV_X1 U5360 ( .A(n8879), .ZN(n4965) );
  NAND2_X1 U5361 ( .A1(n6573), .A2(n4968), .ZN(n4958) );
  NAND2_X1 U5362 ( .A1(n4950), .A2(n6533), .ZN(n4947) );
  OR2_X1 U5363 ( .A1(n6566), .A2(n6565), .ZN(n4421) );
  NAND2_X1 U5364 ( .A1(n4969), .A2(n4968), .ZN(n4967) );
  OR2_X1 U5365 ( .A1(n6626), .A2(n7206), .ZN(n6629) );
  NAND2_X1 U5366 ( .A1(n8792), .A2(n8791), .ZN(n4923) );
  AND2_X1 U5367 ( .A1(n10339), .A2(n6605), .ZN(n6623) );
  XNOR2_X1 U5368 ( .A(n9389), .B(n8915), .ZN(n6459) );
  INV_X1 U5369 ( .A(n7768), .ZN(n6466) );
  AOI21_X1 U5370 ( .B1(n8948), .B2(n7268), .A(n7267), .ZN(n7283) );
  AND2_X1 U5371 ( .A1(n4723), .A2(n7288), .ZN(n4717) );
  NAND2_X1 U5372 ( .A1(n4709), .A2(n9050), .ZN(n9053) );
  OR2_X1 U5373 ( .A1(n9068), .A2(n9083), .ZN(n4725) );
  AND2_X1 U5374 ( .A1(n6471), .A2(n6466), .ZN(n7029) );
  AOI21_X1 U5375 ( .B1(n4734), .B2(n9137), .A(n4453), .ZN(n4733) );
  NAND2_X1 U5376 ( .A1(n4815), .A2(n6418), .ZN(n9113) );
  INV_X1 U5377 ( .A(n6459), .ZN(n9120) );
  NOR2_X1 U5378 ( .A1(n9120), .A2(n4814), .ZN(n4813) );
  INV_X1 U5379 ( .A(n6418), .ZN(n4814) );
  INV_X1 U5380 ( .A(n8890), .ZN(n9139) );
  NAND2_X1 U5381 ( .A1(n4785), .A2(n9152), .ZN(n4784) );
  NAND2_X1 U5382 ( .A1(n9185), .A2(n9184), .ZN(n9183) );
  AND2_X1 U5383 ( .A1(n9180), .A2(n6388), .ZN(n4804) );
  AND2_X1 U5384 ( .A1(n6392), .A2(n6285), .ZN(n9180) );
  NAND2_X1 U5385 ( .A1(n9229), .A2(n4403), .ZN(n9212) );
  AND2_X1 U5386 ( .A1(n9274), .A2(n9270), .ZN(n9265) );
  INV_X1 U5387 ( .A(n9241), .ZN(n9230) );
  NAND2_X1 U5388 ( .A1(n4486), .A2(n4741), .ZN(n9229) );
  INV_X1 U5389 ( .A(n4742), .ZN(n4741) );
  NAND2_X1 U5390 ( .A1(n4405), .A2(n4487), .ZN(n4486) );
  OAI21_X1 U5391 ( .B1(n4743), .B2(n9255), .A(n9230), .ZN(n4742) );
  INV_X1 U5392 ( .A(n4487), .ZN(n4745) );
  NAND2_X1 U5393 ( .A1(n9291), .A2(n4840), .ZN(n9294) );
  NAND2_X1 U5394 ( .A1(n4797), .A2(n6350), .ZN(n4794) );
  OAI22_X1 U5395 ( .A1(n9365), .A2(n6453), .B1(n9334), .B2(n9455), .ZN(n9342)
         );
  NAND3_X1 U5396 ( .A1(n8371), .A2(n7821), .A3(n4522), .ZN(n4827) );
  AND2_X1 U5397 ( .A1(n5930), .A2(n5909), .ZN(n4522) );
  AND4_X1 U5398 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n8785)
         );
  NAND2_X1 U5399 ( .A1(n4493), .A2(n4438), .ZN(n7930) );
  NAND2_X1 U5400 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5861) );
  NOR2_X1 U5401 ( .A1(n5807), .A2(n7720), .ZN(n4776) );
  NAND2_X1 U5402 ( .A1(n10311), .A2(n10309), .ZN(n7707) );
  NAND2_X1 U5403 ( .A1(n9503), .A2(n7029), .ZN(n9312) );
  NAND2_X1 U5404 ( .A1(n6099), .A2(n6098), .ZN(n6617) );
  NAND2_X1 U5405 ( .A1(n6024), .A2(n6023), .ZN(n9432) );
  NAND2_X1 U5406 ( .A1(n9318), .A2(n10402), .ZN(n10393) );
  NAND2_X1 U5407 ( .A1(n6141), .A2(n6140), .ZN(n10338) );
  AND2_X1 U5408 ( .A1(n4429), .A2(n4736), .ZN(n4735) );
  INV_X1 U5409 ( .A(n5772), .ZN(n4736) );
  OR2_X1 U5410 ( .A1(n5936), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5949) );
  INV_X1 U5411 ( .A(n5852), .ZN(n5854) );
  INV_X1 U5412 ( .A(n6703), .ZN(n4555) );
  NAND2_X1 U5413 ( .A1(n5223), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5246) );
  INV_X1 U5414 ( .A(n5225), .ZN(n5223) );
  NAND2_X1 U5415 ( .A1(n8442), .A2(n6871), .ZN(n6639) );
  NAND2_X1 U5416 ( .A1(n4889), .A2(n4888), .ZN(n9592) );
  INV_X1 U5417 ( .A(n9595), .ZN(n4888) );
  INV_X1 U5418 ( .A(n9594), .ZN(n4889) );
  NAND2_X1 U5419 ( .A1(n6706), .A2(n6705), .ZN(n4531) );
  NAND2_X1 U5420 ( .A1(n4566), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5287) );
  INV_X1 U5421 ( .A(n5263), .ZN(n4566) );
  NAND2_X1 U5422 ( .A1(n5330), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5345) );
  INV_X1 U5423 ( .A(n5331), .ZN(n5330) );
  INV_X1 U5424 ( .A(n4569), .ZN(n5365) );
  OR2_X1 U5425 ( .A1(n5607), .A2(n9640), .ZN(n5629) );
  NAND2_X1 U5426 ( .A1(n5589), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5607) );
  INV_X1 U5427 ( .A(n5590), .ZN(n5589) );
  OR2_X1 U5428 ( .A1(n8717), .A2(n6871), .ZN(n6884) );
  NAND2_X1 U5429 ( .A1(n4660), .A2(n4661), .ZN(n5101) );
  AND2_X1 U5430 ( .A1(n5664), .A2(n4658), .ZN(n4661) );
  INV_X1 U5431 ( .A(n5101), .ZN(n4537) );
  NOR2_X1 U5432 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4536) );
  INV_X1 U5433 ( .A(n5190), .ZN(n4659) );
  AND2_X1 U5434 ( .A1(n5574), .A2(n5573), .ZN(n9562) );
  OR2_X1 U5435 ( .A1(n9859), .A2(n5631), .ZN(n5574) );
  AND4_X1 U5436 ( .A1(n5230), .A2(n5229), .A3(n5228), .A4(n5227), .ZN(n7649)
         );
  OR2_X1 U5437 ( .A1(n5631), .A2(n4571), .ZN(n5230) );
  AND2_X1 U5438 ( .A1(n5156), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5089) );
  AND2_X1 U5439 ( .A1(n7063), .A2(n6917), .ZN(n4671) );
  AND2_X1 U5440 ( .A1(n7197), .A2(n6926), .ZN(n7233) );
  NAND2_X1 U5441 ( .A1(n7233), .A2(n7234), .ZN(n7232) );
  NAND2_X1 U5442 ( .A1(n4667), .A2(n4666), .ZN(n7544) );
  INV_X1 U5443 ( .A(n7547), .ZN(n4666) );
  INV_X1 U5444 ( .A(n7546), .ZN(n4667) );
  NOR2_X1 U5445 ( .A1(n9727), .A2(n4678), .ZN(n9729) );
  AND2_X1 U5446 ( .A1(n9728), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4678) );
  NAND2_X1 U5447 ( .A1(n9813), .A2(n5038), .ZN(n9774) );
  INV_X1 U5448 ( .A(n5040), .ZN(n5038) );
  NAND2_X1 U5449 ( .A1(n9807), .A2(n10041), .ZN(n5722) );
  NAND2_X1 U5450 ( .A1(n8694), .A2(n8695), .ZN(n9798) );
  OAI21_X1 U5451 ( .B1(n8547), .B2(n4994), .A(n4998), .ZN(n4993) );
  INV_X1 U5452 ( .A(n5597), .ZN(n9842) );
  NAND2_X1 U5453 ( .A1(n4984), .A2(n5540), .ZN(n9871) );
  NAND2_X1 U5454 ( .A1(n4985), .A2(n4402), .ZN(n4984) );
  INV_X1 U5455 ( .A(n9885), .ZN(n4985) );
  INV_X1 U5456 ( .A(n9891), .ZN(n9889) );
  OR2_X1 U5457 ( .A1(n9949), .A2(n10133), .ZN(n9934) );
  AND2_X1 U5458 ( .A1(n5486), .A2(n5485), .ZN(n9909) );
  NAND2_X1 U5459 ( .A1(n9929), .A2(n9930), .ZN(n9928) );
  AOI21_X1 U5460 ( .B1(n9956), .B2(n4656), .A(n4452), .ZN(n4655) );
  INV_X1 U5461 ( .A(n5445), .ZN(n4656) );
  INV_X1 U5462 ( .A(n9956), .ZN(n4657) );
  AND2_X1 U5463 ( .A1(n8656), .A2(n8657), .ZN(n9930) );
  INV_X1 U5464 ( .A(n5007), .ZN(n5006) );
  OAI21_X1 U5465 ( .B1(n4424), .B2(n5008), .A(n8650), .ZN(n5007) );
  NAND2_X1 U5466 ( .A1(n4693), .A2(n4694), .ZN(n10011) );
  NAND3_X1 U5467 ( .A1(n4650), .A2(n4649), .A3(n5269), .ZN(n8284) );
  NAND2_X1 U5468 ( .A1(n4431), .A2(n4651), .ZN(n4649) );
  NAND2_X1 U5469 ( .A1(n8287), .A2(n8642), .ZN(n8291) );
  NAND2_X1 U5470 ( .A1(n5285), .A2(n5284), .ZN(n8399) );
  AND2_X1 U5471 ( .A1(n8615), .A2(n8613), .ZN(n8484) );
  NAND2_X1 U5472 ( .A1(n4978), .A2(n5253), .ZN(n7579) );
  NAND2_X1 U5473 ( .A1(n4409), .A2(n7591), .ZN(n4978) );
  AND4_X1 U5474 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n7849)
         );
  AND4_X1 U5475 ( .A1(n5211), .A2(n5210), .A3(n5209), .A4(n5208), .ZN(n7632)
         );
  NAND2_X1 U5476 ( .A1(n5704), .A2(n8482), .ZN(n7628) );
  OR2_X1 U5477 ( .A1(n4689), .A2(n4687), .ZN(n4682) );
  AOI21_X1 U5478 ( .B1(n4689), .B2(n4688), .A(n4687), .ZN(n4684) );
  INV_X1 U5479 ( .A(n4689), .ZN(n4685) );
  NAND2_X1 U5480 ( .A1(n7591), .A2(n4979), .ZN(n7594) );
  AND2_X1 U5481 ( .A1(n5194), .A2(n5193), .ZN(n6679) );
  AND2_X1 U5482 ( .A1(n8725), .A2(n6847), .ZN(n7252) );
  INV_X1 U5483 ( .A(n10017), .ZN(n10043) );
  AND2_X1 U5484 ( .A1(n10081), .A2(n10080), .ZN(n10082) );
  NOR2_X1 U5485 ( .A1(n10078), .A2(n10295), .ZN(n10079) );
  NAND2_X1 U5486 ( .A1(n8704), .A2(n8703), .ZN(n10076) );
  INV_X1 U5487 ( .A(n4392), .ZN(n5727) );
  INV_X1 U5488 ( .A(n10295), .ZN(n10180) );
  NAND2_X1 U5489 ( .A1(n6884), .A2(n6979), .ZN(n7245) );
  NAND2_X1 U5490 ( .A1(n5326), .A2(n10234), .ZN(n4526) );
  OAI22_X1 U5491 ( .A1(n6264), .A2(n6263), .B1(SI_30_), .B2(n6262), .ZN(n6267)
         );
  XNOR2_X1 U5492 ( .A(n6264), .B(n6247), .ZN(n8731) );
  NAND2_X1 U5493 ( .A1(n5673), .A2(n10215), .ZN(n4510) );
  XNOR2_X1 U5494 ( .A(n5272), .B(n5271), .ZN(n7019) );
  NAND2_X1 U5495 ( .A1(n4953), .A2(n4952), .ZN(n4949) );
  INV_X1 U5496 ( .A(n7610), .ZN(n4953) );
  INV_X1 U5497 ( .A(n4950), .ZN(n4948) );
  OR2_X1 U5498 ( .A1(n5841), .A2(n7010), .ZN(n5815) );
  OR2_X1 U5499 ( .A1(n5840), .A2(n7017), .ZN(n5816) );
  INV_X1 U5500 ( .A(n8902), .ZN(n8862) );
  NAND2_X1 U5501 ( .A1(n7024), .A2(n6056), .ZN(n5916) );
  INV_X1 U5502 ( .A(n8874), .ZN(n8906) );
  AND2_X1 U5503 ( .A1(n7312), .A2(n6610), .ZN(n8908) );
  NAND2_X1 U5504 ( .A1(n6079), .A2(n6078), .ZN(n9165) );
  OR2_X1 U5505 ( .A1(n9155), .A2(n6073), .ZN(n6079) );
  NAND2_X1 U5506 ( .A1(n4719), .A2(n4723), .ZN(n4718) );
  AOI21_X1 U5507 ( .B1(n7288), .B2(n9018), .A(n4722), .ZN(n4721) );
  INV_X1 U5508 ( .A(n7291), .ZN(n4722) );
  INV_X1 U5509 ( .A(n9097), .ZN(n9056) );
  OAI21_X1 U5510 ( .B1(n9091), .B2(n9094), .A(n4443), .ZN(n4714) );
  OAI22_X1 U5511 ( .A1(n9095), .A2(n9094), .B1(n9093), .B2(n9092), .ZN(n4712)
         );
  XNOR2_X1 U5512 ( .A(n4492), .B(n9377), .ZN(n4491) );
  NAND2_X1 U5513 ( .A1(n9387), .A2(n9385), .ZN(n4492) );
  AND2_X1 U5514 ( .A1(n6178), .A2(n6105), .ZN(n9105) );
  INV_X1 U5515 ( .A(n9300), .ZN(n9356) );
  AND2_X1 U5516 ( .A1(n10335), .A2(n10322), .ZN(n9196) );
  INV_X1 U5517 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n4819) );
  NAND2_X1 U5518 ( .A1(n6222), .A2(n4447), .ZN(n9384) );
  NOR2_X1 U5519 ( .A1(n10405), .A2(n9351), .ZN(n4817) );
  NAND2_X1 U5520 ( .A1(n4519), .A2(n10407), .ZN(n4518) );
  INV_X1 U5521 ( .A(n9383), .ZN(n4519) );
  AND2_X1 U5522 ( .A1(n5057), .A2(n4429), .ZN(n4791) );
  OR2_X1 U5523 ( .A1(n6019), .A2(n6127), .ZN(n6020) );
  NAND2_X1 U5524 ( .A1(n5627), .A2(n5626), .ZN(n10089) );
  NAND2_X1 U5525 ( .A1(n5326), .A2(n4698), .ZN(n5151) );
  NOR2_X1 U5526 ( .A1(n4393), .A2(n6985), .ZN(n4698) );
  OAI21_X1 U5527 ( .B1(n6896), .B2(n6895), .A(n6894), .ZN(n6897) );
  NAND2_X1 U5528 ( .A1(n6999), .A2(n8464), .ZN(n5243) );
  AND2_X1 U5529 ( .A1(n5443), .A2(n5442), .ZN(n9628) );
  AND3_X1 U5530 ( .A1(n5371), .A2(n5370), .A3(n5369), .ZN(n9656) );
  AND2_X1 U5531 ( .A1(n5520), .A2(n5519), .ZN(n9910) );
  INV_X1 U5532 ( .A(n7424), .ZN(n7258) );
  OAI22_X1 U5533 ( .A1(n8722), .A2(n5052), .B1(n8558), .B2(n4607), .ZN(n4606)
         );
  OR3_X1 U5534 ( .A1(n8720), .A2(n8718), .A3(n8717), .ZN(n5052) );
  INV_X1 U5535 ( .A(n9562), .ZN(n9864) );
  INV_X1 U5536 ( .A(n9628), .ZN(n9979) );
  INV_X1 U5537 ( .A(n7849), .ZN(n9670) );
  XNOR2_X1 U5538 ( .A(n7093), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n7090) );
  NAND2_X1 U5539 ( .A1(n4639), .A2(n4645), .ZN(n9820) );
  NAND2_X1 U5540 ( .A1(n9810), .A2(n9809), .ZN(n9811) );
  NAND2_X1 U5541 ( .A1(n9808), .A2(n10041), .ZN(n9809) );
  NAND2_X1 U5542 ( .A1(n4663), .A2(n5372), .ZN(n9995) );
  OR2_X1 U5543 ( .A1(n5326), .A2(n7093), .ZN(n5111) );
  NOR2_X1 U5544 ( .A1(n10464), .A2(n10463), .ZN(n10462) );
  INV_X1 U5545 ( .A(n8613), .ZN(n4748) );
  AND2_X1 U5546 ( .A1(n9975), .A2(n8714), .ZN(n8622) );
  AOI21_X1 U5547 ( .B1(n6344), .B2(n6343), .A(n6342), .ZN(n6351) );
  AOI21_X1 U5548 ( .B1(n4622), .B2(n4440), .A(n6382), .ZN(n6400) );
  NAND2_X1 U5549 ( .A1(n4553), .A2(n4552), .ZN(n8672) );
  NAND2_X1 U5550 ( .A1(n6310), .A2(n6287), .ZN(n6307) );
  NAND2_X1 U5551 ( .A1(n4635), .A2(n4877), .ZN(n4550) );
  NOR2_X1 U5552 ( .A1(n6411), .A2(n4878), .ZN(n4877) );
  AND2_X1 U5553 ( .A1(n6409), .A2(n4583), .ZN(n4878) );
  NOR2_X1 U5554 ( .A1(n4549), .A2(n6412), .ZN(n4548) );
  NAND2_X1 U5555 ( .A1(n4764), .A2(n4767), .ZN(n4763) );
  AND2_X1 U5556 ( .A1(n4762), .A2(n4760), .ZN(n4759) );
  OAI21_X1 U5557 ( .B1(n8680), .B2(n8714), .A(n4384), .ZN(n4761) );
  INV_X1 U5558 ( .A(n4596), .ZN(n4592) );
  NAND2_X1 U5559 ( .A1(n4488), .A2(n4490), .ZN(n4489) );
  NAND2_X1 U5560 ( .A1(n6986), .A2(n5257), .ZN(n4488) );
  OAI21_X1 U5561 ( .B1(n6461), .B2(n6426), .A(n6284), .ZN(n5020) );
  AND3_X1 U5562 ( .A1(n9259), .A2(n9238), .A3(n6398), .ZN(n6198) );
  INV_X1 U5563 ( .A(n7873), .ZN(n6187) );
  NAND2_X1 U5564 ( .A1(n7709), .A2(n6488), .ZN(n6302) );
  INV_X1 U5565 ( .A(SI_19_), .ZN(n8069) );
  INV_X1 U5566 ( .A(SI_16_), .ZN(n8057) );
  NOR2_X1 U5567 ( .A1(n9851), .A2(n5003), .ZN(n5002) );
  INV_X1 U5568 ( .A(n8595), .ZN(n5003) );
  INV_X1 U5569 ( .A(n5640), .ZN(n4876) );
  INV_X1 U5570 ( .A(n4875), .ZN(n4874) );
  OAI21_X1 U5571 ( .B1(n5638), .B2(n4876), .A(n6109), .ZN(n4875) );
  INV_X1 U5572 ( .A(n5582), .ZN(n4904) );
  INV_X1 U5573 ( .A(n4594), .ZN(n4593) );
  INV_X1 U5574 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5072) );
  NOR2_X1 U5575 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4914) );
  AOI21_X1 U5576 ( .B1(n4869), .B2(n4867), .A(n4461), .ZN(n4866) );
  NAND2_X1 U5577 ( .A1(n5490), .A2(n7963), .ZN(n5509) );
  NAND2_X1 U5578 ( .A1(n5339), .A2(SI_13_), .ZN(n5375) );
  NAND2_X1 U5579 ( .A1(n5320), .A2(n5319), .ZN(n5373) );
  NAND2_X1 U5580 ( .A1(n4427), .A2(n4627), .ZN(n5215) );
  AOI21_X1 U5581 ( .B1(n4398), .B2(n8845), .A(n4458), .ZN(n4932) );
  NOR2_X1 U5582 ( .A1(n8805), .A2(n6557), .ZN(n6553) );
  AOI21_X1 U5583 ( .B1(n4894), .B2(n4629), .A(n4892), .ZN(n4631) );
  NAND2_X1 U5584 ( .A1(n6428), .A2(n6426), .ZN(n4629) );
  NAND2_X1 U5585 ( .A1(n4634), .A2(n6428), .ZN(n4633) );
  INV_X1 U5586 ( .A(n4892), .ZN(n4634) );
  OR2_X1 U5587 ( .A1(n9378), .A2(n6617), .ZN(n4782) );
  INV_X1 U5588 ( .A(n6080), .ZN(n4734) );
  NOR2_X1 U5589 ( .A1(n9162), .A2(n4835), .ZN(n4833) );
  AND2_X1 U5590 ( .A1(n9404), .A2(n6066), .ZN(n6411) );
  NOR2_X1 U5591 ( .A1(n4786), .A2(n9192), .ZN(n4785) );
  NAND2_X1 U5592 ( .A1(n9172), .A2(n4787), .ZN(n4786) );
  OAI21_X1 U5593 ( .B1(n4840), .B2(n4839), .A(n6016), .ZN(n4838) );
  NOR2_X1 U5594 ( .A1(n9292), .A2(n6196), .ZN(n6197) );
  NOR2_X1 U5595 ( .A1(n4798), .A2(n6194), .ZN(n4797) );
  NOR2_X1 U5596 ( .A1(n8229), .A2(n9470), .ZN(n4773) );
  OR2_X1 U5597 ( .A1(n5901), .A2(n5758), .ZN(n5923) );
  NOR2_X1 U5598 ( .A1(n7826), .A2(n7915), .ZN(n7825) );
  AND2_X1 U5599 ( .A1(n7873), .A2(n7867), .ZN(n5892) );
  OR2_X1 U5600 ( .A1(n6168), .A2(n7768), .ZN(n6487) );
  NOR2_X1 U5601 ( .A1(n7724), .A2(n7701), .ZN(n7621) );
  OR2_X1 U5602 ( .A1(n7622), .A2(n7876), .ZN(n6318) );
  NAND2_X1 U5603 ( .A1(n7875), .A2(n6320), .ZN(n7830) );
  NAND3_X1 U5604 ( .A1(n6171), .A2(n4776), .A3(n4775), .ZN(n7724) );
  NOR2_X1 U5605 ( .A1(n7688), .A2(n7738), .ZN(n4775) );
  NAND2_X1 U5606 ( .A1(n5771), .A2(n4413), .ZN(n6208) );
  INV_X1 U5607 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6162) );
  OAI21_X1 U5608 ( .B1(n10282), .B2(n6873), .A(n6648), .ZN(n6649) );
  INV_X1 U5609 ( .A(n8244), .ZN(n4896) );
  INV_X1 U5610 ( .A(n6749), .ZN(n4899) );
  NOR2_X1 U5611 ( .A1(n5345), .A2(n5344), .ZN(n4569) );
  AND2_X1 U5612 ( .A1(n8708), .A2(n8504), .ZN(n8715) );
  INV_X1 U5613 ( .A(n7639), .ZN(n4571) );
  NAND2_X1 U5614 ( .A1(n6876), .A2(n9796), .ZN(n5040) );
  NOR2_X1 U5615 ( .A1(n4642), .A2(n4641), .ZN(n4640) );
  INV_X1 U5616 ( .A(n8689), .ZN(n4641) );
  INV_X1 U5617 ( .A(n4646), .ZN(n4642) );
  NAND2_X1 U5618 ( .A1(n5628), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5644) );
  INV_X1 U5619 ( .A(n5629), .ZN(n5628) );
  AOI21_X1 U5620 ( .B1(n5004), .B2(n8599), .A(n4999), .ZN(n4998) );
  INV_X1 U5621 ( .A(n8549), .ZN(n4999) );
  NAND2_X1 U5622 ( .A1(n5002), .A2(n8682), .ZN(n4994) );
  NOR2_X1 U5623 ( .A1(n8547), .A2(n4997), .ZN(n4996) );
  INV_X1 U5624 ( .A(n5002), .ZN(n4997) );
  INV_X1 U5625 ( .A(n5575), .ZN(n4981) );
  NOR2_X1 U5626 ( .A1(n5576), .A2(n4983), .ZN(n4982) );
  INV_X1 U5627 ( .A(n5540), .ZN(n4983) );
  OR2_X1 U5628 ( .A1(n10106), .A2(n9562), .ZN(n8597) );
  NAND2_X1 U5629 ( .A1(n5034), .A2(n9869), .ZN(n5033) );
  INV_X1 U5630 ( .A(n5036), .ZN(n5034) );
  NAND2_X1 U5631 ( .A1(n9883), .A2(n5037), .ZN(n5036) );
  INV_X1 U5632 ( .A(n10118), .ZN(n5037) );
  OR2_X1 U5633 ( .A1(n10118), .A2(n9910), .ZN(n8675) );
  NAND2_X1 U5634 ( .A1(n8321), .A2(n8627), .ZN(n5014) );
  NOR2_X1 U5635 ( .A1(n8399), .A2(n8411), .ZN(n5030) );
  INV_X1 U5636 ( .A(n5253), .ZN(n4651) );
  AND2_X1 U5637 ( .A1(n5024), .A2(n5027), .ZN(n7584) );
  NOR2_X1 U5638 ( .A1(n5025), .A2(n7452), .ZN(n5024) );
  NAND2_X1 U5639 ( .A1(n7597), .A2(n5026), .ZN(n5025) );
  NOR2_X1 U5640 ( .A1(n4688), .A2(n4687), .ZN(n4686) );
  NAND2_X1 U5641 ( .A1(n7454), .A2(n6679), .ZN(n5028) );
  INV_X1 U5642 ( .A(n5028), .ZN(n5027) );
  AND2_X1 U5643 ( .A1(n8479), .A2(n7590), .ZN(n4979) );
  INV_X1 U5644 ( .A(n8519), .ZN(n8574) );
  INV_X1 U5645 ( .A(n7408), .ZN(n8475) );
  NOR2_X1 U5646 ( .A1(n7368), .A2(n7179), .ZN(n7256) );
  NOR2_X1 U5647 ( .A1(n5578), .A2(n4907), .ZN(n4906) );
  INV_X1 U5648 ( .A(n5562), .ZN(n4907) );
  AOI21_X1 U5649 ( .B1(n4596), .B2(n5527), .A(n4595), .ZN(n4594) );
  INV_X1 U5650 ( .A(n5541), .ZN(n4595) );
  NAND2_X1 U5651 ( .A1(n5525), .A2(SI_21_), .ZN(n5526) );
  NAND2_X1 U5652 ( .A1(n5541), .A2(n5532), .ZN(n5542) );
  INV_X1 U5653 ( .A(n5523), .ZN(n5527) );
  OR2_X1 U5654 ( .A1(n5412), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5413) );
  AND2_X1 U5655 ( .A1(n5361), .A2(n5360), .ZN(n5390) );
  NOR2_X1 U5656 ( .A1(n5323), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5361) );
  AND2_X1 U5657 ( .A1(n5300), .A2(n5314), .ZN(n4883) );
  NAND2_X1 U5658 ( .A1(n4479), .A2(n5294), .ZN(n4478) );
  INV_X1 U5659 ( .A(n5271), .ZN(n4479) );
  AOI21_X1 U5660 ( .B1(n4619), .B2(n5255), .A(n4618), .ZN(n4617) );
  NOR2_X1 U5661 ( .A1(n4621), .A2(n4620), .ZN(n4619) );
  NOR2_X1 U5662 ( .A1(n4620), .A2(n4621), .ZN(n4618) );
  NAND2_X1 U5663 ( .A1(n5255), .A2(n5295), .ZN(n4616) );
  NAND2_X1 U5664 ( .A1(n4611), .A2(n4609), .ZN(n5297) );
  NOR2_X1 U5665 ( .A1(n5255), .A2(n4610), .ZN(n4609) );
  INV_X1 U5666 ( .A(n5234), .ZN(n4610) );
  XNOR2_X1 U5667 ( .A(n5215), .B(SI_6_), .ZN(n5212) );
  NAND2_X1 U5668 ( .A1(n4497), .A2(n5199), .ZN(n5213) );
  OAI21_X1 U5669 ( .B1(n5752), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n5141), .ZN(
        n5162) );
  NOR2_X2 U5670 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .ZN(
        n4821) );
  NAND2_X1 U5671 ( .A1(n5761), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5977) );
  INV_X1 U5672 ( .A(n5956), .ZN(n5761) );
  NAND2_X1 U5673 ( .A1(n8889), .A2(n6597), .ZN(n8734) );
  AND2_X1 U5674 ( .A1(n6600), .A2(n6599), .ZN(n6622) );
  INV_X1 U5675 ( .A(n6058), .ZN(n6057) );
  NOR2_X1 U5676 ( .A1(n4411), .A2(n6586), .ZN(n4940) );
  NOR2_X1 U5677 ( .A1(n4945), .A2(n6591), .ZN(n4944) );
  OR2_X1 U5678 ( .A1(n5923), .A2(n7784), .ZN(n5942) );
  AND2_X1 U5679 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5755) );
  OAI21_X1 U5680 ( .B1(n6257), .B2(n6256), .A(n6255), .ZN(n6258) );
  INV_X1 U5681 ( .A(n8447), .ZN(n6471) );
  INV_X1 U5682 ( .A(n6229), .ZN(n6485) );
  INV_X1 U5683 ( .A(n4386), .ZN(n6120) );
  AND3_X1 U5684 ( .A1(n6038), .A2(n6037), .A3(n6036), .ZN(n8774) );
  AND4_X1 U5685 ( .A1(n5947), .A2(n5946), .A3(n5945), .A4(n5944), .ZN(n6539)
         );
  AND4_X1 U5686 ( .A1(n5880), .A2(n5879), .A3(n5878), .A4(n5877), .ZN(n7832)
         );
  AND4_X1 U5687 ( .A1(n5821), .A2(n5822), .A3(n5820), .A4(n5819), .ZN(n7315)
         );
  OAI21_X1 U5688 ( .B1(n7283), .B2(n8959), .A(n7282), .ZN(n8976) );
  NAND2_X1 U5689 ( .A1(n4720), .A2(n7288), .ZN(n9021) );
  OR2_X1 U5690 ( .A1(n9023), .A2(n9018), .ZN(n4720) );
  AOI21_X1 U5691 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7378), .A(n7377), .ZN(
        n7379) );
  NOR2_X1 U5692 ( .A1(n7805), .A2(n8259), .ZN(n8254) );
  AND2_X1 U5693 ( .A1(n9133), .A2(n4779), .ZN(n9099) );
  NOR2_X1 U5694 ( .A1(n4782), .A2(n4780), .ZN(n4779) );
  NAND2_X1 U5695 ( .A1(n4781), .A2(n9127), .ZN(n4780) );
  NAND2_X1 U5696 ( .A1(n9130), .A2(n4813), .ZN(n4807) );
  INV_X1 U5697 ( .A(n4812), .ZN(n4811) );
  AOI21_X1 U5698 ( .B1(n4812), .B2(n4810), .A(n4809), .ZN(n4808) );
  INV_X1 U5699 ( .A(n4813), .ZN(n4810) );
  OR2_X1 U5700 ( .A1(n6083), .A2(n8049), .ZN(n6104) );
  OR2_X1 U5701 ( .A1(n9131), .A2(n6215), .ZN(n4541) );
  XNOR2_X1 U5702 ( .A(n9130), .B(n9137), .ZN(n4543) );
  AND2_X1 U5703 ( .A1(n6069), .A2(n6068), .ZN(n9152) );
  INV_X1 U5704 ( .A(n4833), .ZN(n4832) );
  NOR2_X1 U5705 ( .A1(n9214), .A2(n4783), .ZN(n9168) );
  INV_X1 U5706 ( .A(n4785), .ZN(n4783) );
  NOR3_X1 U5707 ( .A1(n9214), .A2(n9192), .A3(n9415), .ZN(n9187) );
  INV_X1 U5708 ( .A(n9199), .ZN(n9205) );
  NOR2_X1 U5709 ( .A1(n9214), .A2(n9415), .ZN(n9201) );
  AND2_X1 U5710 ( .A1(n6388), .A2(n6394), .ZN(n9199) );
  OR2_X1 U5711 ( .A1(n9232), .A2(n9420), .ZN(n9214) );
  CLKBUF_X1 U5712 ( .A(n9243), .Z(n9244) );
  OR2_X1 U5713 ( .A1(n6009), .A2(n5764), .ZN(n6026) );
  NAND2_X1 U5714 ( .A1(n5765), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6034) );
  INV_X1 U5715 ( .A(n6026), .ZN(n5765) );
  AND2_X1 U5716 ( .A1(n9355), .A2(n4465), .ZN(n9274) );
  NAND2_X1 U5717 ( .A1(n9355), .A2(n4410), .ZN(n9302) );
  NAND2_X1 U5718 ( .A1(n9310), .A2(n9315), .ZN(n9309) );
  AND4_X1 U5719 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n9313)
         );
  AND2_X1 U5720 ( .A1(n9355), .A2(n9341), .ZN(n9337) );
  NAND2_X1 U5721 ( .A1(n4482), .A2(n4481), .ZN(n9365) );
  NAND2_X1 U5722 ( .A1(n4731), .A2(n4824), .ZN(n4481) );
  INV_X1 U5723 ( .A(n4823), .ZN(n4731) );
  NAND2_X1 U5724 ( .A1(n4799), .A2(n4801), .ZN(n8381) );
  INV_X1 U5725 ( .A(n4798), .ZN(n4801) );
  NAND2_X1 U5726 ( .A1(n4800), .A2(n6188), .ZN(n4799) );
  INV_X1 U5727 ( .A(n5930), .ZN(n7924) );
  NAND2_X1 U5728 ( .A1(n7822), .A2(n5909), .ZN(n7925) );
  NAND2_X1 U5729 ( .A1(n4493), .A2(n4792), .ZN(n7927) );
  NAND2_X1 U5730 ( .A1(n7825), .A2(n6172), .ZN(n8375) );
  AND2_X1 U5731 ( .A1(n6328), .A2(n6329), .ZN(n7829) );
  CLKBUF_X1 U5732 ( .A(n7821), .Z(n7822) );
  NAND2_X1 U5733 ( .A1(n6322), .A2(n6320), .ZN(n7873) );
  NAND2_X1 U5734 ( .A1(n5021), .A2(n4406), .ZN(n7875) );
  AND2_X1 U5735 ( .A1(n7621), .A2(n7861), .ZN(n7882) );
  NOR2_X1 U5736 ( .A1(n7681), .A2(n6441), .ZN(n6182) );
  NAND2_X1 U5737 ( .A1(n6171), .A2(n10365), .ZN(n7741) );
  NAND2_X1 U5738 ( .A1(n7718), .A2(n5829), .ZN(n7750) );
  INV_X1 U5739 ( .A(n7707), .ZN(n4544) );
  NAND2_X1 U5740 ( .A1(n6625), .A2(n6166), .ZN(n7657) );
  NOR2_X1 U5741 ( .A1(n10402), .A2(n6466), .ZN(n6607) );
  AND2_X1 U5742 ( .A1(n9377), .A2(n10393), .ZN(n4730) );
  NAND2_X1 U5743 ( .A1(n6082), .A2(n6081), .ZN(n9394) );
  INV_X1 U5744 ( .A(n10393), .ZN(n9475) );
  INV_X1 U5745 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5749) );
  AND4_X1 U5746 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n6128)
         );
  AND2_X1 U5747 ( .A1(n4938), .A2(n6125), .ZN(n4937) );
  NAND2_X1 U5748 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  INV_X1 U5749 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4915) );
  NAND2_X1 U5750 ( .A1(n4524), .A2(n4523), .ZN(n5852) );
  NOR2_X1 U5751 ( .A1(n6750), .A2(n4902), .ZN(n4901) );
  INV_X1 U5752 ( .A(n6742), .ZN(n4902) );
  XNOR2_X1 U5753 ( .A(n4557), .B(n6847), .ZN(n8423) );
  NAND2_X1 U5754 ( .A1(n4585), .A2(n4584), .ZN(n9584) );
  OR2_X1 U5755 ( .A1(n9568), .A2(n6781), .ZN(n4585) );
  OAI22_X1 U5756 ( .A1(n7445), .A2(n6875), .B1(n10286), .B2(n6873), .ZN(n6662)
         );
  NAND2_X1 U5757 ( .A1(n6712), .A2(n6711), .ZN(n6713) );
  INV_X1 U5758 ( .A(n5246), .ZN(n5244) );
  NAND2_X1 U5759 ( .A1(n8245), .A2(n8244), .ZN(n4516) );
  INV_X1 U5760 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5344) );
  INV_X1 U5761 ( .A(n6825), .ZN(n4856) );
  NAND2_X1 U5762 ( .A1(n6826), .A2(n6825), .ZN(n9613) );
  INV_X1 U5763 ( .A(n5308), .ZN(n5306) );
  XNOR2_X1 U5764 ( .A(n4558), .B(n6847), .ZN(n6683) );
  NAND2_X1 U5765 ( .A1(n7553), .A2(n6863), .ZN(n4559) );
  AOI21_X1 U5766 ( .B1(n4886), .B2(n4885), .A(n4450), .ZN(n4884) );
  INV_X1 U5767 ( .A(n6844), .ZN(n4885) );
  OAI211_X1 U5768 ( .C1(n8245), .C2(n4897), .A(n4898), .B(n4895), .ZN(n9570)
         );
  NOR2_X1 U5769 ( .A1(n4899), .A2(n6768), .ZN(n4898) );
  NAND2_X1 U5770 ( .A1(n4901), .A2(n4896), .ZN(n4895) );
  INV_X1 U5771 ( .A(n4901), .ZN(n4897) );
  OR2_X1 U5772 ( .A1(n6888), .A2(n10213), .ZN(n6882) );
  NAND2_X1 U5773 ( .A1(n4569), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U5774 ( .A1(n8559), .A2(n8716), .ZN(n4608) );
  NAND2_X1 U5775 ( .A1(n5656), .A2(n5654), .ZN(n5658) );
  AND2_X1 U5776 ( .A1(n5504), .A2(n5503), .ZN(n9543) );
  AND4_X1 U5777 ( .A1(n5336), .A2(n5335), .A3(n5334), .A4(n5333), .ZN(n7909)
         );
  AND4_X1 U5778 ( .A1(n5313), .A2(n5312), .A3(n5311), .A4(n5310), .ZN(n7948)
         );
  AND4_X1 U5779 ( .A1(n5292), .A2(n5291), .A3(n5290), .A4(n5289), .ZN(n8270)
         );
  AND4_X1 U5780 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n7946)
         );
  OR2_X1 U5781 ( .A1(n5174), .A2(n5115), .ZN(n5118) );
  NAND2_X1 U5782 ( .A1(n5090), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5117) );
  OR2_X1 U5783 ( .A1(n9678), .A2(n9677), .ZN(n9680) );
  NAND2_X1 U5784 ( .A1(n4576), .A2(n4575), .ZN(n7070) );
  INV_X1 U5785 ( .A(n7073), .ZN(n4575) );
  INV_X1 U5786 ( .A(n7072), .ZN(n4576) );
  OAI21_X1 U5787 ( .B1(n7079), .B2(n4670), .A(n4668), .ZN(n6922) );
  AND2_X1 U5788 ( .A1(n4669), .A2(n7037), .ZN(n4668) );
  OR2_X1 U5789 ( .A1(n7164), .A2(n7165), .ZN(n7162) );
  NAND2_X1 U5790 ( .A1(n4578), .A2(n4577), .ZN(n7157) );
  INV_X1 U5791 ( .A(n7160), .ZN(n4577) );
  INV_X1 U5792 ( .A(n7159), .ZN(n4578) );
  NAND2_X1 U5793 ( .A1(n7232), .A2(n6928), .ZN(n7546) );
  NAND2_X1 U5794 ( .A1(n7544), .A2(n6930), .ZN(n7669) );
  AND2_X1 U5795 ( .A1(n7894), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7895) );
  NAND2_X1 U5796 ( .A1(n4675), .A2(n4432), .ZN(n4674) );
  NAND2_X1 U5797 ( .A1(n7771), .A2(n7772), .ZN(n4675) );
  NOR2_X1 U5798 ( .A1(n9729), .A2(n9730), .ZN(n9738) );
  XNOR2_X1 U5799 ( .A(n4579), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U5800 ( .A1(n9736), .A2(n4580), .ZN(n4579) );
  OR2_X1 U5801 ( .A1(n9739), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4580) );
  XNOR2_X1 U5802 ( .A(n4676), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9747) );
  OR2_X1 U5803 ( .A1(n9738), .A2(n4677), .ZN(n4676) );
  AND2_X1 U5804 ( .A1(n9739), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4677) );
  INV_X1 U5805 ( .A(n10073), .ZN(n10072) );
  NAND2_X1 U5806 ( .A1(n9813), .A2(n9796), .ZN(n9790) );
  NAND2_X1 U5807 ( .A1(n4646), .A2(n4422), .ZN(n4645) );
  NAND2_X1 U5808 ( .A1(n9807), .A2(n10043), .ZN(n9810) );
  NAND2_X1 U5809 ( .A1(n4638), .A2(n4980), .ZN(n9816) );
  NOR2_X2 U5810 ( .A1(n5032), .A2(n9917), .ZN(n9855) );
  OR2_X1 U5811 ( .A1(n10106), .A2(n5033), .ZN(n5032) );
  INV_X1 U5812 ( .A(n5567), .ZN(n5566) );
  AND2_X1 U5813 ( .A1(n5559), .A2(n5558), .ZN(n9852) );
  NAND2_X1 U5814 ( .A1(n5001), .A2(n4707), .ZN(n4706) );
  NAND2_X1 U5815 ( .A1(n9850), .A2(n9851), .ZN(n4707) );
  NAND2_X1 U5816 ( .A1(n5005), .A2(n8595), .ZN(n9850) );
  NOR2_X1 U5817 ( .A1(n9917), .A2(n5033), .ZN(n9866) );
  OR2_X1 U5818 ( .A1(n8544), .A2(n8471), .ZN(n9884) );
  INV_X1 U5819 ( .A(n4570), .ZN(n5514) );
  AOI21_X1 U5820 ( .B1(n4989), .B2(n4987), .A(n5710), .ZN(n4986) );
  INV_X1 U5821 ( .A(n4989), .ZN(n4988) );
  AND2_X1 U5822 ( .A1(n8675), .A2(n8673), .ZN(n9891) );
  NAND2_X1 U5823 ( .A1(n4653), .A2(n4652), .ZN(n9915) );
  AOI21_X1 U5824 ( .B1(n4407), .B2(n4657), .A(n4455), .ZN(n4652) );
  INV_X1 U5825 ( .A(n5043), .ZN(n5041) );
  NOR2_X1 U5826 ( .A1(n5043), .A2(n10020), .ZN(n9964) );
  AND2_X1 U5827 ( .A1(n9943), .A2(n9945), .ZN(n9969) );
  NOR2_X1 U5828 ( .A1(n10020), .A2(n5044), .ZN(n9981) );
  NOR2_X1 U5829 ( .A1(n4454), .A2(n4665), .ZN(n4664) );
  INV_X1 U5830 ( .A(n5353), .ZN(n4665) );
  AND4_X1 U5831 ( .A1(n5350), .A2(n5349), .A3(n5348), .A4(n5347), .ZN(n10015)
         );
  AND3_X1 U5832 ( .A1(n5399), .A2(n5398), .A3(n5397), .ZN(n10016) );
  NAND2_X1 U5833 ( .A1(n5014), .A2(n5012), .ZN(n10036) );
  NAND2_X1 U5834 ( .A1(n5014), .A2(n8638), .ZN(n10038) );
  INV_X1 U5835 ( .A(n8489), .ZN(n8325) );
  AND2_X1 U5836 ( .A1(n8638), .A2(n8618), .ZN(n8489) );
  NAND2_X1 U5837 ( .A1(n7796), .A2(n5030), .ZN(n5060) );
  NAND2_X1 U5838 ( .A1(n7796), .A2(n8286), .ZN(n8285) );
  NOR2_X1 U5839 ( .A1(n5011), .A2(n5010), .ZN(n5009) );
  INV_X1 U5840 ( .A(n8607), .ZN(n5010) );
  NAND2_X1 U5841 ( .A1(n7584), .A2(n5726), .ZN(n7797) );
  INV_X1 U5842 ( .A(n7584), .ZN(n7637) );
  NOR2_X1 U5843 ( .A1(n5028), .A2(n7452), .ZN(n7596) );
  NAND2_X1 U5844 ( .A1(n5027), .A2(n5023), .ZN(n7636) );
  NOR2_X1 U5845 ( .A1(n7452), .A2(n7758), .ZN(n5023) );
  NAND2_X1 U5846 ( .A1(n4691), .A2(n8575), .ZN(n8605) );
  NAND2_X1 U5847 ( .A1(n7511), .A2(n8521), .ZN(n4691) );
  NOR2_X1 U5848 ( .A1(n7452), .A2(n7466), .ZN(n7514) );
  NAND2_X1 U5849 ( .A1(n8513), .A2(n8518), .ZN(n7408) );
  CLKBUF_X1 U5850 ( .A(n7248), .Z(n8473) );
  OR2_X1 U5851 ( .A1(n7245), .A2(n5697), .ZN(n5729) );
  INV_X1 U5852 ( .A(n6650), .ZN(n7051) );
  NOR2_X1 U5853 ( .A1(n10071), .A2(n4975), .ZN(n4974) );
  NAND2_X1 U5854 ( .A1(n10075), .A2(n4976), .ZN(n4975) );
  AND2_X1 U5855 ( .A1(n10106), .A2(n10180), .ZN(n4701) );
  AND2_X1 U5856 ( .A1(n4435), .A2(n5077), .ZN(n4756) );
  INV_X1 U5857 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5077) );
  XNOR2_X1 U5858 ( .A(n6244), .B(n6114), .ZN(n8465) );
  XNOR2_X1 U5859 ( .A(n6110), .B(n6109), .ZN(n9501) );
  NAND2_X1 U5860 ( .A1(n4873), .A2(n5640), .ZN(n6110) );
  AND2_X1 U5861 ( .A1(n5562), .A2(n5548), .ZN(n5560) );
  XNOR2_X1 U5862 ( .A(n5489), .B(n5488), .ZN(n7402) );
  AOI21_X1 U5863 ( .B1(n4869), .B2(n4867), .A(n4446), .ZN(n4862) );
  OAI21_X1 U5864 ( .B1(n5450), .B2(n4870), .A(n5449), .ZN(n5465) );
  AND2_X1 U5865 ( .A1(n5451), .A2(n5431), .ZN(n9728) );
  XNOR2_X1 U5866 ( .A(n5318), .B(n5314), .ZN(n7024) );
  AND2_X1 U5867 ( .A1(n5283), .A2(n5323), .ZN(n6950) );
  XNOR2_X1 U5868 ( .A(n4476), .B(n5054), .ZN(n7026) );
  OAI21_X1 U5869 ( .B1(n4480), .B2(n5256), .A(n4477), .ZN(n4476) );
  NAND2_X1 U5870 ( .A1(n5271), .A2(n4616), .ZN(n4480) );
  NAND2_X1 U5871 ( .A1(n4617), .A2(n4478), .ZN(n4477) );
  AND2_X1 U5872 ( .A1(n5192), .A2(n5191), .ZN(n9697) );
  AND2_X1 U5873 ( .A1(n7532), .A2(n6515), .ZN(n7503) );
  NAND2_X1 U5874 ( .A1(n6090), .A2(n6089), .ZN(n9389) );
  AND2_X1 U5875 ( .A1(n4933), .A2(n4430), .ZN(n8740) );
  OR2_X1 U5876 ( .A1(n5841), .A2(n7009), .ZN(n5805) );
  AND4_X1 U5877 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n7731)
         );
  OR2_X1 U5878 ( .A1(n6628), .A2(n6627), .ZN(n8797) );
  NAND2_X1 U5879 ( .A1(n4956), .A2(n4962), .ZN(n8756) );
  NAND2_X1 U5880 ( .A1(n4960), .A2(n4959), .ZN(n8758) );
  NAND2_X1 U5881 ( .A1(n4969), .A2(n4957), .ZN(n4956) );
  NAND2_X1 U5882 ( .A1(n8734), .A2(n8735), .ZN(n8733) );
  AOI21_X1 U5883 ( .B1(n4930), .B2(n7535), .A(n4929), .ZN(n4927) );
  INV_X1 U5884 ( .A(n6521), .ZN(n4929) );
  NAND2_X1 U5885 ( .A1(n6999), .A2(n6056), .ZN(n4841) );
  AND4_X1 U5886 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n9311)
         );
  OR2_X1 U5887 ( .A1(n6507), .A2(n6506), .ZN(n6508) );
  AND4_X1 U5888 ( .A1(n5929), .A2(n5928), .A3(n5927), .A4(n5926), .ZN(n7831)
         );
  INV_X1 U5889 ( .A(n7828), .ZN(n7915) );
  AND3_X1 U5890 ( .A1(n6046), .A2(n6045), .A3(n6044), .ZN(n9248) );
  NAND2_X1 U5891 ( .A1(n4554), .A2(n6573), .ZN(n4955) );
  NAND2_X1 U5892 ( .A1(n6033), .A2(n6032), .ZN(n9425) );
  NOR2_X1 U5893 ( .A1(n8797), .A2(n9312), .ZN(n8874) );
  AND4_X1 U5894 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n9247)
         );
  NAND2_X1 U5895 ( .A1(n4967), .A2(n4421), .ZN(n8880) );
  NAND2_X1 U5896 ( .A1(n4922), .A2(n4920), .ZN(n8889) );
  NOR2_X1 U5897 ( .A1(n8885), .A2(n4921), .ZN(n4920) );
  INV_X1 U5898 ( .A(n4923), .ZN(n4921) );
  NAND2_X1 U5899 ( .A1(n4922), .A2(n4923), .ZN(n8886) );
  AND4_X1 U5900 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n9290)
         );
  INV_X1 U5901 ( .A(n8888), .ZN(n8910) );
  NOR2_X1 U5902 ( .A1(n6439), .A2(n6168), .ZN(n6474) );
  AND2_X1 U5903 ( .A1(n6437), .A2(n4583), .ZN(n4890) );
  INV_X1 U5904 ( .A(P2_U3966), .ZN(n8917) );
  AND2_X1 U5905 ( .A1(n4716), .A2(n4715), .ZN(n9035) );
  OR2_X1 U5906 ( .A1(n7326), .A2(n7327), .ZN(n7373) );
  AND2_X1 U5907 ( .A1(n5965), .A2(n5972), .ZN(n7812) );
  NAND2_X1 U5908 ( .A1(n4725), .A2(n4724), .ZN(n9069) );
  NAND2_X1 U5909 ( .A1(n9068), .A2(n9083), .ZN(n4724) );
  NOR2_X1 U5910 ( .A1(n9069), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U5911 ( .A1(n6270), .A2(n6269), .ZN(n9369) );
  INV_X1 U5912 ( .A(n9389), .ZN(n9127) );
  NAND2_X1 U5913 ( .A1(n4815), .A2(n4813), .ZN(n9117) );
  NAND2_X1 U5914 ( .A1(n4542), .A2(n4539), .ZN(n9135) );
  INV_X1 U5915 ( .A(n4540), .ZN(n4539) );
  NAND2_X1 U5916 ( .A1(n4543), .A2(n10313), .ZN(n4542) );
  OAI21_X1 U5917 ( .B1(n9132), .B2(n9312), .A(n4541), .ZN(n4540) );
  NAND2_X1 U5918 ( .A1(n9138), .A2(n9137), .ZN(n9136) );
  NAND2_X1 U5919 ( .A1(n9150), .A2(n6080), .ZN(n9138) );
  INV_X1 U5920 ( .A(n9152), .ZN(n9400) );
  NAND2_X1 U5921 ( .A1(n9183), .A2(n4834), .ZN(n9174) );
  AND2_X1 U5922 ( .A1(n4806), .A2(n6388), .ZN(n9179) );
  NAND2_X1 U5923 ( .A1(n4740), .A2(n4739), .ZN(n9231) );
  AOI21_X1 U5924 ( .B1(n4744), .B2(n9255), .A(n4743), .ZN(n4739) );
  NAND2_X1 U5925 ( .A1(n4745), .A2(n9255), .ZN(n4740) );
  NAND2_X1 U5926 ( .A1(n9256), .A2(n9255), .ZN(n9254) );
  OR2_X1 U5927 ( .A1(n4744), .A2(n4745), .ZN(n9256) );
  NAND2_X1 U5928 ( .A1(n9294), .A2(n6005), .ZN(n9273) );
  NAND2_X1 U5929 ( .A1(n4825), .A2(n4472), .ZN(n8383) );
  INV_X1 U5930 ( .A(n4826), .ZN(n4828) );
  NAND2_X1 U5931 ( .A1(n6345), .A2(n8372), .ZN(n8310) );
  AND2_X1 U5932 ( .A1(n6171), .A2(n4776), .ZN(n7683) );
  OR2_X1 U5933 ( .A1(n5841), .A2(n6990), .ZN(n5787) );
  AND2_X1 U5934 ( .A1(n10335), .A2(n6176), .ZN(n9300) );
  INV_X1 U5935 ( .A(n9359), .ZN(n10330) );
  NAND2_X1 U5936 ( .A1(n10339), .A2(n6607), .ZN(n9359) );
  NAND2_X1 U5937 ( .A1(n6233), .A2(n6232), .ZN(n6480) );
  AND2_X1 U5938 ( .A1(n9112), .A2(n6231), .ZN(n6232) );
  NAND2_X1 U5939 ( .A1(n4738), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5770) );
  XNOR2_X1 U5940 ( .A(n6139), .B(n6138), .ZN(n9512) );
  INV_X1 U5941 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8408) );
  XNOR2_X1 U5942 ( .A(n6132), .B(n6131), .ZN(n8410) );
  NAND2_X1 U5943 ( .A1(n6147), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6132) );
  INV_X1 U5944 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8449) );
  BUF_X1 U5945 ( .A(n6202), .Z(n8447) );
  INV_X1 U5946 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7770) );
  INV_X1 U5947 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7607) );
  INV_X1 U5948 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7403) );
  INV_X1 U5949 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7243) );
  INV_X1 U5950 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n8191) );
  INV_X1 U5951 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n8140) );
  INV_X1 U5952 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7059) );
  XNOR2_X1 U5953 ( .A(n5914), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9042) );
  INV_X1 U5954 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7034) );
  XNOR2_X1 U5955 ( .A(n5910), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9029) );
  INV_X1 U5956 ( .A(n5874), .ZN(n5888) );
  NAND2_X1 U5957 ( .A1(n9497), .A2(n4727), .ZN(n4726) );
  XNOR2_X1 U5958 ( .A(n6866), .B(n6690), .ZN(n9515) );
  AOI21_X1 U5959 ( .B1(n10089), .B2(n6868), .A(n6867), .ZN(n9514) );
  NAND2_X1 U5960 ( .A1(n7561), .A2(n7562), .ZN(n4849) );
  NAND2_X1 U5961 ( .A1(n9602), .A2(n9603), .ZN(n9550) );
  NAND2_X1 U5962 ( .A1(n9592), .A2(n6844), .ZN(n9559) );
  AND2_X1 U5963 ( .A1(n5463), .A2(n5462), .ZN(n9588) );
  AND2_X1 U5964 ( .A1(n5457), .A2(n5437), .ZN(n9966) );
  NAND2_X1 U5965 ( .A1(n6837), .A2(n9526), .ZN(n9594) );
  NAND2_X1 U5966 ( .A1(n7019), .A2(n8464), .ZN(n4532) );
  NAND2_X1 U5967 ( .A1(n6803), .A2(n6802), .ZN(n9602) );
  NAND2_X1 U5968 ( .A1(n9538), .A2(n6797), .ZN(n6803) );
  INV_X1 U5969 ( .A(n9657), .ZN(n9604) );
  XNOR2_X1 U5970 ( .A(n6696), .B(n6694), .ZN(n7459) );
  INV_X1 U5971 ( .A(n9654), .ZN(n9632) );
  OR2_X1 U5972 ( .A1(n9836), .A2(n5631), .ZN(n5596) );
  AND2_X1 U5973 ( .A1(n5629), .A2(n5608), .ZN(n9814) );
  AND3_X1 U5974 ( .A1(n5422), .A2(n5421), .A3(n5420), .ZN(n9653) );
  AND2_X1 U5975 ( .A1(n9570), .A2(n9569), .ZN(n9651) );
  NAND2_X1 U5976 ( .A1(n6889), .A2(n7133), .ZN(n9660) );
  AND2_X1 U5977 ( .A1(n8722), .A2(n8721), .ZN(n4755) );
  NAND2_X1 U5978 ( .A1(n4538), .A2(n4535), .ZN(n8724) );
  NOR2_X1 U5979 ( .A1(n4758), .A2(n10215), .ZN(n4525) );
  INV_X1 U5980 ( .A(n9853), .ZN(n9808) );
  NAND2_X1 U5981 ( .A1(n5539), .A2(n5538), .ZN(n9894) );
  INV_X1 U5982 ( .A(n9910), .ZN(n9876) );
  INV_X1 U5983 ( .A(n9543), .ZN(n9931) );
  INV_X1 U5984 ( .A(n9909), .ZN(n9947) );
  INV_X1 U5985 ( .A(n9588), .ZN(n9962) );
  INV_X1 U5986 ( .A(n10016), .ZN(n9978) );
  INV_X1 U5987 ( .A(n7909), .ZN(n10040) );
  INV_X1 U5988 ( .A(n7948), .ZN(n9667) );
  INV_X1 U5989 ( .A(n7946), .ZN(n9669) );
  OR2_X1 U5990 ( .A1(n5159), .A2(n5158), .ZN(n9674) );
  OAI22_X1 U5991 ( .A1(n5154), .A2(n6642), .B1(n5174), .B2(n8211), .ZN(n5088)
         );
  OR2_X1 U5992 ( .A1(n7077), .A2(n7076), .ZN(n7079) );
  NAND2_X1 U5993 ( .A1(n7079), .A2(n4671), .ZN(n7062) );
  NAND2_X1 U5994 ( .A1(n7062), .A2(n6919), .ZN(n7036) );
  XNOR2_X1 U5995 ( .A(n4674), .B(n7154), .ZN(n7893) );
  AND2_X1 U5996 ( .A1(n7893), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7902) );
  NOR2_X1 U5997 ( .A1(n7902), .A2(n4672), .ZN(n6935) );
  NOR2_X1 U5998 ( .A1(n4674), .A2(n4673), .ZN(n4672) );
  AOI21_X1 U5999 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9711), .A(n9710), .ZN(
        n9713) );
  OR2_X1 U6000 ( .A1(n6972), .A2(n10226), .ZN(n9741) );
  NAND2_X1 U6001 ( .A1(n8455), .A2(n5326), .ZN(n9756) );
  MUX2_X1 U6002 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9495), .S(n4394), .Z(n8455) );
  NAND2_X1 U6003 ( .A1(n8462), .A2(n8461), .ZN(n10067) );
  NAND2_X1 U6004 ( .A1(n9776), .A2(n9775), .ZN(n10081) );
  INV_X1 U6005 ( .A(n10076), .ZN(n10071) );
  AOI21_X1 U6006 ( .B1(n9786), .B2(n10041), .A(n9771), .ZN(n9772) );
  NOR2_X1 U6007 ( .A1(n9770), .A2(n9769), .ZN(n9771) );
  AOI21_X1 U6008 ( .B1(n5725), .B2(n4705), .A(n5724), .ZN(n10087) );
  NAND2_X1 U6009 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  NAND2_X1 U6010 ( .A1(n9665), .A2(n10043), .ZN(n5723) );
  AOI21_X1 U6011 ( .B1(n9789), .B2(n4705), .A(n9788), .ZN(n10092) );
  INV_X1 U6012 ( .A(n9830), .ZN(n9831) );
  XNOR2_X1 U6013 ( .A(n5048), .B(n9842), .ZN(n9832) );
  AOI22_X1 U6014 ( .A1(n9829), .A2(n10043), .B1(n10041), .B2(n9864), .ZN(n9830) );
  NAND2_X1 U6015 ( .A1(n4704), .A2(n4702), .ZN(n10104) );
  INV_X1 U6016 ( .A(n4703), .ZN(n4702) );
  NAND2_X1 U6017 ( .A1(n4706), .A2(n4705), .ZN(n4704) );
  OAI22_X1 U6018 ( .A1(n9853), .A2(n10017), .B1(n10014), .B2(n9852), .ZN(n4703) );
  NAND2_X1 U6019 ( .A1(n9928), .A2(n8657), .ZN(n9908) );
  NAND2_X1 U6020 ( .A1(n4654), .A2(n4655), .ZN(n9927) );
  OR2_X1 U6021 ( .A1(n4971), .A2(n4657), .ZN(n4654) );
  NAND2_X1 U6022 ( .A1(n4971), .A2(n5445), .ZN(n9957) );
  AND2_X1 U6023 ( .A1(n10011), .A2(n8619), .ZN(n9993) );
  NAND2_X1 U6024 ( .A1(n5354), .A2(n5353), .ZN(n10027) );
  NAND2_X1 U6025 ( .A1(n7579), .A2(n5254), .ZN(n7792) );
  OAI21_X1 U6026 ( .B1(n7511), .B2(n4685), .A(n4684), .ZN(n7630) );
  OR2_X1 U6027 ( .A1(n5166), .A2(n6991), .ZN(n4648) );
  INV_X1 U6028 ( .A(n9920), .ZN(n10054) );
  AND2_X1 U6029 ( .A1(n9940), .A2(n5730), .ZN(n9920) );
  NAND2_X1 U6030 ( .A1(n5729), .A2(n9898), .ZN(n9940) );
  AND2_X2 U6031 ( .A1(n7247), .A2(n7246), .ZN(n10308) );
  NAND2_X1 U6032 ( .A1(n10097), .A2(n4561), .ZN(n10193) );
  INV_X1 U6033 ( .A(n4562), .ZN(n4561) );
  OAI21_X1 U6034 ( .B1(n10098), .B2(n10163), .A(n10096), .ZN(n4562) );
  NAND2_X1 U6035 ( .A1(n4708), .A2(n4699), .ZN(n10195) );
  NOR2_X1 U6036 ( .A1(n10104), .A2(n4700), .ZN(n4699) );
  OR2_X1 U6037 ( .A1(n10107), .A2(n10163), .ZN(n4708) );
  OR2_X1 U6038 ( .A1(n10105), .A2(n4701), .ZN(n4700) );
  OR2_X1 U6039 ( .A1(n10123), .A2(n10122), .ZN(n10198) );
  AND2_X2 U6040 ( .A1(n7247), .A2(n7050), .ZN(n10301) );
  INV_X1 U6042 ( .A(n5083), .ZN(n10223) );
  NAND2_X1 U6043 ( .A1(n5670), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U6044 ( .A1(n5071), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4527) );
  INV_X1 U6045 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8443) );
  INV_X1 U6046 ( .A(n8726), .ZN(n8442) );
  INV_X1 U6047 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7767) );
  CLKBUF_X1 U6048 ( .A(n5700), .Z(n8561) );
  INV_X1 U6049 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8161) );
  INV_X1 U6050 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7405) );
  OAI21_X1 U6051 ( .B1(n5476), .B2(n5475), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5477) );
  INV_X1 U6052 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n8034) );
  INV_X1 U6053 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7185) );
  INV_X1 U6054 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7146) );
  INV_X1 U6055 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7057) );
  INV_X1 U6056 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8178) );
  INV_X1 U6057 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U6058 ( .A1(n5110), .A2(n10215), .ZN(n4679) );
  OAI21_X1 U6059 ( .B1(n10469), .B2(n10472), .A(n8356), .ZN(n10466) );
  NOR2_X1 U6060 ( .A1(n8360), .A2(n10462), .ZN(n10452) );
  AOI21_X1 U6061 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10450), .ZN(n10449) );
  NOR2_X1 U6062 ( .A1(n10449), .A2(n10448), .ZN(n10447) );
  NAND2_X1 U6063 ( .A1(n4949), .A2(n4948), .ZN(n7781) );
  NAND2_X1 U6064 ( .A1(n4716), .A2(n4718), .ZN(n7330) );
  AOI21_X1 U6065 ( .B1(n4712), .B2(n9154), .A(n4711), .ZN(n4710) );
  NAND2_X1 U6066 ( .A1(n4714), .A2(n6278), .ZN(n4713) );
  OAI21_X1 U6067 ( .B1(n9097), .B2(n9098), .A(n9096), .ZN(n4711) );
  NAND2_X1 U6068 ( .A1(n4491), .A2(n9196), .ZN(n6221) );
  NAND2_X1 U6069 ( .A1(n4499), .A2(n4746), .ZN(P2_U3549) );
  OR2_X1 U6070 ( .A1(n10423), .A2(n6119), .ZN(n4746) );
  NAND2_X1 U6071 ( .A1(n4500), .A2(n10423), .ZN(n4499) );
  NAND2_X1 U6072 ( .A1(n4520), .A2(n4436), .ZN(P2_U3517) );
  AOI21_X1 U6073 ( .B1(n6216), .B2(n10407), .A(n4473), .ZN(n4818) );
  NAND2_X1 U6074 ( .A1(n4574), .A2(n4572), .ZN(P1_U3260) );
  AOI21_X1 U6075 ( .B1(n9749), .B2(n8502), .A(n4573), .ZN(n4572) );
  NAND2_X1 U6076 ( .A1(n9748), .A2(n9857), .ZN(n4574) );
  OAI21_X1 U6077 ( .B1(n10245), .B2(n9751), .A(n9750), .ZN(n4573) );
  NAND3_X1 U6078 ( .A1(n7825), .A2(n8790), .A3(n4414), .ZN(n4397) );
  AND2_X1 U6079 ( .A1(n8741), .A2(n4430), .ZN(n4398) );
  OR4_X1 U6080 ( .A1(n8559), .A2(n8502), .A3(n4560), .A4(n4392), .ZN(n4399) );
  OAI21_X1 U6081 ( .B1(n9115), .B2(n6215), .A(n6214), .ZN(n6216) );
  OR3_X1 U6082 ( .A1(n10073), .A2(n10163), .A3(n10076), .ZN(n4400) );
  INV_X1 U6083 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9497) );
  INV_X1 U6084 ( .A(n5818), .ZN(n6093) );
  OR2_X1 U6085 ( .A1(n9270), .A2(n9247), .ZN(n4401) );
  INV_X1 U6086 ( .A(n6458), .ZN(n4549) );
  NAND2_X1 U6087 ( .A1(n10113), .A2(n9894), .ZN(n4402) );
  NAND2_X1 U6088 ( .A1(n10011), .A2(n4424), .ZN(n9974) );
  OR2_X1 U6089 ( .A1(n9237), .A2(n8774), .ZN(n4403) );
  INV_X1 U6090 ( .A(n8505), .ZN(n5711) );
  NAND2_X1 U6091 ( .A1(n5773), .A2(n5774), .ZN(n8445) );
  XNOR2_X1 U6092 ( .A(n5447), .B(SI_17_), .ZN(n5446) );
  AND2_X1 U6093 ( .A1(n5534), .A2(n5533), .ZN(n9883) );
  INV_X1 U6094 ( .A(n9883), .ZN(n10113) );
  AND2_X1 U6095 ( .A1(n4939), .A2(n4463), .ZN(n4404) );
  AND2_X1 U6096 ( .A1(n4836), .A2(n4401), .ZN(n4405) );
  AOI21_X1 U6097 ( .B1(n4870), .B2(n5449), .A(n5464), .ZN(n4869) );
  INV_X1 U6098 ( .A(n4869), .ZN(n4868) );
  AND2_X1 U6099 ( .A1(n6187), .A2(n6318), .ZN(n4406) );
  AND2_X1 U6100 ( .A1(n4655), .A2(n4445), .ZN(n4407) );
  INV_X1 U6101 ( .A(n5449), .ZN(n4867) );
  OR2_X1 U6102 ( .A1(n9435), .A2(n6015), .ZN(n4408) );
  AND2_X1 U6103 ( .A1(n4778), .A2(n4777), .ZN(n4410) );
  AND2_X1 U6104 ( .A1(n6593), .A2(n6592), .ZN(n4411) );
  NAND2_X1 U6105 ( .A1(n10397), .A2(n7832), .ZN(n6320) );
  INV_X1 U6106 ( .A(n6320), .ZN(n4793) );
  OR2_X1 U6107 ( .A1(n6617), .A2(n9115), .ZN(n6424) );
  AND3_X1 U6108 ( .A1(n5806), .A2(n5805), .A3(n5804), .ZN(n7482) );
  INV_X1 U6109 ( .A(n7482), .ZN(n5807) );
  INV_X1 U6110 ( .A(n9180), .ZN(n9184) );
  AND2_X1 U6111 ( .A1(n8574), .A2(n8518), .ZN(n4412) );
  AND2_X1 U6112 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4413) );
  AND2_X1 U6113 ( .A1(n10085), .A2(n9786), .ZN(n10074) );
  AND2_X1 U6114 ( .A1(n4773), .A2(n4772), .ZN(n4414) );
  AND2_X1 U6115 ( .A1(n5030), .A2(n5029), .ZN(n4415) );
  AND2_X1 U6116 ( .A1(n6357), .A2(n9331), .ZN(n8382) );
  AND2_X1 U6117 ( .A1(n10083), .A2(n10082), .ZN(n4416) );
  AND3_X1 U6118 ( .A1(n5912), .A2(n4916), .A3(n4915), .ZN(n4417) );
  OR2_X1 U6119 ( .A1(n9214), .A2(n4784), .ZN(n4418) );
  NAND2_X1 U6120 ( .A1(n9343), .A2(n5997), .ZN(n9291) );
  OR2_X1 U6121 ( .A1(n6819), .A2(n9552), .ZN(n4419) );
  INV_X1 U6122 ( .A(n8820), .ZN(n4969) );
  INV_X1 U6123 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5836) );
  AND3_X1 U6124 ( .A1(n5796), .A2(n5795), .A3(n5794), .ZN(n4420) );
  INV_X1 U6125 ( .A(n7535), .ZN(n6511) );
  INV_X1 U6126 ( .A(n9192), .ZN(n9409) );
  NAND2_X1 U6127 ( .A1(n5754), .A2(n5753), .ZN(n9192) );
  NAND2_X1 U6128 ( .A1(n9817), .A2(n9821), .ZN(n4422) );
  OR2_X1 U6129 ( .A1(n4904), .A2(n5599), .ZN(n4423) );
  AND2_X1 U6130 ( .A1(n9994), .A2(n8619), .ZN(n4424) );
  INV_X1 U6131 ( .A(n8547), .ZN(n5004) );
  NAND2_X1 U6132 ( .A1(n5651), .A2(n5650), .ZN(n9786) );
  AND2_X1 U6133 ( .A1(n9460), .A2(n8920), .ZN(n4425) );
  INV_X1 U6134 ( .A(n8657), .ZN(n4990) );
  AND2_X1 U6135 ( .A1(n8478), .A2(n7506), .ZN(n4426) );
  OR2_X1 U6136 ( .A1(n6986), .A2(n4628), .ZN(n4427) );
  OR2_X1 U6137 ( .A1(n9123), .A2(n6617), .ZN(n4428) );
  INV_X1 U6138 ( .A(n7656), .ZN(n7314) );
  AND2_X1 U6139 ( .A1(n5748), .A2(n6138), .ZN(n4429) );
  NAND2_X1 U6140 ( .A1(n6547), .A2(n6546), .ZN(n4430) );
  INV_X1 U6141 ( .A(n6345), .ZN(n4803) );
  INV_X1 U6142 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4523) );
  NOR2_X1 U6143 ( .A1(n5270), .A2(n4977), .ZN(n4431) );
  INV_X1 U6144 ( .A(n9415), .ZN(n4787) );
  OR2_X1 U6145 ( .A1(n6932), .A2(n6963), .ZN(n4432) );
  OR2_X1 U6146 ( .A1(n6433), .A2(n4583), .ZN(n4433) );
  INV_X1 U6147 ( .A(n5063), .ZN(n5011) );
  INV_X1 U6148 ( .A(n6168), .ZN(n6173) );
  AND2_X1 U6149 ( .A1(n8829), .A2(n8828), .ZN(n4434) );
  INV_X1 U6150 ( .A(n5295), .ZN(n4621) );
  NAND2_X1 U6151 ( .A1(n4830), .A2(n4829), .ZN(n9150) );
  OR2_X1 U6152 ( .A1(n9415), .A2(n8773), .ZN(n6388) );
  NAND2_X1 U6153 ( .A1(n4513), .A2(n4884), .ZN(n9635) );
  NAND2_X1 U6154 ( .A1(n9221), .A2(n6395), .ZN(n9204) );
  AND2_X1 U6155 ( .A1(n5102), .A2(n4758), .ZN(n4435) );
  OAI21_X1 U6156 ( .B1(n6164), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U6157 ( .A1(n5606), .A2(n5605), .ZN(n10094) );
  INV_X1 U6158 ( .A(n10094), .ZN(n4568) );
  AND3_X1 U6159 ( .A1(n4816), .A2(n4518), .A3(n4818), .ZN(n4436) );
  INV_X2 U6160 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10215) );
  AND2_X1 U6161 ( .A1(n9569), .A2(n9580), .ZN(n4437) );
  INV_X1 U6162 ( .A(n6863), .ZN(n6873) );
  NAND2_X1 U6163 ( .A1(n5939), .A2(n5938), .ZN(n9465) );
  AND2_X1 U6164 ( .A1(n7924), .A2(n4792), .ZN(n4438) );
  NOR2_X1 U6165 ( .A1(n5799), .A2(n7265), .ZN(n4439) );
  AND2_X1 U6166 ( .A1(n4855), .A2(n4854), .ZN(n4440) );
  OR2_X1 U6167 ( .A1(n9123), .A2(n4782), .ZN(n4441) );
  AND2_X1 U6168 ( .A1(n4419), .A2(n4514), .ZN(n4442) );
  INV_X1 U6169 ( .A(n6347), .ZN(n4802) );
  NAND2_X1 U6170 ( .A1(n5975), .A2(n5974), .ZN(n9450) );
  AND2_X1 U6171 ( .A1(n9089), .A2(n9090), .ZN(n4443) );
  NAND2_X1 U6172 ( .A1(n5788), .A2(n5787), .ZN(n7720) );
  AND2_X1 U6173 ( .A1(n6682), .A2(n6677), .ZN(n4444) );
  NAND2_X1 U6174 ( .A1(n10133), .A2(n9947), .ZN(n4445) );
  INV_X1 U6175 ( .A(n4835), .ZN(n4834) );
  INV_X1 U6176 ( .A(n5294), .ZN(n4620) );
  NAND2_X1 U6177 ( .A1(n4489), .A2(n5258), .ZN(n5294) );
  XNOR2_X1 U6178 ( .A(n9400), .B(n9165), .ZN(n6458) );
  AND2_X1 U6179 ( .A1(n5466), .A2(SI_18_), .ZN(n4446) );
  AND2_X1 U6180 ( .A1(n4809), .A2(n4730), .ZN(n4447) );
  AND2_X1 U6181 ( .A1(n4946), .A2(n4944), .ZN(n4448) );
  NAND2_X1 U6182 ( .A1(n9470), .A2(n8922), .ZN(n4449) );
  INV_X1 U6183 ( .A(n4401), .ZN(n4743) );
  INV_X1 U6184 ( .A(n6440), .ZN(n4545) );
  INV_X1 U6185 ( .A(n5931), .ZN(n4524) );
  INV_X1 U6186 ( .A(n6005), .ZN(n4839) );
  OR2_X1 U6187 ( .A1(n9442), .A2(n9280), .ZN(n6005) );
  INV_X1 U6188 ( .A(n8599), .ZN(n5000) );
  AND2_X1 U6189 ( .A1(n6852), .A2(n6851), .ZN(n4450) );
  OR2_X1 U6190 ( .A1(n9378), .A2(n6225), .ZN(n6432) );
  INV_X1 U6191 ( .A(n6432), .ZN(n5018) );
  AND2_X1 U6192 ( .A1(n4603), .A2(n4605), .ZN(n4451) );
  AND2_X1 U6193 ( .A1(n10138), .A2(n9962), .ZN(n4452) );
  NOR2_X1 U6194 ( .A1(n9394), .A2(n8916), .ZN(n4453) );
  INV_X1 U6195 ( .A(n5035), .ZN(n9879) );
  NOR2_X1 U6196 ( .A1(n9917), .A2(n5036), .ZN(n5035) );
  INV_X1 U6197 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8150) );
  AND2_X1 U6198 ( .A1(n10159), .A2(n10042), .ZN(n4454) );
  NOR2_X1 U6199 ( .A1(n10133), .A2(n9947), .ZN(n4455) );
  OR2_X1 U6200 ( .A1(n5896), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n4456) );
  INV_X1 U6201 ( .A(n6585), .ZN(n6586) );
  OR2_X1 U6202 ( .A1(n4958), .A2(n4965), .ZN(n4457) );
  INV_X1 U6203 ( .A(n7454), .ZN(n7466) );
  AND2_X1 U6204 ( .A1(n5173), .A2(n5172), .ZN(n7454) );
  INV_X1 U6205 ( .A(n6876), .ZN(n10085) );
  AND2_X1 U6206 ( .A1(n5643), .A2(n5642), .ZN(n6876) );
  OAI21_X1 U6207 ( .B1(n4906), .B2(n4423), .A(n5598), .ZN(n4903) );
  OR2_X1 U6208 ( .A1(n6554), .A2(n6553), .ZN(n4458) );
  NAND2_X1 U6209 ( .A1(n6533), .A2(n4952), .ZN(n4459) );
  AND2_X1 U6210 ( .A1(n9172), .A2(n6066), .ZN(n4460) );
  OR2_X1 U6211 ( .A1(n5488), .A2(n4446), .ZN(n4461) );
  INV_X1 U6212 ( .A(n9603), .ZN(n4861) );
  AND3_X1 U6213 ( .A1(n5279), .A2(n5278), .A3(n5277), .ZN(n5280) );
  INV_X1 U6214 ( .A(n5001), .ZN(n9827) );
  NAND2_X1 U6215 ( .A1(n5005), .A2(n5002), .ZN(n5001) );
  INV_X1 U6216 ( .A(n4836), .ZN(n4744) );
  NAND2_X1 U6217 ( .A1(n4838), .A2(n4408), .ZN(n4836) );
  AND2_X1 U6218 ( .A1(n6424), .A2(n6422), .ZN(n6461) );
  INV_X1 U6219 ( .A(n6461), .ZN(n4809) );
  INV_X1 U6220 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4916) );
  INV_X1 U6221 ( .A(n5154), .ZN(n5087) );
  XNOR2_X1 U6222 ( .A(n5315), .B(SI_11_), .ZN(n5314) );
  NAND2_X1 U6223 ( .A1(n6116), .A2(n6115), .ZN(n9378) );
  AND2_X1 U6224 ( .A1(n6422), .A2(n6421), .ZN(n4462) );
  OR2_X1 U6225 ( .A1(n4941), .A2(n4411), .ZN(n4463) );
  AND2_X1 U6226 ( .A1(n5575), .A2(n4402), .ZN(n4464) );
  AND2_X1 U6227 ( .A1(n4410), .A2(n9277), .ZN(n4465) );
  NAND2_X1 U6228 ( .A1(n7331), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4466) );
  AND2_X1 U6229 ( .A1(n8715), .A2(n8705), .ZN(n4467) );
  INV_X1 U6230 ( .A(n5013), .ZN(n5012) );
  AND2_X1 U6231 ( .A1(n4715), .A2(n9036), .ZN(n4468) );
  AND2_X1 U6232 ( .A1(n4858), .A2(n4856), .ZN(n4469) );
  INV_X1 U6233 ( .A(n5708), .ZN(n5008) );
  AND2_X1 U6234 ( .A1(n5062), .A2(n9241), .ZN(n4470) );
  NAND2_X1 U6235 ( .A1(n10073), .A2(n4974), .ZN(n4471) );
  AND2_X1 U6236 ( .A1(n9558), .A2(n4887), .ZN(n4886) );
  INV_X1 U6237 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U6238 ( .A1(n5373), .A2(n5322), .ZN(n5338) );
  NAND2_X1 U6239 ( .A1(n6704), .A2(n4849), .ZN(n7646) );
  NAND2_X1 U6240 ( .A1(n4509), .A2(n6697), .ZN(n7561) );
  AND4_X1 U6241 ( .A1(n6014), .A2(n6013), .A3(n6012), .A4(n6011), .ZN(n9289)
         );
  NAND2_X1 U6242 ( .A1(n9355), .A2(n4778), .ZN(n9301) );
  NAND2_X1 U6243 ( .A1(n4737), .A2(n5748), .ZN(n6135) );
  INV_X2 U6244 ( .A(n10405), .ZN(n10407) );
  NAND2_X1 U6245 ( .A1(n6250), .A2(n6249), .ZN(n9100) );
  INV_X1 U6246 ( .A(n9100), .ZN(n4781) );
  NAND2_X1 U6247 ( .A1(n7411), .A2(n8518), .ZN(n7446) );
  NAND2_X1 U6248 ( .A1(n7628), .A2(n8607), .ZN(n7572) );
  NAND2_X1 U6249 ( .A1(n4827), .A2(n4828), .ZN(n8315) );
  NAND2_X1 U6250 ( .A1(n6432), .A2(n6284), .ZN(n9377) );
  INV_X1 U6251 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5912) );
  INV_X1 U6252 ( .A(n8819), .ZN(n4968) );
  INV_X1 U6253 ( .A(n4949), .ZN(n7609) );
  OR2_X1 U6254 ( .A1(n9465), .A2(n8921), .ZN(n4472) );
  NAND2_X1 U6255 ( .A1(n5021), .A2(n6318), .ZN(n7872) );
  NAND2_X1 U6256 ( .A1(n7825), .A2(n4773), .ZN(n4774) );
  NAND2_X1 U6257 ( .A1(n6568), .A2(n6569), .ZN(n4970) );
  NOR2_X1 U6258 ( .A1(n10020), .A2(n10154), .ZN(n5045) );
  NOR2_X1 U6259 ( .A1(n10407), .A2(n4819), .ZN(n4473) );
  AND2_X1 U6260 ( .A1(n6112), .A2(n6111), .ZN(n4474) );
  INV_X1 U6261 ( .A(n6279), .ZN(n10398) );
  INV_X1 U6262 ( .A(n10163), .ZN(n4976) );
  INV_X1 U6263 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U6264 ( .A1(n4545), .A2(n4544), .ZN(n7705) );
  AND2_X1 U6265 ( .A1(n7502), .A2(n6515), .ZN(n4930) );
  INV_X1 U6266 ( .A(n7640), .ZN(n5026) );
  AND2_X1 U6267 ( .A1(n8442), .A2(n8502), .ZN(n8702) );
  INV_X1 U6268 ( .A(n10313), .ZN(n9351) );
  OR2_X1 U6269 ( .A1(n6280), .A2(n6203), .ZN(n10313) );
  INV_X1 U6270 ( .A(n7709), .ZN(n7313) );
  INV_X1 U6271 ( .A(n7173), .ZN(n7134) );
  INV_X1 U6272 ( .A(n9460), .ZN(n4772) );
  NAND2_X1 U6273 ( .A1(n5329), .A2(n5328), .ZN(n10170) );
  INV_X1 U6274 ( .A(n10170), .ZN(n5029) );
  NAND2_X1 U6275 ( .A1(n7532), .A2(n4930), .ZN(n7501) );
  OR2_X1 U6276 ( .A1(n9154), .A2(n6202), .ZN(n6484) );
  AND2_X1 U6277 ( .A1(n5713), .A2(n8719), .ZN(n10045) );
  NAND2_X1 U6278 ( .A1(n6512), .A2(n6511), .ZN(n7532) );
  AND2_X1 U6279 ( .A1(n7079), .A2(n6917), .ZN(n4475) );
  INV_X1 U6280 ( .A(n7154), .ZN(n4673) );
  INV_X1 U6281 ( .A(n9857), .ZN(n8502) );
  INV_X1 U6282 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U6283 ( .A1(n4393), .A2(n7022), .ZN(n4490) );
  NAND3_X1 U6284 ( .A1(n5021), .A2(n6328), .A3(n4406), .ZN(n4493) );
  NAND2_X1 U6285 ( .A1(n4494), .A2(n5188), .ZN(n5197) );
  NAND2_X1 U6286 ( .A1(n5185), .A2(n5184), .ZN(n4494) );
  OAI211_X1 U6287 ( .C1(n5185), .C2(n4496), .A(n4495), .B(n5196), .ZN(n4497)
         );
  NAND2_X1 U6288 ( .A1(n4390), .A2(n5188), .ZN(n4495) );
  INV_X1 U6289 ( .A(n5188), .ZN(n4496) );
  NAND3_X1 U6290 ( .A1(n4789), .A2(n4470), .A3(n4498), .ZN(n9243) );
  NAND3_X1 U6291 ( .A1(n9310), .A2(n6198), .A3(n9315), .ZN(n4498) );
  AND2_X2 U6292 ( .A1(n9243), .A2(n6404), .ZN(n9220) );
  NAND3_X1 U6293 ( .A1(n4820), .A2(n9383), .A3(n9382), .ZN(n4500) );
  NAND3_X1 U6294 ( .A1(n4850), .A2(n6714), .A3(n4501), .ZN(n4504) );
  OR2_X1 U6295 ( .A1(n4505), .A2(n4851), .ZN(n4501) );
  AND2_X1 U6296 ( .A1(n4508), .A2(n4507), .ZN(n4503) );
  INV_X1 U6297 ( .A(n6697), .ZN(n4505) );
  NAND2_X1 U6298 ( .A1(n4850), .A2(n6714), .ZN(n4506) );
  INV_X1 U6299 ( .A(n7841), .ZN(n7840) );
  NAND4_X1 U6300 ( .A1(n5667), .A2(n5664), .A3(n5668), .A4(n5673), .ZN(n4511)
         );
  NAND3_X1 U6301 ( .A1(n5667), .A2(n5664), .A3(n5668), .ZN(n5670) );
  NAND3_X1 U6302 ( .A1(n6837), .A2(n9526), .A3(n4886), .ZN(n4513) );
  INV_X1 U6303 ( .A(n9635), .ZN(n4512) );
  NAND2_X2 U6304 ( .A1(n9584), .A2(n6785), .ZN(n9538) );
  NAND2_X2 U6305 ( .A1(n6674), .A2(n6673), .ZN(n4515) );
  NAND2_X1 U6306 ( .A1(n4515), .A2(n6677), .ZN(n7395) );
  NAND2_X1 U6307 ( .A1(n7190), .A2(n4515), .ZN(n7193) );
  NAND2_X1 U6308 ( .A1(n4516), .A2(n4901), .ZN(n4900) );
  NAND2_X1 U6309 ( .A1(n4516), .A2(n6742), .ZN(n8302) );
  INV_X1 U6310 ( .A(n4771), .ZN(n4768) );
  NAND2_X1 U6311 ( .A1(n5659), .A2(n5658), .ZN(n5700) );
  AOI21_X2 U6312 ( .B1(n9961), .B2(n8603), .A(n5709), .ZN(n9929) );
  NAND2_X2 U6313 ( .A1(n4697), .A2(n5006), .ZN(n9961) );
  NAND3_X1 U6314 ( .A1(n4400), .A2(n4416), .A3(n4471), .ZN(n10190) );
  NAND2_X2 U6315 ( .A1(n7411), .A2(n4412), .ZN(n7511) );
  NAND4_X1 U6316 ( .A1(n5067), .A2(n5066), .A3(n5065), .A4(n5068), .ZN(n5666)
         );
  AND2_X2 U6317 ( .A1(n10220), .A2(n5083), .ZN(n5156) );
  NOR2_X1 U6318 ( .A1(n5677), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4529) );
  XNOR2_X1 U6319 ( .A(n4517), .B(n6847), .ZN(n6660) );
  OAI22_X1 U6320 ( .A1(n6875), .A2(n7173), .B1(n7424), .B2(n6873), .ZN(n4517)
         );
  NAND2_X2 U6321 ( .A1(n5081), .A2(n5083), .ZN(n5611) );
  NAND2_X1 U6322 ( .A1(n6678), .A2(n4559), .ZN(n4558) );
  NAND2_X2 U6323 ( .A1(n9185), .A2(n4831), .ZN(n4830) );
  NAND2_X1 U6324 ( .A1(n9121), .A2(n9120), .ZN(n9119) );
  AOI22_X2 U6325 ( .A1(n9212), .A2(n6047), .B1(n9420), .B2(n8918), .ZN(n9200)
         );
  NAND2_X2 U6326 ( .A1(n4420), .A2(n5798), .ZN(n8930) );
  NAND2_X1 U6327 ( .A1(n9387), .A2(n5047), .ZN(n4521) );
  INV_X1 U6328 ( .A(n7745), .ZN(n4729) );
  AOI21_X1 U6329 ( .B1(n7676), .B2(n5844), .A(n4728), .ZN(n7736) );
  NAND2_X1 U6330 ( .A1(n4716), .A2(n4468), .ZN(n9034) );
  INV_X1 U6331 ( .A(n4721), .ZN(n4719) );
  NAND2_X1 U6332 ( .A1(n4713), .A2(n4710), .ZN(P2_U3264) );
  NAND2_X1 U6333 ( .A1(n4857), .A2(n4858), .ZN(n6826) );
  NAND2_X2 U6334 ( .A1(n5720), .A2(n8724), .ZN(n5326) );
  NAND2_X1 U6335 ( .A1(n5100), .A2(n4525), .ZN(n4538) );
  NAND2_X1 U6336 ( .A1(n4528), .A2(n4527), .ZN(n5669) );
  OAI21_X1 U6337 ( .B1(n4529), .B2(n10215), .A(P1_IR_REG_24__SCAN_IN), .ZN(
        n4528) );
  OR2_X2 U6338 ( .A1(n8706), .A2(n10076), .ZN(n4752) );
  NAND2_X1 U6339 ( .A1(n5561), .A2(n5560), .ZN(n5563) );
  NAND2_X1 U6340 ( .A1(n8713), .A2(n4753), .ZN(n8722) );
  NOR2_X1 U6341 ( .A1(n4755), .A2(n4606), .ZN(n8730) );
  NAND2_X1 U6342 ( .A1(n4905), .A2(n5582), .ZN(n5600) );
  NAND2_X1 U6343 ( .A1(n4644), .A2(n8689), .ZN(n4643) );
  NAND2_X1 U6344 ( .A1(n9804), .A2(n8687), .ZN(n5597) );
  INV_X1 U6345 ( .A(n4993), .ZN(n4992) );
  NAND2_X1 U6346 ( .A1(n9178), .A2(n6285), .ZN(n9163) );
  NAND2_X1 U6347 ( .A1(n6218), .A2(n10335), .ZN(n6219) );
  OAI21_X1 U6348 ( .B1(n5528), .B2(n5527), .A(n5526), .ZN(n5543) );
  NAND3_X1 U6349 ( .A1(n4530), .A2(n6476), .A3(n6475), .ZN(P2_U3244) );
  NAND2_X1 U6350 ( .A1(n6283), .A2(n6282), .ZN(n4530) );
  NAND2_X1 U6351 ( .A1(n4807), .A2(n4812), .ZN(n6224) );
  NAND2_X1 U6352 ( .A1(n6198), .A2(n4790), .ZN(n4789) );
  NAND2_X1 U6353 ( .A1(n5156), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5084) );
  XNOR2_X1 U6354 ( .A(n4531), .B(n6847), .ZN(n7846) );
  NAND2_X1 U6355 ( .A1(n4534), .A2(n4556), .ZN(n6641) );
  NAND2_X1 U6356 ( .A1(n4395), .A2(n7179), .ZN(n4534) );
  OAI21_X2 U6357 ( .B1(n9163), .B2(n9173), .A(n6200), .ZN(n9145) );
  NAND2_X1 U6358 ( .A1(n6752), .A2(n6751), .ZN(n4557) );
  NOR2_X1 U6359 ( .A1(n5475), .A2(n4913), .ZN(n4911) );
  OAI21_X1 U6360 ( .B1(n9567), .B2(n9647), .A(n9571), .ZN(n6777) );
  NAND2_X1 U6361 ( .A1(n6778), .A2(n9581), .ZN(n4564) );
  NOR2_X1 U6362 ( .A1(n5658), .A2(n5655), .ZN(n4845) );
  NAND2_X2 U6363 ( .A1(n7930), .A2(n6337), .ZN(n8372) );
  NAND2_X1 U6364 ( .A1(n4788), .A2(n7745), .ZN(n7678) );
  NOR2_X2 U6365 ( .A1(n5746), .A2(n5745), .ZN(n5747) );
  NOR4_X2 U6366 ( .A1(n6464), .A2(n6463), .A3(n9377), .A4(n6462), .ZN(n6465)
         );
  NOR4_X1 U6367 ( .A1(n6449), .A2(n7617), .A3(n6448), .A4(n6447), .ZN(n6450)
         );
  NAND2_X1 U6368 ( .A1(n4546), .A2(n4462), .ZN(n6423) );
  NAND2_X1 U6369 ( .A1(n6420), .A2(n6419), .ZN(n4546) );
  AOI21_X1 U6370 ( .B1(n4550), .B2(n4548), .A(n4547), .ZN(n6417) );
  AND3_X2 U6371 ( .A1(n6278), .A2(n6466), .A3(n8447), .ZN(n6435) );
  OR2_X1 U6372 ( .A1(n4851), .A2(n7562), .ZN(n4850) );
  NAND2_X1 U6373 ( .A1(n8425), .A2(n6779), .ZN(n9568) );
  NAND2_X1 U6374 ( .A1(n8672), .A2(n8671), .ZN(n8674) );
  NAND2_X1 U6375 ( .A1(n8665), .A2(n8714), .ZN(n4552) );
  NAND2_X1 U6376 ( .A1(n8666), .A2(n8702), .ZN(n4553) );
  AND4_X1 U6377 ( .A1(n8632), .A2(n8633), .A3(n9976), .A4(n8631), .ZN(n8647)
         );
  NAND2_X1 U6378 ( .A1(n4882), .A2(n4880), .ZN(n5381) );
  INV_X1 U6379 ( .A(n4970), .ZN(n4966) );
  INV_X1 U6380 ( .A(n4962), .ZN(n4554) );
  OAI21_X2 U6381 ( .B1(n8855), .B2(n4943), .A(n6585), .ZN(n6589) );
  XNOR2_X1 U6382 ( .A(n6713), .B(n6847), .ZN(n7841) );
  AOI21_X2 U6383 ( .B1(n7904), .B2(n6734), .A(n5059), .ZN(n8245) );
  INV_X1 U6384 ( .A(n5700), .ZN(n4560) );
  NAND2_X1 U6385 ( .A1(n6653), .A2(n6654), .ZN(n7127) );
  NAND2_X1 U6386 ( .A1(n6647), .A2(n7117), .ZN(n6653) );
  OR2_X1 U6387 ( .A1(n6702), .A2(n4555), .ZN(n6704) );
  NOR2_X2 U6388 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5074) );
  INV_X1 U6389 ( .A(n5470), .ZN(n5474) );
  NAND2_X1 U6390 ( .A1(n7943), .A2(n7944), .ZN(n7904) );
  AOI21_X1 U6391 ( .B1(n9517), .B2(n9515), .A(n9514), .ZN(n6901) );
  INV_X1 U6392 ( .A(n5100), .ZN(n4757) );
  INV_X1 U6393 ( .A(n5471), .ZN(n5473) );
  NAND2_X1 U6394 ( .A1(n4900), .A2(n6749), .ZN(n8425) );
  NOR2_X2 U6395 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5073) );
  INV_X1 U6396 ( .A(n7118), .ZN(n6646) );
  NAND2_X1 U6397 ( .A1(n6644), .A2(n6645), .ZN(n7118) );
  NOR2_X2 U6398 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5068) );
  AOI21_X2 U6399 ( .B1(n9812), .B2(n4705), .A(n9811), .ZN(n10097) );
  NAND2_X1 U6400 ( .A1(n7360), .A2(n5702), .ZN(n8564) );
  AOI21_X2 U6401 ( .B1(n9892), .B2(n9891), .A(n4563), .ZN(n9875) );
  NAND2_X1 U6402 ( .A1(n4752), .A2(n4467), .ZN(n4751) );
  NAND2_X1 U6403 ( .A1(n4751), .A2(n8707), .ZN(n8712) );
  INV_X1 U6404 ( .A(n6197), .ZN(n4790) );
  NOR2_X1 U6405 ( .A1(n6991), .A2(n5840), .ZN(n5786) );
  NAND2_X1 U6406 ( .A1(n6833), .A2(n6834), .ZN(n9525) );
  NAND2_X1 U6407 ( .A1(n4821), .A2(n9751), .ZN(n5095) );
  NAND2_X1 U6408 ( .A1(n4586), .A2(n5144), .ZN(n5147) );
  NAND2_X1 U6409 ( .A1(n5128), .A2(n5129), .ZN(n4586) );
  INV_X1 U6410 ( .A(n6833), .ZN(n6836) );
  AOI21_X1 U6411 ( .B1(n9570), .B2(n4437), .A(n4564), .ZN(n4584) );
  NAND2_X1 U6412 ( .A1(n9614), .A2(n9612), .ZN(n9611) );
  NAND2_X1 U6413 ( .A1(n5204), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5225) );
  NAND3_X1 U6414 ( .A1(n4640), .A2(n4647), .A3(n4980), .ZN(n4565) );
  NOR2_X2 U6415 ( .A1(n5436), .A2(n4567), .ZN(n5455) );
  NOR2_X2 U6416 ( .A1(n5498), .A2(n5497), .ZN(n4570) );
  NAND2_X1 U6417 ( .A1(n4757), .A2(n4435), .ZN(n5078) );
  NAND2_X1 U6418 ( .A1(n4857), .A2(n4469), .ZN(n9614) );
  OAI21_X1 U6419 ( .B1(n6423), .B2(n4633), .A(n4630), .ZN(n4632) );
  OAI21_X1 U6420 ( .B1(n6400), .B2(n6383), .A(n4852), .ZN(n6385) );
  NAND2_X1 U6421 ( .A1(n4582), .A2(n4581), .ZN(n6311) );
  INV_X2 U6422 ( .A(n6435), .ZN(n4583) );
  NAND2_X1 U6423 ( .A1(n5213), .A2(n5214), .ZN(n5217) );
  NAND2_X1 U6424 ( .A1(n5012), .A2(n4696), .ZN(n4695) );
  NAND2_X1 U6425 ( .A1(n5705), .A2(n8638), .ZN(n5013) );
  OAI21_X2 U6426 ( .B1(n5381), .B2(n5380), .A(n5379), .ZN(n5406) );
  NAND2_X1 U6427 ( .A1(n4806), .A2(n4804), .ZN(n9178) );
  INV_X1 U6428 ( .A(n6704), .ZN(n4851) );
  NAND2_X1 U6429 ( .A1(n5281), .A2(n4912), .ZN(n5660) );
  XNOR2_X1 U6430 ( .A(n4586), .B(n5142), .ZN(n5131) );
  NAND2_X1 U6431 ( .A1(n5528), .A2(n4590), .ZN(n4588) );
  NAND2_X1 U6432 ( .A1(n5528), .A2(n4596), .ZN(n4589) );
  NAND2_X1 U6433 ( .A1(n5408), .A2(n4603), .ZN(n4600) );
  NAND2_X1 U6434 ( .A1(n4600), .A2(n4601), .ZN(n4865) );
  NAND3_X1 U6435 ( .A1(n8723), .A2(n4399), .A3(n4608), .ZN(n4607) );
  NAND2_X1 U6436 ( .A1(n5297), .A2(n5296), .ZN(n5299) );
  XNOR2_X1 U6437 ( .A(n4612), .B(n5231), .ZN(n6995) );
  NAND2_X1 U6438 ( .A1(n6328), .A2(n6337), .ZN(n6331) );
  NAND2_X1 U6439 ( .A1(n5297), .A2(n5295), .ZN(n5272) );
  NAND2_X1 U6440 ( .A1(n4625), .A2(n4623), .ZN(n4622) );
  NAND2_X1 U6441 ( .A1(n4624), .A2(n6364), .ZN(n4623) );
  OAI21_X1 U6442 ( .B1(n6351), .B2(n4803), .A(n6346), .ZN(n4624) );
  NAND2_X1 U6443 ( .A1(n4626), .A2(n6363), .ZN(n4625) );
  OAI21_X1 U6444 ( .B1(n6351), .B2(n6350), .A(n6349), .ZN(n4626) );
  NAND2_X1 U6445 ( .A1(n6986), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4627) );
  NOR2_X1 U6446 ( .A1(n4631), .A2(n6463), .ZN(n4630) );
  NAND2_X1 U6447 ( .A1(n4632), .A2(n4433), .ZN(n4891) );
  NAND2_X1 U6448 ( .A1(n4636), .A2(n4879), .ZN(n4635) );
  NAND2_X1 U6449 ( .A1(n4637), .A2(n6408), .ZN(n4636) );
  NAND2_X1 U6450 ( .A1(n6391), .A2(n6390), .ZN(n4637) );
  NAND3_X1 U6451 ( .A1(n4464), .A2(n5522), .A3(n5521), .ZN(n4647) );
  INV_X1 U6452 ( .A(n4645), .ZN(n4644) );
  CLKBUF_X1 U6453 ( .A(n4647), .Z(n4638) );
  NAND3_X1 U6454 ( .A1(n4638), .A2(n4980), .A3(n4646), .ZN(n4639) );
  NAND3_X1 U6455 ( .A1(n4431), .A2(n4409), .A3(n7591), .ZN(n4650) );
  AOI21_X1 U6456 ( .B1(n8284), .B2(n8472), .A(n5293), .ZN(n8267) );
  NAND2_X1 U6457 ( .A1(n4971), .A2(n4407), .ZN(n4653) );
  NAND4_X1 U6458 ( .A1(n5663), .A2(n4658), .A3(n4681), .A4(n4659), .ZN(n5100)
         );
  INV_X1 U6459 ( .A(n5190), .ZN(n5664) );
  NAND2_X1 U6460 ( .A1(n5354), .A2(n4664), .ZN(n4663) );
  NAND3_X1 U6461 ( .A1(n4680), .A2(n5170), .A3(n4679), .ZN(n7093) );
  NAND3_X1 U6462 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4680) );
  OAI21_X2 U6463 ( .B1(n9875), .B2(n8544), .A(n8678), .ZN(n9863) );
  NOR2_X2 U6464 ( .A1(n5076), .A2(n5665), .ZN(n4681) );
  NAND2_X1 U6465 ( .A1(n7511), .A2(n4686), .ZN(n4683) );
  NAND2_X1 U6466 ( .A1(n4683), .A2(n4682), .ZN(n5704) );
  INV_X1 U6467 ( .A(n8575), .ZN(n4690) );
  OR2_X2 U6468 ( .A1(n8321), .A2(n5013), .ZN(n4693) );
  INV_X2 U6469 ( .A(n5432), .ZN(n8466) );
  NAND2_X2 U6470 ( .A1(n5326), .A2(n6986), .ZN(n5432) );
  NAND2_X1 U6471 ( .A1(n9053), .A2(n9052), .ZN(n9066) );
  NAND2_X1 U6472 ( .A1(n9049), .A2(n9048), .ZN(n4709) );
  NOR2_X1 U6473 ( .A1(n8253), .A2(n8254), .ZN(n9049) );
  NAND2_X1 U6474 ( .A1(n9023), .A2(n4717), .ZN(n4716) );
  MUX2_X1 U6475 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10334), .S(n8931), .Z(n7220)
         );
  NOR2_X1 U6476 ( .A1(n7681), .A2(n5846), .ZN(n4728) );
  NAND3_X1 U6477 ( .A1(n7751), .A2(n7750), .A3(n4729), .ZN(n7676) );
  NAND2_X2 U6478 ( .A1(n9119), .A2(n6097), .ZN(n6222) );
  NAND2_X1 U6479 ( .A1(n4825), .A2(n4824), .ZN(n8385) );
  NAND2_X1 U6480 ( .A1(n4823), .A2(n4827), .ZN(n4825) );
  NAND2_X1 U6481 ( .A1(n4732), .A2(n4733), .ZN(n9121) );
  NAND3_X1 U6482 ( .A1(n4830), .A2(n4829), .A3(n9137), .ZN(n4732) );
  NAND3_X1 U6483 ( .A1(n5952), .A2(n5747), .A3(n4429), .ZN(n5771) );
  NAND3_X1 U6484 ( .A1(n5952), .A2(n5747), .A3(n4735), .ZN(n4738) );
  CLKBUF_X1 U6485 ( .A(n5015), .Z(n4737) );
  INV_X1 U6486 ( .A(n4737), .ZN(n6133) );
  NAND2_X2 U6487 ( .A1(n7628), .A2(n5009), .ZN(n7789) );
  NAND2_X1 U6488 ( .A1(n4757), .A2(n4756), .ZN(n5080) );
  INV_X1 U6489 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4758) );
  OAI21_X1 U6490 ( .B1(n4763), .B2(n4761), .A(n4759), .ZN(n8698) );
  NAND2_X1 U6491 ( .A1(n4766), .A2(n4764), .ZN(n4760) );
  NAND2_X1 U6492 ( .A1(n8693), .A2(n4765), .ZN(n4764) );
  INV_X1 U6493 ( .A(n8686), .ZN(n4766) );
  AND2_X1 U6494 ( .A1(n8684), .A2(n8685), .ZN(n4767) );
  XNOR2_X1 U6495 ( .A(n6650), .B(n7368), .ZN(n7248) );
  NAND2_X2 U6496 ( .A1(n4769), .A2(n4768), .ZN(n6650) );
  AND2_X1 U6497 ( .A1(n4770), .A2(n5085), .ZN(n4769) );
  NAND2_X1 U6498 ( .A1(n5087), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4770) );
  OAI21_X1 U6499 ( .B1(n5086), .B2(n5174), .A(n5084), .ZN(n4771) );
  NAND2_X1 U6500 ( .A1(n5771), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6205) );
  NAND3_X1 U6501 ( .A1(n7825), .A2(n8790), .A3(n4773), .ZN(n8389) );
  INV_X1 U6502 ( .A(n4774), .ZN(n8374) );
  NAND3_X1 U6503 ( .A1(n6171), .A2(n4776), .A3(n6497), .ZN(n7723) );
  NAND2_X1 U6504 ( .A1(n9133), .A2(n9127), .ZN(n9123) );
  NAND2_X1 U6505 ( .A1(n7705), .A2(n7746), .ZN(n4788) );
  NAND2_X1 U6506 ( .A1(n9309), .A2(n6197), .ZN(n9239) );
  NAND2_X1 U6507 ( .A1(n5015), .A2(n4791), .ZN(n5774) );
  NAND2_X1 U6508 ( .A1(n8372), .A2(n4797), .ZN(n4795) );
  INV_X1 U6509 ( .A(n8372), .ZN(n4800) );
  NAND3_X1 U6510 ( .A1(n4795), .A2(n6193), .A3(n4794), .ZN(n6195) );
  NAND2_X1 U6511 ( .A1(n9221), .A2(n4805), .ZN(n4806) );
  AOI21_X1 U6512 ( .B1(n6217), .B2(n10313), .A(n6216), .ZN(n9382) );
  NAND2_X1 U6513 ( .A1(n6217), .A2(n4817), .ZN(n4816) );
  OAI211_X2 U6514 ( .C1(n5799), .C2(n8931), .A(n5816), .B(n5815), .ZN(n6488)
         );
  XNOR2_X1 U6515 ( .A(n5109), .B(n5108), .ZN(n7017) );
  MUX2_X1 U6516 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9513), .S(n5799), .Z(n10353)
         );
  NAND4_X1 U6517 ( .A1(n4821), .A2(n8147), .A3(n8345), .A4(
        P1_ADDR_REG_4__SCAN_IN), .ZN(n8157) );
  OAI21_X1 U6518 ( .B1(n9185), .B2(n4832), .A(n4831), .ZN(n9151) );
  NOR2_X1 U6519 ( .A1(n9409), .A2(n9206), .ZN(n4835) );
  OAI21_X2 U6520 ( .B1(n7138), .B2(n7139), .A(n4843), .ZN(n7171) );
  NAND2_X1 U6521 ( .A1(n4843), .A2(n4842), .ZN(n7139) );
  NAND2_X1 U6522 ( .A1(n6660), .A2(n6661), .ZN(n4842) );
  OR2_X1 U6523 ( .A1(n6660), .A2(n6661), .ZN(n4843) );
  NAND2_X1 U6524 ( .A1(n6657), .A2(n7128), .ZN(n7138) );
  NAND2_X1 U6525 ( .A1(n4844), .A2(n6667), .ZN(n7188) );
  NAND2_X1 U6526 ( .A1(n7171), .A2(n7170), .ZN(n4844) );
  XNOR2_X1 U6527 ( .A(n6664), .B(n6665), .ZN(n7170) );
  XNOR2_X1 U6528 ( .A(n6662), .B(n6847), .ZN(n6664) );
  AOI21_X1 U6529 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(n10215), .A(n4845), .ZN(
        n4848) );
  NAND2_X1 U6530 ( .A1(n5658), .A2(n4847), .ZN(n4846) );
  NOR2_X1 U6531 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n10215), .ZN(n4847) );
  NAND2_X1 U6532 ( .A1(n8726), .A2(n9857), .ZN(n5701) );
  OAI21_X1 U6533 ( .B1(n5450), .B2(n4868), .A(n4862), .ZN(n5489) );
  NAND2_X1 U6534 ( .A1(n5639), .A2(n5638), .ZN(n4873) );
  NAND2_X1 U6535 ( .A1(n5301), .A2(n4883), .ZN(n4882) );
  NAND2_X1 U6536 ( .A1(n4882), .A2(n5317), .ZN(n5337) );
  NAND2_X1 U6537 ( .A1(n5301), .A2(n5300), .ZN(n5318) );
  AOI21_X1 U6538 ( .B1(n4891), .B2(n6438), .A(n4890), .ZN(n6439) );
  NOR2_X1 U6539 ( .A1(n9377), .A2(n6427), .ZN(n4894) );
  NAND2_X1 U6540 ( .A1(n5563), .A2(n4906), .ZN(n4905) );
  NAND2_X1 U6541 ( .A1(n5563), .A2(n5562), .ZN(n5579) );
  NAND2_X1 U6542 ( .A1(n5281), .A2(n5280), .ZN(n5476) );
  NAND2_X1 U6543 ( .A1(n5281), .A2(n4911), .ZN(n4910) );
  NAND2_X1 U6544 ( .A1(n8794), .A2(n4924), .ZN(n4922) );
  OAI21_X2 U6545 ( .B1(n6512), .B2(n4928), .A(n4927), .ZN(n7476) );
  INV_X1 U6546 ( .A(n4930), .ZN(n4928) );
  INV_X1 U6547 ( .A(n8846), .ZN(n4934) );
  NAND2_X1 U6548 ( .A1(n4931), .A2(n4932), .ZN(n6560) );
  NAND2_X1 U6549 ( .A1(n8846), .A2(n4398), .ZN(n4931) );
  INV_X1 U6550 ( .A(n8845), .ZN(n4935) );
  NAND2_X1 U6551 ( .A1(n5984), .A2(n4938), .ZN(n6123) );
  NAND2_X1 U6552 ( .A1(n5984), .A2(n4937), .ZN(n4936) );
  NAND2_X1 U6553 ( .A1(n8855), .A2(n6585), .ZN(n4946) );
  NAND2_X1 U6554 ( .A1(n8855), .A2(n4940), .ZN(n4939) );
  NOR2_X1 U6555 ( .A1(n6586), .A2(n6587), .ZN(n4945) );
  NOR2_X1 U6556 ( .A1(n7609), .A2(n5061), .ZN(n7783) );
  INV_X1 U6557 ( .A(n4954), .ZN(n8838) );
  INV_X1 U6558 ( .A(n4421), .ZN(n4964) );
  OR2_X4 U6559 ( .A1(n5083), .A2(n10220), .ZN(n5154) );
  XNOR2_X2 U6560 ( .A(n4972), .B(P1_IR_REG_30__SCAN_IN), .ZN(n10220) );
  NAND2_X2 U6561 ( .A1(n5652), .A2(n8470), .ZN(n10073) );
  AND2_X2 U6562 ( .A1(n9797), .A2(n5637), .ZN(n5652) );
  OAI21_X2 U6563 ( .B1(n9915), .B2(n5505), .A(n5506), .ZN(n9890) );
  OAI21_X1 U6564 ( .B1(n9929), .B2(n4988), .A(n4986), .ZN(n4991) );
  INV_X1 U6565 ( .A(n4991), .ZN(n9892) );
  NAND2_X1 U6566 ( .A1(n9863), .A2(n4996), .ZN(n4995) );
  NAND2_X1 U6567 ( .A1(n6224), .A2(n5019), .ZN(n5016) );
  NAND2_X1 U6568 ( .A1(n5016), .A2(n5017), .ZN(n6257) );
  AND2_X2 U6569 ( .A1(n5022), .A2(n5777), .ZN(n5831) );
  NAND3_X1 U6570 ( .A1(n5022), .A2(n5777), .A3(P2_REG3_REG_1__SCAN_IN), .ZN(
        n5812) );
  XNOR2_X2 U6571 ( .A(n5776), .B(n5775), .ZN(n5778) );
  NAND2_X1 U6572 ( .A1(n4415), .A2(n7796), .ZN(n5031) );
  INV_X1 U6573 ( .A(n5031), .ZN(n10049) );
  NOR2_X1 U6574 ( .A1(n9917), .A2(n10118), .ZN(n9901) );
  INV_X1 U6575 ( .A(n10020), .ZN(n5042) );
  NAND3_X1 U6576 ( .A1(n5042), .A2(n9955), .A3(n5041), .ZN(n9949) );
  INV_X1 U6577 ( .A(n5045), .ZN(n10003) );
  OR2_X1 U6578 ( .A1(n6488), .A2(n10353), .ZN(n10329) );
  XNOR2_X1 U6579 ( .A(n5049), .B(n9821), .ZN(n9812) );
  NAND2_X2 U6580 ( .A1(n5751), .A2(n5750), .ZN(n5799) );
  NAND2_X1 U6581 ( .A1(n6208), .A2(n5772), .ZN(n5751) );
  XOR2_X1 U6582 ( .A(n9369), .B(n9099), .Z(n9371) );
  NAND2_X1 U6583 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  OR2_X1 U6584 ( .A1(n9538), .A2(n9539), .ZN(n9623) );
  NOR2_X1 U6585 ( .A1(n5786), .A2(n4439), .ZN(n5788) );
  AND2_X4 U6586 ( .A1(n6904), .A2(n7358), .ZN(n6863) );
  XNOR2_X1 U6587 ( .A(n5561), .B(n5560), .ZN(n8240) );
  XNOR2_X1 U6588 ( .A(n5618), .B(n5617), .ZN(n8438) );
  NAND2_X1 U6589 ( .A1(n5752), .A2(n6985), .ZN(n5141) );
  NAND2_X1 U6590 ( .A1(n8733), .A2(n6621), .ZN(n6637) );
  INV_X1 U6591 ( .A(n9382), .ZN(n6218) );
  INV_X1 U6592 ( .A(n6123), .ZN(n6129) );
  OAI21_X1 U6593 ( .B1(n10087), .B2(n10062), .A(n5733), .ZN(n5734) );
  NAND2_X1 U6594 ( .A1(n9855), .A2(n9839), .ZN(n9833) );
  INV_X1 U6595 ( .A(n7737), .ZN(n6184) );
  OR2_X1 U6596 ( .A1(n5432), .A2(n5132), .ZN(n5134) );
  OR2_X1 U6597 ( .A1(n5611), .A2(n5082), .ZN(n5085) );
  NAND2_X1 U6598 ( .A1(n7693), .A2(n7694), .ZN(n7692) );
  NAND2_X1 U6599 ( .A1(n9676), .A2(n7179), .ZN(n7249) );
  XNOR2_X1 U6600 ( .A(n9785), .B(n9784), .ZN(n9789) );
  AOI22_X2 U6601 ( .A1(n9200), .A2(n9205), .B1(n8773), .B2(n4787), .ZN(n9185)
         );
  INV_X2 U6602 ( .A(n10335), .ZN(n10337) );
  OR2_X1 U6603 ( .A1(n8717), .A2(n4391), .ZN(n10014) );
  AND2_X1 U6604 ( .A1(n6220), .A2(n6219), .ZN(n5046) );
  AND2_X1 U6605 ( .A1(n9386), .A2(n5056), .ZN(n5047) );
  OR2_X1 U6606 ( .A1(n9827), .A2(n9828), .ZN(n5048) );
  OR2_X1 U6607 ( .A1(n9806), .A2(n9805), .ZN(n5049) );
  OR2_X1 U6608 ( .A1(n6222), .A2(n4809), .ZN(n5050) );
  AND3_X1 U6609 ( .A1(n6484), .A2(n6485), .A3(n7032), .ZN(n5051) );
  NOR3_X1 U6610 ( .A1(n10076), .A2(n10163), .A3(n10075), .ZN(n5053) );
  AND2_X1 U6611 ( .A1(n10124), .A2(n9543), .ZN(n8505) );
  AND2_X1 U6612 ( .A1(n5300), .A2(n5276), .ZN(n5054) );
  AND2_X1 U6613 ( .A1(n5425), .A2(n5411), .ZN(n5055) );
  INV_X1 U6614 ( .A(n7829), .ZN(n5907) );
  NAND2_X1 U6615 ( .A1(n5721), .A2(n4391), .ZN(n10017) );
  INV_X1 U6616 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5748) );
  AND2_X1 U6617 ( .A1(n9385), .A2(n10393), .ZN(n5056) );
  AOI21_X1 U6618 ( .B1(n9105), .B2(n5831), .A(n6108), .ZN(n9115) );
  NOR2_X1 U6619 ( .A1(n5772), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5057) );
  INV_X1 U6620 ( .A(n8229), .ZN(n6172) );
  OR2_X1 U6621 ( .A1(n6418), .A2(n4583), .ZN(n5058) );
  AND2_X1 U6622 ( .A1(n7029), .A2(n7222), .ZN(n10317) );
  INV_X1 U6623 ( .A(n10317), .ZN(n6215) );
  INV_X4 U6624 ( .A(n6496), .ZN(n7656) );
  NOR2_X1 U6625 ( .A1(n6733), .A2(n7906), .ZN(n5059) );
  AND2_X1 U6626 ( .A1(n6529), .A2(n6528), .ZN(n5061) );
  AND2_X1 U6627 ( .A1(n6199), .A2(n9242), .ZN(n5062) );
  INV_X1 U6628 ( .A(n5827), .ZN(n10320) );
  NAND2_X1 U6629 ( .A1(n10179), .A2(n7849), .ZN(n5063) );
  INV_X1 U6630 ( .A(n10179), .ZN(n5726) );
  OR2_X1 U6631 ( .A1(n10088), .A2(n10028), .ZN(n5064) );
  INV_X1 U6632 ( .A(n10039), .ZN(n5705) );
  AND2_X1 U6633 ( .A1(n6404), .A2(n6398), .ZN(n6384) );
  AND2_X1 U6634 ( .A1(n9180), .A2(n6389), .ZN(n6390) );
  AND2_X1 U6635 ( .A1(n6459), .A2(n5058), .ZN(n6419) );
  INV_X1 U6636 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5075) );
  AND2_X1 U6637 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5759) );
  NAND2_X1 U6638 ( .A1(n8710), .A2(n8709), .ZN(n8711) );
  INV_X1 U6639 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6640 ( .A1(n8805), .A2(n6557), .ZN(n6558) );
  OR2_X1 U6641 ( .A1(n10338), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6159) );
  INV_X1 U6642 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5286) );
  AND2_X1 U6643 ( .A1(n10109), .A2(n9852), .ZN(n8682) );
  NOR2_X1 U6644 ( .A1(n5053), .A2(n10079), .ZN(n10080) );
  INV_X1 U6645 ( .A(n8537), .ZN(n8649) );
  AND2_X1 U6646 ( .A1(n8617), .A2(n8613), .ZN(n8642) );
  INV_X1 U6647 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5071) );
  INV_X1 U6648 ( .A(SI_20_), .ZN(n7963) );
  INV_X1 U6649 ( .A(n5375), .ZN(n5380) );
  INV_X1 U6650 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6651 ( .A1(n6163), .A2(n6162), .ZN(n6130) );
  AND2_X1 U6652 ( .A1(n6503), .A2(n7484), .ZN(n6498) );
  INV_X1 U6653 ( .A(n6493), .ZN(n7340) );
  OR2_X1 U6654 ( .A1(n6071), .A2(n6070), .ZN(n6083) );
  NAND2_X1 U6655 ( .A1(n6057), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6071) );
  INV_X1 U6656 ( .A(n7825), .ZN(n7934) );
  OR2_X1 U6657 ( .A1(n10338), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6143) );
  INV_X1 U6658 ( .A(n9786), .ZN(n9768) );
  INV_X1 U6659 ( .A(n7396), .ZN(n6682) );
  INV_X1 U6660 ( .A(n5206), .ZN(n5204) );
  INV_X1 U6661 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5102) );
  INV_X1 U6662 ( .A(n9994), .ZN(n5400) );
  NAND2_X1 U6663 ( .A1(n8726), .A2(n4560), .ZN(n8717) );
  INV_X1 U6664 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6665 ( .A1(n5385), .A2(n5384), .ZN(n5407) );
  NAND2_X1 U6666 ( .A1(n6130), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6145) );
  INV_X1 U6667 ( .A(n9334), .ZN(n8850) );
  INV_X1 U6668 ( .A(n8903), .ZN(n8863) );
  INV_X1 U6669 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7784) );
  AND2_X1 U6670 ( .A1(n6623), .A2(n6629), .ZN(n6166) );
  INV_X1 U6671 ( .A(n7189), .ZN(n6673) );
  AND2_X1 U6672 ( .A1(n9568), .A2(n9567), .ZN(n9648) );
  OR2_X1 U6673 ( .A1(n9793), .A2(n5631), .ZN(n5636) );
  OR2_X1 U6674 ( .A1(n5631), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5140) );
  AOI22_X1 U6675 ( .A1(n9786), .A2(n10043), .B1(n10041), .B2(n9829), .ZN(n9787) );
  NAND2_X1 U6676 ( .A1(n10106), .A2(n9562), .ZN(n8594) );
  AND2_X1 U6677 ( .A1(n5711), .A2(n8671), .ZN(n9913) );
  INV_X1 U6678 ( .A(n10287), .ZN(n10181) );
  INV_X1 U6679 ( .A(n7368), .ZN(n10282) );
  XNOR2_X1 U6680 ( .A(n5524), .B(SI_21_), .ZN(n5523) );
  XNOR2_X1 U6681 ( .A(n5466), .B(SI_18_), .ZN(n5464) );
  XNOR2_X1 U6682 ( .A(n5382), .B(SI_14_), .ZN(n5377) );
  NAND2_X1 U6683 ( .A1(n6145), .A2(n6144), .ZN(n6147) );
  AND2_X1 U6684 ( .A1(n6631), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8902) );
  AOI21_X1 U6685 ( .B1(n6474), .B2(n5051), .A(n6473), .ZN(n6475) );
  OR2_X1 U6686 ( .A1(n9169), .A2(n6073), .ZN(n6065) );
  AND4_X1 U6687 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n5958), .ZN(n8743)
         );
  INV_X1 U6688 ( .A(n9094), .ZN(n9051) );
  AND2_X1 U6689 ( .A1(n7213), .A2(n7212), .ZN(n9088) );
  INV_X1 U6690 ( .A(n9090), .ZN(n9077) );
  INV_X1 U6691 ( .A(n9312), .ZN(n10316) );
  INV_X1 U6692 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6238) );
  INV_X1 U6693 ( .A(n10396), .ZN(n10390) );
  OR2_X1 U6694 ( .A1(n6168), .A2(n6167), .ZN(n10402) );
  OR3_X1 U6695 ( .A1(n6236), .A2(n6607), .A3(n6235), .ZN(n6479) );
  AND2_X1 U6696 ( .A1(n5636), .A2(n5635), .ZN(n9641) );
  OR2_X1 U6697 ( .A1(n5631), .A2(n5178), .ZN(n5183) );
  INV_X1 U6698 ( .A(n10245), .ZN(n9733) );
  INV_X1 U6699 ( .A(n9787), .ZN(n9788) );
  NAND2_X1 U6700 ( .A1(n10292), .A2(n5698), .ZN(n9898) );
  OR2_X1 U6701 ( .A1(n7054), .A2(n5727), .ZN(n10287) );
  AND2_X1 U6702 ( .A1(n10000), .A2(n10186), .ZN(n10163) );
  INV_X1 U6703 ( .A(n10292), .ZN(n10186) );
  AND2_X1 U6704 ( .A1(n8702), .A2(n4392), .ZN(n10292) );
  AND2_X1 U6705 ( .A1(n5683), .A2(n5682), .ZN(n10212) );
  AND2_X1 U6706 ( .A1(n5241), .A2(n5260), .ZN(n7014) );
  OAI21_X1 U6707 ( .B1(n8454), .B2(n6990), .A(n5143), .ZN(n5130) );
  INV_X1 U6708 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8345) );
  INV_X1 U6709 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n8354) );
  NOR2_X1 U6710 ( .A1(n6903), .A2(P2_U3152), .ZN(n7207) );
  INV_X1 U6711 ( .A(n9432), .ZN(n9270) );
  INV_X1 U6712 ( .A(n8908), .ZN(n8897) );
  NAND2_X1 U6713 ( .A1(n6096), .A2(n6095), .ZN(n8915) );
  INV_X1 U6714 ( .A(n9313), .ZN(n9280) );
  NAND2_X1 U6715 ( .A1(n7224), .A2(n7223), .ZN(n9094) );
  INV_X1 U6716 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n9098) );
  INV_X1 U6717 ( .A(n9196), .ZN(n9366) );
  OR2_X1 U6718 ( .A1(n6479), .A2(n6237), .ZN(n10420) );
  INV_X2 U6719 ( .A(n10420), .ZN(n10423) );
  OR2_X1 U6720 ( .A1(n6479), .A2(n6478), .ZN(n10405) );
  NAND2_X1 U6721 ( .A1(n10339), .A2(n10338), .ZN(n10346) );
  INV_X1 U6722 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8243) );
  INV_X1 U6723 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7153) );
  INV_X1 U6724 ( .A(n9660), .ZN(n9629) );
  INV_X1 U6725 ( .A(n9650), .ZN(n9636) );
  INV_X1 U6726 ( .A(n9852), .ZN(n9877) );
  INV_X1 U6727 ( .A(n9653), .ZN(n9998) );
  OR2_X1 U6728 ( .A1(n6972), .A2(n4391), .ZN(n9746) );
  OR2_X1 U6729 ( .A1(n10243), .A2(n10239), .ZN(n9745) );
  INV_X1 U6730 ( .A(n5734), .ZN(n5735) );
  INV_X1 U6731 ( .A(n10308), .ZN(n10306) );
  INV_X1 U6732 ( .A(n10301), .ZN(n10299) );
  NOR2_X1 U6733 ( .A1(n10213), .A2(n10212), .ZN(n10265) );
  AND2_X1 U6734 ( .A1(n6904), .A2(n5680), .ZN(n6979) );
  INV_X1 U6735 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7156) );
  INV_X1 U6736 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8199) );
  OAI21_X1 U6737 ( .B1(n8355), .B2(n8354), .A(n8353), .ZN(n10472) );
  NOR2_X1 U6738 ( .A1(n10452), .A2(n10451), .ZN(n10450) );
  AND2_X2 U6739 ( .A1(n7207), .A2(n10345), .ZN(P2_U3966) );
  NAND2_X1 U6740 ( .A1(n5064), .A2(n5735), .ZN(P1_U3263) );
  NOR2_X1 U6741 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5067) );
  NAND2_X1 U6742 ( .A1(n5070), .A2(n5069), .ZN(n5471) );
  NAND3_X1 U6743 ( .A1(n5072), .A2(n5678), .A3(n5071), .ZN(n5665) );
  NAND2_X1 U6744 ( .A1(n5074), .A2(n5073), .ZN(n5470) );
  NAND3_X1 U6745 ( .A1(n5472), .A2(n5673), .A3(n5075), .ZN(n5076) );
  NAND2_X1 U6746 ( .A1(n5078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6747 ( .A1(n10223), .A2(n10220), .ZN(n5174) );
  INV_X1 U6748 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5086) );
  INV_X1 U6749 ( .A(n10220), .ZN(n5081) );
  INV_X1 U6750 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5082) );
  INV_X1 U6751 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6642) );
  INV_X1 U6752 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8211) );
  INV_X1 U6753 ( .A(n5088), .ZN(n5092) );
  INV_X1 U6754 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5093) );
  NAND3_X1 U6755 ( .A1(n5093), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5094) );
  NAND2_X4 U6756 ( .A1(n5095), .A2(n5094), .ZN(n5752) );
  NAND2_X1 U6757 ( .A1(n5752), .A2(SI_0_), .ZN(n5097) );
  INV_X1 U6758 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6759 ( .A1(n5097), .A2(n5096), .ZN(n5099) );
  NAND2_X1 U6760 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5122) );
  INV_X1 U6761 ( .A(n5122), .ZN(n5098) );
  NAND2_X1 U6762 ( .A1(n5752), .A2(n5098), .ZN(n5105) );
  NAND2_X1 U6763 ( .A1(n5099), .A2(n5105), .ZN(n10234) );
  NAND2_X1 U6764 ( .A1(n7249), .A2(n7051), .ZN(n5113) );
  INV_X2 U6765 ( .A(n5752), .ZN(n6986) );
  NAND2_X1 U6766 ( .A1(n5326), .A2(n4394), .ZN(n5166) );
  NAND2_X1 U6767 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5126) );
  INV_X1 U6768 ( .A(n5126), .ZN(n5104) );
  NAND2_X1 U6769 ( .A1(n6986), .A2(n5104), .ZN(n5825) );
  NAND2_X1 U6770 ( .A1(n5105), .A2(n5825), .ZN(n5107) );
  INV_X1 U6771 ( .A(SI_1_), .ZN(n5106) );
  XNOR2_X1 U6772 ( .A(n5107), .B(n5106), .ZN(n5109) );
  MUX2_X1 U6773 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5752), .Z(n5108) );
  OAI211_X2 U6774 ( .C1(n5166), .C2(n7017), .A(n5112), .B(n5111), .ZN(n7368)
         );
  NAND2_X1 U6775 ( .A1(n5113), .A2(n7368), .ZN(n5114) );
  OAI21_X1 U6776 ( .B1(n7051), .B2(n7249), .A(n5114), .ZN(n5136) );
  NAND2_X1 U6777 ( .A1(n5179), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5119) );
  INV_X1 U6778 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6779 ( .A1(n5156), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5116) );
  AND4_X2 U6780 ( .A1(n5119), .A2(n5118), .A3(n5117), .A4(n5116), .ZN(n7173)
         );
  INV_X1 U6781 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7018) );
  NAND2_X1 U6782 ( .A1(n5122), .A2(n7018), .ZN(n5120) );
  NAND2_X1 U6783 ( .A1(n5120), .A2(SI_1_), .ZN(n5121) );
  OAI21_X1 U6784 ( .B1(n7018), .B2(n5122), .A(n5121), .ZN(n5123) );
  NAND2_X1 U6785 ( .A1(n5752), .A2(n5123), .ZN(n5129) );
  INV_X1 U6786 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7010) );
  NAND2_X1 U6787 ( .A1(n5126), .A2(n7010), .ZN(n5124) );
  NAND2_X1 U6788 ( .A1(n5124), .A2(SI_1_), .ZN(n5125) );
  OAI21_X1 U6789 ( .B1(n5126), .B2(n7010), .A(n5125), .ZN(n5127) );
  NAND2_X1 U6790 ( .A1(n6986), .A2(n5127), .ZN(n5128) );
  INV_X1 U6791 ( .A(SI_2_), .ZN(n5142) );
  NAND2_X1 U6792 ( .A1(n5752), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5143) );
  INV_X1 U6793 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6794 ( .A1(n5170), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5148) );
  XNOR2_X1 U6795 ( .A(n5148), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U6796 ( .A1(n5479), .A2(n6983), .ZN(n5133) );
  NAND2_X1 U6797 ( .A1(n7173), .A2(n7424), .ZN(n5135) );
  NAND2_X1 U6798 ( .A1(n5179), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6799 ( .A1(n5090), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6800 ( .A1(n8456), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5137) );
  INV_X1 U6801 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7009) );
  INV_X1 U6802 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6985) );
  INV_X1 U6803 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6990) );
  OAI211_X1 U6804 ( .C1(n5752), .C2(n6990), .A(n5143), .B(n5142), .ZN(n5144)
         );
  NAND2_X1 U6805 ( .A1(n5752), .A2(n5132), .ZN(n5145) );
  OAI211_X1 U6806 ( .C1(n5752), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5145), .B(
        SI_2_), .ZN(n5146) );
  NAND2_X1 U6807 ( .A1(n5147), .A2(n5146), .ZN(n5160) );
  XNOR2_X1 U6808 ( .A(n5161), .B(n5160), .ZN(n7008) );
  INV_X1 U6809 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6810 ( .A1(n5148), .A2(n5168), .ZN(n5149) );
  NAND2_X1 U6811 ( .A1(n5149), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6812 ( .A1(n5479), .A2(n6984), .ZN(n5152) );
  NAND2_X1 U6813 ( .A1(n9675), .A2(n10286), .ZN(n8513) );
  NAND2_X1 U6814 ( .A1(n7445), .A2(n7176), .ZN(n8518) );
  NAND2_X1 U6815 ( .A1(n7409), .A2(n7408), .ZN(n7407) );
  NAND2_X1 U6816 ( .A1(n7445), .A2(n10286), .ZN(n5153) );
  NAND2_X1 U6817 ( .A1(n7407), .A2(n5153), .ZN(n7444) );
  INV_X1 U6818 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5155) );
  XNOR2_X1 U6819 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7453) );
  OAI22_X1 U6820 ( .A1(n5154), .A2(n5155), .B1(n5631), .B2(n7453), .ZN(n5159)
         );
  INV_X1 U6821 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7451) );
  INV_X1 U6822 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5157) );
  OAI22_X1 U6823 ( .A1(n5716), .A2(n7451), .B1(n5611), .B2(n5157), .ZN(n5158)
         );
  NAND2_X1 U6824 ( .A1(n5161), .A2(n5160), .ZN(n5165) );
  INV_X1 U6825 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6826 ( .A1(n5163), .A2(SI_3_), .ZN(n5164) );
  INV_X1 U6827 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6988) );
  INV_X1 U6828 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6982) );
  MUX2_X1 U6829 ( .A(n6988), .B(n6982), .S(n5752), .Z(n5186) );
  XNOR2_X1 U6830 ( .A(n5186), .B(SI_4_), .ZN(n5184) );
  XNOR2_X1 U6831 ( .A(n5185), .B(n4390), .ZN(n6980) );
  NAND2_X1 U6832 ( .A1(n6980), .A2(n5218), .ZN(n5173) );
  NAND2_X1 U6833 ( .A1(n5168), .A2(n5167), .ZN(n5169) );
  OAI21_X1 U6834 ( .B1(n5170), .B2(n5169), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5171) );
  XNOR2_X1 U6835 ( .A(n5171), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9688) );
  AOI22_X1 U6836 ( .A1(n8466), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n5479), .B2(
        n9688), .ZN(n5172) );
  NOR2_X1 U6837 ( .A1(n9674), .A2(n7454), .ZN(n8519) );
  NAND2_X1 U6838 ( .A1(n9674), .A2(n7454), .ZN(n8514) );
  NAND2_X1 U6839 ( .A1(n8574), .A2(n8514), .ZN(n8477) );
  INV_X1 U6840 ( .A(n9674), .ZN(n7397) );
  NAND2_X1 U6841 ( .A1(n7397), .A2(n7454), .ZN(n7506) );
  INV_X1 U6842 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6843 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5175) );
  NAND2_X1 U6844 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  AND2_X1 U6845 ( .A1(n5206), .A2(n5177), .ZN(n7516) );
  INV_X1 U6846 ( .A(n7516), .ZN(n5178) );
  NAND2_X1 U6847 ( .A1(n8457), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6848 ( .A1(n7002), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6849 ( .A1(n8456), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5180) );
  INV_X1 U6850 ( .A(n5186), .ZN(n5187) );
  NAND2_X1 U6851 ( .A1(n5187), .A2(SI_4_), .ZN(n5188) );
  MUX2_X1 U6852 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5752), .Z(n5198) );
  XNOR2_X1 U6853 ( .A(n5198), .B(SI_5_), .ZN(n5195) );
  XNOR2_X1 U6854 ( .A(n5197), .B(n5195), .ZN(n6989) );
  NAND2_X1 U6855 ( .A1(n6989), .A2(n5218), .ZN(n5194) );
  NAND2_X1 U6856 ( .A1(n5190), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5189) );
  MUX2_X1 U6857 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5189), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5192) );
  NOR2_X2 U6858 ( .A1(n5190), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5220) );
  INV_X1 U6859 ( .A(n5220), .ZN(n5191) );
  AOI22_X1 U6860 ( .A1(n8466), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5479), .B2(
        n9697), .ZN(n5193) );
  NAND2_X1 U6861 ( .A1(n7461), .A2(n7553), .ZN(n8575) );
  NAND2_X1 U6862 ( .A1(n6679), .A2(n9673), .ZN(n8516) );
  NAND2_X1 U6863 ( .A1(n8575), .A2(n8516), .ZN(n8478) );
  INV_X1 U6864 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U6865 ( .A1(n5198), .A2(SI_5_), .ZN(n5199) );
  XNOR2_X1 U6866 ( .A(n5213), .B(n5212), .ZN(n6992) );
  NAND2_X1 U6867 ( .A1(n6992), .A2(n8464), .ZN(n5203) );
  OR2_X1 U6868 ( .A1(n5220), .A2(n10215), .ZN(n5201) );
  XNOR2_X1 U6869 ( .A(n5201), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6993) );
  AOI22_X1 U6870 ( .A1(n8466), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5479), .B2(
        n6993), .ZN(n5202) );
  NAND2_X1 U6871 ( .A1(n5203), .A2(n5202), .ZN(n7758) );
  NAND2_X1 U6872 ( .A1(n8457), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5211) );
  INV_X1 U6873 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6874 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  AND2_X1 U6875 ( .A1(n5225), .A2(n5207), .ZN(n7757) );
  NAND2_X1 U6876 ( .A1(n5718), .A2(n7757), .ZN(n5210) );
  NAND2_X1 U6877 ( .A1(n7002), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6878 ( .A1(n7001), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5208) );
  OR2_X1 U6879 ( .A1(n7758), .A2(n7632), .ZN(n8604) );
  INV_X1 U6880 ( .A(n8578), .ZN(n8606) );
  NAND2_X1 U6881 ( .A1(n8604), .A2(n8606), .ZN(n8479) );
  NAND2_X1 U6882 ( .A1(n7553), .A2(n9673), .ZN(n7590) );
  INV_X1 U6883 ( .A(n5212), .ZN(n5214) );
  NAND2_X1 U6884 ( .A1(n5215), .A2(SI_6_), .ZN(n5216) );
  MUX2_X1 U6885 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8454), .Z(n5233) );
  XNOR2_X1 U6886 ( .A(n5233), .B(SI_7_), .ZN(n5231) );
  NAND2_X1 U6887 ( .A1(n6995), .A2(n8464), .ZN(n5222) );
  OR2_X1 U6888 ( .A1(n5281), .A2(n10215), .ZN(n5238) );
  XNOR2_X1 U6889 ( .A(n5238), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7064) );
  AOI22_X1 U6890 ( .A1(n8466), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5479), .B2(
        n7064), .ZN(n5221) );
  INV_X1 U6891 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6892 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  AND2_X1 U6893 ( .A1(n5246), .A2(n5226), .ZN(n7639) );
  NAND2_X1 U6894 ( .A1(n8457), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6895 ( .A1(n7002), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6896 ( .A1(n8456), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5227) );
  OR2_X1 U6897 ( .A1(n7640), .A2(n7649), .ZN(n8609) );
  NAND2_X1 U6898 ( .A1(n7640), .A2(n7649), .ZN(n8607) );
  NAND2_X1 U6899 ( .A1(n8609), .A2(n8607), .ZN(n7634) );
  INV_X1 U6900 ( .A(n7634), .ZN(n8482) );
  INV_X1 U6901 ( .A(n7632), .ZN(n9672) );
  NOR2_X1 U6902 ( .A1(n7758), .A2(n9672), .ZN(n7574) );
  NOR2_X1 U6903 ( .A1(n7640), .A2(n9671), .ZN(n7576) );
  AOI21_X1 U6904 ( .B1(n7574), .B2(n7634), .A(n7576), .ZN(n5252) );
  INV_X1 U6905 ( .A(n5231), .ZN(n5232) );
  NAND2_X1 U6906 ( .A1(n5233), .A2(SI_7_), .ZN(n5234) );
  INV_X1 U6907 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7000) );
  INV_X1 U6908 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7016) );
  MUX2_X1 U6909 ( .A(n7000), .B(n7016), .S(n8454), .Z(n5235) );
  INV_X1 U6910 ( .A(SI_8_), .ZN(n8198) );
  INV_X1 U6911 ( .A(n5235), .ZN(n5236) );
  NAND2_X1 U6912 ( .A1(n5236), .A2(SI_8_), .ZN(n5237) );
  AOI21_X1 U6913 ( .B1(n5238), .B2(n5279), .A(n10215), .ZN(n5239) );
  NAND2_X1 U6914 ( .A1(n5239), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5241) );
  INV_X1 U6915 ( .A(n5239), .ZN(n5240) );
  NAND2_X1 U6916 ( .A1(n5240), .A2(n5278), .ZN(n5260) );
  AOI22_X1 U6917 ( .A1(n8466), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7014), .B2(
        n5479), .ZN(n5242) );
  INV_X1 U6918 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6919 ( .A1(n5246), .A2(n5245), .ZN(n5247) );
  AND2_X1 U6920 ( .A1(n5263), .A2(n5247), .ZN(n7652) );
  NAND2_X1 U6921 ( .A1(n5718), .A2(n7652), .ZN(n5251) );
  NAND2_X1 U6922 ( .A1(n8457), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6923 ( .A1(n7002), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6924 ( .A1(n7001), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5248) );
  OR2_X1 U6925 ( .A1(n10179), .A2(n7849), .ZN(n8612) );
  NAND2_X1 U6926 ( .A1(n8612), .A2(n5063), .ZN(n7573) );
  NAND2_X1 U6927 ( .A1(n10179), .A2(n9670), .ZN(n5254) );
  INV_X1 U6928 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5257) );
  INV_X1 U6929 ( .A(SI_9_), .ZN(n5258) );
  NAND2_X1 U6930 ( .A1(n5259), .A2(SI_9_), .ZN(n5298) );
  AND2_X1 U6931 ( .A1(n5294), .A2(n5298), .ZN(n5271) );
  NAND2_X1 U6932 ( .A1(n5260), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5261) );
  XNOR2_X1 U6933 ( .A(n5261), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7021) );
  AOI22_X1 U6934 ( .A1(n7021), .A2(n5479), .B1(n8466), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6935 ( .A1(n5263), .A2(n8150), .ZN(n5264) );
  AND2_X1 U6936 ( .A1(n5287), .A2(n5264), .ZN(n7853) );
  NAND2_X1 U6937 ( .A1(n5718), .A2(n7853), .ZN(n5268) );
  NAND2_X1 U6938 ( .A1(n5179), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6939 ( .A1(n7002), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6940 ( .A1(n8456), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5265) );
  AND2_X1 U6941 ( .A1(n10174), .A2(n9669), .ZN(n5270) );
  OR2_X1 U6942 ( .A1(n10174), .A2(n9669), .ZN(n5269) );
  MUX2_X1 U6943 ( .A(n7034), .B(n8199), .S(n4394), .Z(n5274) );
  INV_X1 U6944 ( .A(SI_10_), .ZN(n5273) );
  INV_X1 U6945 ( .A(n5274), .ZN(n5275) );
  NAND2_X1 U6946 ( .A1(n5275), .A2(SI_10_), .ZN(n5276) );
  NAND2_X1 U6947 ( .A1(n7026), .A2(n8464), .ZN(n5285) );
  NAND2_X1 U6948 ( .A1(n5476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5282) );
  MUX2_X1 U6949 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5282), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5283) );
  AOI22_X1 U6950 ( .A1(n8466), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5479), .B2(
        n6950), .ZN(n5284) );
  OR2_X2 U6951 ( .A1(n5287), .A2(n5286), .ZN(n5308) );
  NAND2_X1 U6952 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  AND2_X1 U6953 ( .A1(n5308), .A2(n5288), .ZN(n8398) );
  NAND2_X1 U6954 ( .A1(n5718), .A2(n8398), .ZN(n5292) );
  NAND2_X1 U6955 ( .A1(n8457), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6956 ( .A1(n7001), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6957 ( .A1(n7002), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6958 ( .A1(n8399), .A2(n8270), .ZN(n8617) );
  NAND2_X1 U6959 ( .A1(n8636), .A2(n8617), .ZN(n8472) );
  INV_X1 U6960 ( .A(n8270), .ZN(n9668) );
  NOR2_X1 U6961 ( .A1(n8399), .A2(n9668), .ZN(n5293) );
  AND2_X1 U6962 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  NAND3_X1 U6963 ( .A1(n5299), .A2(n5054), .A3(n5298), .ZN(n5301) );
  INV_X1 U6964 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5302) );
  MUX2_X1 U6965 ( .A(n5302), .B(n8178), .S(n4393), .Z(n5315) );
  NAND2_X1 U6966 ( .A1(n7024), .A2(n8464), .ZN(n5305) );
  NAND2_X1 U6967 ( .A1(n5323), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5303) );
  XNOR2_X1 U6968 ( .A(n5303), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7027) );
  AOI22_X1 U6969 ( .A1(n8466), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7027), .B2(
        n5479), .ZN(n5304) );
  NAND2_X1 U6970 ( .A1(n8457), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5313) );
  INV_X1 U6971 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6972 ( .A1(n5308), .A2(n5307), .ZN(n5309) );
  AND2_X1 U6973 ( .A1(n5331), .A2(n5309), .ZN(n8278) );
  NAND2_X1 U6974 ( .A1(n5718), .A2(n8278), .ZN(n5312) );
  NAND2_X1 U6975 ( .A1(n7002), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6976 ( .A1(n7001), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6977 ( .A1(n8411), .A2(n7948), .ZN(n8320) );
  NAND2_X1 U6978 ( .A1(n8527), .A2(n8320), .ZN(n8486) );
  NAND2_X1 U6979 ( .A1(n8267), .A2(n8486), .ZN(n8324) );
  NAND2_X1 U6980 ( .A1(n8411), .A2(n9667), .ZN(n8323) );
  INV_X1 U6981 ( .A(n5315), .ZN(n5316) );
  NAND2_X1 U6982 ( .A1(n5316), .A2(SI_11_), .ZN(n5317) );
  MUX2_X1 U6983 ( .A(n7059), .B(n7057), .S(n4393), .Z(n5320) );
  INV_X1 U6984 ( .A(SI_12_), .ZN(n5319) );
  INV_X1 U6985 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6986 ( .A1(n5321), .A2(SI_12_), .ZN(n5322) );
  XNOR2_X1 U6987 ( .A(n5337), .B(n5338), .ZN(n7056) );
  NAND2_X1 U6988 ( .A1(n7056), .A2(n8464), .ZN(n5329) );
  OR2_X1 U6989 ( .A1(n5361), .A2(n10215), .ZN(n5325) );
  INV_X1 U6990 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6991 ( .A1(n5325), .A2(n5324), .ZN(n5340) );
  OAI21_X1 U6992 ( .B1(n5325), .B2(n5324), .A(n5340), .ZN(n7543) );
  OAI22_X1 U6993 ( .A1(n7543), .A2(n5326), .B1(n5432), .B2(n7057), .ZN(n5327)
         );
  INV_X1 U6994 ( .A(n5327), .ZN(n5328) );
  INV_X1 U6995 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U6996 ( .A1(n5331), .A2(n8036), .ZN(n5332) );
  AND2_X1 U6997 ( .A1(n5345), .A2(n5332), .ZN(n8330) );
  NAND2_X1 U6998 ( .A1(n5718), .A2(n8330), .ZN(n5336) );
  NAND2_X1 U6999 ( .A1(n5179), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U7000 ( .A1(n7002), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U7001 ( .A1(n8456), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U7002 ( .A1(n10170), .A2(n10040), .ZN(n10033) );
  NAND3_X1 U7003 ( .A1(n8324), .A2(n8323), .A3(n10033), .ZN(n5352) );
  MUX2_X1 U7004 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4394), .Z(n5339) );
  NOR2_X1 U7005 ( .A1(n5339), .A2(SI_13_), .ZN(n5374) );
  INV_X1 U7006 ( .A(n5374), .ZN(n5357) );
  AND2_X1 U7007 ( .A1(n5375), .A2(n5357), .ZN(n5355) );
  NAND2_X1 U7008 ( .A1(n7125), .A2(n8464), .ZN(n5343) );
  NAND2_X1 U7009 ( .A1(n5340), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5341) );
  XNOR2_X1 U7010 ( .A(n5341), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7126) );
  AOI22_X1 U7011 ( .A1(n7126), .A2(n5479), .B1(n8466), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5342) );
  NAND2_X2 U7012 ( .A1(n5343), .A2(n5342), .ZN(n10164) );
  INV_X1 U7013 ( .A(n10164), .ZN(n10055) );
  NAND2_X1 U7014 ( .A1(n5345), .A2(n5344), .ZN(n5346) );
  AND2_X1 U7015 ( .A1(n5365), .A2(n5346), .ZN(n10052) );
  NAND2_X1 U7016 ( .A1(n5718), .A2(n10052), .ZN(n5350) );
  NAND2_X1 U7017 ( .A1(n5179), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U7018 ( .A1(n7001), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U7019 ( .A1(n7002), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U7020 ( .A1(n10170), .A2(n7909), .ZN(n8618) );
  AOI22_X1 U7021 ( .A1(n10055), .A2(n10015), .B1(n8489), .B2(n10033), .ZN(
        n5351) );
  NAND2_X1 U7022 ( .A1(n5352), .A2(n5351), .ZN(n5354) );
  INV_X1 U7023 ( .A(n10015), .ZN(n9666) );
  NAND2_X1 U7024 ( .A1(n10164), .A2(n9666), .ZN(n5353) );
  NAND2_X1 U7025 ( .A1(n5356), .A2(n5355), .ZN(n5358) );
  NAND2_X1 U7026 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  MUX2_X1 U7027 ( .A(n8140), .B(n7146), .S(n4393), .Z(n5382) );
  NAND2_X1 U7028 ( .A1(n7145), .A2(n8464), .ZN(n5364) );
  NOR2_X1 U7029 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5360) );
  OR2_X1 U7030 ( .A1(n5390), .A2(n10215), .ZN(n5362) );
  XNOR2_X1 U7031 ( .A(n5362), .B(P1_IR_REG_14__SCAN_IN), .ZN(n6963) );
  AOI22_X1 U7032 ( .A1(n6963), .A2(n5479), .B1(n8466), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5363) );
  NAND2_X2 U7033 ( .A1(n5364), .A2(n5363), .ZN(n10159) );
  INV_X1 U7034 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U7035 ( .A1(n5365), .A2(n8165), .ZN(n5366) );
  NAND2_X1 U7036 ( .A1(n5395), .A2(n5366), .ZN(n10022) );
  OR2_X1 U7037 ( .A1(n5631), .A2(n10022), .ZN(n5371) );
  NAND2_X1 U7038 ( .A1(n7001), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U7039 ( .A1(n7002), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5367) );
  AND2_X1 U7040 ( .A1(n5368), .A2(n5367), .ZN(n5370) );
  NAND2_X1 U7041 ( .A1(n8457), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5369) );
  OR2_X1 U7042 ( .A1(n10159), .A2(n10042), .ZN(n5372) );
  INV_X1 U7043 ( .A(n5373), .ZN(n5376) );
  AOI21_X1 U7044 ( .B1(n5376), .B2(n5375), .A(n5374), .ZN(n5378) );
  INV_X1 U7045 ( .A(n5382), .ZN(n5383) );
  NAND2_X1 U7046 ( .A1(n5383), .A2(SI_14_), .ZN(n5404) );
  NAND2_X1 U7047 ( .A1(n5406), .A2(n5404), .ZN(n5388) );
  MUX2_X1 U7048 ( .A(n7153), .B(n7156), .S(n4393), .Z(n5385) );
  INV_X1 U7049 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U7050 ( .A1(n5386), .A2(SI_15_), .ZN(n5387) );
  NAND2_X1 U7051 ( .A1(n5407), .A2(n5387), .ZN(n5402) );
  NAND2_X1 U7052 ( .A1(n7152), .A2(n8464), .ZN(n5393) );
  INV_X1 U7053 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U7054 ( .A1(n5390), .A2(n5389), .ZN(n5412) );
  NAND2_X1 U7055 ( .A1(n5412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5391) );
  XNOR2_X1 U7056 ( .A(n5391), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7154) );
  AOI22_X1 U7057 ( .A1(n7154), .A2(n5479), .B1(n8466), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5392) );
  INV_X1 U7058 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5394) );
  OR2_X2 U7059 ( .A1(n5395), .A2(n5394), .ZN(n5418) );
  NAND2_X1 U7060 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  AND2_X1 U7061 ( .A1(n5418), .A2(n5396), .ZN(n10004) );
  NAND2_X1 U7062 ( .A1(n10004), .A2(n5718), .ZN(n5399) );
  AOI22_X1 U7063 ( .A1(n8456), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7002), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U7064 ( .A1(n5179), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U7065 ( .A1(n10154), .A2(n9978), .ZN(n5401) );
  NAND2_X1 U7066 ( .A1(n9997), .A2(n5401), .ZN(n9987) );
  INV_X1 U7067 ( .A(n5402), .ZN(n5403) );
  MUX2_X1 U7068 ( .A(n8191), .B(n7185), .S(n4393), .Z(n5409) );
  INV_X1 U7069 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U7070 ( .A1(n5410), .A2(SI_16_), .ZN(n5411) );
  NAND2_X1 U7071 ( .A1(n7184), .A2(n8464), .ZN(n5415) );
  NAND2_X1 U7072 ( .A1(n5413), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5427) );
  XNOR2_X1 U7073 ( .A(n5427), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9711) );
  AOI22_X1 U7074 ( .A1(n9711), .A2(n5479), .B1(n8466), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5414) );
  INV_X1 U7075 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U7076 ( .A1(n5418), .A2(n5417), .ZN(n5419) );
  NAND2_X1 U7077 ( .A1(n5436), .A2(n5419), .ZN(n9982) );
  OR2_X1 U7078 ( .A1(n9982), .A2(n5631), .ZN(n5422) );
  AOI22_X1 U7079 ( .A1(n8456), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7002), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U7080 ( .A1(n5179), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5420) );
  AND2_X2 U7081 ( .A1(n10149), .A2(n9653), .ZN(n8537) );
  NAND2_X1 U7082 ( .A1(n8650), .A2(n8649), .ZN(n9986) );
  NAND2_X1 U7083 ( .A1(n9987), .A2(n9986), .ZN(n9989) );
  NAND2_X1 U7084 ( .A1(n10149), .A2(n9998), .ZN(n5423) );
  MUX2_X1 U7085 ( .A(n7243), .B(n8034), .S(n4394), .Z(n5447) );
  XNOR2_X1 U7086 ( .A(n5450), .B(n5446), .ZN(n7205) );
  NAND2_X1 U7087 ( .A1(n7205), .A2(n8464), .ZN(n5435) );
  INV_X1 U7088 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U7089 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  NAND2_X1 U7090 ( .A1(n5428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5430) );
  INV_X1 U7091 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U7092 ( .A1(n5430), .A2(n5429), .ZN(n5451) );
  OR2_X1 U7093 ( .A1(n5430), .A2(n5429), .ZN(n5431) );
  NOR2_X1 U7094 ( .A1(n5432), .A2(n8034), .ZN(n5433) );
  AOI21_X1 U7095 ( .B1(n9728), .B2(n5479), .A(n5433), .ZN(n5434) );
  INV_X1 U7096 ( .A(n5455), .ZN(n5457) );
  NAND2_X1 U7097 ( .A1(n5436), .A2(n4567), .ZN(n5437) );
  NAND2_X1 U7098 ( .A1(n9966), .A2(n5718), .ZN(n5443) );
  INV_X1 U7099 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U7100 ( .A1(n7002), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U7101 ( .A1(n8456), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5438) );
  OAI211_X1 U7102 ( .C1(n5440), .C2(n5154), .A(n5439), .B(n5438), .ZN(n5441)
         );
  INV_X1 U7103 ( .A(n5441), .ZN(n5442) );
  OR2_X1 U7104 ( .A1(n10144), .A2(n9979), .ZN(n5444) );
  NAND2_X1 U7105 ( .A1(n10144), .A2(n9979), .ZN(n5445) );
  INV_X1 U7106 ( .A(n5447), .ZN(n5448) );
  NAND2_X1 U7107 ( .A1(n5448), .A2(SI_17_), .ZN(n5449) );
  MUX2_X1 U7108 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4393), .Z(n5466) );
  NAND2_X1 U7109 ( .A1(n7351), .A2(n8464), .ZN(n5454) );
  NAND2_X1 U7110 ( .A1(n5451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5452) );
  XNOR2_X1 U7111 ( .A(n5452), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9739) );
  AOI22_X1 U7112 ( .A1(n9739), .A2(n5479), .B1(n8466), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5453) );
  INV_X1 U7113 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U7114 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  NAND2_X1 U7115 ( .A1(n5498), .A2(n5458), .ZN(n9952) );
  OR2_X1 U7116 ( .A1(n9952), .A2(n5631), .ZN(n5463) );
  INV_X1 U7117 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U7118 ( .A1(n7002), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U7119 ( .A1(n7001), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5459) );
  OAI211_X1 U7120 ( .C1(n9720), .C2(n5154), .A(n5460), .B(n5459), .ZN(n5461)
         );
  INV_X1 U7121 ( .A(n5461), .ZN(n5462) );
  OR2_X1 U7122 ( .A1(n10138), .A2(n9588), .ZN(n8655) );
  NAND2_X1 U7123 ( .A1(n10138), .A2(n9588), .ZN(n8540) );
  NAND2_X1 U7124 ( .A1(n8655), .A2(n8540), .ZN(n9956) );
  MUX2_X1 U7125 ( .A(n7403), .B(n7405), .S(n4394), .Z(n5467) );
  INV_X1 U7126 ( .A(n5467), .ZN(n5468) );
  NAND2_X1 U7127 ( .A1(n5468), .A2(SI_19_), .ZN(n5469) );
  NAND2_X1 U7128 ( .A1(n7402), .A2(n8464), .ZN(n5481) );
  AOI22_X1 U7129 ( .A1(n8502), .A2(n5479), .B1(n8466), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n5480) );
  XNOR2_X1 U7130 ( .A(n5498), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9935) );
  NAND2_X1 U7131 ( .A1(n9935), .A2(n5718), .ZN(n5486) );
  INV_X1 U7132 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9737) );
  NAND2_X1 U7133 ( .A1(n7002), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7134 ( .A1(n7001), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5482) );
  OAI211_X1 U7135 ( .C1(n5154), .C2(n9737), .A(n5483), .B(n5482), .ZN(n5484)
         );
  INV_X1 U7136 ( .A(n5484), .ZN(n5485) );
  MUX2_X1 U7137 ( .A(n7607), .B(n8161), .S(n4393), .Z(n5490) );
  INV_X1 U7138 ( .A(n5490), .ZN(n5491) );
  NAND2_X1 U7139 ( .A1(n5491), .A2(SI_20_), .ZN(n5492) );
  XNOR2_X1 U7140 ( .A(n5508), .B(n5507), .ZN(n7571) );
  NAND2_X1 U7141 ( .A1(n7571), .A2(n8464), .ZN(n5494) );
  NAND2_X1 U7142 ( .A1(n8466), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5493) );
  INV_X1 U7143 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5496) );
  INV_X1 U7144 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5495) );
  OAI21_X1 U7145 ( .B1(n5498), .B2(n5496), .A(n5495), .ZN(n5499) );
  NAND2_X1 U7146 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5497) );
  NAND2_X1 U7147 ( .A1(n5499), .A2(n5514), .ZN(n9918) );
  OR2_X1 U7148 ( .A1(n9918), .A2(n5631), .ZN(n5504) );
  INV_X1 U7149 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U7150 ( .A1(n8457), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7151 ( .A1(n8456), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5500) );
  OAI211_X1 U7152 ( .C1(n5611), .C2(n10200), .A(n5501), .B(n5500), .ZN(n5502)
         );
  INV_X1 U7153 ( .A(n5502), .ZN(n5503) );
  NOR2_X1 U7154 ( .A1(n10124), .A2(n9931), .ZN(n5505) );
  NAND2_X1 U7155 ( .A1(n10124), .A2(n9931), .ZN(n5506) );
  NAND2_X1 U7156 ( .A1(n5508), .A2(n5507), .ZN(n5510) );
  MUX2_X1 U7157 ( .A(n7770), .B(n7767), .S(n4394), .Z(n5524) );
  XNOR2_X1 U7158 ( .A(n5528), .B(n5523), .ZN(n7766) );
  NAND2_X1 U7159 ( .A1(n7766), .A2(n8464), .ZN(n5512) );
  NAND2_X1 U7160 ( .A1(n8466), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5511) );
  INV_X1 U7161 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7162 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  NAND2_X1 U7163 ( .A1(n5553), .A2(n5515), .ZN(n9899) );
  OR2_X1 U7164 ( .A1(n9899), .A2(n5631), .ZN(n5520) );
  INV_X1 U7165 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8104) );
  NAND2_X1 U7166 ( .A1(n5179), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7167 ( .A1(n7001), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5516) );
  OAI211_X1 U7168 ( .C1(n5611), .C2(n8104), .A(n5517), .B(n5516), .ZN(n5518)
         );
  INV_X1 U7169 ( .A(n5518), .ZN(n5519) );
  NAND2_X1 U7170 ( .A1(n10118), .A2(n9910), .ZN(n8673) );
  NAND2_X1 U7171 ( .A1(n10118), .A2(n9876), .ZN(n5521) );
  INV_X1 U7172 ( .A(n5524), .ZN(n5525) );
  MUX2_X1 U7173 ( .A(n8449), .B(n8443), .S(n4393), .Z(n5530) );
  INV_X1 U7174 ( .A(SI_22_), .ZN(n5529) );
  INV_X1 U7175 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7176 ( .A1(n5531), .A2(SI_22_), .ZN(n5532) );
  XNOR2_X1 U7177 ( .A(n5543), .B(n5542), .ZN(n8441) );
  NAND2_X1 U7178 ( .A1(n8441), .A2(n8464), .ZN(n5534) );
  NAND2_X1 U7179 ( .A1(n8466), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5533) );
  XNOR2_X1 U7180 ( .A(n5553), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U7181 ( .A1(n9881), .A2(n5718), .ZN(n5539) );
  INV_X1 U7182 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U7183 ( .A1(n5179), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7184 ( .A1(n7001), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5535) );
  OAI211_X1 U7185 ( .C1(n5611), .C2(n8180), .A(n5536), .B(n5535), .ZN(n5537)
         );
  INV_X1 U7186 ( .A(n5537), .ZN(n5538) );
  OR2_X1 U7187 ( .A1(n10113), .A2(n9894), .ZN(n5540) );
  INV_X1 U7188 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5544) );
  MUX2_X1 U7189 ( .A(n8243), .B(n5544), .S(n4394), .Z(n5546) );
  INV_X1 U7190 ( .A(SI_23_), .ZN(n5545) );
  NAND2_X1 U7191 ( .A1(n5546), .A2(n5545), .ZN(n5562) );
  INV_X1 U7192 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U7193 ( .A1(n5547), .A2(SI_23_), .ZN(n5548) );
  NAND2_X1 U7194 ( .A1(n8240), .A2(n8464), .ZN(n5550) );
  NAND2_X1 U7195 ( .A1(n8466), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5549) );
  INV_X1 U7196 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5552) );
  INV_X1 U7197 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5551) );
  OAI21_X1 U7198 ( .B1(n5553), .B2(n5552), .A(n5551), .ZN(n5554) );
  OR3_X2 U7199 ( .A1(n5553), .A2(n5552), .A3(n5551), .ZN(n5567) );
  AND2_X1 U7200 ( .A1(n5554), .A2(n5567), .ZN(n9867) );
  NAND2_X1 U7201 ( .A1(n9867), .A2(n5718), .ZN(n5559) );
  INV_X1 U7202 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U7203 ( .A1(n8457), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7204 ( .A1(n7002), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5555) );
  OAI211_X1 U7205 ( .C1(n8189), .C2(n5716), .A(n5556), .B(n5555), .ZN(n5557)
         );
  INV_X1 U7206 ( .A(n5557), .ZN(n5558) );
  NOR2_X1 U7207 ( .A1(n10109), .A2(n9877), .ZN(n9846) );
  INV_X1 U7208 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8396) );
  MUX2_X1 U7209 ( .A(n8408), .B(n8396), .S(n4394), .Z(n5580) );
  XNOR2_X1 U7210 ( .A(n5580), .B(SI_24_), .ZN(n5577) );
  NAND2_X1 U7211 ( .A1(n8395), .A2(n8464), .ZN(n5565) );
  NAND2_X1 U7212 ( .A1(n8466), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5564) );
  NAND2_X2 U7213 ( .A1(n5565), .A2(n5564), .ZN(n10106) );
  INV_X1 U7214 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U7215 ( .A1(n5567), .A2(n9596), .ZN(n5568) );
  NAND2_X1 U7216 ( .A1(n5590), .A2(n5568), .ZN(n9859) );
  INV_X1 U7217 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7218 ( .A1(n7002), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7219 ( .A1(n8456), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5569) );
  OAI211_X1 U7220 ( .C1(n5571), .C2(n5154), .A(n5570), .B(n5569), .ZN(n5572)
         );
  INV_X1 U7221 ( .A(n5572), .ZN(n5573) );
  INV_X1 U7222 ( .A(n9851), .ZN(n8685) );
  OR2_X1 U7223 ( .A1(n9846), .A2(n8685), .ZN(n5576) );
  NAND2_X1 U7224 ( .A1(n10109), .A2(n9877), .ZN(n9847) );
  OR2_X1 U7225 ( .A1(n8685), .A2(n9847), .ZN(n5575) );
  NAND2_X1 U7226 ( .A1(n10106), .A2(n9864), .ZN(n9840) );
  INV_X1 U7227 ( .A(n5577), .ZN(n5578) );
  INV_X1 U7228 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U7229 ( .A1(n5581), .A2(SI_24_), .ZN(n5582) );
  INV_X1 U7230 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8437) );
  INV_X1 U7231 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8434) );
  MUX2_X1 U7232 ( .A(n8437), .B(n8434), .S(n4393), .Z(n5584) );
  INV_X1 U7233 ( .A(SI_25_), .ZN(n5583) );
  NAND2_X1 U7234 ( .A1(n5584), .A2(n5583), .ZN(n5598) );
  INV_X1 U7235 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7236 ( .A1(n5585), .A2(SI_25_), .ZN(n5586) );
  NAND2_X1 U7237 ( .A1(n5598), .A2(n5586), .ZN(n5599) );
  XNOR2_X1 U7238 ( .A(n5600), .B(n5599), .ZN(n8432) );
  NAND2_X1 U7239 ( .A1(n8432), .A2(n8464), .ZN(n5588) );
  NAND2_X1 U7240 ( .A1(n8466), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5587) );
  INV_X1 U7241 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U7242 ( .A1(n5590), .A2(n9561), .ZN(n5591) );
  NAND2_X1 U7243 ( .A1(n5607), .A2(n5591), .ZN(n9836) );
  INV_X1 U7244 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U7245 ( .A1(n7002), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7246 ( .A1(n7001), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5592) );
  OAI211_X1 U7247 ( .C1(n8179), .C2(n5154), .A(n5593), .B(n5592), .ZN(n5594)
         );
  INV_X1 U7248 ( .A(n5594), .ZN(n5595) );
  NAND2_X1 U7249 ( .A1(n10099), .A2(n9853), .ZN(n8687) );
  AND2_X1 U7250 ( .A1(n9840), .A2(n5597), .ZN(n9817) );
  INV_X1 U7251 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9509) );
  INV_X1 U7252 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8439) );
  MUX2_X1 U7253 ( .A(n9509), .B(n8439), .S(n4393), .Z(n5602) );
  INV_X1 U7254 ( .A(SI_26_), .ZN(n5601) );
  NAND2_X1 U7255 ( .A1(n5602), .A2(n5601), .ZN(n5619) );
  INV_X1 U7256 ( .A(n5602), .ZN(n5603) );
  NAND2_X1 U7257 ( .A1(n5603), .A2(SI_26_), .ZN(n5604) );
  NAND2_X1 U7258 ( .A1(n8438), .A2(n8464), .ZN(n5606) );
  NAND2_X1 U7259 ( .A1(n8466), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5605) );
  INV_X1 U7260 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U7261 ( .A1(n5607), .A2(n9640), .ZN(n5608) );
  NAND2_X1 U7262 ( .A1(n9814), .A2(n5718), .ZN(n5614) );
  INV_X1 U7263 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U7264 ( .A1(n5179), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7265 ( .A1(n7001), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5609) );
  OAI211_X1 U7266 ( .C1(n5611), .C2(n8137), .A(n5610), .B(n5609), .ZN(n5612)
         );
  INV_X1 U7267 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7268 ( .A1(n10094), .A2(n9829), .ZN(n5615) );
  AND2_X2 U7269 ( .A1(n8689), .A2(n5615), .ZN(n9821) );
  INV_X1 U7270 ( .A(n9821), .ZN(n5616) );
  OR2_X1 U7271 ( .A1(n10099), .A2(n9808), .ZN(n9818) );
  NAND2_X1 U7272 ( .A1(n5618), .A2(n5617), .ZN(n5620) );
  INV_X1 U7273 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9505) );
  INV_X1 U7274 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5621) );
  MUX2_X1 U7275 ( .A(n9505), .B(n5621), .S(n4394), .Z(n5623) );
  INV_X1 U7276 ( .A(SI_27_), .ZN(n5622) );
  NAND2_X1 U7277 ( .A1(n5623), .A2(n5622), .ZN(n5640) );
  INV_X1 U7278 ( .A(n5623), .ZN(n5624) );
  NAND2_X1 U7279 ( .A1(n5624), .A2(SI_27_), .ZN(n5625) );
  NAND2_X1 U7280 ( .A1(n9504), .A2(n8464), .ZN(n5627) );
  NAND2_X1 U7281 ( .A1(n8466), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5626) );
  INV_X1 U7282 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9518) );
  NAND2_X1 U7283 ( .A1(n5629), .A2(n9518), .ZN(n5630) );
  NAND2_X1 U7284 ( .A1(n5644), .A2(n5630), .ZN(n9793) );
  INV_X1 U7285 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U7286 ( .A1(n8456), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7287 ( .A1(n7002), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5632) );
  OAI211_X1 U7288 ( .C1(n8210), .C2(n5154), .A(n5633), .B(n5632), .ZN(n5634)
         );
  INV_X1 U7289 ( .A(n5634), .ZN(n5635) );
  NAND2_X1 U7290 ( .A1(n10089), .A2(n9641), .ZN(n8695) );
  NAND2_X1 U7291 ( .A1(n9799), .A2(n9798), .ZN(n9797) );
  OR2_X1 U7292 ( .A1(n10089), .A2(n9807), .ZN(n5637) );
  INV_X1 U7293 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9502) );
  INV_X1 U7294 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5641) );
  MUX2_X1 U7295 ( .A(n9502), .B(n5641), .S(n4394), .Z(n6112) );
  XNOR2_X1 U7296 ( .A(n6112), .B(SI_28_), .ZN(n6109) );
  NAND2_X1 U7297 ( .A1(n9501), .A2(n8464), .ZN(n5643) );
  NAND2_X1 U7298 ( .A1(n8466), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5642) );
  INV_X1 U7299 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U7300 ( .A1(n5644), .A2(n8047), .ZN(n5645) );
  NAND2_X1 U7301 ( .A1(n6890), .A2(n5718), .ZN(n5651) );
  INV_X1 U7302 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7303 ( .A1(n7002), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7304 ( .A1(n7001), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5646) );
  OAI211_X1 U7305 ( .C1(n5154), .C2(n5648), .A(n5647), .B(n5646), .ZN(n5649)
         );
  INV_X1 U7306 ( .A(n5649), .ZN(n5650) );
  NOR2_X1 U7307 ( .A1(n5652), .A2(n8470), .ZN(n5653) );
  OR2_X2 U7308 ( .A1(n10072), .A2(n5653), .ZN(n10088) );
  INV_X1 U7309 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5654) );
  INV_X1 U7310 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5655) );
  INV_X1 U7311 ( .A(n5656), .ZN(n5657) );
  NAND2_X1 U7312 ( .A1(n5657), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5659) );
  INV_X1 U7313 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5661) );
  NAND3_X1 U7314 ( .A1(n5668), .A2(n5220), .A3(n5663), .ZN(n5677) );
  NOR2_X1 U7315 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  NAND2_X1 U7316 ( .A1(n5669), .A2(n5670), .ZN(n8397) );
  INV_X1 U7317 ( .A(n8397), .ZN(n5676) );
  INV_X1 U7318 ( .A(n8433), .ZN(n5675) );
  NAND3_X2 U7319 ( .A1(n5676), .A2(n5683), .A3(n5675), .ZN(n6904) );
  NAND2_X1 U7320 ( .A1(n5677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5679) );
  XNOR2_X1 U7321 ( .A(n5679), .B(n5678), .ZN(n8236) );
  AND2_X1 U7322 ( .A1(n8236), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7323 ( .A1(n8433), .A2(P1_B_REG_SCAN_IN), .ZN(n5681) );
  MUX2_X1 U7324 ( .A(P1_B_REG_SCAN_IN), .B(n5681), .S(n8397), .Z(n5682) );
  INV_X1 U7325 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U7326 ( .A1(n10212), .A2(n8207), .ZN(n5685) );
  INV_X1 U7327 ( .A(n5683), .ZN(n8440) );
  NAND2_X1 U7328 ( .A1(n8440), .A2(n8433), .ZN(n5684) );
  NAND2_X1 U7329 ( .A1(n5685), .A2(n5684), .ZN(n7047) );
  INV_X1 U7330 ( .A(n7047), .ZN(n6977) );
  NOR4_X1 U7331 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8159) );
  NOR2_X1 U7332 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .ZN(
        n5688) );
  NOR4_X1 U7333 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5687) );
  NOR4_X1 U7334 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5686) );
  NAND4_X1 U7335 ( .A1(n8159), .A2(n5688), .A3(n5687), .A4(n5686), .ZN(n5694)
         );
  NOR4_X1 U7336 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5692) );
  NOR4_X1 U7337 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5691) );
  NOR4_X1 U7338 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n5690) );
  NOR4_X1 U7339 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5689) );
  NAND4_X1 U7340 ( .A1(n5692), .A2(n5691), .A3(n5690), .A4(n5689), .ZN(n5693)
         );
  OAI21_X1 U7341 ( .B1(n5694), .B2(n5693), .A(n10212), .ZN(n7046) );
  INV_X1 U7342 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7343 ( .A1(n10212), .A2(n5695), .ZN(n5696) );
  NAND2_X1 U7344 ( .A1(n8440), .A2(n8397), .ZN(n10214) );
  NAND2_X1 U7345 ( .A1(n5696), .A2(n10214), .ZN(n7244) );
  NAND3_X1 U7346 ( .A1(n6977), .A2(n7046), .A3(n7244), .ZN(n5697) );
  AND2_X1 U7347 ( .A1(n8561), .A2(n6979), .ZN(n5698) );
  OR2_X1 U7348 ( .A1(n7358), .A2(n5701), .ZN(n8725) );
  NAND2_X4 U7349 ( .A1(n5701), .A2(n7358), .ZN(n6847) );
  NAND2_X1 U7350 ( .A1(n9940), .A2(n7252), .ZN(n10028) );
  NAND2_X1 U7351 ( .A1(n7248), .A2(n7361), .ZN(n7360) );
  NAND2_X1 U7352 ( .A1(n7051), .A2(n7368), .ZN(n5702) );
  NAND2_X1 U7353 ( .A1(n8564), .A2(n8474), .ZN(n5703) );
  NAND2_X1 U7354 ( .A1(n5703), .A2(n8563), .ZN(n7410) );
  NAND2_X1 U7355 ( .A1(n7410), .A2(n8475), .ZN(n7411) );
  AND2_X1 U7356 ( .A1(n8516), .A2(n8514), .ZN(n8521) );
  OR2_X1 U7357 ( .A1(n10174), .A2(n7946), .ZN(n8615) );
  AND2_X1 U7358 ( .A1(n8615), .A2(n8612), .ZN(n8634) );
  NAND2_X1 U7359 ( .A1(n7789), .A2(n8634), .ZN(n8287) );
  NAND2_X1 U7360 ( .A1(n10174), .A2(n7946), .ZN(n8613) );
  AND2_X2 U7361 ( .A1(n8291), .A2(n8636), .ZN(n8273) );
  NAND2_X1 U7362 ( .A1(n8273), .A2(n8527), .ZN(n8321) );
  NAND2_X1 U7363 ( .A1(n10164), .A2(n10015), .ZN(n10010) );
  NAND2_X1 U7364 ( .A1(n8531), .A2(n10010), .ZN(n10039) );
  NAND2_X1 U7365 ( .A1(n8619), .A2(n8532), .ZN(n10026) );
  INV_X1 U7366 ( .A(n10010), .ZN(n5706) );
  NOR2_X1 U7367 ( .A1(n10026), .A2(n5706), .ZN(n5707) );
  AND2_X1 U7368 ( .A1(n8649), .A2(n9975), .ZN(n5708) );
  NAND2_X1 U7369 ( .A1(n10144), .A2(n9628), .ZN(n9945) );
  AND2_X1 U7370 ( .A1(n8540), .A2(n9945), .ZN(n8603) );
  OR2_X1 U7371 ( .A1(n10144), .A2(n9628), .ZN(n9943) );
  NAND2_X1 U7372 ( .A1(n8655), .A2(n9943), .ZN(n8541) );
  AND2_X1 U7373 ( .A1(n8541), .A2(n8540), .ZN(n5709) );
  OR2_X1 U7374 ( .A1(n10133), .A2(n9909), .ZN(n8656) );
  NAND2_X1 U7375 ( .A1(n10133), .A2(n9909), .ZN(n8657) );
  INV_X1 U7376 ( .A(n8671), .ZN(n5710) );
  INV_X1 U7377 ( .A(n9894), .ZN(n9531) );
  NAND2_X1 U7378 ( .A1(n10113), .A2(n9531), .ZN(n8678) );
  INV_X1 U7379 ( .A(n10109), .ZN(n9869) );
  NAND2_X1 U7380 ( .A1(n9869), .A2(n9877), .ZN(n8595) );
  NAND2_X1 U7381 ( .A1(n8687), .A2(n8594), .ZN(n8599) );
  OR2_X1 U7382 ( .A1(n10094), .A2(n9519), .ZN(n5712) );
  NAND2_X1 U7383 ( .A1(n5712), .A2(n9804), .ZN(n8547) );
  NAND2_X1 U7384 ( .A1(n10094), .A2(n9519), .ZN(n8549) );
  OAI21_X1 U7385 ( .B1(n9785), .B2(n9798), .A(n8694), .ZN(n9766) );
  XNOR2_X1 U7386 ( .A(n9766), .B(n8470), .ZN(n5725) );
  NAND2_X1 U7387 ( .A1(n8726), .A2(n8502), .ZN(n5713) );
  OR2_X1 U7388 ( .A1(n8561), .A2(n4392), .ZN(n8719) );
  INV_X1 U7389 ( .A(n9778), .ZN(n5719) );
  INV_X1 U7390 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U7391 ( .A1(n8457), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7392 ( .A1(n7002), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5714) );
  OAI211_X1 U7393 ( .C1(n5716), .C2(n9777), .A(n5715), .B(n5714), .ZN(n5717)
         );
  AOI21_X1 U7394 ( .B1(n5719), .B2(n5718), .A(n5717), .ZN(n8469) );
  INV_X1 U7395 ( .A(n8469), .ZN(n9665) );
  INV_X1 U7396 ( .A(n8717), .ZN(n5721) );
  NAND2_X1 U7397 ( .A1(n7256), .A2(n7424), .ZN(n7257) );
  INV_X1 U7398 ( .A(n7758), .ZN(n7597) );
  INV_X1 U7399 ( .A(n8399), .ZN(n8286) );
  INV_X1 U7400 ( .A(n10159), .ZN(n10025) );
  NAND2_X1 U7401 ( .A1(n10050), .A2(n10025), .ZN(n10020) );
  INV_X1 U7402 ( .A(n10144), .ZN(n9968) );
  INV_X1 U7403 ( .A(n10138), .ZN(n9955) );
  INV_X1 U7404 ( .A(n10106), .ZN(n9854) );
  INV_X1 U7405 ( .A(n10099), .ZN(n9839) );
  NOR2_X2 U7406 ( .A1(n9833), .A2(n10094), .ZN(n9813) );
  INV_X1 U7407 ( .A(n10089), .ZN(n9796) );
  NAND2_X1 U7408 ( .A1(n8442), .A2(n8561), .ZN(n7054) );
  INV_X1 U7409 ( .A(n9774), .ZN(n5728) );
  AOI211_X1 U7410 ( .C1(n10085), .C2(n9790), .A(n10287), .B(n5728), .ZN(n10084) );
  NOR2_X1 U7411 ( .A1(n5729), .A2(n8502), .ZN(n10031) );
  INV_X1 U7412 ( .A(n10031), .ZN(n9903) );
  OR2_X1 U7413 ( .A1(n7054), .A2(n4392), .ZN(n6887) );
  INV_X1 U7414 ( .A(n6887), .ZN(n5730) );
  INV_X2 U7415 ( .A(n9898), .ZN(n10051) );
  AOI22_X1 U7416 ( .A1(n6890), .A2(n10051), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n10062), .ZN(n5731) );
  OAI21_X1 U7417 ( .B1(n6876), .B2(n10054), .A(n5731), .ZN(n5732) );
  AOI21_X1 U7418 ( .B1(n10084), .B2(n10031), .A(n5732), .ZN(n5733) );
  AND3_X2 U7419 ( .A1(n5740), .A2(n5739), .A3(n5933), .ZN(n5952) );
  NOR2_X1 U7420 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5743) );
  NOR2_X1 U7421 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5742) );
  NAND4_X1 U7422 ( .A1(n5743), .A2(n5742), .A3(n5741), .A4(n6127), .ZN(n5746)
         );
  INV_X2 U7423 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8163) );
  NAND4_X1 U7424 ( .A1(n8163), .A2(n5744), .A3(n6144), .A4(n6131), .ZN(n5745)
         );
  NAND2_X1 U7425 ( .A1(n6204), .A2(n5749), .ZN(n5772) );
  NAND2_X1 U7426 ( .A1(n8240), .A2(n6056), .ZN(n5754) );
  OR2_X1 U7427 ( .A1(n5841), .A2(n8243), .ZN(n5753) );
  INV_X1 U7428 ( .A(n5861), .ZN(n5756) );
  NAND2_X1 U7429 ( .A1(n5756), .A2(n5755), .ZN(n5882) );
  INV_X1 U7430 ( .A(n5882), .ZN(n5757) );
  NAND2_X1 U7431 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5758) );
  NAND2_X1 U7432 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n5762) );
  NAND2_X1 U7433 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5764) );
  INV_X1 U7434 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8839) );
  INV_X1 U7435 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8860) );
  INV_X1 U7436 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5767) );
  OAI21_X1 U7437 ( .B1(n6050), .B2(n8860), .A(n5767), .ZN(n5769) );
  NAND2_X1 U7438 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5768) );
  AND2_X1 U7439 ( .A1(n5769), .A2(n6058), .ZN(n9188) );
  INV_X1 U7440 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U7441 ( .A1(n9188), .A2(n5831), .ZN(n5784) );
  INV_X1 U7442 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n5781) );
  NOR2_X2 U7443 ( .A1(n5778), .A2(n5777), .ZN(n5817) );
  INV_X1 U7444 ( .A(n5817), .ZN(n5797) );
  INV_X2 U7445 ( .A(n5797), .ZN(n6210) );
  NAND2_X1 U7446 ( .A1(n6210), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5780) );
  INV_X4 U7447 ( .A(n6093), .ZN(n6251) );
  NAND2_X1 U7448 ( .A1(n6251), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5779) );
  OAI211_X1 U7449 ( .C1(n6120), .C2(n5781), .A(n5780), .B(n5779), .ZN(n5782)
         );
  INV_X1 U7450 ( .A(n5782), .ZN(n5783) );
  NAND2_X1 U7451 ( .A1(n5784), .A2(n5783), .ZN(n9164) );
  INV_X1 U7452 ( .A(n9164), .ZN(n9206) );
  OR2_X1 U7453 ( .A1(n5838), .A2(n9497), .ZN(n5800) );
  XNOR2_X1 U7454 ( .A(n5800), .B(n5836), .ZN(n7265) );
  NAND2_X1 U7455 ( .A1(n5831), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7456 ( .A1(n5817), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7457 ( .A1(n4385), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7458 ( .A1(n5818), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7459 ( .A1(n10365), .A2(n10315), .ZN(n6303) );
  NAND2_X1 U7460 ( .A1(n6303), .A2(n7746), .ZN(n6440) );
  NAND2_X1 U7461 ( .A1(n5793), .A2(n10365), .ZN(n5828) );
  NAND2_X1 U7462 ( .A1(n4545), .A2(n5828), .ZN(n7751) );
  NAND2_X1 U7463 ( .A1(n4385), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7464 ( .A1(n5818), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5795) );
  INV_X1 U7465 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U7466 ( .A1(n5831), .A2(n7753), .ZN(n5794) );
  NAND2_X1 U7467 ( .A1(n5817), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5798) );
  OR2_X1 U7468 ( .A1(n7008), .A2(n5840), .ZN(n5806) );
  NAND2_X1 U7469 ( .A1(n5800), .A2(n5836), .ZN(n5801) );
  NAND2_X1 U7470 ( .A1(n5801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5803) );
  INV_X1 U7471 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5802) );
  XNOR2_X1 U7472 ( .A(n5803), .B(n5802), .ZN(n8944) );
  OR2_X1 U7473 ( .A1(n5799), .A2(n8944), .ZN(n5804) );
  NAND2_X1 U7474 ( .A1(n5808), .A2(n5807), .ZN(n7679) );
  NAND2_X1 U7475 ( .A1(n8930), .A2(n7482), .ZN(n6308) );
  NAND2_X1 U7476 ( .A1(n4385), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7477 ( .A1(n5817), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7478 ( .A1(n5818), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5809) );
  AND4_X2 U7479 ( .A1(n5812), .A2(n5811), .A3(n5810), .A4(n5809), .ZN(n7709)
         );
  NAND2_X1 U7480 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5813) );
  INV_X1 U7481 ( .A(n5838), .ZN(n5814) );
  NAND2_X1 U7482 ( .A1(n10309), .A2(n6302), .ZN(n6443) );
  NAND2_X1 U7483 ( .A1(n4385), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7484 ( .A1(n5831), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7485 ( .A1(n5817), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7486 ( .A1(n5818), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7487 ( .A1(n6986), .A2(SI_0_), .ZN(n5824) );
  INV_X1 U7488 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7489 ( .A1(n5824), .A2(n5823), .ZN(n5826) );
  AND2_X1 U7490 ( .A1(n5826), .A2(n5825), .ZN(n9513) );
  NAND2_X1 U7491 ( .A1(n6293), .A2(n10353), .ZN(n5827) );
  NAND2_X1 U7492 ( .A1(n6443), .A2(n5827), .ZN(n7718) );
  NAND2_X1 U7493 ( .A1(n7709), .A2(n10326), .ZN(n7717) );
  AND2_X1 U7494 ( .A1(n7717), .A2(n5828), .ZN(n5829) );
  NAND2_X1 U7495 ( .A1(n5808), .A2(n7482), .ZN(n7675) );
  NAND2_X1 U7496 ( .A1(n4386), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5835) );
  INV_X1 U7497 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U7498 ( .A1(n7753), .A2(n8200), .ZN(n5830) );
  AND2_X1 U7499 ( .A1(n5830), .A2(n5861), .ZN(n7685) );
  NAND2_X1 U7500 ( .A1(n5831), .A2(n7685), .ZN(n5834) );
  NAND2_X1 U7501 ( .A1(n5818), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7502 ( .A1(n5817), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5832) );
  NOR2_X1 U7503 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5837) );
  NAND2_X1 U7504 ( .A1(n5838), .A2(n5837), .ZN(n5931) );
  NAND2_X1 U7505 ( .A1(n5931), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5839) );
  XNOR2_X1 U7506 ( .A(n5839), .B(n4523), .ZN(n7296) );
  NAND2_X1 U7507 ( .A1(n6056), .A2(n6980), .ZN(n5843) );
  OR2_X1 U7508 ( .A1(n5841), .A2(n6988), .ZN(n5842) );
  OAI211_X1 U7509 ( .C1(n5799), .C2(n7296), .A(n5843), .B(n5842), .ZN(n7688)
         );
  NAND2_X1 U7510 ( .A1(n7731), .A2(n6497), .ZN(n5845) );
  AND2_X1 U7511 ( .A1(n7675), .A2(n5845), .ZN(n5844) );
  INV_X1 U7512 ( .A(n5845), .ZN(n5846) );
  INV_X1 U7513 ( .A(n7731), .ZN(n8929) );
  NAND2_X1 U7514 ( .A1(n7731), .A2(n7688), .ZN(n6288) );
  NAND2_X1 U7515 ( .A1(n4386), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5850) );
  XNOR2_X1 U7516 ( .A(n5861), .B(P2_REG3_REG_5__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U7517 ( .A1(n6043), .A2(n7733), .ZN(n5849) );
  NAND2_X1 U7518 ( .A1(n5818), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7519 ( .A1(n5817), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5847) );
  AND4_X2 U7520 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n7536)
         );
  NAND2_X1 U7521 ( .A1(n5852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5851) );
  MUX2_X1 U7522 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5851), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5855) );
  INV_X1 U7523 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7524 ( .A1(n5854), .A2(n5853), .ZN(n5872) );
  NAND2_X1 U7525 ( .A1(n5855), .A2(n5872), .ZN(n8960) );
  INV_X1 U7526 ( .A(n8960), .ZN(n8965) );
  AOI22_X1 U7527 ( .A1(n6022), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6021), .B2(
        n8965), .ZN(n5857) );
  NAND2_X1 U7528 ( .A1(n6989), .A2(n6056), .ZN(n5856) );
  INV_X1 U7529 ( .A(n7738), .ZN(n10383) );
  AND2_X1 U7530 ( .A1(n7536), .A2(n10383), .ZN(n5858) );
  NAND2_X1 U7531 ( .A1(n7536), .A2(n7738), .ZN(n6290) );
  INV_X1 U7532 ( .A(n7536), .ZN(n8928) );
  NAND2_X1 U7533 ( .A1(n8928), .A2(n10383), .ZN(n6310) );
  NAND2_X1 U7534 ( .A1(n6290), .A2(n6310), .ZN(n7737) );
  OAI22_X1 U7535 ( .A1(n7736), .A2(n5858), .B1(n10383), .B2(n7737), .ZN(n7691)
         );
  NAND2_X1 U7536 ( .A1(n4386), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5866) );
  INV_X1 U7537 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5860) );
  INV_X1 U7538 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5859) );
  OAI21_X1 U7539 ( .B1(n5861), .B2(n5860), .A(n5859), .ZN(n5862) );
  AND2_X1 U7540 ( .A1(n5882), .A2(n5862), .ZN(n7698) );
  NAND2_X1 U7541 ( .A1(n6043), .A2(n7698), .ZN(n5865) );
  NAND2_X1 U7542 ( .A1(n6251), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7543 ( .A1(n6210), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7544 ( .A1(n6992), .A2(n6056), .ZN(n5869) );
  NAND2_X1 U7545 ( .A1(n5872), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5867) );
  XNOR2_X1 U7546 ( .A(n5867), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8979) );
  AOI22_X1 U7547 ( .A1(n6022), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6021), .B2(
        n8979), .ZN(n5868) );
  NAND2_X1 U7548 ( .A1(n5869), .A2(n5868), .ZN(n7701) );
  AND2_X1 U7549 ( .A1(n7730), .A2(n7701), .ZN(n6291) );
  INV_X1 U7550 ( .A(n6291), .ZN(n7618) );
  INV_X1 U7551 ( .A(n7701), .ZN(n10391) );
  INV_X1 U7552 ( .A(n7730), .ZN(n8927) );
  NAND2_X1 U7553 ( .A1(n10391), .A2(n8927), .ZN(n6312) );
  NAND2_X1 U7554 ( .A1(n7618), .A2(n6312), .ZN(n6448) );
  NAND2_X1 U7555 ( .A1(n7691), .A2(n6448), .ZN(n5871) );
  OR2_X1 U7556 ( .A1(n7730), .A2(n10391), .ZN(n5870) );
  NAND2_X1 U7557 ( .A1(n5871), .A2(n5870), .ZN(n7616) );
  INV_X1 U7558 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U7559 ( .A1(n5874), .A2(n5873), .ZN(n5896) );
  NAND2_X1 U7560 ( .A1(n5896), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5875) );
  XNOR2_X1 U7561 ( .A(n5875), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7303) );
  AOI22_X1 U7562 ( .A1(n6022), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6021), .B2(
        n7303), .ZN(n5876) );
  NAND2_X1 U7563 ( .A1(n4386), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5880) );
  XNOR2_X1 U7564 ( .A(n5901), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n7477) );
  NAND2_X1 U7565 ( .A1(n6043), .A2(n7477), .ZN(n5879) );
  NAND2_X1 U7566 ( .A1(n6251), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7567 ( .A1(n6210), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7568 ( .A1(n4386), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5887) );
  INV_X1 U7569 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7570 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  AND2_X1 U7571 ( .A1(n5901), .A2(n5883), .ZN(n7859) );
  NAND2_X1 U7572 ( .A1(n6043), .A2(n7859), .ZN(n5886) );
  NAND2_X1 U7573 ( .A1(n6251), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7574 ( .A1(n6210), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5884) );
  INV_X1 U7575 ( .A(n7876), .ZN(n8926) );
  NAND2_X1 U7576 ( .A1(n6995), .A2(n6056), .ZN(n5891) );
  NAND2_X1 U7577 ( .A1(n5888), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U7578 ( .A(n5889), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8995) );
  AOI22_X1 U7579 ( .A1(n6022), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6021), .B2(
        n8995), .ZN(n5890) );
  OR2_X1 U7580 ( .A1(n8926), .A2(n7622), .ZN(n7867) );
  NAND2_X1 U7581 ( .A1(n7616), .A2(n5892), .ZN(n5895) );
  NAND2_X1 U7582 ( .A1(n7622), .A2(n7876), .ZN(n6336) );
  AND2_X2 U7583 ( .A1(n6318), .A2(n6336), .ZN(n7868) );
  AND2_X1 U7584 ( .A1(n7868), .A2(n7867), .ZN(n5893) );
  INV_X1 U7585 ( .A(n7832), .ZN(n8925) );
  AOI22_X1 U7586 ( .A1(n5893), .A2(n7873), .B1(n10397), .B2(n8925), .ZN(n5894)
         );
  NAND2_X1 U7587 ( .A1(n5895), .A2(n5894), .ZN(n7823) );
  INV_X1 U7588 ( .A(n7823), .ZN(n5908) );
  NAND2_X1 U7589 ( .A1(n7019), .A2(n6056), .ZN(n5898) );
  NAND2_X1 U7590 ( .A1(n4456), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5910) );
  AOI22_X1 U7591 ( .A1(n6022), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6021), .B2(
        n9029), .ZN(n5897) );
  NAND2_X1 U7592 ( .A1(n4386), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5906) );
  INV_X1 U7593 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5900) );
  INV_X1 U7594 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5899) );
  OAI21_X1 U7595 ( .B1(n5901), .B2(n5900), .A(n5899), .ZN(n5902) );
  AND2_X1 U7596 ( .A1(n5902), .A2(n5923), .ZN(n7914) );
  NAND2_X1 U7597 ( .A1(n6043), .A2(n7914), .ZN(n5905) );
  NAND2_X1 U7598 ( .A1(n6251), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7599 ( .A1(n6210), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5903) );
  NAND4_X1 U7600 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n8924)
         );
  AND2_X1 U7601 ( .A1(n7828), .A2(n8924), .ZN(n6324) );
  INV_X1 U7602 ( .A(n8924), .ZN(n7877) );
  NAND2_X1 U7603 ( .A1(n7915), .A2(n7877), .ZN(n6329) );
  NAND2_X1 U7604 ( .A1(n5908), .A2(n5907), .ZN(n7821) );
  NAND2_X1 U7605 ( .A1(n7828), .A2(n7877), .ZN(n5909) );
  NAND2_X1 U7606 ( .A1(n5910), .A2(n4916), .ZN(n5911) );
  NAND2_X1 U7607 ( .A1(n5911), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7608 ( .A1(n5921), .A2(n5912), .ZN(n5913) );
  NAND2_X1 U7609 ( .A1(n5913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5914) );
  AOI22_X1 U7610 ( .A1(n9042), .A2(n6021), .B1(n6022), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7611 ( .A1(n4386), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U7612 ( .A(n5942), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U7613 ( .A1(n6043), .A2(n8873), .ZN(n5919) );
  NAND2_X1 U7614 ( .A1(n6251), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7615 ( .A1(n6210), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7616 ( .A1(n9470), .A2(n8785), .ZN(n6345) );
  NAND2_X1 U7617 ( .A1(n8309), .A2(n6345), .ZN(n8371) );
  INV_X1 U7618 ( .A(n8371), .ZN(n8369) );
  XNOR2_X1 U7619 ( .A(n5921), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7331) );
  AOI22_X1 U7620 ( .A1(n6022), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7331), .B2(
        n6021), .ZN(n5922) );
  NAND2_X1 U7621 ( .A1(n4386), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7622 ( .A1(n5923), .A2(n7784), .ZN(n5924) );
  NAND2_X1 U7623 ( .A1(n5942), .A2(n5924), .ZN(n8230) );
  INV_X1 U7624 ( .A(n8230), .ZN(n5925) );
  NAND2_X1 U7625 ( .A1(n6043), .A2(n5925), .ZN(n5928) );
  NAND2_X1 U7626 ( .A1(n6251), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7627 ( .A1(n6210), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5926) );
  INV_X1 U7628 ( .A(n7831), .ZN(n8923) );
  AND2_X1 U7629 ( .A1(n8229), .A2(n8923), .ZN(n8367) );
  INV_X1 U7630 ( .A(n8785), .ZN(n8922) );
  NAND2_X1 U7631 ( .A1(n7056), .A2(n6056), .ZN(n5939) );
  INV_X1 U7632 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5932) );
  NAND4_X1 U7633 ( .A1(n4524), .A2(n4417), .A3(n5933), .A4(n5932), .ZN(n5936)
         );
  NAND2_X1 U7634 ( .A1(n5936), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5935) );
  INV_X1 U7635 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5934) );
  MUX2_X1 U7636 ( .A(n5935), .B(P2_IR_REG_31__SCAN_IN), .S(n5934), .Z(n5937)
         );
  NAND2_X1 U7637 ( .A1(n5937), .A2(n5949), .ZN(n7371) );
  INV_X1 U7638 ( .A(n7371), .ZN(n7378) );
  AOI22_X1 U7639 ( .A1(n6022), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6021), .B2(
        n7378), .ZN(n5938) );
  NAND2_X1 U7640 ( .A1(n4386), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5947) );
  INV_X1 U7641 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5941) );
  INV_X1 U7642 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5940) );
  OAI21_X1 U7643 ( .B1(n5942), .B2(n5941), .A(n5940), .ZN(n5943) );
  AND2_X1 U7644 ( .A1(n5956), .A2(n5943), .ZN(n8783) );
  NAND2_X1 U7645 ( .A1(n5831), .A2(n8783), .ZN(n5946) );
  NAND2_X1 U7646 ( .A1(n6251), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7647 ( .A1(n6210), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7648 ( .A1(n9465), .A2(n6539), .ZN(n6346) );
  NAND2_X1 U7649 ( .A1(n9465), .A2(n6539), .ZN(n6347) );
  NAND2_X1 U7650 ( .A1(n6346), .A2(n6347), .ZN(n8316) );
  INV_X1 U7651 ( .A(n8316), .ZN(n5948) );
  INV_X1 U7652 ( .A(n6539), .ZN(n8921) );
  NAND2_X1 U7653 ( .A1(n7125), .A2(n6056), .ZN(n5955) );
  NAND2_X1 U7654 ( .A1(n5949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5950) );
  MUX2_X1 U7655 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5950), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n5951) );
  INV_X1 U7656 ( .A(n5951), .ZN(n5953) );
  NOR2_X1 U7657 ( .A1(n5953), .A2(n5984), .ZN(n7375) );
  AOI22_X1 U7658 ( .A1(n6022), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6021), .B2(
        n7375), .ZN(n5954) );
  NAND2_X1 U7659 ( .A1(n4386), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5961) );
  INV_X1 U7660 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U7661 ( .A1(n5956), .A2(n8162), .ZN(n5957) );
  AND2_X1 U7662 ( .A1(n5977), .A2(n5957), .ZN(n8847) );
  NAND2_X1 U7663 ( .A1(n6043), .A2(n8847), .ZN(n5960) );
  NAND2_X1 U7664 ( .A1(n6210), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7665 ( .A1(n6251), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5958) );
  OR2_X2 U7666 ( .A1(n9460), .A2(n8743), .ZN(n6357) );
  NAND2_X1 U7667 ( .A1(n9460), .A2(n8743), .ZN(n9331) );
  INV_X1 U7668 ( .A(n8743), .ZN(n8920) );
  NAND2_X1 U7669 ( .A1(n7145), .A2(n6056), .ZN(n5967) );
  OR2_X1 U7670 ( .A1(n5984), .A2(n9497), .ZN(n5964) );
  INV_X1 U7671 ( .A(n5964), .ZN(n5962) );
  NAND2_X1 U7672 ( .A1(n5962), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5965) );
  INV_X1 U7673 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U7674 ( .A1(n5964), .A2(n5963), .ZN(n5972) );
  AOI22_X1 U7675 ( .A1(n6022), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6021), .B2(
        n7812), .ZN(n5966) );
  NAND2_X1 U7676 ( .A1(n4386), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5971) );
  XNOR2_X1 U7677 ( .A(n5977), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U7678 ( .A1(n6043), .A2(n9358), .ZN(n5970) );
  NAND2_X1 U7679 ( .A1(n6210), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7680 ( .A1(n6251), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5968) );
  NAND4_X1 U7681 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(n9334)
         );
  XNOR2_X1 U7682 ( .A(n9455), .B(n8850), .ZN(n9364) );
  INV_X1 U7683 ( .A(n9364), .ZN(n6453) );
  NAND2_X1 U7684 ( .A1(n7152), .A2(n6056), .ZN(n5975) );
  NAND2_X1 U7685 ( .A1(n5972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U7686 ( .A(n5973), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8259) );
  AOI22_X1 U7687 ( .A1(n6022), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6021), .B2(
        n8259), .ZN(n5974) );
  NAND2_X1 U7688 ( .A1(n4386), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5982) );
  INV_X1 U7689 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5976) );
  INV_X1 U7690 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7957) );
  OAI21_X1 U7691 ( .B1(n5977), .B2(n5976), .A(n7957), .ZN(n5978) );
  AND2_X1 U7692 ( .A1(n5978), .A2(n5990), .ZN(n9339) );
  NAND2_X1 U7693 ( .A1(n5831), .A2(n9339), .ZN(n5981) );
  NAND2_X1 U7694 ( .A1(n6251), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7695 ( .A1(n6210), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5979) );
  OR2_X1 U7696 ( .A1(n9450), .A2(n9311), .ZN(n6365) );
  NAND2_X1 U7697 ( .A1(n9450), .A2(n9311), .ZN(n6368) );
  NAND2_X1 U7698 ( .A1(n6365), .A2(n6368), .ZN(n6360) );
  NAND2_X1 U7699 ( .A1(n9342), .A2(n6360), .ZN(n9343) );
  NAND2_X1 U7700 ( .A1(n7184), .A2(n6056), .ZN(n5989) );
  NAND2_X1 U7701 ( .A1(n5985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5986) );
  MUX2_X1 U7702 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5986), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5987) );
  AND2_X1 U7703 ( .A1(n6123), .A2(n5987), .ZN(n9061) );
  AOI22_X1 U7704 ( .A1(n6022), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6021), .B2(
        n9061), .ZN(n5988) );
  NAND2_X1 U7705 ( .A1(n4386), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5995) );
  INV_X1 U7706 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8255) );
  NAND2_X1 U7707 ( .A1(n5990), .A2(n8255), .ZN(n5991) );
  AND2_X1 U7708 ( .A1(n6009), .A2(n5991), .ZN(n9324) );
  NAND2_X1 U7709 ( .A1(n5831), .A2(n9324), .ZN(n5994) );
  NAND2_X1 U7710 ( .A1(n6210), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7711 ( .A1(n6251), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7712 ( .A1(n9445), .A2(n9290), .ZN(n9286) );
  OR2_X1 U7713 ( .A1(n9445), .A2(n9290), .ZN(n5996) );
  NAND2_X1 U7714 ( .A1(n9286), .A2(n5996), .ZN(n6370) );
  INV_X1 U7715 ( .A(n9311), .ZN(n8919) );
  OR2_X1 U7716 ( .A1(n9450), .A2(n8919), .ZN(n9314) );
  AND2_X1 U7717 ( .A1(n6370), .A2(n9314), .ZN(n5997) );
  NAND2_X1 U7718 ( .A1(n7205), .A2(n6056), .ZN(n6000) );
  NAND2_X1 U7719 ( .A1(n6123), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5998) );
  XNOR2_X1 U7720 ( .A(n5998), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9072) );
  AOI22_X1 U7721 ( .A1(n6022), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6021), .B2(
        n9072), .ZN(n5999) );
  NAND2_X1 U7722 ( .A1(n4386), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6004) );
  XNOR2_X1 U7723 ( .A(n6009), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U7724 ( .A1(n5831), .A2(n8821), .ZN(n6003) );
  NAND2_X1 U7725 ( .A1(n6210), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7726 ( .A1(n6251), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7727 ( .A1(n9442), .A2(n9313), .ZN(n6371) );
  INV_X1 U7728 ( .A(n9290), .ZN(n9335) );
  NAND2_X1 U7729 ( .A1(n9445), .A2(n9335), .ZN(n9293) );
  NAND2_X1 U7730 ( .A1(n7351), .A2(n6056), .ZN(n6007) );
  XNOR2_X1 U7731 ( .A(n6017), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9083) );
  AOI22_X1 U7732 ( .A1(n6022), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6021), .B2(
        n9083), .ZN(n6006) );
  NAND2_X2 U7733 ( .A1(n6007), .A2(n6006), .ZN(n9435) );
  NAND2_X1 U7734 ( .A1(n4385), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6014) );
  INV_X1 U7735 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9054) );
  INV_X1 U7736 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6008) );
  OAI21_X1 U7737 ( .B1(n6009), .B2(n9054), .A(n6008), .ZN(n6010) );
  AND2_X1 U7738 ( .A1(n6010), .A2(n6026), .ZN(n9275) );
  NAND2_X1 U7739 ( .A1(n5831), .A2(n9275), .ZN(n6013) );
  NAND2_X1 U7740 ( .A1(n6251), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7741 ( .A1(n6210), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7742 ( .A1(n9435), .A2(n6015), .ZN(n6016) );
  INV_X1 U7743 ( .A(n9435), .ZN(n9277) );
  INV_X1 U7744 ( .A(n9289), .ZN(n6015) );
  NAND2_X1 U7745 ( .A1(n7402), .A2(n6056), .ZN(n6024) );
  NAND2_X1 U7746 ( .A1(n6017), .A2(n6126), .ZN(n6018) );
  AOI22_X1 U7747 ( .A1(n6022), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6278), .B2(
        n6021), .ZN(n6023) );
  INV_X1 U7748 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U7749 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  AND2_X1 U7750 ( .A1(n6034), .A2(n6027), .ZN(n9267) );
  NAND2_X1 U7751 ( .A1(n9267), .A2(n5831), .ZN(n6031) );
  NAND2_X1 U7752 ( .A1(n6251), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7753 ( .A1(n4386), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7754 ( .A1(n6210), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7755 ( .A1(n9432), .A2(n9247), .ZN(n9242) );
  NAND2_X1 U7756 ( .A1(n6398), .A2(n9242), .ZN(n9255) );
  NAND2_X1 U7757 ( .A1(n7571), .A2(n6056), .ZN(n6033) );
  OR2_X1 U7758 ( .A1(n6248), .A2(n7607), .ZN(n6032) );
  NAND2_X1 U7759 ( .A1(n6034), .A2(n8839), .ZN(n6035) );
  AND2_X1 U7760 ( .A1(n6041), .A2(n6035), .ZN(n9235) );
  NAND2_X1 U7761 ( .A1(n9235), .A2(n5831), .ZN(n6038) );
  AOI22_X1 U7762 ( .A1(n4386), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6251), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7763 ( .A1(n6210), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7764 ( .A1(n9425), .A2(n8774), .ZN(n6401) );
  INV_X1 U7765 ( .A(n9425), .ZN(n9237) );
  NAND2_X1 U7766 ( .A1(n7766), .A2(n6056), .ZN(n6040) );
  OR2_X1 U7767 ( .A1(n5841), .A2(n7770), .ZN(n6039) );
  INV_X1 U7768 ( .A(n9420), .ZN(n9219) );
  INV_X1 U7769 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U7770 ( .A1(n6041), .A2(n8772), .ZN(n6042) );
  NAND2_X1 U7771 ( .A1(n6050), .A2(n6042), .ZN(n9216) );
  INV_X1 U7772 ( .A(n6043), .ZN(n6073) );
  OR2_X1 U7773 ( .A1(n9216), .A2(n6073), .ZN(n6046) );
  AOI22_X1 U7774 ( .A1(n4386), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6251), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7775 ( .A1(n6210), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7776 ( .A1(n9219), .A2(n9248), .ZN(n6047) );
  INV_X1 U7777 ( .A(n9248), .ZN(n8918) );
  NAND2_X1 U7778 ( .A1(n8441), .A2(n6056), .ZN(n6049) );
  OR2_X1 U7779 ( .A1(n6248), .A2(n8449), .ZN(n6048) );
  XNOR2_X1 U7780 ( .A(n6050), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n9202) );
  INV_X1 U7781 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7782 ( .A1(n6210), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7783 ( .A1(n6251), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7784 ( .C1(n6120), .C2(n6053), .A(n6052), .B(n6051), .ZN(n6054)
         );
  AOI21_X1 U7785 ( .B1(n9202), .B2(n5831), .A(n6054), .ZN(n8773) );
  NAND2_X1 U7786 ( .A1(n9415), .A2(n8773), .ZN(n6394) );
  NAND2_X1 U7787 ( .A1(n9409), .A2(n9164), .ZN(n6392) );
  NAND2_X1 U7788 ( .A1(n9192), .A2(n9206), .ZN(n6285) );
  NOR2_X1 U7789 ( .A1(n6248), .A2(n8408), .ZN(n6055) );
  AOI21_X2 U7790 ( .B1(n8395), .B2(n6056), .A(n6055), .ZN(n9172) );
  INV_X1 U7791 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U7792 ( .A1(n6058), .A2(n8832), .ZN(n6059) );
  NAND2_X1 U7793 ( .A1(n6071), .A2(n6059), .ZN(n9169) );
  INV_X1 U7794 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7795 ( .A1(n4386), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7796 ( .A1(n6251), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6060) );
  OAI211_X1 U7797 ( .C1(n6062), .C2(n5797), .A(n6061), .B(n6060), .ZN(n6063)
         );
  INV_X1 U7798 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7799 ( .A1(n6065), .A2(n6064), .ZN(n9181) );
  AND2_X1 U7800 ( .A1(n9172), .A2(n9181), .ZN(n6410) );
  INV_X1 U7801 ( .A(n6410), .ZN(n6200) );
  INV_X1 U7802 ( .A(n9172), .ZN(n9404) );
  INV_X1 U7803 ( .A(n9181), .ZN(n6066) );
  INV_X1 U7804 ( .A(n6411), .ZN(n6067) );
  NAND2_X1 U7805 ( .A1(n6200), .A2(n6067), .ZN(n9173) );
  INV_X1 U7806 ( .A(n9173), .ZN(n9162) );
  NAND2_X1 U7807 ( .A1(n8432), .A2(n6056), .ZN(n6069) );
  OR2_X1 U7808 ( .A1(n6248), .A2(n8437), .ZN(n6068) );
  INV_X1 U7809 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7810 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  NAND2_X1 U7811 ( .A1(n6083), .A2(n6072), .ZN(n9155) );
  INV_X1 U7812 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7813 ( .A1(n6251), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7814 ( .A1(n6210), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6074) );
  OAI211_X1 U7815 ( .C1(n6120), .C2(n6076), .A(n6075), .B(n6074), .ZN(n6077)
         );
  INV_X1 U7816 ( .A(n6077), .ZN(n6078) );
  NAND2_X1 U7817 ( .A1(n8438), .A2(n6056), .ZN(n6082) );
  OR2_X1 U7818 ( .A1(n5841), .A2(n9509), .ZN(n6081) );
  INV_X1 U7819 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U7820 ( .A1(n6083), .A2(n8049), .ZN(n6084) );
  NAND2_X1 U7821 ( .A1(n6104), .A2(n6084), .ZN(n8890) );
  INV_X1 U7822 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8188) );
  NAND2_X1 U7823 ( .A1(n6251), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7824 ( .A1(n6210), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6085) );
  OAI211_X1 U7825 ( .C1(n6120), .C2(n8188), .A(n6086), .B(n6085), .ZN(n6087)
         );
  AOI21_X1 U7826 ( .B1(n9139), .B2(n5831), .A(n6087), .ZN(n9114) );
  NOR2_X1 U7827 ( .A1(n9394), .A2(n9114), .ZN(n6416) );
  INV_X1 U7828 ( .A(n6416), .ZN(n6088) );
  NAND2_X1 U7829 ( .A1(n9394), .A2(n9114), .ZN(n6418) );
  INV_X1 U7830 ( .A(n9114), .ZN(n8916) );
  NAND2_X1 U7831 ( .A1(n9504), .A2(n6056), .ZN(n6090) );
  OR2_X1 U7832 ( .A1(n6248), .A2(n9505), .ZN(n6089) );
  XNOR2_X1 U7833 ( .A(n6104), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U7834 ( .A1(n9124), .A2(n5831), .ZN(n6096) );
  INV_X1 U7835 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U7836 ( .A1(n4386), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7837 ( .A1(n6210), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6091) );
  OAI211_X1 U7838 ( .C1(n6093), .C2(n8026), .A(n6092), .B(n6091), .ZN(n6094)
         );
  INV_X1 U7839 ( .A(n6094), .ZN(n6095) );
  NAND2_X1 U7840 ( .A1(n9501), .A2(n6056), .ZN(n6099) );
  OR2_X1 U7841 ( .A1(n5841), .A2(n9502), .ZN(n6098) );
  INV_X1 U7842 ( .A(n6104), .ZN(n6101) );
  AND2_X1 U7843 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6100) );
  NAND2_X1 U7844 ( .A1(n6101), .A2(n6100), .ZN(n6178) );
  INV_X1 U7845 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6103) );
  INV_X1 U7846 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6102) );
  OAI21_X1 U7847 ( .B1(n6104), .B2(n6103), .A(n6102), .ZN(n6105) );
  NAND2_X1 U7848 ( .A1(n6251), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7849 ( .A1(n6210), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6106) );
  OAI211_X1 U7850 ( .C1(n6120), .C2(n6238), .A(n6107), .B(n6106), .ZN(n6108)
         );
  NAND2_X1 U7851 ( .A1(n6617), .A2(n9115), .ZN(n6422) );
  INV_X1 U7852 ( .A(n9115), .ZN(n8914) );
  OR2_X1 U7853 ( .A1(n6617), .A2(n8914), .ZN(n9385) );
  INV_X1 U7854 ( .A(n9385), .ZN(n9376) );
  INV_X1 U7855 ( .A(SI_28_), .ZN(n6111) );
  INV_X1 U7856 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8446) );
  INV_X1 U7857 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6113) );
  MUX2_X1 U7858 ( .A(n8446), .B(n6113), .S(n4393), .Z(n6242) );
  XNOR2_X1 U7859 ( .A(n6242), .B(SI_29_), .ZN(n6114) );
  NAND2_X1 U7860 ( .A1(n8465), .A2(n6056), .ZN(n6116) );
  OR2_X1 U7861 ( .A1(n6248), .A2(n8446), .ZN(n6115) );
  INV_X1 U7862 ( .A(n6178), .ZN(n6122) );
  INV_X1 U7863 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7864 ( .A1(n6210), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7865 ( .A1(n6251), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6117) );
  OAI211_X1 U7866 ( .C1(n6120), .C2(n6119), .A(n6118), .B(n6117), .ZN(n6121)
         );
  AOI21_X1 U7867 ( .B1(n6122), .B2(n6043), .A(n6121), .ZN(n6225) );
  NAND2_X1 U7868 ( .A1(n9378), .A2(n6225), .ZN(n6284) );
  INV_X1 U7869 ( .A(n9377), .ZN(n9386) );
  INV_X1 U7870 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6125) );
  INV_X1 U7871 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7872 ( .A1(n6129), .A2(n6128), .ZN(n6164) );
  XNOR2_X1 U7873 ( .A(n8410), .B(P2_B_REG_SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7874 ( .A1(n6133), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6134) );
  MUX2_X1 U7875 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6134), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6136) );
  NAND2_X1 U7876 ( .A1(n6136), .A2(n6135), .ZN(n8435) );
  NAND2_X1 U7877 ( .A1(n6137), .A2(n8435), .ZN(n6141) );
  NAND2_X1 U7878 ( .A1(n6135), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6139) );
  INV_X1 U7879 ( .A(n9512), .ZN(n6140) );
  AND2_X1 U7880 ( .A1(n8410), .A2(n9512), .ZN(n10348) );
  INV_X1 U7881 ( .A(n10348), .ZN(n6142) );
  OR2_X1 U7882 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  NAND2_X1 U7883 ( .A1(n6147), .A2(n6146), .ZN(n10345) );
  AND2_X1 U7884 ( .A1(n10345), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6148) );
  NOR4_X1 U7885 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6157) );
  NOR4_X1 U7886 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6156) );
  INV_X1 U7887 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10343) );
  INV_X1 U7888 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10341) );
  INV_X1 U7889 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10342) );
  INV_X1 U7890 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10344) );
  NAND4_X1 U7891 ( .A1(n10343), .A2(n10341), .A3(n10342), .A4(n10344), .ZN(
        n6154) );
  NOR4_X1 U7892 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6152) );
  NOR4_X1 U7893 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6151) );
  NOR4_X1 U7894 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6150) );
  NOR4_X1 U7895 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6149) );
  NAND4_X1 U7896 ( .A1(n6152), .A2(n6151), .A3(n6150), .A4(n6149), .ZN(n6153)
         );
  NOR4_X1 U7897 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6154), .A4(n6153), .ZN(n6155) );
  AND3_X1 U7898 ( .A1(n6157), .A2(n6156), .A3(n6155), .ZN(n6158) );
  NOR2_X1 U7899 ( .A1(n10338), .A2(n6158), .ZN(n6235) );
  NAND2_X1 U7900 ( .A1(n9512), .A2(n8435), .ZN(n10351) );
  NAND2_X1 U7901 ( .A1(n6159), .A2(n10351), .ZN(n6234) );
  NOR2_X1 U7902 ( .A1(n6235), .A2(n6234), .ZN(n6605) );
  XNOR2_X1 U7903 ( .A(n6163), .B(n6162), .ZN(n6202) );
  NAND2_X1 U7904 ( .A1(n6164), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6165) );
  INV_X1 U7905 ( .A(n7029), .ZN(n7206) );
  NAND2_X1 U7906 ( .A1(n6278), .A2(n8447), .ZN(n6167) );
  NAND2_X1 U7907 ( .A1(n6487), .A2(n8447), .ZN(n6170) );
  NOR2_X1 U7908 ( .A1(n7029), .A2(n6278), .ZN(n6169) );
  NAND2_X1 U7909 ( .A1(n6170), .A2(n6169), .ZN(n9318) );
  OR2_X1 U7910 ( .A1(n6487), .A2(n9154), .ZN(n7870) );
  NAND2_X1 U7911 ( .A1(n9318), .A2(n7870), .ZN(n10322) );
  INV_X1 U7912 ( .A(n10329), .ZN(n6171) );
  INV_X1 U7913 ( .A(n7622), .ZN(n7861) );
  INV_X1 U7914 ( .A(n10397), .ZN(n7886) );
  NAND2_X1 U7915 ( .A1(n7882), .A2(n7886), .ZN(n7826) );
  INV_X1 U7916 ( .A(n9465), .ZN(n8790) );
  INV_X1 U7917 ( .A(n9450), .ZN(n9341) );
  INV_X1 U7918 ( .A(n9445), .ZN(n9326) );
  NAND2_X1 U7919 ( .A1(n9265), .A2(n9237), .ZN(n9232) );
  AND2_X2 U7920 ( .A1(n6202), .A2(n7768), .ZN(n6229) );
  NAND2_X1 U7921 ( .A1(n9378), .A2(n4428), .ZN(n6174) );
  NAND3_X1 U7922 ( .A1(n4441), .A2(n10398), .A3(n6174), .ZN(n9380) );
  INV_X1 U7923 ( .A(n7657), .ZN(n6175) );
  NAND2_X1 U7924 ( .A1(n6175), .A2(n9154), .ZN(n7714) );
  NAND2_X1 U7925 ( .A1(n6168), .A2(n6229), .ZN(n10325) );
  INV_X1 U7926 ( .A(n10325), .ZN(n6176) );
  INV_X1 U7927 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6177) );
  OAI22_X1 U7928 ( .A1(n6178), .A2(n9359), .B1(n10335), .B2(n6177), .ZN(n6179)
         );
  AOI21_X1 U7929 ( .B1(n9378), .B2(n9300), .A(n6179), .ZN(n6180) );
  OAI21_X1 U7930 ( .B1(n9380), .B2(n7714), .A(n6180), .ZN(n6181) );
  INV_X1 U7931 ( .A(n6181), .ZN(n6220) );
  NAND2_X1 U7932 ( .A1(n7315), .A2(n10353), .ZN(n10314) );
  NAND2_X1 U7933 ( .A1(n6302), .A2(n10314), .ZN(n10311) );
  NAND2_X1 U7934 ( .A1(n7678), .A2(n6182), .ZN(n6183) );
  NAND2_X1 U7935 ( .A1(n6183), .A2(n6287), .ZN(n7726) );
  INV_X1 U7936 ( .A(n7726), .ZN(n6185) );
  NAND2_X1 U7937 ( .A1(n6185), .A2(n6184), .ZN(n7727) );
  NAND2_X1 U7938 ( .A1(n7727), .A2(n6290), .ZN(n7693) );
  INV_X1 U7939 ( .A(n6448), .ZN(n7694) );
  INV_X1 U7940 ( .A(n7868), .ZN(n7617) );
  NOR2_X1 U7941 ( .A1(n7617), .A2(n6291), .ZN(n6186) );
  NAND2_X1 U7942 ( .A1(n6346), .A2(n8309), .ZN(n6350) );
  INV_X1 U7943 ( .A(n6350), .ZN(n6188) );
  NAND2_X1 U7944 ( .A1(n9455), .A2(n8850), .ZN(n6189) );
  NAND2_X1 U7945 ( .A1(n6189), .A2(n9331), .ZN(n6194) );
  AND2_X1 U7946 ( .A1(n6357), .A2(n8850), .ZN(n6359) );
  INV_X1 U7947 ( .A(n6359), .ZN(n6190) );
  NAND2_X1 U7948 ( .A1(n6190), .A2(n9357), .ZN(n6191) );
  OAI211_X1 U7949 ( .C1(n8850), .C2(n6357), .A(n6365), .B(n6191), .ZN(n6192)
         );
  INV_X1 U7950 ( .A(n6192), .ZN(n6193) );
  NAND2_X1 U7951 ( .A1(n6195), .A2(n6368), .ZN(n9310) );
  INV_X1 U7952 ( .A(n6370), .ZN(n9315) );
  INV_X1 U7953 ( .A(n9286), .ZN(n6196) );
  OR2_X1 U7954 ( .A1(n9435), .A2(n9289), .ZN(n9259) );
  NAND2_X1 U7955 ( .A1(n9435), .A2(n9289), .ZN(n9240) );
  INV_X1 U7956 ( .A(n9240), .ZN(n6399) );
  NAND2_X1 U7957 ( .A1(n6398), .A2(n6399), .ZN(n6199) );
  XNOR2_X1 U7958 ( .A(n9420), .B(n8918), .ZN(n9222) );
  INV_X1 U7959 ( .A(n9222), .ZN(n9213) );
  NAND2_X1 U7960 ( .A1(n9420), .A2(n9248), .ZN(n6395) );
  NAND2_X1 U7961 ( .A1(n9145), .A2(n6458), .ZN(n9148) );
  INV_X1 U7962 ( .A(n9165), .ZN(n9131) );
  NOR2_X1 U7963 ( .A1(n9400), .A2(n9131), .ZN(n6414) );
  INV_X1 U7964 ( .A(n6414), .ZN(n6201) );
  INV_X1 U7965 ( .A(n8915), .ZN(n9132) );
  NOR2_X1 U7966 ( .A1(n9389), .A2(n9132), .ZN(n6425) );
  XNOR2_X1 U7967 ( .A(n6241), .B(n9377), .ZN(n6217) );
  AND2_X1 U7968 ( .A1(n6168), .A2(n6466), .ZN(n6280) );
  INV_X1 U7969 ( .A(n6484), .ZN(n6203) );
  NAND2_X1 U7970 ( .A1(n6205), .A2(n6204), .ZN(n6207) );
  NAND2_X1 U7971 ( .A1(n6207), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6206) );
  XNOR2_X1 U7972 ( .A(n6206), .B(P2_IR_REG_28__SCAN_IN), .ZN(n7222) );
  INV_X1 U7973 ( .A(n7222), .ZN(n9503) );
  AND2_X1 U7974 ( .A1(n6208), .A2(n6207), .ZN(n7221) );
  AND2_X1 U7975 ( .A1(n7221), .A2(P2_B_REG_SCAN_IN), .ZN(n6209) );
  NOR2_X1 U7976 ( .A1(n9312), .A2(n6209), .ZN(n8450) );
  NAND2_X1 U7977 ( .A1(n4385), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7978 ( .A1(n6251), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7979 ( .A1(n6210), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6211) );
  AND3_X1 U7980 ( .A1(n6213), .A2(n6212), .A3(n6211), .ZN(n6271) );
  INV_X1 U7981 ( .A(n6271), .ZN(n8912) );
  NAND2_X1 U7982 ( .A1(n8450), .A2(n8912), .ZN(n6214) );
  NAND2_X1 U7983 ( .A1(n6221), .A2(n5046), .ZN(P2_U3267) );
  NAND2_X1 U7984 ( .A1(n9387), .A2(n5050), .ZN(n9110) );
  NAND2_X1 U7985 ( .A1(n9110), .A2(n10393), .ZN(n6233) );
  OAI211_X1 U7986 ( .C1(n6224), .C2(n6461), .A(n6223), .B(n10313), .ZN(n6227)
         );
  INV_X1 U7987 ( .A(n6225), .ZN(n8913) );
  AOI22_X1 U7988 ( .A1(n8913), .A2(n10316), .B1(n10317), .B2(n8915), .ZN(n6226) );
  AND2_X1 U7989 ( .A1(n6227), .A2(n6226), .ZN(n9112) );
  NAND2_X1 U7990 ( .A1(n9123), .A2(n6617), .ZN(n6228) );
  AND2_X1 U7991 ( .A1(n4428), .A2(n6228), .ZN(n9104) );
  OR2_X1 U7992 ( .A1(n9154), .A2(n6485), .ZN(n6230) );
  NAND2_X2 U7993 ( .A1(n10325), .A2(n6230), .ZN(n10396) );
  AOI22_X1 U7994 ( .A1(n9104), .A2(n10398), .B1(n6617), .B2(n10396), .ZN(n6231) );
  INV_X1 U7995 ( .A(n6234), .ZN(n6236) );
  NAND2_X1 U7996 ( .A1(n10339), .A2(n6629), .ZN(n6477) );
  OR2_X1 U7997 ( .A1(n6625), .A2(n6477), .ZN(n6237) );
  NAND2_X1 U7998 ( .A1(n6480), .A2(n10423), .ZN(n6240) );
  OR2_X1 U7999 ( .A1(n10423), .A2(n6238), .ZN(n6239) );
  NAND2_X1 U8000 ( .A1(n6240), .A2(n6239), .ZN(P2_U3548) );
  INV_X1 U8001 ( .A(n6257), .ZN(n6259) );
  INV_X1 U8002 ( .A(n6242), .ZN(n6245) );
  NOR2_X1 U8003 ( .A1(n6245), .A2(SI_29_), .ZN(n6243) );
  NAND2_X1 U8004 ( .A1(n6245), .A2(SI_29_), .ZN(n6246) );
  MUX2_X1 U8005 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4394), .Z(n6262) );
  XNOR2_X1 U8006 ( .A(n6262), .B(SI_30_), .ZN(n6247) );
  NAND2_X1 U8007 ( .A1(n8731), .A2(n6056), .ZN(n6250) );
  INV_X1 U8008 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8732) );
  OR2_X1 U8009 ( .A1(n6248), .A2(n8732), .ZN(n6249) );
  OR2_X1 U8010 ( .A1(n9100), .A2(n6271), .ZN(n6431) );
  INV_X1 U8011 ( .A(n6431), .ZN(n6256) );
  NAND2_X1 U8012 ( .A1(n4386), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U8013 ( .A1(n6210), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U8014 ( .A1(n6251), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6252) );
  AND3_X1 U8015 ( .A1(n6254), .A2(n6253), .A3(n6252), .ZN(n6273) );
  INV_X1 U8016 ( .A(n6273), .ZN(n8451) );
  OR2_X1 U8017 ( .A1(n8451), .A2(n7768), .ZN(n6255) );
  OAI21_X1 U8018 ( .B1(n6259), .B2(n9100), .A(n6258), .ZN(n6276) );
  INV_X1 U8019 ( .A(n6262), .ZN(n6261) );
  INV_X1 U8020 ( .A(SI_30_), .ZN(n6260) );
  NOR2_X1 U8021 ( .A1(n6261), .A2(n6260), .ZN(n6263) );
  MUX2_X1 U8022 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4393), .Z(n6265) );
  INV_X1 U8023 ( .A(SI_31_), .ZN(n8102) );
  XNOR2_X1 U8024 ( .A(n6265), .B(n8102), .ZN(n6266) );
  XNOR2_X1 U8025 ( .A(n6267), .B(n6266), .ZN(n9495) );
  NAND2_X1 U8026 ( .A1(n9495), .A2(n6056), .ZN(n6270) );
  INV_X1 U8027 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6268) );
  OR2_X1 U8028 ( .A1(n5841), .A2(n6268), .ZN(n6269) );
  OR2_X1 U8029 ( .A1(n9369), .A2(n6273), .ZN(n6436) );
  AND2_X1 U8030 ( .A1(n9100), .A2(n6271), .ZN(n6429) );
  INV_X1 U8031 ( .A(n6429), .ZN(n6272) );
  NAND2_X1 U8032 ( .A1(n6436), .A2(n6272), .ZN(n6464) );
  INV_X1 U8033 ( .A(n6464), .ZN(n6275) );
  NAND2_X1 U8034 ( .A1(n9369), .A2(n6273), .ZN(n6434) );
  INV_X1 U8035 ( .A(n6434), .ZN(n6274) );
  AOI21_X1 U8036 ( .B1(n6276), .B2(n6275), .A(n6274), .ZN(n6277) );
  XNOR2_X1 U8037 ( .A(n6277), .B(n9154), .ZN(n6283) );
  NOR2_X1 U8038 ( .A1(n10345), .A2(P2_U3152), .ZN(n7032) );
  OAI21_X1 U8039 ( .B1(n7314), .B2(n6280), .A(n7032), .ZN(n6281) );
  INV_X1 U8040 ( .A(n6281), .ZN(n6282) );
  INV_X1 U8041 ( .A(n6284), .ZN(n6430) );
  INV_X1 U8042 ( .A(n6285), .ZN(n6409) );
  INV_X1 U8043 ( .A(n9331), .ZN(n6286) );
  NOR4_X1 U8044 ( .A1(n9364), .A2(n4802), .A3(n6286), .A4(n6435), .ZN(n6364)
         );
  NAND2_X1 U8045 ( .A1(n6290), .A2(n6288), .ZN(n6442) );
  NOR2_X1 U8046 ( .A1(n6442), .A2(n6441), .ZN(n6289) );
  AOI21_X1 U8047 ( .B1(n6311), .B2(n6290), .A(n6289), .ZN(n6292) );
  OAI21_X1 U8048 ( .B1(n6292), .B2(n6291), .A(n4583), .ZN(n6299) );
  INV_X1 U8049 ( .A(n6311), .ZN(n6297) );
  INV_X1 U8050 ( .A(n10353), .ZN(n7663) );
  NAND2_X1 U8051 ( .A1(n6293), .A2(n7663), .ZN(n6300) );
  AND2_X1 U8052 ( .A1(n6300), .A2(n6466), .ZN(n6294) );
  OAI211_X1 U8053 ( .C1(n10311), .C2(n6294), .A(n6303), .B(n10309), .ZN(n6295)
         );
  NAND3_X1 U8054 ( .A1(n6295), .A2(n7746), .A3(n4583), .ZN(n6296) );
  NAND3_X1 U8055 ( .A1(n6297), .A2(n7745), .A3(n6296), .ZN(n6298) );
  NAND2_X1 U8056 ( .A1(n6299), .A2(n6298), .ZN(n6306) );
  NAND2_X1 U8057 ( .A1(n10309), .A2(n6300), .ZN(n6301) );
  NAND3_X1 U8058 ( .A1(n7746), .A2(n6302), .A3(n6301), .ZN(n6304) );
  NAND3_X1 U8059 ( .A1(n6304), .A2(n6435), .A3(n6303), .ZN(n6305) );
  NAND3_X1 U8060 ( .A1(n6306), .A2(n6312), .A3(n6305), .ZN(n6317) );
  INV_X1 U8061 ( .A(n6307), .ZN(n6309) );
  AND2_X1 U8062 ( .A1(n6309), .A2(n6308), .ZN(n6446) );
  AOI21_X1 U8063 ( .B1(n6311), .B2(n6310), .A(n6446), .ZN(n6314) );
  INV_X1 U8064 ( .A(n6312), .ZN(n6313) );
  OAI21_X1 U8065 ( .B1(n6314), .B2(n6313), .A(n6435), .ZN(n6316) );
  OAI21_X1 U8066 ( .B1(n7618), .B2(n4583), .A(n7868), .ZN(n6315) );
  INV_X1 U8067 ( .A(n6318), .ZN(n6319) );
  NOR3_X1 U8068 ( .A1(n6334), .A2(n6319), .A3(n7873), .ZN(n6321) );
  NOR2_X1 U8069 ( .A1(n6321), .A2(n4793), .ZN(n6326) );
  INV_X1 U8070 ( .A(n6322), .ZN(n6323) );
  NOR2_X1 U8071 ( .A1(n6324), .A2(n6323), .ZN(n6325) );
  MUX2_X1 U8072 ( .A(n6326), .B(n6325), .S(n4583), .Z(n6327) );
  NAND2_X1 U8073 ( .A1(n6327), .A2(n6329), .ZN(n6344) );
  INV_X1 U8074 ( .A(n6329), .ZN(n6330) );
  MUX2_X1 U8075 ( .A(n6331), .B(n6330), .S(n4583), .Z(n6333) );
  NOR2_X1 U8076 ( .A1(n6333), .A2(n6332), .ZN(n6343) );
  INV_X1 U8077 ( .A(n6334), .ZN(n6335) );
  NAND4_X1 U8078 ( .A1(n6343), .A2(n6187), .A3(n6336), .A4(n6335), .ZN(n6338)
         );
  NAND3_X1 U8079 ( .A1(n6338), .A2(n8309), .A3(n6337), .ZN(n6341) );
  NAND2_X1 U8080 ( .A1(n6345), .A2(n6339), .ZN(n6340) );
  MUX2_X1 U8081 ( .A(n6341), .B(n6340), .S(n6435), .Z(n6342) );
  NOR2_X1 U8082 ( .A1(n9334), .A2(n4583), .ZN(n6354) );
  NAND2_X1 U8083 ( .A1(n9334), .A2(n4583), .ZN(n6356) );
  NAND3_X1 U8084 ( .A1(n8382), .A2(n6347), .A3(n6356), .ZN(n6348) );
  AOI211_X1 U8085 ( .C1(n6354), .C2(n9455), .A(n6348), .B(n6360), .ZN(n6349)
         );
  INV_X1 U8086 ( .A(n6356), .ZN(n6353) );
  INV_X1 U8087 ( .A(n6357), .ZN(n6352) );
  MUX2_X1 U8088 ( .A(n6435), .B(n6353), .S(n6352), .Z(n6355) );
  NOR3_X1 U8089 ( .A1(n6355), .A2(n9357), .A3(n6354), .ZN(n6362) );
  OAI211_X1 U8090 ( .C1(n6357), .C2(n6435), .A(n9357), .B(n6356), .ZN(n6358)
         );
  AOI21_X1 U8091 ( .B1(n6359), .B2(n6435), .A(n6358), .ZN(n6361) );
  INV_X1 U8092 ( .A(n6360), .ZN(n9345) );
  OAI21_X1 U8093 ( .B1(n6362), .B2(n6361), .A(n9345), .ZN(n6363) );
  INV_X1 U8094 ( .A(n6365), .ZN(n6366) );
  NAND2_X1 U8095 ( .A1(n6366), .A2(n6435), .ZN(n6367) );
  OAI21_X1 U8096 ( .B1(n6435), .B2(n6368), .A(n6367), .ZN(n6369) );
  INV_X1 U8097 ( .A(n6371), .ZN(n6381) );
  NOR2_X1 U8098 ( .A1(n9335), .A2(n4583), .ZN(n6372) );
  AND2_X1 U8099 ( .A1(n9445), .A2(n6372), .ZN(n6376) );
  OAI21_X1 U8100 ( .B1(n9290), .B2(n6435), .A(n9326), .ZN(n6375) );
  INV_X1 U8101 ( .A(n6372), .ZN(n6373) );
  OAI21_X1 U8102 ( .B1(n9280), .B2(n6373), .A(n9445), .ZN(n6374) );
  AOI22_X1 U8103 ( .A1(n6376), .A2(n9442), .B1(n6375), .B2(n6374), .ZN(n6380)
         );
  AND2_X1 U8104 ( .A1(n9280), .A2(n4583), .ZN(n6378) );
  OAI21_X1 U8105 ( .B1(n9280), .B2(n4583), .A(n9442), .ZN(n6377) );
  OAI21_X1 U8106 ( .B1(n6378), .B2(n9442), .A(n6377), .ZN(n6379) );
  OAI211_X1 U8107 ( .C1(n6381), .C2(n6380), .A(n9259), .B(n6379), .ZN(n6382)
         );
  INV_X1 U8108 ( .A(n9259), .ZN(n6383) );
  NAND2_X1 U8109 ( .A1(n6385), .A2(n6384), .ZN(n6386) );
  NAND3_X1 U8110 ( .A1(n6386), .A2(n6395), .A3(n6401), .ZN(n6387) );
  NAND2_X1 U8111 ( .A1(n9219), .A2(n8918), .ZN(n6403) );
  NAND4_X1 U8112 ( .A1(n6387), .A2(n6435), .A3(n6388), .A4(n6403), .ZN(n6391)
         );
  MUX2_X1 U8113 ( .A(n6394), .B(n6388), .S(n4583), .Z(n6389) );
  INV_X1 U8114 ( .A(n6392), .ZN(n6393) );
  OAI21_X1 U8115 ( .B1(n6410), .B2(n6393), .A(n6435), .ZN(n6408) );
  INV_X1 U8116 ( .A(n6394), .ZN(n6397) );
  INV_X1 U8117 ( .A(n6395), .ZN(n6396) );
  NOR3_X1 U8118 ( .A1(n6397), .A2(n6396), .A3(n6435), .ZN(n6407) );
  OAI21_X1 U8119 ( .B1(n6400), .B2(n6399), .A(n6398), .ZN(n6402) );
  NAND3_X1 U8120 ( .A1(n6402), .A2(n6401), .A3(n9242), .ZN(n6405) );
  NAND3_X1 U8121 ( .A1(n6405), .A2(n6404), .A3(n6403), .ZN(n6406) );
  MUX2_X1 U8122 ( .A(n6411), .B(n6410), .S(n4583), .Z(n6412) );
  OAI21_X1 U8123 ( .B1(n9152), .B2(n9165), .A(n6418), .ZN(n6413) );
  NOR2_X1 U8124 ( .A1(n6416), .A2(n6414), .ZN(n6415) );
  OAI22_X1 U8125 ( .A1(n6417), .A2(n6416), .B1(n4583), .B2(n6415), .ZN(n6420)
         );
  NAND3_X1 U8126 ( .A1(n9389), .A2(n9132), .A3(n4583), .ZN(n6421) );
  INV_X1 U8127 ( .A(n6424), .ZN(n6426) );
  OAI21_X1 U8128 ( .B1(n6426), .B2(n6425), .A(n6435), .ZN(n6428) );
  INV_X1 U8129 ( .A(n6617), .ZN(n9108) );
  NOR3_X1 U8130 ( .A1(n9108), .A2(n8914), .A3(n4583), .ZN(n6427) );
  NAND2_X1 U8131 ( .A1(n6434), .A2(n6431), .ZN(n6463) );
  NOR2_X1 U8132 ( .A1(n6463), .A2(n5018), .ZN(n6433) );
  NAND3_X1 U8133 ( .A1(n6464), .A2(n6435), .A3(n6434), .ZN(n6438) );
  INV_X1 U8134 ( .A(n6436), .ZN(n6437) );
  INV_X1 U8135 ( .A(n6474), .ZN(n6469) );
  NAND2_X1 U8136 ( .A1(n9259), .A2(n9240), .ZN(n9278) );
  INV_X1 U8137 ( .A(n8382), .ZN(n6452) );
  NOR3_X1 U8138 ( .A1(n6440), .A2(n6441), .A3(n6173), .ZN(n6445) );
  INV_X1 U8139 ( .A(n6442), .ZN(n6444) );
  INV_X1 U8140 ( .A(n6443), .ZN(n10321) );
  OAI21_X1 U8141 ( .B1(n6293), .B2(n10353), .A(n5827), .ZN(n7659) );
  NAND4_X1 U8142 ( .A1(n6445), .A2(n6444), .A3(n10321), .A4(n7659), .ZN(n6449)
         );
  INV_X1 U8143 ( .A(n6446), .ZN(n6447) );
  NAND4_X1 U8144 ( .A1(n7924), .A2(n6187), .A3(n7829), .A4(n6450), .ZN(n6451)
         );
  NAND4_X1 U8145 ( .A1(n9315), .A2(n9345), .A3(n6454), .A4(n6453), .ZN(n6455)
         );
  NOR4_X1 U8146 ( .A1(n9255), .A2(n9278), .A3(n9292), .A4(n6455), .ZN(n6456)
         );
  NAND4_X1 U8147 ( .A1(n6456), .A2(n9241), .A3(n9199), .A4(n9222), .ZN(n6457)
         );
  NOR4_X1 U8148 ( .A1(n9137), .A2(n9184), .A3(n9173), .A4(n6457), .ZN(n6460)
         );
  NAND4_X1 U8149 ( .A1(n6461), .A2(n6460), .A3(n6459), .A4(n6458), .ZN(n6462)
         );
  XOR2_X1 U8150 ( .A(n9154), .B(n6465), .Z(n6467) );
  OAI22_X1 U8151 ( .A1(n6467), .A2(n6466), .B1(n6168), .B2(n6484), .ZN(n6468)
         );
  NAND3_X1 U8152 ( .A1(n6469), .A2(n6468), .A3(n7032), .ZN(n6476) );
  INV_X1 U8153 ( .A(n7032), .ZN(n8241) );
  NAND4_X1 U8154 ( .A1(n10339), .A2(n6626), .A3(n7221), .A4(n10317), .ZN(n6470) );
  OAI211_X1 U8155 ( .C1(n6471), .C2(n8241), .A(n6470), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6472) );
  INV_X1 U8156 ( .A(n6472), .ZN(n6473) );
  INV_X1 U8157 ( .A(n6477), .ZN(n7311) );
  NAND2_X1 U8158 ( .A1(n6625), .A2(n7311), .ZN(n6478) );
  NAND2_X1 U8159 ( .A1(n6480), .A2(n10407), .ZN(n6483) );
  INV_X1 U8160 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6481) );
  OR2_X1 U8161 ( .A1(n10407), .A2(n6481), .ZN(n6482) );
  NAND2_X1 U8162 ( .A1(n6483), .A2(n6482), .ZN(P2_U3516) );
  NOR2_X1 U8163 ( .A1(n7709), .A2(n6496), .ZN(n7341) );
  INV_X1 U8164 ( .A(n7341), .ZN(n6489) );
  XNOR2_X1 U8165 ( .A(n4388), .B(n6488), .ZN(n6493) );
  NAND2_X1 U8166 ( .A1(n6489), .A2(n7340), .ZN(n7343) );
  NAND2_X1 U8167 ( .A1(n10320), .A2(n7656), .ZN(n7317) );
  OR2_X1 U8168 ( .A1(n6588), .A2(n10353), .ZN(n6490) );
  NAND2_X1 U8169 ( .A1(n7317), .A2(n6490), .ZN(n7342) );
  INV_X2 U8170 ( .A(n5793), .ZN(n10315) );
  NAND2_X1 U8171 ( .A1(n7656), .A2(n10315), .ZN(n6492) );
  XNOR2_X1 U8172 ( .A(n4389), .B(n10365), .ZN(n6491) );
  NAND2_X1 U8173 ( .A1(n6492), .A2(n6491), .ZN(n7344) );
  NAND3_X1 U8174 ( .A1(n7343), .A2(n7342), .A3(n7344), .ZN(n6495) );
  OR2_X1 U8175 ( .A1(n6492), .A2(n6491), .ZN(n7345) );
  NAND3_X1 U8176 ( .A1(n7344), .A2(n7341), .A3(n6493), .ZN(n6494) );
  NAND3_X1 U8177 ( .A1(n6495), .A2(n7345), .A3(n6494), .ZN(n7483) );
  OR2_X1 U8178 ( .A1(n7731), .A2(n6496), .ZN(n7524) );
  XNOR2_X1 U8179 ( .A(n4389), .B(n6497), .ZN(n7523) );
  NAND2_X1 U8180 ( .A1(n7524), .A2(n7523), .ZN(n6503) );
  NAND2_X1 U8181 ( .A1(n7656), .A2(n8930), .ZN(n6500) );
  XNOR2_X1 U8182 ( .A(n6588), .B(n7482), .ZN(n6499) );
  NAND2_X1 U8183 ( .A1(n6500), .A2(n6499), .ZN(n7484) );
  NAND2_X1 U8184 ( .A1(n7483), .A2(n6498), .ZN(n6505) );
  NOR2_X1 U8185 ( .A1(n6500), .A2(n6499), .ZN(n7521) );
  INV_X1 U8186 ( .A(n7523), .ZN(n6502) );
  INV_X1 U8187 ( .A(n7524), .ZN(n6501) );
  AOI22_X1 U8188 ( .A1(n6503), .A2(n7521), .B1(n6502), .B2(n6501), .ZN(n6504)
         );
  NAND2_X1 U8189 ( .A1(n6505), .A2(n6504), .ZN(n7496) );
  INV_X1 U8190 ( .A(n7656), .ZN(n6510) );
  NOR2_X1 U8191 ( .A1(n7536), .A2(n6510), .ZN(n6507) );
  XNOR2_X1 U8192 ( .A(n6588), .B(n7738), .ZN(n6506) );
  NAND2_X1 U8193 ( .A1(n6507), .A2(n6506), .ZN(n6509) );
  AND2_X1 U8194 ( .A1(n6509), .A2(n6508), .ZN(n7495) );
  NAND2_X1 U8195 ( .A1(n7496), .A2(n7495), .ZN(n7494) );
  NAND2_X1 U8196 ( .A1(n7494), .A2(n6509), .ZN(n7534) );
  INV_X1 U8197 ( .A(n7534), .ZN(n6512) );
  XNOR2_X1 U8198 ( .A(n7701), .B(n6603), .ZN(n6514) );
  OR2_X1 U8199 ( .A1(n7730), .A2(n6510), .ZN(n6513) );
  XNOR2_X1 U8200 ( .A(n6514), .B(n6513), .ZN(n7535) );
  NAND2_X1 U8201 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  XNOR2_X1 U8202 ( .A(n7622), .B(n4389), .ZN(n6516) );
  NOR2_X1 U8203 ( .A1(n7876), .A2(n6510), .ZN(n6517) );
  NAND2_X1 U8204 ( .A1(n6516), .A2(n6517), .ZN(n6521) );
  INV_X1 U8205 ( .A(n6516), .ZN(n6519) );
  INV_X1 U8206 ( .A(n6517), .ZN(n6518) );
  NAND2_X1 U8207 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  AND2_X1 U8208 ( .A1(n6521), .A2(n6520), .ZN(n7502) );
  XNOR2_X1 U8209 ( .A(n10397), .B(n6598), .ZN(n6522) );
  NOR2_X1 U8210 ( .A1(n7832), .A2(n7314), .ZN(n6523) );
  NAND2_X1 U8211 ( .A1(n6522), .A2(n6523), .ZN(n6527) );
  INV_X1 U8212 ( .A(n6522), .ZN(n6525) );
  INV_X1 U8213 ( .A(n6523), .ZN(n6524) );
  NAND2_X1 U8214 ( .A1(n6525), .A2(n6524), .ZN(n6526) );
  AND2_X1 U8215 ( .A1(n6527), .A2(n6526), .ZN(n7475) );
  NAND2_X1 U8216 ( .A1(n7476), .A2(n7475), .ZN(n7474) );
  NAND2_X1 U8217 ( .A1(n7474), .A2(n6527), .ZN(n7610) );
  XNOR2_X1 U8218 ( .A(n7828), .B(n6598), .ZN(n6529) );
  NAND2_X1 U8219 ( .A1(n7656), .A2(n8924), .ZN(n6528) );
  XNOR2_X1 U8220 ( .A(n6529), .B(n6528), .ZN(n7611) );
  XNOR2_X1 U8221 ( .A(n8229), .B(n6603), .ZN(n6530) );
  NOR2_X1 U8222 ( .A1(n7831), .A2(n7314), .ZN(n6531) );
  XNOR2_X1 U8223 ( .A(n6530), .B(n6531), .ZN(n7782) );
  INV_X1 U8224 ( .A(n6530), .ZN(n6532) );
  NAND2_X1 U8225 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  XNOR2_X1 U8226 ( .A(n9470), .B(n6598), .ZN(n6534) );
  NOR2_X1 U8227 ( .A1(n8785), .A2(n7314), .ZN(n6535) );
  NAND2_X1 U8228 ( .A1(n6534), .A2(n6535), .ZN(n8868) );
  NAND2_X1 U8229 ( .A1(n8870), .A2(n8868), .ZN(n6538) );
  INV_X1 U8230 ( .A(n6534), .ZN(n6537) );
  INV_X1 U8231 ( .A(n6535), .ZN(n6536) );
  NAND2_X1 U8232 ( .A1(n6537), .A2(n6536), .ZN(n8869) );
  NAND2_X1 U8233 ( .A1(n6538), .A2(n8869), .ZN(n8780) );
  XNOR2_X1 U8234 ( .A(n9465), .B(n6603), .ZN(n6540) );
  OR2_X1 U8235 ( .A1(n6539), .A2(n7314), .ZN(n6541) );
  NAND2_X1 U8236 ( .A1(n6540), .A2(n6541), .ZN(n6545) );
  INV_X1 U8237 ( .A(n6540), .ZN(n6543) );
  INV_X1 U8238 ( .A(n6541), .ZN(n6542) );
  NAND2_X1 U8239 ( .A1(n6543), .A2(n6542), .ZN(n6544) );
  AND2_X1 U8240 ( .A1(n6545), .A2(n6544), .ZN(n8781) );
  NAND2_X1 U8241 ( .A1(n8780), .A2(n8781), .ZN(n8779) );
  NAND2_X1 U8242 ( .A1(n8779), .A2(n6545), .ZN(n8846) );
  XNOR2_X1 U8243 ( .A(n9460), .B(n6598), .ZN(n6547) );
  NOR2_X1 U8244 ( .A1(n8743), .A2(n7314), .ZN(n6546) );
  XNOR2_X1 U8245 ( .A(n6547), .B(n6546), .ZN(n8845) );
  XNOR2_X1 U8246 ( .A(n9455), .B(n6603), .ZN(n6548) );
  NAND2_X1 U8247 ( .A1(n7656), .A2(n9334), .ZN(n6549) );
  NAND2_X1 U8248 ( .A1(n6548), .A2(n6549), .ZN(n8803) );
  INV_X1 U8249 ( .A(n6548), .ZN(n6551) );
  INV_X1 U8250 ( .A(n6549), .ZN(n6550) );
  NAND2_X1 U8251 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  AND2_X1 U8252 ( .A1(n8803), .A2(n6552), .ZN(n8741) );
  INV_X1 U8253 ( .A(n8803), .ZN(n6554) );
  XNOR2_X1 U8254 ( .A(n9450), .B(n6598), .ZN(n8805) );
  NOR2_X1 U8255 ( .A1(n9311), .A2(n7314), .ZN(n6557) );
  NOR2_X1 U8256 ( .A1(n9290), .A2(n7314), .ZN(n6556) );
  XNOR2_X1 U8257 ( .A(n9445), .B(n6598), .ZN(n6555) );
  NOR2_X1 U8258 ( .A1(n6555), .A2(n6556), .ZN(n6561) );
  AOI21_X1 U8259 ( .B1(n6556), .B2(n6555), .A(n6561), .ZN(n8810) );
  INV_X1 U8260 ( .A(n8805), .ZN(n8807) );
  INV_X1 U8261 ( .A(n6557), .ZN(n8900) );
  NAND2_X1 U8262 ( .A1(n6560), .A2(n6559), .ZN(n8811) );
  INV_X1 U8263 ( .A(n6561), .ZN(n6562) );
  XNOR2_X1 U8264 ( .A(n9442), .B(n6598), .ZN(n6563) );
  NOR2_X1 U8265 ( .A1(n9313), .A2(n7314), .ZN(n6564) );
  XNOR2_X1 U8266 ( .A(n6563), .B(n6564), .ZN(n8819) );
  INV_X1 U8267 ( .A(n6563), .ZN(n6566) );
  INV_X1 U8268 ( .A(n6564), .ZN(n6565) );
  XNOR2_X1 U8269 ( .A(n9435), .B(n6603), .ZN(n6567) );
  NOR2_X1 U8270 ( .A1(n9289), .A2(n7314), .ZN(n6569) );
  XNOR2_X1 U8271 ( .A(n6567), .B(n6569), .ZN(n8879) );
  INV_X1 U8272 ( .A(n6567), .ZN(n6568) );
  NOR2_X1 U8273 ( .A1(n9247), .A2(n7314), .ZN(n6571) );
  XNOR2_X1 U8274 ( .A(n9432), .B(n6598), .ZN(n6570) );
  NOR2_X1 U8275 ( .A1(n6570), .A2(n6571), .ZN(n6572) );
  AOI21_X1 U8276 ( .B1(n6571), .B2(n6570), .A(n6572), .ZN(n8757) );
  INV_X1 U8277 ( .A(n6572), .ZN(n6573) );
  XNOR2_X1 U8278 ( .A(n9425), .B(n6598), .ZN(n6574) );
  NOR2_X1 U8279 ( .A1(n8774), .A2(n7314), .ZN(n6575) );
  XNOR2_X1 U8280 ( .A(n6574), .B(n6575), .ZN(n8837) );
  INV_X1 U8281 ( .A(n6574), .ZN(n6577) );
  INV_X1 U8282 ( .A(n6575), .ZN(n6576) );
  XNOR2_X1 U8283 ( .A(n9420), .B(n6603), .ZN(n6582) );
  NOR2_X1 U8284 ( .A1(n9248), .A2(n7314), .ZN(n6580) );
  XNOR2_X1 U8285 ( .A(n6582), .B(n6580), .ZN(n8770) );
  NAND2_X1 U8286 ( .A1(n8771), .A2(n8770), .ZN(n8855) );
  XNOR2_X1 U8287 ( .A(n9415), .B(n6603), .ZN(n6578) );
  INV_X1 U8288 ( .A(n8773), .ZN(n9224) );
  NAND2_X1 U8289 ( .A1(n9224), .A2(n7656), .ZN(n8856) );
  NAND2_X1 U8290 ( .A1(n6578), .A2(n8856), .ZN(n6587) );
  INV_X1 U8291 ( .A(n6578), .ZN(n8857) );
  INV_X1 U8292 ( .A(n6582), .ZN(n6579) );
  NAND2_X1 U8293 ( .A1(n6579), .A2(n6580), .ZN(n8854) );
  NAND2_X1 U8294 ( .A1(n8854), .A2(n8856), .ZN(n6584) );
  INV_X1 U8295 ( .A(n6580), .ZN(n6581) );
  NOR3_X1 U8296 ( .A1(n6582), .A2(n8773), .A3(n6581), .ZN(n6583) );
  AOI21_X2 U8297 ( .B1(n8857), .B2(n6584), .A(n6583), .ZN(n6585) );
  XNOR2_X1 U8298 ( .A(n9409), .B(n6598), .ZN(n6591) );
  XNOR2_X2 U8299 ( .A(n6589), .B(n6591), .ZN(n8827) );
  XNOR2_X1 U8300 ( .A(n9172), .B(n6598), .ZN(n8829) );
  INV_X1 U8301 ( .A(n8829), .ZN(n6593) );
  AND2_X1 U8302 ( .A1(n9164), .A2(n7656), .ZN(n8826) );
  OAI21_X1 U8303 ( .B1(n6593), .B2(n9181), .A(n8826), .ZN(n6590) );
  INV_X1 U8304 ( .A(n6590), .ZN(n6594) );
  NAND2_X1 U8305 ( .A1(n9181), .A2(n7656), .ZN(n8828) );
  INV_X1 U8306 ( .A(n8828), .ZN(n6592) );
  AOI21_X2 U8307 ( .B1(n8827), .B2(n6594), .A(n4404), .ZN(n8794) );
  XNOR2_X1 U8308 ( .A(n9152), .B(n6598), .ZN(n8792) );
  NAND2_X1 U8309 ( .A1(n9165), .A2(n7656), .ZN(n8791) );
  XNOR2_X1 U8310 ( .A(n9394), .B(n6598), .ZN(n6596) );
  NOR2_X1 U8311 ( .A1(n9114), .A2(n7314), .ZN(n6595) );
  NAND2_X1 U8312 ( .A1(n6596), .A2(n6595), .ZN(n6597) );
  OAI21_X1 U8313 ( .B1(n6596), .B2(n6595), .A(n6597), .ZN(n8885) );
  XNOR2_X1 U8314 ( .A(n9389), .B(n6598), .ZN(n6600) );
  INV_X1 U8315 ( .A(n6600), .ZN(n6602) );
  AND2_X1 U8316 ( .A1(n8915), .A2(n7656), .ZN(n6599) );
  INV_X1 U8317 ( .A(n6599), .ZN(n6601) );
  AOI21_X1 U8318 ( .B1(n6602), .B2(n6601), .A(n6622), .ZN(n8735) );
  OR2_X1 U8319 ( .A1(n9115), .A2(n7314), .ZN(n6604) );
  XNOR2_X1 U8320 ( .A(n6604), .B(n6603), .ZN(n6618) );
  INV_X1 U8321 ( .A(n6618), .ZN(n6615) );
  INV_X1 U8322 ( .A(n6605), .ZN(n6606) );
  OR2_X1 U8323 ( .A1(n6625), .A2(n6606), .ZN(n6609) );
  INV_X1 U8324 ( .A(n6607), .ZN(n6608) );
  NAND2_X1 U8325 ( .A1(n6609), .A2(n6608), .ZN(n7312) );
  AND2_X1 U8326 ( .A1(n10339), .A2(n10396), .ZN(n6610) );
  NOR2_X1 U8327 ( .A1(n10396), .A2(n7029), .ZN(n6611) );
  NAND2_X1 U8328 ( .A1(n6623), .A2(n6611), .ZN(n6612) );
  NOR2_X2 U8329 ( .A1(n6625), .A2(n6612), .ZN(n8888) );
  AOI21_X1 U8330 ( .B1(n6617), .B2(n8908), .A(n8888), .ZN(n6620) );
  INV_X1 U8331 ( .A(n6620), .ZN(n6614) );
  NAND3_X1 U8332 ( .A1(n6617), .A2(n10390), .A3(n6615), .ZN(n6613) );
  OAI211_X1 U8333 ( .C1(n6615), .C2(n6617), .A(n6614), .B(n6613), .ZN(n6638)
         );
  NAND3_X1 U8334 ( .A1(n6617), .A2(n10390), .A3(n6618), .ZN(n6616) );
  OAI21_X1 U8335 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(n6619) );
  NOR3_X1 U8336 ( .A1(n6620), .A2(n6622), .A3(n6619), .ZN(n6621) );
  INV_X1 U8337 ( .A(n6622), .ZN(n6634) );
  INV_X1 U8338 ( .A(n6623), .ZN(n6624) );
  OR2_X1 U8339 ( .A1(n6625), .A2(n6624), .ZN(n6628) );
  INV_X1 U8340 ( .A(n6626), .ZN(n6627) );
  NOR2_X2 U8341 ( .A1(n8797), .A2(n6215), .ZN(n8903) );
  AOI22_X1 U8342 ( .A1(n8915), .A2(n8903), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6633) );
  AND3_X1 U8343 ( .A1(n6629), .A2(n10345), .A3(n6903), .ZN(n6630) );
  NAND2_X1 U8344 ( .A1(n7312), .A2(n6630), .ZN(n6631) );
  AOI22_X1 U8345 ( .A1(n8913), .A2(n8874), .B1(n8902), .B2(n9105), .ZN(n6632)
         );
  OAI211_X1 U8346 ( .C1(n6638), .C2(n6634), .A(n6633), .B(n6632), .ZN(n6635)
         );
  INV_X1 U8347 ( .A(n6635), .ZN(n6636) );
  OAI211_X1 U8348 ( .C1(n8733), .C2(n6638), .A(n6637), .B(n6636), .ZN(P2_U3222) );
  AND2_X4 U8349 ( .A1(n6639), .A2(n6863), .ZN(n6830) );
  NOR2_X1 U8350 ( .A1(n6904), .A2(n6642), .ZN(n6643) );
  AOI21_X1 U8351 ( .B1(n6863), .B2(n7179), .A(n6643), .ZN(n6645) );
  NAND2_X1 U8352 ( .A1(n7119), .A2(n7118), .ZN(n7117) );
  NAND2_X1 U8353 ( .A1(n6646), .A2(n6847), .ZN(n6647) );
  NAND2_X1 U8354 ( .A1(n4395), .A2(n6650), .ZN(n6648) );
  XNOR2_X1 U8355 ( .A(n6690), .B(n6649), .ZN(n6654) );
  NAND2_X1 U8356 ( .A1(n6830), .A2(n6650), .ZN(n6652) );
  INV_X2 U8357 ( .A(n4395), .ZN(n6875) );
  NAND2_X1 U8358 ( .A1(n6663), .A2(n7368), .ZN(n6651) );
  NAND2_X1 U8359 ( .A1(n6652), .A2(n6651), .ZN(n7130) );
  NAND2_X1 U8360 ( .A1(n7127), .A2(n7130), .ZN(n6657) );
  INV_X1 U8361 ( .A(n6653), .ZN(n6656) );
  INV_X1 U8362 ( .A(n6654), .ZN(n6655) );
  NAND2_X1 U8363 ( .A1(n6656), .A2(n6655), .ZN(n7128) );
  OAI22_X1 U8365 ( .A1(n7173), .A2(n6659), .B1(n7424), .B2(n6875), .ZN(n6661)
         );
  AOI22_X1 U8366 ( .A1(n9675), .A2(n6830), .B1(n6663), .B2(n7176), .ZN(n6665)
         );
  INV_X1 U8367 ( .A(n6664), .ZN(n6666) );
  NAND2_X1 U8368 ( .A1(n6666), .A2(n6665), .ZN(n6667) );
  INV_X1 U8369 ( .A(n7188), .ZN(n6674) );
  NAND2_X1 U8370 ( .A1(n6663), .A2(n9674), .ZN(n6669) );
  NAND2_X1 U8371 ( .A1(n7466), .A2(n6863), .ZN(n6668) );
  NAND2_X1 U8372 ( .A1(n6669), .A2(n6668), .ZN(n6670) );
  XNOR2_X1 U8373 ( .A(n6670), .B(n6847), .ZN(n6675) );
  NAND2_X1 U8374 ( .A1(n6830), .A2(n9674), .ZN(n6672) );
  NAND2_X1 U8375 ( .A1(n6868), .A2(n7466), .ZN(n6671) );
  NAND2_X1 U8376 ( .A1(n6672), .A2(n6671), .ZN(n6676) );
  XNOR2_X1 U8377 ( .A(n6675), .B(n6676), .ZN(n7189) );
  NAND2_X1 U8378 ( .A1(n6675), .A2(n6676), .ZN(n6677) );
  NAND2_X1 U8379 ( .A1(n6663), .A2(n9673), .ZN(n6678) );
  NAND2_X1 U8380 ( .A1(n6830), .A2(n9673), .ZN(n6681) );
  OR2_X1 U8381 ( .A1(n6875), .A2(n6679), .ZN(n6680) );
  NAND2_X1 U8382 ( .A1(n6681), .A2(n6680), .ZN(n6684) );
  XNOR2_X1 U8383 ( .A(n6683), .B(n6684), .ZN(n7396) );
  INV_X1 U8384 ( .A(n6683), .ZN(n6686) );
  INV_X1 U8385 ( .A(n6684), .ZN(n6685) );
  NAND2_X1 U8386 ( .A1(n6686), .A2(n6685), .ZN(n6687) );
  NAND2_X1 U8387 ( .A1(n7758), .A2(n6863), .ZN(n6689) );
  NAND2_X1 U8388 ( .A1(n9672), .A2(n6868), .ZN(n6688) );
  NAND2_X1 U8389 ( .A1(n6689), .A2(n6688), .ZN(n6691) );
  XNOR2_X1 U8390 ( .A(n6691), .B(n6690), .ZN(n6696) );
  NAND2_X1 U8391 ( .A1(n7758), .A2(n6868), .ZN(n6693) );
  NAND2_X1 U8392 ( .A1(n9672), .A2(n6830), .ZN(n6692) );
  NAND2_X1 U8393 ( .A1(n6693), .A2(n6692), .ZN(n6694) );
  INV_X1 U8394 ( .A(n6694), .ZN(n6695) );
  NAND2_X1 U8395 ( .A1(n6696), .A2(n6695), .ZN(n6697) );
  NAND2_X1 U8396 ( .A1(n7640), .A2(n6863), .ZN(n6699) );
  NAND2_X1 U8397 ( .A1(n9671), .A2(n6663), .ZN(n6698) );
  NAND2_X1 U8398 ( .A1(n6699), .A2(n6698), .ZN(n6700) );
  NOR2_X1 U8399 ( .A1(n7649), .A2(n4396), .ZN(n6701) );
  AOI21_X1 U8400 ( .B1(n7640), .B2(n6868), .A(n6701), .ZN(n6703) );
  XNOR2_X1 U8401 ( .A(n6702), .B(n6703), .ZN(n7562) );
  NAND2_X1 U8402 ( .A1(n10174), .A2(n6863), .ZN(n6706) );
  NAND2_X1 U8403 ( .A1(n9669), .A2(n6868), .ZN(n6705) );
  NAND2_X1 U8404 ( .A1(n10174), .A2(n6868), .ZN(n6708) );
  NAND2_X1 U8405 ( .A1(n9669), .A2(n6830), .ZN(n6707) );
  NAND2_X1 U8406 ( .A1(n6708), .A2(n6707), .ZN(n7845) );
  NAND2_X1 U8407 ( .A1(n10179), .A2(n6663), .ZN(n6710) );
  NAND2_X1 U8408 ( .A1(n9670), .A2(n6830), .ZN(n6709) );
  NAND2_X1 U8409 ( .A1(n6710), .A2(n6709), .ZN(n7843) );
  NAND2_X1 U8410 ( .A1(n10179), .A2(n6863), .ZN(n6712) );
  NAND2_X1 U8411 ( .A1(n9670), .A2(n6868), .ZN(n6711) );
  AOI22_X1 U8412 ( .A1(n7846), .A2(n7845), .B1(n7843), .B2(n7841), .ZN(n6714)
         );
  INV_X1 U8413 ( .A(n7846), .ZN(n6717) );
  OAI21_X1 U8414 ( .B1(n7841), .B2(n7843), .A(n7845), .ZN(n6716) );
  NOR2_X1 U8415 ( .A1(n7845), .A2(n7843), .ZN(n6715) );
  NAND2_X1 U8416 ( .A1(n8399), .A2(n6863), .ZN(n6719) );
  NAND2_X1 U8417 ( .A1(n9668), .A2(n6868), .ZN(n6718) );
  NAND2_X1 U8418 ( .A1(n6719), .A2(n6718), .ZN(n6720) );
  XNOR2_X1 U8419 ( .A(n6720), .B(n6847), .ZN(n6722) );
  NOR2_X1 U8420 ( .A1(n8270), .A2(n4396), .ZN(n6721) );
  AOI21_X1 U8421 ( .B1(n8399), .B2(n4395), .A(n6721), .ZN(n6723) );
  XNOR2_X1 U8422 ( .A(n6722), .B(n6723), .ZN(n7944) );
  INV_X1 U8423 ( .A(n6722), .ZN(n6724) );
  NAND2_X1 U8424 ( .A1(n6724), .A2(n6723), .ZN(n7903) );
  NAND2_X1 U8425 ( .A1(n8411), .A2(n6863), .ZN(n6726) );
  NAND2_X1 U8426 ( .A1(n9667), .A2(n6868), .ZN(n6725) );
  NAND2_X1 U8427 ( .A1(n6726), .A2(n6725), .ZN(n6727) );
  XNOR2_X1 U8428 ( .A(n6727), .B(n6847), .ZN(n6732) );
  INV_X1 U8429 ( .A(n6732), .ZN(n6729) );
  NOR2_X1 U8430 ( .A1(n7948), .A2(n4396), .ZN(n6728) );
  AOI21_X1 U8431 ( .B1(n8411), .B2(n6663), .A(n6728), .ZN(n6731) );
  NAND2_X1 U8432 ( .A1(n6729), .A2(n6731), .ZN(n6730) );
  AND2_X1 U8433 ( .A1(n7903), .A2(n6730), .ZN(n6734) );
  INV_X1 U8434 ( .A(n6730), .ZN(n6733) );
  XNOR2_X1 U8435 ( .A(n6732), .B(n6731), .ZN(n7906) );
  NAND2_X1 U8436 ( .A1(n10170), .A2(n6863), .ZN(n6736) );
  NAND2_X1 U8437 ( .A1(n10040), .A2(n6868), .ZN(n6735) );
  NAND2_X1 U8438 ( .A1(n6736), .A2(n6735), .ZN(n6737) );
  XNOR2_X1 U8439 ( .A(n6737), .B(n6847), .ZN(n6739) );
  NOR2_X1 U8440 ( .A1(n7909), .A2(n4396), .ZN(n6738) );
  AOI21_X1 U8441 ( .B1(n10170), .B2(n6663), .A(n6738), .ZN(n6740) );
  XNOR2_X1 U8442 ( .A(n6739), .B(n6740), .ZN(n8244) );
  INV_X1 U8443 ( .A(n6739), .ZN(n6741) );
  NAND2_X1 U8444 ( .A1(n6741), .A2(n6740), .ZN(n6742) );
  NAND2_X1 U8445 ( .A1(n10164), .A2(n6863), .ZN(n6744) );
  NAND2_X1 U8446 ( .A1(n9666), .A2(n6868), .ZN(n6743) );
  NAND2_X1 U8447 ( .A1(n6744), .A2(n6743), .ZN(n6745) );
  XNOR2_X1 U8448 ( .A(n6745), .B(n6690), .ZN(n8300) );
  NOR2_X1 U8449 ( .A1(n10015), .A2(n4396), .ZN(n6746) );
  AOI21_X1 U8450 ( .B1(n10164), .B2(n6868), .A(n6746), .ZN(n8299) );
  AND2_X1 U8451 ( .A1(n8300), .A2(n8299), .ZN(n6750) );
  INV_X1 U8452 ( .A(n8300), .ZN(n6748) );
  INV_X1 U8453 ( .A(n8299), .ZN(n6747) );
  NAND2_X1 U8454 ( .A1(n6748), .A2(n6747), .ZN(n6749) );
  NAND2_X1 U8455 ( .A1(n10159), .A2(n6863), .ZN(n6752) );
  NAND2_X1 U8456 ( .A1(n10042), .A2(n6868), .ZN(n6751) );
  NAND2_X1 U8457 ( .A1(n10159), .A2(n6868), .ZN(n6754) );
  NAND2_X1 U8458 ( .A1(n10042), .A2(n6830), .ZN(n6753) );
  NAND2_X1 U8459 ( .A1(n6754), .A2(n6753), .ZN(n6755) );
  AND2_X1 U8460 ( .A1(n8423), .A2(n6755), .ZN(n6768) );
  INV_X1 U8461 ( .A(n8423), .ZN(n6756) );
  INV_X1 U8462 ( .A(n6755), .ZN(n8422) );
  NAND2_X1 U8463 ( .A1(n6756), .A2(n8422), .ZN(n6779) );
  NAND2_X1 U8464 ( .A1(n10154), .A2(n6863), .ZN(n6758) );
  NAND2_X1 U8465 ( .A1(n9978), .A2(n4395), .ZN(n6757) );
  NAND2_X1 U8466 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  XNOR2_X1 U8467 ( .A(n6759), .B(n6847), .ZN(n6769) );
  AND2_X1 U8468 ( .A1(n6779), .A2(n6769), .ZN(n9569) );
  NAND2_X1 U8469 ( .A1(n10149), .A2(n6863), .ZN(n6761) );
  NAND2_X1 U8470 ( .A1(n9998), .A2(n6868), .ZN(n6760) );
  NAND2_X1 U8471 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  XNOR2_X1 U8472 ( .A(n6762), .B(n6690), .ZN(n6773) );
  NOR2_X1 U8473 ( .A1(n9653), .A2(n4396), .ZN(n6763) );
  AOI21_X1 U8474 ( .B1(n10149), .B2(n6663), .A(n6763), .ZN(n6774) );
  NAND2_X1 U8475 ( .A1(n6773), .A2(n6774), .ZN(n9580) );
  NAND2_X1 U8476 ( .A1(n10144), .A2(n6863), .ZN(n6765) );
  NAND2_X1 U8477 ( .A1(n9979), .A2(n6868), .ZN(n6764) );
  NAND2_X1 U8478 ( .A1(n6765), .A2(n6764), .ZN(n6766) );
  XNOR2_X1 U8479 ( .A(n6766), .B(n6847), .ZN(n6782) );
  NOR2_X1 U8480 ( .A1(n9628), .A2(n4396), .ZN(n6767) );
  AOI21_X1 U8481 ( .B1(n10144), .B2(n6868), .A(n6767), .ZN(n6783) );
  XNOR2_X1 U8482 ( .A(n6782), .B(n6783), .ZN(n9581) );
  INV_X1 U8483 ( .A(n6768), .ZN(n6771) );
  INV_X1 U8484 ( .A(n6769), .ZN(n6770) );
  AND2_X1 U8485 ( .A1(n6771), .A2(n6770), .ZN(n9567) );
  NOR2_X1 U8486 ( .A1(n10016), .A2(n4396), .ZN(n6772) );
  AOI21_X1 U8487 ( .B1(n10154), .B2(n6868), .A(n6772), .ZN(n9647) );
  INV_X1 U8488 ( .A(n6773), .ZN(n6776) );
  INV_X1 U8489 ( .A(n6774), .ZN(n6775) );
  NAND2_X1 U8490 ( .A1(n6776), .A2(n6775), .ZN(n9571) );
  NAND2_X1 U8491 ( .A1(n6777), .A2(n9580), .ZN(n6778) );
  INV_X1 U8492 ( .A(n9647), .ZN(n6780) );
  NAND2_X1 U8493 ( .A1(n9580), .A2(n6780), .ZN(n6781) );
  INV_X1 U8494 ( .A(n6782), .ZN(n6784) );
  NAND2_X1 U8495 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  NAND2_X1 U8496 ( .A1(n10133), .A2(n6863), .ZN(n6787) );
  OR2_X1 U8497 ( .A1(n9909), .A2(n6875), .ZN(n6786) );
  NAND2_X1 U8498 ( .A1(n6787), .A2(n6786), .ZN(n6788) );
  XNOR2_X1 U8499 ( .A(n6788), .B(n6847), .ZN(n9537) );
  NAND2_X1 U8500 ( .A1(n10133), .A2(n6868), .ZN(n6790) );
  OR2_X1 U8501 ( .A1(n9909), .A2(n4396), .ZN(n6789) );
  NAND2_X1 U8502 ( .A1(n6790), .A2(n6789), .ZN(n9536) );
  NAND2_X1 U8503 ( .A1(n9537), .A2(n9536), .ZN(n9535) );
  NAND2_X1 U8504 ( .A1(n10138), .A2(n6863), .ZN(n6792) );
  NAND2_X1 U8505 ( .A1(n9962), .A2(n6868), .ZN(n6791) );
  NAND2_X1 U8506 ( .A1(n6792), .A2(n6791), .ZN(n6793) );
  XNOR2_X1 U8507 ( .A(n6793), .B(n6847), .ZN(n6798) );
  NAND2_X1 U8508 ( .A1(n10138), .A2(n6868), .ZN(n6795) );
  NAND2_X1 U8509 ( .A1(n9962), .A2(n6830), .ZN(n6794) );
  NAND2_X1 U8510 ( .A1(n6795), .A2(n6794), .ZN(n9621) );
  NAND2_X1 U8511 ( .A1(n6798), .A2(n9621), .ZN(n6796) );
  AND2_X1 U8512 ( .A1(n9535), .A2(n6796), .ZN(n6797) );
  OAI21_X1 U8513 ( .B1(n6798), .B2(n9621), .A(n9536), .ZN(n6801) );
  INV_X1 U8514 ( .A(n9537), .ZN(n6800) );
  INV_X1 U8515 ( .A(n6798), .ZN(n9539) );
  NOR2_X1 U8516 ( .A1(n9536), .A2(n9621), .ZN(n6799) );
  AOI22_X1 U8517 ( .A1(n6801), .A2(n6800), .B1(n9539), .B2(n6799), .ZN(n6802)
         );
  NAND2_X1 U8518 ( .A1(n10124), .A2(n6863), .ZN(n6805) );
  NAND2_X1 U8519 ( .A1(n9931), .A2(n6868), .ZN(n6804) );
  NAND2_X1 U8520 ( .A1(n6805), .A2(n6804), .ZN(n6806) );
  XNOR2_X1 U8521 ( .A(n6806), .B(n6847), .ZN(n6808) );
  NOR2_X1 U8522 ( .A1(n9543), .A2(n4396), .ZN(n6807) );
  AOI21_X1 U8523 ( .B1(n10124), .B2(n4395), .A(n6807), .ZN(n6809) );
  XNOR2_X1 U8524 ( .A(n6808), .B(n6809), .ZN(n9603) );
  INV_X1 U8525 ( .A(n6808), .ZN(n6810) );
  NAND2_X1 U8526 ( .A1(n6810), .A2(n6809), .ZN(n9549) );
  NAND2_X1 U8527 ( .A1(n10118), .A2(n6863), .ZN(n6812) );
  NAND2_X1 U8528 ( .A1(n9876), .A2(n6868), .ZN(n6811) );
  NAND2_X1 U8529 ( .A1(n6812), .A2(n6811), .ZN(n6813) );
  XNOR2_X1 U8530 ( .A(n6813), .B(n6847), .ZN(n6818) );
  INV_X1 U8531 ( .A(n6818), .ZN(n6815) );
  NOR2_X1 U8532 ( .A1(n9910), .A2(n4396), .ZN(n6814) );
  AOI21_X1 U8533 ( .B1(n10118), .B2(n6868), .A(n6814), .ZN(n6817) );
  NAND2_X1 U8534 ( .A1(n6815), .A2(n6817), .ZN(n6816) );
  AND2_X1 U8535 ( .A1(n9549), .A2(n6816), .ZN(n6820) );
  INV_X1 U8536 ( .A(n6816), .ZN(n6819) );
  XNOR2_X1 U8537 ( .A(n6818), .B(n6817), .ZN(n9552) );
  OR2_X1 U8538 ( .A1(n9883), .A2(n6875), .ZN(n6822) );
  NAND2_X1 U8539 ( .A1(n9894), .A2(n6830), .ZN(n6821) );
  AND2_X1 U8540 ( .A1(n6822), .A2(n6821), .ZN(n6825) );
  OAI22_X1 U8541 ( .A1(n9883), .A2(n6873), .B1(n9531), .B2(n6875), .ZN(n6824)
         );
  XNOR2_X1 U8542 ( .A(n6824), .B(n6690), .ZN(n9612) );
  NAND2_X1 U8543 ( .A1(n10109), .A2(n6863), .ZN(n6828) );
  NAND2_X1 U8544 ( .A1(n9877), .A2(n6868), .ZN(n6827) );
  NAND2_X1 U8545 ( .A1(n6828), .A2(n6827), .ZN(n6829) );
  XNOR2_X1 U8546 ( .A(n6829), .B(n6690), .ZN(n6834) );
  NAND2_X1 U8547 ( .A1(n10109), .A2(n6868), .ZN(n6832) );
  NAND2_X1 U8548 ( .A1(n9877), .A2(n6830), .ZN(n6831) );
  NAND2_X1 U8549 ( .A1(n6832), .A2(n6831), .ZN(n9528) );
  INV_X1 U8550 ( .A(n6834), .ZN(n6835) );
  NAND2_X1 U8551 ( .A1(n10106), .A2(n6863), .ZN(n6839) );
  NAND2_X1 U8552 ( .A1(n9864), .A2(n6663), .ZN(n6838) );
  NAND2_X1 U8553 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  XNOR2_X1 U8554 ( .A(n6840), .B(n6690), .ZN(n6843) );
  NOR2_X1 U8555 ( .A1(n9562), .A2(n4396), .ZN(n6841) );
  AOI21_X1 U8556 ( .B1(n10106), .B2(n6868), .A(n6841), .ZN(n6842) );
  XNOR2_X1 U8557 ( .A(n6843), .B(n6842), .ZN(n9595) );
  NAND2_X1 U8558 ( .A1(n6843), .A2(n6842), .ZN(n6844) );
  NAND2_X1 U8559 ( .A1(n10099), .A2(n6863), .ZN(n6846) );
  NAND2_X1 U8560 ( .A1(n9808), .A2(n4395), .ZN(n6845) );
  NAND2_X1 U8561 ( .A1(n6846), .A2(n6845), .ZN(n6848) );
  XNOR2_X1 U8562 ( .A(n6848), .B(n6847), .ZN(n6850) );
  NOR2_X1 U8563 ( .A1(n9853), .A2(n4396), .ZN(n6849) );
  AOI21_X1 U8564 ( .B1(n10099), .B2(n6868), .A(n6849), .ZN(n6851) );
  XNOR2_X1 U8565 ( .A(n6850), .B(n6851), .ZN(n9558) );
  INV_X1 U8566 ( .A(n6850), .ZN(n6852) );
  NAND2_X1 U8567 ( .A1(n10094), .A2(n6863), .ZN(n6854) );
  NAND2_X1 U8568 ( .A1(n9829), .A2(n6868), .ZN(n6853) );
  NAND2_X1 U8569 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  XNOR2_X1 U8570 ( .A(n6855), .B(n6690), .ZN(n6858) );
  NOR2_X1 U8571 ( .A1(n9519), .A2(n4396), .ZN(n6856) );
  AOI21_X1 U8572 ( .B1(n10094), .B2(n4395), .A(n6856), .ZN(n6859) );
  XNOR2_X1 U8573 ( .A(n6858), .B(n6859), .ZN(n9637) );
  INV_X1 U8574 ( .A(n9637), .ZN(n6857) );
  INV_X1 U8575 ( .A(n6858), .ZN(n6861) );
  INV_X1 U8576 ( .A(n6859), .ZN(n6860) );
  NAND2_X1 U8577 ( .A1(n6861), .A2(n6860), .ZN(n6862) );
  NAND2_X1 U8578 ( .A1(n9638), .A2(n6862), .ZN(n6870) );
  NAND2_X1 U8579 ( .A1(n10089), .A2(n6863), .ZN(n6865) );
  NAND2_X1 U8580 ( .A1(n9807), .A2(n4395), .ZN(n6864) );
  NAND2_X1 U8581 ( .A1(n6865), .A2(n6864), .ZN(n6866) );
  NOR2_X1 U8582 ( .A1(n9641), .A2(n4396), .ZN(n6867) );
  INV_X1 U8583 ( .A(n9515), .ZN(n6869) );
  NAND2_X1 U8584 ( .A1(n6870), .A2(n6869), .ZN(n6896) );
  INV_X1 U8585 ( .A(n7244), .ZN(n7049) );
  NAND3_X1 U8586 ( .A1(n6977), .A2(n7049), .A3(n7046), .ZN(n6888) );
  INV_X1 U8587 ( .A(n6979), .ZN(n10213) );
  OR2_X1 U8588 ( .A1(n7054), .A2(n6871), .ZN(n10295) );
  NAND2_X1 U8589 ( .A1(n10295), .A2(n8717), .ZN(n6872) );
  OAI22_X1 U8590 ( .A1(n6876), .A2(n6873), .B1(n9768), .B2(n6875), .ZN(n6874)
         );
  XNOR2_X1 U8591 ( .A(n6874), .B(n6690), .ZN(n6878) );
  OAI22_X1 U8592 ( .A1(n6876), .A2(n6875), .B1(n9768), .B2(n4396), .ZN(n6877)
         );
  XNOR2_X1 U8593 ( .A(n6878), .B(n6877), .ZN(n6879) );
  NAND3_X1 U8594 ( .A1(n6896), .A2(n9650), .A3(n6879), .ZN(n6900) );
  INV_X1 U8595 ( .A(n6879), .ZN(n6880) );
  NAND2_X1 U8596 ( .A1(n6880), .A2(n9650), .ZN(n6895) );
  INV_X1 U8597 ( .A(n6895), .ZN(n6881) );
  NAND2_X1 U8598 ( .A1(n6901), .A2(n6881), .ZN(n6899) );
  NOR2_X1 U8599 ( .A1(n6882), .A2(n8725), .ZN(n6883) );
  INV_X1 U8600 ( .A(n4391), .ZN(n10226) );
  NAND2_X1 U8601 ( .A1(n6883), .A2(n10226), .ZN(n9657) );
  NAND2_X1 U8602 ( .A1(n6883), .A2(n4391), .ZN(n9654) );
  OR2_X1 U8603 ( .A1(n8469), .A2(n9654), .ZN(n6892) );
  AND3_X1 U8604 ( .A1(n6904), .A2(n6884), .A3(n8236), .ZN(n6885) );
  NAND2_X1 U8605 ( .A1(n6888), .A2(n10295), .ZN(n7131) );
  NAND2_X1 U8606 ( .A1(n6885), .A2(n7131), .ZN(n6886) );
  NAND2_X1 U8607 ( .A1(n6886), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6889) );
  NAND3_X1 U8608 ( .A1(n5730), .A2(n6888), .A3(n6979), .ZN(n7133) );
  AOI22_X1 U8609 ( .A1(n6890), .A2(n9660), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6891) );
  OAI211_X1 U8610 ( .C1(n9641), .C2(n9657), .A(n6892), .B(n6891), .ZN(n6893)
         );
  AOI21_X1 U8611 ( .B1(n10085), .B2(n4380), .A(n6893), .ZN(n6894) );
  INV_X1 U8612 ( .A(n6897), .ZN(n6898) );
  OAI211_X1 U8613 ( .C1(n6901), .C2(n6900), .A(n6899), .B(n6898), .ZN(P1_U3218) );
  INV_X1 U8614 ( .A(n8236), .ZN(n6902) );
  NOR2_X1 U8615 ( .A1(n6904), .A2(n6902), .ZN(n6970) );
  AND2_X2 U8616 ( .A1(n6970), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND2_X1 U8617 ( .A1(n8717), .A2(n6904), .ZN(n6905) );
  NAND2_X1 U8618 ( .A1(n6905), .A2(n8236), .ZN(n6967) );
  NAND2_X1 U8619 ( .A1(n6967), .A2(n5326), .ZN(n6906) );
  NAND2_X1 U8620 ( .A1(n6906), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U8621 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7120) );
  INV_X1 U8622 ( .A(n7120), .ZN(n7089) );
  NAND2_X1 U8623 ( .A1(n7090), .A2(n7089), .ZN(n7088) );
  INV_X1 U8624 ( .A(n7093), .ZN(n6936) );
  NAND2_X1 U8625 ( .A1(n6936), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U8626 ( .A1(n7088), .A2(n6907), .ZN(n7111) );
  INV_X1 U8627 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6908) );
  XNOR2_X1 U8628 ( .A(n6983), .B(n6908), .ZN(n7112) );
  NAND2_X1 U8629 ( .A1(n7111), .A2(n7112), .ZN(n7110) );
  NAND2_X1 U8630 ( .A1(n6983), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U8631 ( .A1(n7110), .A2(n6909), .ZN(n7101) );
  INV_X1 U8632 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6910) );
  XNOR2_X1 U8633 ( .A(n6984), .B(n6910), .ZN(n7102) );
  NAND2_X1 U8634 ( .A1(n7101), .A2(n7102), .ZN(n7100) );
  NAND2_X1 U8635 ( .A1(n6984), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U8636 ( .A1(n7100), .A2(n6911), .ZN(n9684) );
  MUX2_X1 U8637 ( .A(n7451), .B(P1_REG2_REG_4__SCAN_IN), .S(n9688), .Z(n9683)
         );
  OR2_X1 U8638 ( .A1(n9684), .A2(n9683), .ZN(n9686) );
  OR2_X1 U8639 ( .A1(n9688), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8640 ( .A1(n9686), .A2(n6912), .ZN(n9693) );
  INV_X1 U8641 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6913) );
  XNOR2_X1 U8642 ( .A(n9697), .B(n6913), .ZN(n9692) );
  NAND2_X1 U8643 ( .A1(n9693), .A2(n9692), .ZN(n6915) );
  INV_X1 U8644 ( .A(n9697), .ZN(n7011) );
  NAND2_X1 U8645 ( .A1(n7011), .A2(n6913), .ZN(n6914) );
  NAND2_X1 U8646 ( .A1(n6915), .A2(n6914), .ZN(n7077) );
  INV_X1 U8647 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6916) );
  MUX2_X1 U8648 ( .A(n6916), .B(P1_REG2_REG_6__SCAN_IN), .S(n6993), .Z(n7076)
         );
  NAND2_X1 U8649 ( .A1(n6993), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6917) );
  INV_X1 U8650 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6918) );
  XNOR2_X1 U8651 ( .A(n7064), .B(n6918), .ZN(n7063) );
  OR2_X1 U8652 ( .A1(n7064), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6919) );
  INV_X1 U8653 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6920) );
  XNOR2_X1 U8654 ( .A(n7014), .B(n6920), .ZN(n7037) );
  OR2_X1 U8655 ( .A1(n7014), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U8656 ( .A1(n6922), .A2(n6921), .ZN(n7164) );
  INV_X1 U8657 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6923) );
  MUX2_X1 U8658 ( .A(n6923), .B(P1_REG2_REG_9__SCAN_IN), .S(n7021), .Z(n7165)
         );
  NAND2_X1 U8659 ( .A1(n7021), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U8660 ( .A1(n7162), .A2(n6924), .ZN(n7199) );
  INV_X1 U8661 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6925) );
  MUX2_X1 U8662 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n6925), .S(n6950), .Z(n7198)
         );
  NAND2_X1 U8663 ( .A1(n7199), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U8664 ( .A1(n6950), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6926) );
  INV_X1 U8665 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6927) );
  XNOR2_X1 U8666 ( .A(n7027), .B(n6927), .ZN(n7234) );
  OR2_X1 U8667 ( .A1(n7027), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6928) );
  INV_X1 U8668 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6929) );
  XNOR2_X1 U8669 ( .A(n7543), .B(n6929), .ZN(n7547) );
  OR2_X1 U8670 ( .A1(n7543), .A2(n6929), .ZN(n6930) );
  INV_X1 U8671 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8063) );
  MUX2_X1 U8672 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n8063), .S(n7126), .Z(n7668)
         );
  NAND2_X1 U8673 ( .A1(n7669), .A2(n7668), .ZN(n7667) );
  NAND2_X1 U8674 ( .A1(n7126), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U8675 ( .A1(n7667), .A2(n6931), .ZN(n6932) );
  INV_X1 U8676 ( .A(n6963), .ZN(n7773) );
  XNOR2_X1 U8677 ( .A(n6932), .B(n7773), .ZN(n7771) );
  INV_X1 U8678 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U8679 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9711), .ZN(n6933) );
  OAI21_X1 U8680 ( .B1(n9711), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6933), .ZN(
        n6934) );
  NOR2_X1 U8681 ( .A1(n8724), .A2(P1_U3084), .ZN(n10229) );
  AND2_X1 U8682 ( .A1(n6967), .A2(n10229), .ZN(n9740) );
  INV_X1 U8683 ( .A(n9740), .ZN(n6972) );
  NOR2_X1 U8684 ( .A1(n6935), .A2(n6934), .ZN(n9707) );
  AOI211_X1 U8685 ( .C1(n6935), .C2(n6934), .A(n9746), .B(n9707), .ZN(n6976)
         );
  XNOR2_X1 U8686 ( .A(n7093), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n7085) );
  AND2_X1 U8687 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7084) );
  NAND2_X1 U8688 ( .A1(n7085), .A2(n7084), .ZN(n7083) );
  NAND2_X1 U8689 ( .A1(n6936), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6937) );
  NAND2_X1 U8690 ( .A1(n7083), .A2(n6937), .ZN(n7107) );
  INV_X1 U8691 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6938) );
  XNOR2_X1 U8692 ( .A(n6983), .B(n6938), .ZN(n7108) );
  NAND2_X1 U8693 ( .A1(n7107), .A2(n7108), .ZN(n7106) );
  NAND2_X1 U8694 ( .A1(n6983), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6939) );
  NAND2_X1 U8695 ( .A1(n7106), .A2(n6939), .ZN(n7095) );
  INV_X1 U8696 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10304) );
  MUX2_X1 U8697 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10304), .S(n6984), .Z(n7096)
         );
  NAND2_X1 U8698 ( .A1(n7095), .A2(n7096), .ZN(n7094) );
  NAND2_X1 U8699 ( .A1(n6984), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U8700 ( .A1(n7094), .A2(n6940), .ZN(n9678) );
  MUX2_X1 U8701 ( .A(n5155), .B(P1_REG1_REG_4__SCAN_IN), .S(n9688), .Z(n9677)
         );
  OR2_X1 U8702 ( .A1(n9688), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6941) );
  AND2_X1 U8703 ( .A1(n9680), .A2(n6941), .ZN(n9700) );
  INV_X1 U8704 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6942) );
  XNOR2_X1 U8705 ( .A(n9697), .B(n6942), .ZN(n9701) );
  NAND2_X1 U8706 ( .A1(n9700), .A2(n9701), .ZN(n9698) );
  NAND2_X1 U8707 ( .A1(n9697), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U8708 ( .A1(n9698), .A2(n6943), .ZN(n7072) );
  XNOR2_X1 U8709 ( .A(n6993), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n7073) );
  OR2_X1 U8710 ( .A1(n6993), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U8711 ( .A1(n7070), .A2(n6944), .ZN(n7060) );
  INV_X1 U8712 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6945) );
  XNOR2_X1 U8713 ( .A(n7064), .B(n6945), .ZN(n7061) );
  NOR2_X1 U8714 ( .A1(n7064), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6946) );
  AOI21_X1 U8715 ( .B1(n7060), .B2(n7061), .A(n6946), .ZN(n7042) );
  INV_X1 U8716 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6947) );
  XNOR2_X1 U8717 ( .A(n7014), .B(n6947), .ZN(n7041) );
  NAND2_X1 U8718 ( .A1(n7042), .A2(n7041), .ZN(n7040) );
  NAND2_X1 U8719 ( .A1(n7014), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6948) );
  NAND2_X1 U8720 ( .A1(n7040), .A2(n6948), .ZN(n7159) );
  XNOR2_X1 U8721 ( .A(n7021), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7160) );
  OR2_X1 U8722 ( .A1(n7021), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8723 ( .A1(n7157), .A2(n6949), .ZN(n7194) );
  INV_X1 U8724 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6951) );
  XNOR2_X1 U8725 ( .A(n6950), .B(n6951), .ZN(n7195) );
  NAND2_X1 U8726 ( .A1(n7194), .A2(n7195), .ZN(n6953) );
  INV_X1 U8727 ( .A(n6950), .ZN(n7196) );
  NAND2_X1 U8728 ( .A1(n7196), .A2(n6951), .ZN(n6952) );
  NAND2_X1 U8729 ( .A1(n6953), .A2(n6952), .ZN(n7230) );
  INV_X1 U8730 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8417) );
  XNOR2_X1 U8731 ( .A(n7027), .B(n8417), .ZN(n7231) );
  NAND2_X1 U8732 ( .A1(n7230), .A2(n7231), .ZN(n6955) );
  OR2_X1 U8733 ( .A1(n7027), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8734 ( .A1(n6955), .A2(n6954), .ZN(n7541) );
  XNOR2_X1 U8735 ( .A(n7543), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7542) );
  NAND2_X1 U8736 ( .A1(n7541), .A2(n7542), .ZN(n6958) );
  INV_X1 U8737 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U8738 ( .A1(n7543), .A2(n6956), .ZN(n6957) );
  NAND2_X1 U8739 ( .A1(n6958), .A2(n6957), .ZN(n7664) );
  INV_X1 U8740 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6959) );
  XNOR2_X1 U8741 ( .A(n7126), .B(n6959), .ZN(n7665) );
  NAND2_X1 U8742 ( .A1(n7664), .A2(n7665), .ZN(n6961) );
  OR2_X1 U8743 ( .A1(n7126), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6960) );
  NAND2_X1 U8744 ( .A1(n6961), .A2(n6960), .ZN(n7774) );
  INV_X1 U8745 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6962) );
  XNOR2_X1 U8746 ( .A(n6963), .B(n6962), .ZN(n7775) );
  NOR2_X1 U8747 ( .A1(n6963), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6964) );
  AOI21_X1 U8748 ( .B1(n7774), .B2(n7775), .A(n6964), .ZN(n6965) );
  XOR2_X1 U8749 ( .A(n7154), .B(n6965), .Z(n7894) );
  AOI21_X1 U8750 ( .B1(n6965), .B2(n7154), .A(n7895), .ZN(n6969) );
  XNOR2_X1 U8751 ( .A(n9711), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n6968) );
  AND2_X1 U8752 ( .A1(n5326), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6966) );
  NAND2_X1 U8753 ( .A1(n6967), .A2(n6966), .ZN(n10243) );
  INV_X1 U8754 ( .A(n8724), .ZN(n10239) );
  NOR2_X1 U8755 ( .A1(n6969), .A2(n6968), .ZN(n9710) );
  AOI211_X1 U8756 ( .C1(n6969), .C2(n6968), .A(n9745), .B(n9710), .ZN(n6975)
         );
  OR2_X1 U8757 ( .A1(P1_U3083), .A2(n6970), .ZN(n10245) );
  INV_X1 U8758 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n6971) );
  NOR2_X1 U8759 ( .A1(n10245), .A2(n6971), .ZN(n6974) );
  INV_X1 U8760 ( .A(n9711), .ZN(n7186) );
  NAND2_X1 U8761 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9575) );
  OAI21_X1 U8762 ( .B1(n9741), .B2(n7186), .A(n9575), .ZN(n6973) );
  OR4_X1 U8763 ( .A1(n6976), .A2(n6975), .A3(n6974), .A4(n6973), .ZN(P1_U3257)
         );
  NAND2_X1 U8764 ( .A1(n6977), .A2(n6979), .ZN(n6978) );
  OAI21_X1 U8765 ( .B1(n6979), .B2(n8207), .A(n6978), .ZN(P1_U3441) );
  NOR2_X1 U8766 ( .A1(n4393), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10230) );
  INV_X1 U8767 ( .A(n10230), .ZN(n8444) );
  INV_X1 U8768 ( .A(n6980), .ZN(n6987) );
  INV_X1 U8769 ( .A(n9688), .ZN(n6981) );
  OAI222_X1 U8770 ( .A1(n8444), .A2(n6982), .B1(n10232), .B2(n6987), .C1(
        P1_U3084), .C2(n6981), .ZN(P1_U3349) );
  INV_X1 U8771 ( .A(n6983), .ZN(n7114) );
  OAI222_X1 U8772 ( .A1(n8444), .A2(n5132), .B1(n10232), .B2(n6991), .C1(
        P1_U3084), .C2(n7114), .ZN(P1_U3351) );
  INV_X1 U8773 ( .A(n6984), .ZN(n7105) );
  OAI222_X1 U8774 ( .A1(n8444), .A2(n6985), .B1(n10232), .B2(n7008), .C1(
        P1_U3084), .C2(n7105), .ZN(P1_U3350) );
  AND2_X1 U8775 ( .A1(n4393), .A2(P2_U3152), .ZN(n9499) );
  INV_X2 U8776 ( .A(n9499), .ZN(n9508) );
  NAND2_X1 U8777 ( .A1(n6986), .A2(P2_U3152), .ZN(n9506) );
  OAI222_X1 U8778 ( .A1(n9508), .A2(n6988), .B1(n9506), .B2(n6987), .C1(
        P2_U3152), .C2(n7296), .ZN(P2_U3354) );
  INV_X1 U8779 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8197) );
  INV_X1 U8780 ( .A(n6989), .ZN(n7012) );
  OAI222_X1 U8781 ( .A1(n9508), .A2(n8197), .B1(n9506), .B2(n7012), .C1(
        P2_U3152), .C2(n8960), .ZN(P2_U3353) );
  OAI222_X1 U8782 ( .A1(n7265), .A2(P2_U3152), .B1(n9506), .B2(n6991), .C1(
        n6990), .C2(n9508), .ZN(P2_U3356) );
  INV_X1 U8783 ( .A(n6992), .ZN(n6994) );
  INV_X1 U8784 ( .A(n6993), .ZN(n7074) );
  OAI222_X1 U8785 ( .A1(n8444), .A2(n4628), .B1(n10232), .B2(n6994), .C1(
        P1_U3084), .C2(n7074), .ZN(P1_U3347) );
  INV_X1 U8786 ( .A(n8979), .ZN(n7285) );
  OAI222_X1 U8787 ( .A1(n9508), .A2(n5200), .B1(n9506), .B2(n6994), .C1(
        P2_U3152), .C2(n7285), .ZN(P2_U3352) );
  INV_X1 U8788 ( .A(n6995), .ZN(n6998) );
  AOI22_X1 U8789 ( .A1(n7064), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10230), .ZN(n6996) );
  OAI21_X1 U8790 ( .B1(n6998), .B2(n10232), .A(n6996), .ZN(P1_U3346) );
  AOI22_X1 U8791 ( .A1(n8995), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n9499), .ZN(n6997) );
  OAI21_X1 U8792 ( .B1(n6998), .B2(n9506), .A(n6997), .ZN(P2_U3351) );
  INV_X1 U8793 ( .A(n6999), .ZN(n7015) );
  INV_X1 U8794 ( .A(n7303), .ZN(n9009) );
  OAI222_X1 U8795 ( .A1(n9508), .A2(n7000), .B1(n9506), .B2(n7015), .C1(
        P2_U3152), .C2(n9009), .ZN(P2_U3350) );
  NAND2_X1 U8796 ( .A1(n5087), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U8797 ( .A1(n7001), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U8798 ( .A1(n7002), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7003) );
  AND3_X1 U8799 ( .A1(n7005), .A2(n7004), .A3(n7003), .ZN(n9769) );
  INV_X1 U8800 ( .A(P1_U4006), .ZN(n7007) );
  NAND2_X1 U8801 ( .A1(n7007), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7006) );
  OAI21_X1 U8802 ( .B1(n9769), .B2(n7007), .A(n7006), .ZN(P1_U3585) );
  INV_X1 U8803 ( .A(n9506), .ZN(n8239) );
  INV_X1 U8804 ( .A(n8239), .ZN(n9511) );
  OAI222_X1 U8805 ( .A1(n9508), .A2(n7009), .B1(n9511), .B2(n7008), .C1(
        P2_U3152), .C2(n8944), .ZN(P2_U3355) );
  OAI222_X1 U8806 ( .A1(n8931), .A2(P2_U3152), .B1(n9511), .B2(n7017), .C1(
        n7010), .C2(n9508), .ZN(P2_U3357) );
  INV_X1 U8807 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7013) );
  OAI222_X1 U8808 ( .A1(n8444), .A2(n7013), .B1(n10232), .B2(n7012), .C1(
        P1_U3084), .C2(n7011), .ZN(P1_U3348) );
  INV_X1 U8809 ( .A(n7014), .ZN(n7038) );
  OAI222_X1 U8810 ( .A1(n8444), .A2(n7016), .B1(n10232), .B2(n7015), .C1(
        P1_U3084), .C2(n7038), .ZN(P1_U3345) );
  OAI222_X1 U8811 ( .A1(n8444), .A2(n7018), .B1(n10232), .B2(n7017), .C1(
        P1_U3084), .C2(n7093), .ZN(P1_U3352) );
  INV_X1 U8812 ( .A(n7019), .ZN(n7023) );
  AOI22_X1 U8813 ( .A1(n9029), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9499), .ZN(n7020) );
  OAI21_X1 U8814 ( .B1(n7023), .B2(n9506), .A(n7020), .ZN(P2_U3349) );
  INV_X1 U8815 ( .A(n7021), .ZN(n7161) );
  OAI222_X1 U8816 ( .A1(n10232), .A2(n7023), .B1(n7161), .B2(P1_U3084), .C1(
        n7022), .C2(n8444), .ZN(P1_U3344) );
  INV_X1 U8817 ( .A(n7024), .ZN(n7028) );
  AOI22_X1 U8818 ( .A1(n9042), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9499), .ZN(n7025) );
  OAI21_X1 U8819 ( .B1(n7028), .B2(n9506), .A(n7025), .ZN(P2_U3347) );
  INV_X1 U8820 ( .A(n7026), .ZN(n7033) );
  OAI222_X1 U8821 ( .A1(n10232), .A2(n7033), .B1(n7196), .B2(P1_U3084), .C1(
        n8199), .C2(n8444), .ZN(P1_U3343) );
  INV_X1 U8822 ( .A(n7027), .ZN(n7236) );
  OAI222_X1 U8823 ( .A1(n10232), .A2(n7028), .B1(n7236), .B2(P1_U3084), .C1(
        n8178), .C2(n8444), .ZN(P1_U3342) );
  NAND2_X1 U8824 ( .A1(n10339), .A2(n7029), .ZN(n7030) );
  NAND2_X1 U8825 ( .A1(n7030), .A2(n5799), .ZN(n7031) );
  OAI21_X1 U8826 ( .B1(n7032), .B2(n10339), .A(n7031), .ZN(n9097) );
  NOR2_X1 U8827 ( .A1(n9056), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8828 ( .A(n7331), .ZN(n7293) );
  OAI222_X1 U8829 ( .A1(n9508), .A2(n7034), .B1(n9511), .B2(n7033), .C1(n7293), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8830 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U8831 ( .A1(P2_U3966), .A2(n8451), .ZN(n7035) );
  OAI21_X1 U8832 ( .B1(P2_U3966), .B2(n8109), .A(n7035), .ZN(P2_U3583) );
  XOR2_X1 U8833 ( .A(n7037), .B(n7036), .Z(n7045) );
  NAND2_X1 U8834 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7648) );
  OAI21_X1 U8835 ( .B1(n9741), .B2(n7038), .A(n7648), .ZN(n7039) );
  AOI21_X1 U8836 ( .B1(n9733), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7039), .ZN(
        n7044) );
  INV_X1 U8837 ( .A(n9745), .ZN(n9699) );
  OAI211_X1 U8838 ( .C1(n7042), .C2(n7041), .A(n7040), .B(n9699), .ZN(n7043)
         );
  OAI211_X1 U8839 ( .C1(n7045), .C2(n9746), .A(n7044), .B(n7043), .ZN(P1_U3249) );
  NAND2_X1 U8840 ( .A1(n7047), .A2(n7046), .ZN(n7048) );
  AOI21_X1 U8841 ( .B1(n10292), .B2(n8561), .A(n7048), .ZN(n7247) );
  NOR2_X1 U8842 ( .A1(n7245), .A2(n7049), .ZN(n7050) );
  INV_X1 U8843 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8032) );
  AND2_X1 U8844 ( .A1(n7366), .A2(n9676), .ZN(n8562) );
  NOR2_X1 U8845 ( .A1(n7361), .A2(n8562), .ZN(n8476) );
  NAND2_X1 U8846 ( .A1(n8725), .A2(n7054), .ZN(n7052) );
  OAI22_X1 U8847 ( .A1(n8476), .A2(n7052), .B1(n7051), .B2(n10017), .ZN(n7147)
         );
  INV_X1 U8848 ( .A(n7147), .ZN(n7053) );
  OAI21_X1 U8849 ( .B1(n7366), .B2(n7054), .A(n7053), .ZN(n10187) );
  NAND2_X1 U8850 ( .A1(n10187), .A2(n10301), .ZN(n7055) );
  OAI21_X1 U8851 ( .B1(n10301), .B2(n8032), .A(n7055), .ZN(P1_U3454) );
  INV_X1 U8852 ( .A(n7056), .ZN(n7058) );
  OAI222_X1 U8853 ( .A1(n8444), .A2(n7057), .B1(n10232), .B2(n7058), .C1(
        P1_U3084), .C2(n7543), .ZN(P1_U3341) );
  OAI222_X1 U8854 ( .A1(n9508), .A2(n7059), .B1(n9511), .B2(n7058), .C1(
        P2_U3152), .C2(n7371), .ZN(P2_U3346) );
  XOR2_X1 U8855 ( .A(n7061), .B(n7060), .Z(n7069) );
  INV_X1 U8856 ( .A(n9746), .ZN(n9695) );
  OAI21_X1 U8857 ( .B1(n7063), .B2(n4475), .A(n7062), .ZN(n7067) );
  INV_X1 U8858 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8341) );
  INV_X1 U8859 ( .A(n9741), .ZN(n9696) );
  AND2_X1 U8860 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7563) );
  AOI21_X1 U8861 ( .B1(n9696), .B2(n7064), .A(n7563), .ZN(n7065) );
  OAI21_X1 U8862 ( .B1(n8341), .B2(n10245), .A(n7065), .ZN(n7066) );
  AOI21_X1 U8863 ( .B1(n9695), .B2(n7067), .A(n7066), .ZN(n7068) );
  OAI21_X1 U8864 ( .B1(n9745), .B2(n7069), .A(n7068), .ZN(P1_U3248) );
  INV_X1 U8865 ( .A(n7070), .ZN(n7071) );
  AOI21_X1 U8866 ( .B1(n7073), .B2(n7072), .A(n7071), .ZN(n7082) );
  NAND2_X1 U8867 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7460) );
  OAI21_X1 U8868 ( .B1(n9741), .B2(n7074), .A(n7460), .ZN(n7075) );
  AOI21_X1 U8869 ( .B1(n9733), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7075), .ZN(
        n7081) );
  NAND2_X1 U8870 ( .A1(n7077), .A2(n7076), .ZN(n7078) );
  NAND3_X1 U8871 ( .A1(n9695), .A2(n7079), .A3(n7078), .ZN(n7080) );
  OAI211_X1 U8872 ( .C1(n7082), .C2(n9745), .A(n7081), .B(n7080), .ZN(P1_U3247) );
  OAI211_X1 U8873 ( .C1(n7085), .C2(n7084), .A(n9699), .B(n7083), .ZN(n7086)
         );
  OAI21_X1 U8874 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n5086), .A(n7086), .ZN(n7087) );
  AOI21_X1 U8875 ( .B1(n9733), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n7087), .ZN(
        n7092) );
  OAI211_X1 U8876 ( .C1(n7090), .C2(n7089), .A(n9695), .B(n7088), .ZN(n7091)
         );
  OAI211_X1 U8877 ( .C1(n9741), .C2(n7093), .A(n7092), .B(n7091), .ZN(P1_U3242) );
  INV_X1 U8878 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8343) );
  OAI211_X1 U8879 ( .C1(n7096), .C2(n7095), .A(n9699), .B(n7094), .ZN(n7098)
         );
  INV_X1 U8880 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7416) );
  NOR2_X1 U8881 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7416), .ZN(n7175) );
  INV_X1 U8882 ( .A(n7175), .ZN(n7097) );
  OAI211_X1 U8883 ( .C1(n8343), .C2(n10245), .A(n7098), .B(n7097), .ZN(n7099)
         );
  INV_X1 U8884 ( .A(n7099), .ZN(n7104) );
  OAI211_X1 U8885 ( .C1(n7102), .C2(n7101), .A(n9695), .B(n7100), .ZN(n7103)
         );
  OAI211_X1 U8886 ( .C1(n9741), .C2(n7105), .A(n7104), .B(n7103), .ZN(P1_U3244) );
  OAI21_X1 U8887 ( .B1(n7108), .B2(n7107), .A(n7106), .ZN(n7109) );
  OAI22_X1 U8888 ( .A1(n9745), .A2(n7109), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5115), .ZN(n7116) );
  OAI21_X1 U8889 ( .B1(n7112), .B2(n7111), .A(n7110), .ZN(n7113) );
  OAI22_X1 U8890 ( .A1(n7114), .A2(n9741), .B1(n9746), .B2(n7113), .ZN(n7115)
         );
  AOI211_X1 U8891 ( .C1(n9733), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n7116), .B(
        n7115), .ZN(n7124) );
  OAI21_X1 U8892 ( .B1(n7119), .B2(n7118), .A(n7117), .ZN(n7181) );
  MUX2_X1 U8893 ( .A(n7181), .B(n7120), .S(n10239), .Z(n7123) );
  INV_X1 U8894 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U8895 ( .A1(n10239), .A2(n7150), .ZN(n7121) );
  NAND2_X1 U8896 ( .A1(n10226), .A2(n7121), .ZN(n10237) );
  NAND2_X1 U8897 ( .A1(n10237), .A2(n10240), .ZN(n7122) );
  OAI211_X1 U8898 ( .C1(n7123), .C2(n4391), .A(P1_U4006), .B(n7122), .ZN(n9689) );
  NAND2_X1 U8899 ( .A1(n7124), .A2(n9689), .ZN(P1_U3243) );
  INV_X1 U8900 ( .A(n7125), .ZN(n7143) );
  INV_X1 U8901 ( .A(n7126), .ZN(n7666) );
  INV_X1 U8902 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8024) );
  OAI222_X1 U8903 ( .A1(n10232), .A2(n7143), .B1(n7666), .B2(P1_U3084), .C1(
        n8024), .C2(n8444), .ZN(P1_U3340) );
  NAND2_X1 U8904 ( .A1(n7128), .A2(n7127), .ZN(n7129) );
  XOR2_X1 U8905 ( .A(n7130), .B(n7129), .Z(n7137) );
  INV_X1 U8906 ( .A(n7245), .ZN(n7132) );
  NAND3_X1 U8907 ( .A1(n7133), .A2(n7132), .A3(n7131), .ZN(n7180) );
  AOI22_X1 U8908 ( .A1(n4380), .A2(n7368), .B1(n7180), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7136) );
  AOI22_X1 U8909 ( .A1(n9604), .A2(n9676), .B1(n9632), .B2(n7134), .ZN(n7135)
         );
  OAI211_X1 U8910 ( .C1(n7137), .C2(n9636), .A(n7136), .B(n7135), .ZN(P1_U3220) );
  XOR2_X1 U8911 ( .A(n7138), .B(n7139), .Z(n7142) );
  AOI22_X1 U8912 ( .A1(n4380), .A2(n7258), .B1(n7180), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7141) );
  AOI22_X1 U8913 ( .A1(n9604), .A2(n6650), .B1(n9632), .B2(n9675), .ZN(n7140)
         );
  OAI211_X1 U8914 ( .C1(n7142), .C2(n9636), .A(n7141), .B(n7140), .ZN(P1_U3235) );
  INV_X1 U8915 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7144) );
  INV_X1 U8916 ( .A(n7375), .ZN(n7431) );
  OAI222_X1 U8917 ( .A1(n9508), .A2(n7144), .B1(n9511), .B2(n7143), .C1(n7431), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8918 ( .A(n7145), .ZN(n7151) );
  OAI222_X1 U8919 ( .A1(n10232), .A2(n7151), .B1(n7773), .B2(P1_U3084), .C1(
        n7146), .C2(n8444), .ZN(P1_U3339) );
  NOR2_X2 U8920 ( .A1(n9903), .A2(n10287), .ZN(n10060) );
  OAI21_X1 U8921 ( .B1(n10060), .B2(n9920), .A(n7179), .ZN(n7149) );
  AOI22_X1 U8922 ( .A1(n7147), .A2(n9940), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10051), .ZN(n7148) );
  OAI211_X1 U8923 ( .C1(n9940), .C2(n7150), .A(n7149), .B(n7148), .ZN(P1_U3291) );
  INV_X1 U8924 ( .A(n7812), .ZN(n7804) );
  OAI222_X1 U8925 ( .A1(n9508), .A2(n8140), .B1(n9511), .B2(n7151), .C1(n7804), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8926 ( .A(n7152), .ZN(n7155) );
  INV_X1 U8927 ( .A(n8259), .ZN(n7807) );
  OAI222_X1 U8928 ( .A1(n9508), .A2(n7153), .B1(n9511), .B2(n7155), .C1(
        P2_U3152), .C2(n7807), .ZN(P2_U3343) );
  OAI222_X1 U8929 ( .A1(n8444), .A2(n7156), .B1(n10232), .B2(n7155), .C1(
        P1_U3084), .C2(n4673), .ZN(P1_U3338) );
  INV_X1 U8930 ( .A(n7157), .ZN(n7158) );
  AOI21_X1 U8931 ( .B1(n7160), .B2(n7159), .A(n7158), .ZN(n7169) );
  NAND2_X1 U8932 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7850) );
  OAI21_X1 U8933 ( .B1(n9741), .B2(n7161), .A(n7850), .ZN(n7167) );
  INV_X1 U8934 ( .A(n7162), .ZN(n7163) );
  AOI211_X1 U8935 ( .C1(n7165), .C2(n7164), .A(n9746), .B(n7163), .ZN(n7166)
         );
  AOI211_X1 U8936 ( .C1(n9733), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7167), .B(
        n7166), .ZN(n7168) );
  OAI21_X1 U8937 ( .B1(n7169), .B2(n9745), .A(n7168), .ZN(P1_U3250) );
  XNOR2_X1 U8938 ( .A(n7171), .B(n7170), .ZN(n7172) );
  NAND2_X1 U8939 ( .A1(n7172), .A2(n9650), .ZN(n7178) );
  OAI22_X1 U8940 ( .A1(n7173), .A2(n9657), .B1(n9654), .B2(n7397), .ZN(n7174)
         );
  AOI211_X1 U8941 ( .C1(n7176), .C2(n4380), .A(n7175), .B(n7174), .ZN(n7177)
         );
  OAI211_X1 U8942 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9629), .A(n7178), .B(
        n7177), .ZN(P1_U3216) );
  AOI22_X1 U8943 ( .A1(n9632), .A2(n6650), .B1(n7179), .B2(n4380), .ZN(n7183)
         );
  AOI22_X1 U8944 ( .A1(n7181), .A2(n9650), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7180), .ZN(n7182) );
  NAND2_X1 U8945 ( .A1(n7183), .A2(n7182), .ZN(P1_U3230) );
  INV_X1 U8946 ( .A(n7184), .ZN(n7187) );
  OAI222_X1 U8947 ( .A1(n10232), .A2(n7187), .B1(n7186), .B2(P1_U3084), .C1(
        n7185), .C2(n8444), .ZN(P1_U3337) );
  INV_X1 U8948 ( .A(n9061), .ZN(n8256) );
  OAI222_X1 U8949 ( .A1(n9508), .A2(n8191), .B1(n9511), .B2(n7187), .C1(n8256), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  AOI21_X1 U8950 ( .B1(n7188), .B2(n7189), .A(n9636), .ZN(n7190) );
  AND2_X1 U8951 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9682) );
  OAI22_X1 U8952 ( .A1(n7445), .A2(n9657), .B1(n9654), .B2(n7461), .ZN(n7191)
         );
  AOI211_X1 U8953 ( .C1(n7466), .C2(n4380), .A(n9682), .B(n7191), .ZN(n7192)
         );
  OAI211_X1 U8954 ( .C1(n9629), .C2(n7453), .A(n7193), .B(n7192), .ZN(P1_U3228) );
  XOR2_X1 U8955 ( .A(n7195), .B(n7194), .Z(n7204) );
  NAND2_X1 U8956 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7947) );
  OAI21_X1 U8957 ( .B1(n9741), .B2(n7196), .A(n7947), .ZN(n7202) );
  OAI211_X1 U8958 ( .C1(n7199), .C2(n7198), .A(n7197), .B(n9695), .ZN(n7200)
         );
  INV_X1 U8959 ( .A(n7200), .ZN(n7201) );
  AOI211_X1 U8960 ( .C1(n9733), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n7202), .B(
        n7201), .ZN(n7203) );
  OAI21_X1 U8961 ( .B1(n9745), .B2(n7204), .A(n7203), .ZN(P1_U3251) );
  INV_X1 U8962 ( .A(n7205), .ZN(n7242) );
  INV_X1 U8963 ( .A(n9728), .ZN(n9716) );
  OAI222_X1 U8964 ( .A1(n10232), .A2(n7242), .B1(n9716), .B2(P1_U3084), .C1(
        n8034), .C2(n8444), .ZN(P1_U3336) );
  NAND2_X1 U8965 ( .A1(n10339), .A2(n7206), .ZN(n7209) );
  INV_X1 U8966 ( .A(n7207), .ZN(n7208) );
  NAND3_X1 U8967 ( .A1(n7209), .A2(n8241), .A3(n7208), .ZN(n7213) );
  NAND2_X1 U8968 ( .A1(n7213), .A2(n5799), .ZN(n7210) );
  NAND2_X1 U8969 ( .A1(n7210), .A2(n8917), .ZN(n7224) );
  NAND2_X1 U8970 ( .A1(n7224), .A2(n9503), .ZN(n9090) );
  INV_X1 U8971 ( .A(n7265), .ZN(n7270) );
  INV_X1 U8972 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n8346) );
  XNOR2_X1 U8973 ( .A(n7265), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n7215) );
  INV_X1 U8974 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10409) );
  MUX2_X1 U8975 ( .A(n10409), .B(P2_REG1_REG_1__SCAN_IN), .S(n8931), .Z(n8939)
         );
  AND2_X1 U8976 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8938) );
  NAND2_X1 U8977 ( .A1(n8939), .A2(n8938), .ZN(n8937) );
  INV_X1 U8978 ( .A(n8931), .ZN(n8936) );
  NAND2_X1 U8979 ( .A1(n8936), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7211) );
  NAND2_X1 U8980 ( .A1(n8937), .A2(n7211), .ZN(n7214) );
  INV_X1 U8981 ( .A(n7221), .ZN(n9507) );
  AND2_X1 U8982 ( .A1(n9507), .A2(n5799), .ZN(n7212) );
  NAND2_X1 U8983 ( .A1(n7214), .A2(n7215), .ZN(n7272) );
  OAI211_X1 U8984 ( .C1(n7215), .C2(n7214), .A(n9088), .B(n7272), .ZN(n7217)
         );
  INV_X1 U8985 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U8986 ( .A1(P2_U3152), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7216) );
  OAI211_X1 U8987 ( .C1(n8346), .C2(n9097), .A(n7217), .B(n7216), .ZN(n7228)
         );
  INV_X1 U8988 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10334) );
  INV_X1 U8989 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7219) );
  INV_X1 U8990 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7218) );
  NOR3_X1 U8991 ( .A1(n7220), .A2(n7219), .A3(n7218), .ZN(n8932) );
  AOI21_X1 U8992 ( .B1(n8936), .B2(P2_REG2_REG_1__SCAN_IN), .A(n8932), .ZN(
        n7226) );
  INV_X1 U8993 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7710) );
  MUX2_X1 U8994 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7710), .S(n7265), .Z(n7225)
         );
  NOR2_X1 U8995 ( .A1(n7226), .A2(n7225), .ZN(n8950) );
  AND2_X1 U8996 ( .A1(n7222), .A2(n7221), .ZN(n7223) );
  AOI211_X1 U8997 ( .C1(n7226), .C2(n7225), .A(n8950), .B(n9094), .ZN(n7227)
         );
  AOI211_X1 U8998 ( .C1(n9077), .C2(n7270), .A(n7228), .B(n7227), .ZN(n7229)
         );
  INV_X1 U8999 ( .A(n7229), .ZN(P2_U3247) );
  XOR2_X1 U9000 ( .A(n7231), .B(n7230), .Z(n7241) );
  OAI21_X1 U9001 ( .B1(n7234), .B2(n7233), .A(n7232), .ZN(n7239) );
  INV_X1 U9002 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7235) );
  NOR2_X1 U9003 ( .A1(n10245), .A2(n7235), .ZN(n7238) );
  NAND2_X1 U9004 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7907) );
  OAI21_X1 U9005 ( .B1(n9741), .B2(n7236), .A(n7907), .ZN(n7237) );
  AOI211_X1 U9006 ( .C1(n7239), .C2(n9695), .A(n7238), .B(n7237), .ZN(n7240)
         );
  OAI21_X1 U9007 ( .B1(n9745), .B2(n7241), .A(n7240), .ZN(P1_U3252) );
  INV_X1 U9008 ( .A(n9072), .ZN(n9059) );
  OAI222_X1 U9009 ( .A1(n9508), .A2(n7243), .B1(n9511), .B2(n7242), .C1(n9059), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NOR2_X1 U9010 ( .A1(n7245), .A2(n7244), .ZN(n7246) );
  INV_X1 U9011 ( .A(n8473), .ZN(n7357) );
  INV_X1 U9012 ( .A(n7249), .ZN(n7356) );
  NAND2_X1 U9013 ( .A1(n7357), .A2(n7356), .ZN(n7355) );
  NAND2_X1 U9014 ( .A1(n6650), .A2(n7368), .ZN(n7250) );
  NAND2_X1 U9015 ( .A1(n7355), .A2(n7250), .ZN(n7251) );
  XNOR2_X1 U9016 ( .A(n7251), .B(n8474), .ZN(n7426) );
  INV_X1 U9017 ( .A(n7426), .ZN(n7260) );
  NAND2_X1 U9018 ( .A1(n7252), .A2(n9857), .ZN(n10000) );
  INV_X1 U9019 ( .A(n10000), .ZN(n10048) );
  XOR2_X1 U9020 ( .A(n8564), .B(n8474), .Z(n7254) );
  AOI22_X1 U9021 ( .A1(n10043), .A2(n9675), .B1(n10041), .B2(n6650), .ZN(n7253) );
  OAI21_X1 U9022 ( .B1(n7254), .B2(n10045), .A(n7253), .ZN(n7255) );
  AOI21_X1 U9023 ( .B1(n10048), .B2(n7426), .A(n7255), .ZN(n7428) );
  INV_X1 U9024 ( .A(n7256), .ZN(n7365) );
  INV_X1 U9025 ( .A(n7257), .ZN(n7406) );
  AOI21_X1 U9026 ( .B1(n7258), .B2(n7365), .A(n7406), .ZN(n7421) );
  AOI22_X1 U9027 ( .A1(n7421), .A2(n10181), .B1(n10180), .B2(n7258), .ZN(n7259) );
  OAI211_X1 U9028 ( .C1(n10186), .C2(n7260), .A(n7428), .B(n7259), .ZN(n7262)
         );
  NAND2_X1 U9029 ( .A1(n7262), .A2(n10308), .ZN(n7261) );
  OAI21_X1 U9030 ( .B1(n10308), .B2(n6938), .A(n7261), .ZN(P1_U3525) );
  INV_X1 U9031 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U9032 ( .A1(n7262), .A2(n10301), .ZN(n7263) );
  OAI21_X1 U9033 ( .B1(n10301), .B2(n7264), .A(n7263), .ZN(P1_U3460) );
  NOR2_X1 U9034 ( .A1(n7265), .A2(n7710), .ZN(n8945) );
  INV_X1 U9035 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7749) );
  MUX2_X1 U9036 ( .A(n7749), .B(P2_REG2_REG_3__SCAN_IN), .S(n8944), .Z(n7266)
         );
  OAI21_X1 U9037 ( .B1(n8950), .B2(n8945), .A(n7266), .ZN(n8948) );
  INV_X1 U9038 ( .A(n8944), .ZN(n8951) );
  NAND2_X1 U9039 ( .A1(n8951), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7268) );
  INV_X1 U9040 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7281) );
  MUX2_X1 U9041 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7281), .S(n7296), .Z(n7267)
         );
  INV_X1 U9042 ( .A(n7283), .ZN(n8963) );
  NAND3_X1 U9043 ( .A1(n8948), .A2(n7268), .A3(n7267), .ZN(n7269) );
  NAND3_X1 U9044 ( .A1(n9051), .A2(n8963), .A3(n7269), .ZN(n7280) );
  INV_X1 U9045 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7277) );
  INV_X1 U9046 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10415) );
  MUX2_X1 U9047 ( .A(n10415), .B(P2_REG1_REG_4__SCAN_IN), .S(n7296), .Z(n7275)
         );
  NAND2_X1 U9048 ( .A1(n7270), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7271) );
  NAND2_X1 U9049 ( .A1(n7272), .A2(n7271), .ZN(n8953) );
  XNOR2_X1 U9050 ( .A(n8944), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U9051 ( .A1(n8953), .A2(n8954), .ZN(n8952) );
  NAND2_X1 U9052 ( .A1(n8951), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7273) );
  NAND2_X1 U9053 ( .A1(n8952), .A2(n7273), .ZN(n7274) );
  NAND2_X1 U9054 ( .A1(n7274), .A2(n7275), .ZN(n7298) );
  OAI211_X1 U9055 ( .C1(n7275), .C2(n7274), .A(n9088), .B(n7298), .ZN(n7276)
         );
  NAND2_X1 U9056 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7527) );
  OAI211_X1 U9057 ( .C1(n9097), .C2(n7277), .A(n7276), .B(n7527), .ZN(n7278)
         );
  INV_X1 U9058 ( .A(n7278), .ZN(n7279) );
  OAI211_X1 U9059 ( .C1(n9090), .C2(n7296), .A(n7280), .B(n7279), .ZN(P2_U3249) );
  NOR2_X1 U9060 ( .A1(n7296), .A2(n7281), .ZN(n8959) );
  INV_X1 U9061 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7735) );
  MUX2_X1 U9062 ( .A(n7735), .B(P2_REG2_REG_5__SCAN_IN), .S(n8960), .Z(n7282)
         );
  NAND2_X1 U9063 ( .A1(n8965), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8975) );
  INV_X1 U9064 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7284) );
  MUX2_X1 U9065 ( .A(n7284), .B(P2_REG2_REG_6__SCAN_IN), .S(n8979), .Z(n8974)
         );
  NOR2_X1 U9066 ( .A1(n7285), .A2(n7284), .ZN(n8990) );
  INV_X1 U9067 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7858) );
  MUX2_X1 U9068 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7858), .S(n8995), .Z(n8989)
         );
  NAND2_X1 U9069 ( .A1(n8995), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9004) );
  INV_X1 U9070 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7286) );
  MUX2_X1 U9071 ( .A(n7286), .B(P2_REG2_REG_8__SCAN_IN), .S(n7303), .Z(n9003)
         );
  AOI21_X1 U9072 ( .B1(n9005), .B2(n9004), .A(n9003), .ZN(n9023) );
  NOR2_X1 U9073 ( .A1(n9009), .A2(n7286), .ZN(n9018) );
  INV_X1 U9074 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7287) );
  MUX2_X1 U9075 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7287), .S(n9029), .Z(n7288)
         );
  NAND2_X1 U9076 ( .A1(n9029), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7291) );
  INV_X1 U9077 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7289) );
  MUX2_X1 U9078 ( .A(n7289), .B(P2_REG2_REG_10__SCAN_IN), .S(n7331), .Z(n7290)
         );
  NAND3_X1 U9079 ( .A1(n9021), .A2(n7291), .A3(n7290), .ZN(n7292) );
  NAND2_X1 U9080 ( .A1(n7292), .A2(n9051), .ZN(n7310) );
  NOR2_X1 U9081 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7784), .ZN(n7295) );
  NOR2_X1 U9082 ( .A1(n9090), .A2(n7293), .ZN(n7294) );
  AOI211_X1 U9083 ( .C1(n9056), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7295), .B(
        n7294), .ZN(n7309) );
  OR2_X1 U9084 ( .A1(n7296), .A2(n10415), .ZN(n7297) );
  NAND2_X1 U9085 ( .A1(n7298), .A2(n7297), .ZN(n8968) );
  XNOR2_X1 U9086 ( .A(n8960), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U9087 ( .A1(n8968), .A2(n8969), .ZN(n8967) );
  NAND2_X1 U9088 ( .A1(n8965), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7299) );
  NAND2_X1 U9089 ( .A1(n8967), .A2(n7299), .ZN(n8983) );
  INV_X1 U9090 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7300) );
  XNOR2_X1 U9091 ( .A(n8979), .B(n7300), .ZN(n8984) );
  NAND2_X1 U9092 ( .A1(n8983), .A2(n8984), .ZN(n8982) );
  NAND2_X1 U9093 ( .A1(n8979), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7301) );
  NAND2_X1 U9094 ( .A1(n8982), .A2(n7301), .ZN(n8997) );
  INV_X1 U9095 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8091) );
  MUX2_X1 U9096 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8091), .S(n8995), .Z(n8998)
         );
  NAND2_X1 U9097 ( .A1(n8997), .A2(n8998), .ZN(n8996) );
  NAND2_X1 U9098 ( .A1(n8995), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7302) );
  NAND2_X1 U9099 ( .A1(n8996), .A2(n7302), .ZN(n9013) );
  INV_X1 U9100 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10421) );
  MUX2_X1 U9101 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10421), .S(n7303), .Z(n9014)
         );
  NAND2_X1 U9102 ( .A1(n9013), .A2(n9014), .ZN(n9012) );
  NAND2_X1 U9103 ( .A1(n7303), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7304) );
  NAND2_X1 U9104 ( .A1(n9012), .A2(n7304), .ZN(n9028) );
  INV_X1 U9105 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7892) );
  MUX2_X1 U9106 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7892), .S(n9029), .Z(n9027)
         );
  NAND2_X1 U9107 ( .A1(n9028), .A2(n9027), .ZN(n9026) );
  NAND2_X1 U9108 ( .A1(n9029), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7305) );
  NAND2_X1 U9109 ( .A1(n9026), .A2(n7305), .ZN(n7307) );
  INV_X1 U9110 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7941) );
  XNOR2_X1 U9111 ( .A(n7331), .B(n7941), .ZN(n7306) );
  NAND2_X1 U9112 ( .A1(n7307), .A2(n7306), .ZN(n7322) );
  OAI211_X1 U9113 ( .C1(n7307), .C2(n7306), .A(n7322), .B(n9088), .ZN(n7308)
         );
  OAI211_X1 U9114 ( .C1(n7330), .C2(n7310), .A(n7309), .B(n7308), .ZN(P2_U3255) );
  NAND2_X1 U9115 ( .A1(n7312), .A2(n7311), .ZN(n8892) );
  INV_X1 U9116 ( .A(n8892), .ZN(n7320) );
  INV_X1 U9117 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7658) );
  AOI22_X1 U9118 ( .A1(n8874), .A2(n7313), .B1(n10353), .B2(n8908), .ZN(n7319)
         );
  OAI21_X1 U9119 ( .B1(n7315), .B2(n7314), .A(n7663), .ZN(n7316) );
  NAND3_X1 U9120 ( .A1(n8888), .A2(n7317), .A3(n7316), .ZN(n7318) );
  OAI211_X1 U9121 ( .C1(n7320), .C2(n7658), .A(n7319), .B(n7318), .ZN(P2_U3234) );
  INV_X1 U9122 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8164) );
  XNOR2_X1 U9123 ( .A(n7371), .B(n8164), .ZN(n7327) );
  NAND2_X1 U9124 ( .A1(n7331), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7321) );
  NAND2_X1 U9125 ( .A1(n7322), .A2(n7321), .ZN(n9041) );
  INV_X1 U9126 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7323) );
  XNOR2_X1 U9127 ( .A(n9042), .B(n7323), .ZN(n9040) );
  NAND2_X1 U9128 ( .A1(n9041), .A2(n9040), .ZN(n9039) );
  NAND2_X1 U9129 ( .A1(n9042), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U9130 ( .A1(n9039), .A2(n7324), .ZN(n7326) );
  INV_X1 U9131 ( .A(n7373), .ZN(n7325) );
  AOI21_X1 U9132 ( .B1(n7327), .B2(n7326), .A(n7325), .ZN(n7339) );
  INV_X1 U9133 ( .A(n9088), .ZN(n9092) );
  INV_X1 U9134 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7329) );
  AND2_X1 U9135 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8787) );
  INV_X1 U9136 ( .A(n8787), .ZN(n7328) );
  OAI21_X1 U9137 ( .B1(n9097), .B2(n7329), .A(n7328), .ZN(n7337) );
  INV_X1 U9138 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7332) );
  MUX2_X1 U9139 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7332), .S(n9042), .Z(n9036)
         );
  OAI21_X1 U9140 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n9042), .A(n9034), .ZN(
        n7335) );
  INV_X1 U9141 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7333) );
  MUX2_X1 U9142 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7333), .S(n7371), .Z(n7334)
         );
  NOR2_X1 U9143 ( .A1(n7335), .A2(n7334), .ZN(n7377) );
  AOI211_X1 U9144 ( .C1(n7335), .C2(n7334), .A(n9094), .B(n7377), .ZN(n7336)
         );
  AOI211_X1 U9145 ( .C1(n9077), .C2(n7378), .A(n7337), .B(n7336), .ZN(n7338)
         );
  OAI21_X1 U9146 ( .B1(n7339), .B2(n9092), .A(n7338), .ZN(P2_U3257) );
  XNOR2_X1 U9147 ( .A(n7341), .B(n7340), .ZN(n8764) );
  INV_X1 U9148 ( .A(n7342), .ZN(n8765) );
  NAND2_X1 U9149 ( .A1(n8764), .A2(n8765), .ZN(n8763) );
  NAND2_X1 U9150 ( .A1(n8763), .A2(n7343), .ZN(n7347) );
  NAND2_X1 U9151 ( .A1(n7345), .A2(n7344), .ZN(n7346) );
  XNOR2_X1 U9152 ( .A(n7347), .B(n7346), .ZN(n7350) );
  AOI22_X1 U9153 ( .A1(n8903), .A2(n7313), .B1(n8874), .B2(n8930), .ZN(n7349)
         );
  AOI22_X1 U9154 ( .A1(n8908), .A2(n7720), .B1(n8892), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7348) );
  OAI211_X1 U9155 ( .C1(n8910), .C2(n7350), .A(n7349), .B(n7348), .ZN(P2_U3239) );
  INV_X1 U9156 ( .A(n7351), .ZN(n7354) );
  AOI22_X1 U9157 ( .A1(n9083), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9499), .ZN(n7352) );
  OAI21_X1 U9158 ( .B1(n7354), .B2(n9506), .A(n7352), .ZN(P2_U3340) );
  AOI22_X1 U9159 ( .A1(n9739), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10230), .ZN(n7353) );
  OAI21_X1 U9160 ( .B1(n7354), .B2(n10232), .A(n7353), .ZN(P1_U3335) );
  OAI21_X1 U9161 ( .B1(n7357), .B2(n7356), .A(n7355), .ZN(n10280) );
  NOR2_X1 U9162 ( .A1(n7358), .A2(n9857), .ZN(n7359) );
  NAND2_X1 U9163 ( .A1(n9940), .A2(n7359), .ZN(n10057) );
  AOI22_X1 U9164 ( .A1(n10043), .A2(n7134), .B1(n10041), .B2(n9676), .ZN(n7364) );
  OAI21_X1 U9165 ( .B1(n7361), .B2(n8473), .A(n7360), .ZN(n7362) );
  NAND2_X1 U9166 ( .A1(n7362), .A2(n4705), .ZN(n7363) );
  OAI211_X1 U9167 ( .C1(n10280), .C2(n10000), .A(n7364), .B(n7363), .ZN(n10283) );
  OAI211_X1 U9168 ( .C1(n10282), .C2(n7366), .A(n10181), .B(n7365), .ZN(n10281) );
  OAI22_X1 U9169 ( .A1(n10281), .A2(n8502), .B1(n9898), .B2(n5086), .ZN(n7367)
         );
  OAI21_X1 U9170 ( .B1(n10283), .B2(n7367), .A(n9940), .ZN(n7370) );
  AOI22_X1 U9171 ( .A1(n9920), .A2(n7368), .B1(n10062), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7369) );
  OAI211_X1 U9172 ( .C1(n10280), .C2(n10057), .A(n7370), .B(n7369), .ZN(
        P1_U3290) );
  INV_X1 U9173 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8187) );
  XNOR2_X1 U9174 ( .A(n7375), .B(n8187), .ZN(n7429) );
  NAND2_X1 U9175 ( .A1(n7371), .A2(n8164), .ZN(n7372) );
  NAND2_X1 U9176 ( .A1(n7373), .A2(n7372), .ZN(n7430) );
  XOR2_X1 U9177 ( .A(n7429), .B(n7430), .Z(n7385) );
  INV_X1 U9178 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7374) );
  NOR2_X1 U9179 ( .A1(n7431), .A2(n7374), .ZN(n7376) );
  NOR2_X1 U9180 ( .A1(n7375), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7434) );
  NOR2_X1 U9181 ( .A1(n7376), .A2(n7434), .ZN(n7380) );
  NAND2_X1 U9182 ( .A1(n7379), .A2(n7380), .ZN(n7437) );
  OAI21_X1 U9183 ( .B1(n7380), .B2(n7379), .A(n7437), .ZN(n7383) );
  NAND2_X1 U9184 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U9185 ( .A1(n9056), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7381) );
  OAI211_X1 U9186 ( .C1(n9090), .C2(n7431), .A(n8848), .B(n7381), .ZN(n7382)
         );
  AOI21_X1 U9187 ( .B1(n7383), .B2(n9051), .A(n7382), .ZN(n7384) );
  OAI21_X1 U9188 ( .B1(n9092), .B2(n7385), .A(n7384), .ZN(P2_U3258) );
  AOI22_X1 U9189 ( .A1(n9051), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9088), .ZN(n7390) );
  INV_X1 U9190 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U9191 ( .A1(n9088), .A2(n7386), .ZN(n7387) );
  OAI211_X1 U9192 ( .C1(n9094), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7387), .B(
        n9090), .ZN(n7388) );
  INV_X1 U9193 ( .A(n7388), .ZN(n7389) );
  MUX2_X1 U9194 ( .A(n7390), .B(n7389), .S(P2_IR_REG_0__SCAN_IN), .Z(n7392) );
  AOI22_X1 U9195 ( .A1(n9056), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n7391) );
  NAND2_X1 U9196 ( .A1(n7392), .A2(n7391), .ZN(P2_U3245) );
  INV_X1 U9197 ( .A(n7393), .ZN(n7394) );
  AOI21_X1 U9198 ( .B1(n7396), .B2(n7395), .A(n7394), .ZN(n7401) );
  NOR2_X1 U9199 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5176), .ZN(n9702) );
  OAI22_X1 U9200 ( .A1(n7397), .A2(n9657), .B1(n9654), .B2(n7632), .ZN(n7398)
         );
  AOI211_X1 U9201 ( .C1(n7553), .C2(n4380), .A(n9702), .B(n7398), .ZN(n7400)
         );
  NAND2_X1 U9202 ( .A1(n9660), .A2(n7516), .ZN(n7399) );
  OAI211_X1 U9203 ( .C1(n7401), .C2(n9636), .A(n7400), .B(n7399), .ZN(P1_U3225) );
  INV_X1 U9204 ( .A(n7402), .ZN(n7404) );
  OAI222_X1 U9205 ( .A1(n9508), .A2(n7403), .B1(n9511), .B2(n7404), .C1(
        P2_U3152), .C2(n9154), .ZN(P2_U3339) );
  OAI222_X1 U9206 ( .A1(n8444), .A2(n7405), .B1(n10232), .B2(n7404), .C1(n9857), .C2(P1_U3084), .ZN(P1_U3334) );
  INV_X1 U9207 ( .A(n10060), .ZN(n9923) );
  OAI21_X1 U9208 ( .B1(n7406), .B2(n10286), .A(n7452), .ZN(n10288) );
  OAI21_X1 U9209 ( .B1(n7409), .B2(n7408), .A(n7407), .ZN(n10291) );
  INV_X1 U9210 ( .A(n10291), .ZN(n7415) );
  AOI22_X1 U9211 ( .A1(n10041), .A2(n7134), .B1(n10043), .B2(n9674), .ZN(n7414) );
  OAI21_X1 U9212 ( .B1(n8475), .B2(n7410), .A(n7411), .ZN(n7412) );
  NAND2_X1 U9213 ( .A1(n7412), .A2(n4705), .ZN(n7413) );
  OAI211_X1 U9214 ( .C1(n7415), .C2(n10000), .A(n7414), .B(n7413), .ZN(n10289)
         );
  NAND2_X1 U9215 ( .A1(n10289), .A2(n9940), .ZN(n7420) );
  INV_X1 U9216 ( .A(n10057), .ZN(n8406) );
  AOI22_X1 U9217 ( .A1(n10062), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10051), .B2(
        n7416), .ZN(n7417) );
  OAI21_X1 U9218 ( .B1(n10054), .B2(n10286), .A(n7417), .ZN(n7418) );
  AOI21_X1 U9219 ( .B1(n8406), .B2(n10291), .A(n7418), .ZN(n7419) );
  OAI211_X1 U9220 ( .C1(n9923), .C2(n10288), .A(n7420), .B(n7419), .ZN(
        P1_U3288) );
  NAND2_X1 U9221 ( .A1(n10060), .A2(n7421), .ZN(n7423) );
  AOI22_X1 U9222 ( .A1(n10062), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10051), .ZN(n7422) );
  OAI211_X1 U9223 ( .C1(n7424), .C2(n10054), .A(n7423), .B(n7422), .ZN(n7425)
         );
  AOI21_X1 U9224 ( .B1(n8406), .B2(n7426), .A(n7425), .ZN(n7427) );
  OAI21_X1 U9225 ( .B1(n7428), .B2(n10062), .A(n7427), .ZN(P1_U3289) );
  INV_X1 U9226 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8177) );
  XNOR2_X1 U9227 ( .A(n7812), .B(n8177), .ZN(n7814) );
  NAND2_X1 U9228 ( .A1(n7430), .A2(n7429), .ZN(n7433) );
  NAND2_X1 U9229 ( .A1(n7431), .A2(n8187), .ZN(n7432) );
  NAND2_X1 U9230 ( .A1(n7433), .A2(n7432), .ZN(n7815) );
  XOR2_X1 U9231 ( .A(n7814), .B(n7815), .Z(n7443) );
  INV_X1 U9232 ( .A(n7434), .ZN(n7435) );
  INV_X1 U9233 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9361) );
  MUX2_X1 U9234 ( .A(n9361), .B(P2_REG2_REG_14__SCAN_IN), .S(n7812), .Z(n7436)
         );
  AOI21_X1 U9235 ( .B1(n7437), .B2(n7435), .A(n7436), .ZN(n7803) );
  AND3_X1 U9236 ( .A1(n7437), .A2(n7436), .A3(n7435), .ZN(n7438) );
  OAI21_X1 U9237 ( .B1(n7803), .B2(n7438), .A(n9051), .ZN(n7442) );
  INV_X1 U9238 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7439) );
  NAND2_X1 U9239 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8746) );
  OAI21_X1 U9240 ( .B1(n9097), .B2(n7439), .A(n8746), .ZN(n7440) );
  AOI21_X1 U9241 ( .B1(n9077), .B2(n7812), .A(n7440), .ZN(n7441) );
  OAI211_X1 U9242 ( .C1(n7443), .C2(n9092), .A(n7442), .B(n7441), .ZN(P2_U3259) );
  OAI21_X1 U9243 ( .B1(n7444), .B2(n8477), .A(n7507), .ZN(n7450) );
  INV_X1 U9244 ( .A(n7450), .ZN(n7470) );
  OAI22_X1 U9245 ( .A1(n10017), .A2(n7461), .B1(n7445), .B2(n10014), .ZN(n7449) );
  XNOR2_X1 U9246 ( .A(n7446), .B(n8477), .ZN(n7447) );
  NOR2_X1 U9247 ( .A1(n7447), .A2(n10045), .ZN(n7448) );
  AOI211_X1 U9248 ( .C1(n10048), .C2(n7450), .A(n7449), .B(n7448), .ZN(n7469)
         );
  MUX2_X1 U9249 ( .A(n7451), .B(n7469), .S(n9940), .Z(n7457) );
  AOI21_X1 U9250 ( .B1(n7466), .B2(n7452), .A(n7514), .ZN(n7467) );
  OAI22_X1 U9251 ( .A1(n10054), .A2(n7454), .B1(n9898), .B2(n7453), .ZN(n7455)
         );
  AOI21_X1 U9252 ( .B1(n10060), .B2(n7467), .A(n7455), .ZN(n7456) );
  OAI211_X1 U9253 ( .C1(n7470), .C2(n10057), .A(n7457), .B(n7456), .ZN(
        P1_U3287) );
  XOR2_X1 U9254 ( .A(n7458), .B(n7459), .Z(n7465) );
  OAI21_X1 U9255 ( .B1(n9657), .B2(n7461), .A(n7460), .ZN(n7462) );
  AOI21_X1 U9256 ( .B1(n9632), .B2(n9671), .A(n7462), .ZN(n7464) );
  AOI22_X1 U9257 ( .A1(n9660), .A2(n7757), .B1(n4380), .B2(n7758), .ZN(n7463)
         );
  OAI211_X1 U9258 ( .C1(n7465), .C2(n9636), .A(n7464), .B(n7463), .ZN(P1_U3237) );
  AOI22_X1 U9259 ( .A1(n7467), .A2(n10181), .B1(n10180), .B2(n7466), .ZN(n7468) );
  OAI211_X1 U9260 ( .C1(n7470), .C2(n10186), .A(n7469), .B(n7468), .ZN(n7472)
         );
  NAND2_X1 U9261 ( .A1(n7472), .A2(n10301), .ZN(n7471) );
  OAI21_X1 U9262 ( .B1(n10301), .B2(n5157), .A(n7471), .ZN(P1_U3466) );
  NAND2_X1 U9263 ( .A1(n7472), .A2(n10308), .ZN(n7473) );
  OAI21_X1 U9264 ( .B1(n10308), .B2(n5155), .A(n7473), .ZN(P1_U3527) );
  OAI211_X1 U9265 ( .C1(n7476), .C2(n7475), .A(n7474), .B(n8888), .ZN(n7481)
         );
  NAND2_X1 U9266 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n9008) );
  OAI21_X1 U9267 ( .B1(n8906), .B2(n7877), .A(n9008), .ZN(n7479) );
  INV_X1 U9268 ( .A(n7477), .ZN(n7885) );
  OAI22_X1 U9269 ( .A1(n8863), .A2(n7876), .B1(n8862), .B2(n7885), .ZN(n7478)
         );
  AOI211_X1 U9270 ( .C1(n8908), .C2(n10397), .A(n7479), .B(n7478), .ZN(n7480)
         );
  NAND2_X1 U9271 ( .A1(n7481), .A2(n7480), .ZN(P2_U3223) );
  OAI22_X1 U9272 ( .A1(n8906), .A2(n7731), .B1(n7482), .B2(n8897), .ZN(n7489)
         );
  INV_X1 U9273 ( .A(n7483), .ZN(n7487) );
  INV_X1 U9274 ( .A(n7521), .ZN(n7485) );
  NAND2_X1 U9275 ( .A1(n7485), .A2(n7484), .ZN(n7486) );
  NOR2_X1 U9276 ( .A1(n7487), .A2(n7486), .ZN(n7522) );
  AOI211_X1 U9277 ( .C1(n7487), .C2(n7486), .A(n8910), .B(n7522), .ZN(n7488)
         );
  AOI211_X1 U9278 ( .C1(n8903), .C2(n10315), .A(n7489), .B(n7488), .ZN(n7491)
         );
  MUX2_X1 U9279 ( .A(n8862), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n7490) );
  NAND2_X1 U9280 ( .A1(n7491), .A2(n7490), .ZN(P2_U3220) );
  OAI22_X1 U9281 ( .A1(n8897), .A2(n10383), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5860), .ZN(n7493) );
  OAI22_X1 U9282 ( .A1(n7730), .A2(n8906), .B1(n8863), .B2(n7731), .ZN(n7492)
         );
  AOI211_X1 U9283 ( .C1(n7733), .C2(n8902), .A(n7493), .B(n7492), .ZN(n7498)
         );
  OAI211_X1 U9284 ( .C1(n7496), .C2(n7495), .A(n7494), .B(n8888), .ZN(n7497)
         );
  NAND2_X1 U9285 ( .A1(n7498), .A2(n7497), .ZN(P2_U3229) );
  NAND2_X1 U9286 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9001) );
  OAI21_X1 U9287 ( .B1(n8897), .B2(n7861), .A(n9001), .ZN(n7500) );
  OAI22_X1 U9288 ( .A1(n7730), .A2(n8863), .B1(n8906), .B2(n7832), .ZN(n7499)
         );
  AOI211_X1 U9289 ( .C1(n7859), .C2(n8902), .A(n7500), .B(n7499), .ZN(n7505)
         );
  OAI211_X1 U9290 ( .C1(n7503), .C2(n7502), .A(n7501), .B(n8888), .ZN(n7504)
         );
  NAND2_X1 U9291 ( .A1(n7505), .A2(n7504), .ZN(P2_U3215) );
  NAND2_X1 U9292 ( .A1(n7507), .A2(n7506), .ZN(n7509) );
  INV_X1 U9293 ( .A(n8478), .ZN(n7508) );
  NAND2_X1 U9294 ( .A1(n7509), .A2(n7508), .ZN(n7510) );
  NAND2_X1 U9295 ( .A1(n7591), .A2(n7510), .ZN(n7556) );
  NAND2_X1 U9296 ( .A1(n7511), .A2(n8514), .ZN(n7512) );
  XNOR2_X1 U9297 ( .A(n7512), .B(n8478), .ZN(n7513) );
  AOI222_X1 U9298 ( .A1(n4705), .A2(n7513), .B1(n9672), .B2(n10043), .C1(n9674), .C2(n10041), .ZN(n7555) );
  INV_X1 U9299 ( .A(n7514), .ZN(n7515) );
  AOI211_X1 U9300 ( .C1(n7553), .C2(n7515), .A(n10287), .B(n7596), .ZN(n7552)
         );
  AOI22_X1 U9301 ( .A1(n7552), .A2(n9857), .B1(n10051), .B2(n7516), .ZN(n7517)
         );
  AOI21_X1 U9302 ( .B1(n7555), .B2(n7517), .A(n10062), .ZN(n7518) );
  INV_X1 U9303 ( .A(n7518), .ZN(n7520) );
  AOI22_X1 U9304 ( .A1(n9920), .A2(n7553), .B1(n10062), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n7519) );
  OAI211_X1 U9305 ( .C1(n7556), .C2(n10028), .A(n7520), .B(n7519), .ZN(
        P1_U3286) );
  NOR2_X1 U9306 ( .A1(n7522), .A2(n7521), .ZN(n7526) );
  XNOR2_X1 U9307 ( .A(n7524), .B(n7523), .ZN(n7525) );
  XNOR2_X1 U9308 ( .A(n7526), .B(n7525), .ZN(n7531) );
  OAI21_X1 U9309 ( .B1(n8897), .B2(n6497), .A(n7527), .ZN(n7529) );
  OAI22_X1 U9310 ( .A1(n5808), .A2(n8863), .B1(n8906), .B2(n7536), .ZN(n7528)
         );
  AOI211_X1 U9311 ( .C1(n7685), .C2(n8902), .A(n7529), .B(n7528), .ZN(n7530)
         );
  OAI21_X1 U9312 ( .B1(n8910), .B2(n7531), .A(n7530), .ZN(P2_U3232) );
  INV_X1 U9313 ( .A(n7532), .ZN(n7533) );
  AOI21_X1 U9314 ( .B1(n7535), .B2(n7534), .A(n7533), .ZN(n7540) );
  NAND2_X1 U9315 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8980) );
  OAI21_X1 U9316 ( .B1(n8897), .B2(n10391), .A(n8980), .ZN(n7538) );
  OAI22_X1 U9317 ( .A1(n7536), .A2(n8863), .B1(n8906), .B2(n7876), .ZN(n7537)
         );
  AOI211_X1 U9318 ( .C1(n7698), .C2(n8902), .A(n7538), .B(n7537), .ZN(n7539)
         );
  OAI21_X1 U9319 ( .B1(n7540), .B2(n8910), .A(n7539), .ZN(P2_U3241) );
  XOR2_X1 U9320 ( .A(n7542), .B(n7541), .Z(n7551) );
  NAND2_X1 U9321 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8246) );
  OAI21_X1 U9322 ( .B1(n9741), .B2(n7543), .A(n8246), .ZN(n7549) );
  INV_X1 U9323 ( .A(n7544), .ZN(n7545) );
  AOI211_X1 U9324 ( .C1(n7547), .C2(n7546), .A(n9746), .B(n7545), .ZN(n7548)
         );
  AOI211_X1 U9325 ( .C1(n9733), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7549), .B(
        n7548), .ZN(n7550) );
  OAI21_X1 U9326 ( .B1(n9745), .B2(n7551), .A(n7550), .ZN(P1_U3253) );
  AOI21_X1 U9327 ( .B1(n10180), .B2(n7553), .A(n7552), .ZN(n7554) );
  OAI211_X1 U9328 ( .C1(n10163), .C2(n7556), .A(n7555), .B(n7554), .ZN(n7558)
         );
  NAND2_X1 U9329 ( .A1(n7558), .A2(n10308), .ZN(n7557) );
  OAI21_X1 U9330 ( .B1(n10308), .B2(n6942), .A(n7557), .ZN(P1_U3528) );
  INV_X1 U9331 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U9332 ( .A1(n7558), .A2(n10301), .ZN(n7559) );
  OAI21_X1 U9333 ( .B1(n10301), .B2(n7560), .A(n7559), .ZN(P1_U3469) );
  XNOR2_X1 U9334 ( .A(n7562), .B(n7561), .ZN(n7569) );
  AOI21_X1 U9335 ( .B1(n9632), .B2(n9670), .A(n7563), .ZN(n7567) );
  NAND2_X1 U9336 ( .A1(n4380), .A2(n7640), .ZN(n7566) );
  NAND2_X1 U9337 ( .A1(n9660), .A2(n7639), .ZN(n7565) );
  OR2_X1 U9338 ( .A1(n9657), .A2(n7632), .ZN(n7564) );
  NAND4_X1 U9339 ( .A1(n7567), .A2(n7566), .A3(n7565), .A4(n7564), .ZN(n7568)
         );
  AOI21_X1 U9340 ( .B1(n7569), .B2(n9650), .A(n7568), .ZN(n7570) );
  INV_X1 U9341 ( .A(n7570), .ZN(P1_U3211) );
  INV_X1 U9342 ( .A(n7571), .ZN(n7608) );
  OAI222_X1 U9343 ( .A1(n10232), .A2(n7608), .B1(P1_U3084), .B2(n4392), .C1(
        n8161), .C2(n8444), .ZN(P1_U3333) );
  INV_X1 U9344 ( .A(n7573), .ZN(n8483) );
  XNOR2_X1 U9345 ( .A(n7572), .B(n8483), .ZN(n7583) );
  INV_X1 U9346 ( .A(n7574), .ZN(n7575) );
  NAND2_X1 U9347 ( .A1(n7594), .A2(n7575), .ZN(n7635) );
  NAND2_X1 U9348 ( .A1(n7635), .A2(n7634), .ZN(n7633) );
  INV_X1 U9349 ( .A(n7576), .ZN(n7577) );
  NAND2_X1 U9350 ( .A1(n7633), .A2(n7577), .ZN(n7578) );
  NAND2_X1 U9351 ( .A1(n7578), .A2(n8483), .ZN(n7580) );
  NAND2_X1 U9352 ( .A1(n7580), .A2(n7579), .ZN(n10185) );
  AOI22_X1 U9353 ( .A1(n10041), .A2(n9671), .B1(n10043), .B2(n9669), .ZN(n7581) );
  OAI21_X1 U9354 ( .B1(n10185), .B2(n10000), .A(n7581), .ZN(n7582) );
  AOI21_X1 U9355 ( .B1(n7583), .B2(n4705), .A(n7582), .ZN(n10184) );
  INV_X1 U9356 ( .A(n7797), .ZN(n7585) );
  AOI21_X1 U9357 ( .B1(n10179), .B2(n7637), .A(n7585), .ZN(n10182) );
  AOI22_X1 U9358 ( .A1(n10062), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7652), .B2(
        n10051), .ZN(n7586) );
  OAI21_X1 U9359 ( .B1(n10054), .B2(n5726), .A(n7586), .ZN(n7588) );
  NOR2_X1 U9360 ( .A1(n10185), .A2(n10057), .ZN(n7587) );
  AOI211_X1 U9361 ( .C1(n10182), .C2(n10060), .A(n7588), .B(n7587), .ZN(n7589)
         );
  OAI21_X1 U9362 ( .B1(n10062), .B2(n10184), .A(n7589), .ZN(P1_U3283) );
  INV_X1 U9363 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9364 ( .A1(n7591), .A2(n7590), .ZN(n7593) );
  INV_X1 U9365 ( .A(n8479), .ZN(n7592) );
  NAND2_X1 U9366 ( .A1(n7593), .A2(n7592), .ZN(n7595) );
  NAND2_X1 U9367 ( .A1(n7595), .A2(n7594), .ZN(n7764) );
  OAI21_X1 U9368 ( .B1(n7596), .B2(n7597), .A(n7636), .ZN(n7760) );
  OAI22_X1 U9369 ( .A1(n7760), .A2(n10287), .B1(n7597), .B2(n10295), .ZN(n7601) );
  XNOR2_X1 U9370 ( .A(n8605), .B(n8479), .ZN(n7600) );
  NAND2_X1 U9371 ( .A1(n7764), .A2(n10048), .ZN(n7599) );
  AOI22_X1 U9372 ( .A1(n10043), .A2(n9671), .B1(n10041), .B2(n9673), .ZN(n7598) );
  OAI211_X1 U9373 ( .C1(n7600), .C2(n10045), .A(n7599), .B(n7598), .ZN(n7761)
         );
  AOI211_X1 U9374 ( .C1(n10292), .C2(n7764), .A(n7601), .B(n7761), .ZN(n7604)
         );
  OR2_X1 U9375 ( .A1(n7604), .A2(n10306), .ZN(n7602) );
  OAI21_X1 U9376 ( .B1(n10308), .B2(n7603), .A(n7602), .ZN(P1_U3529) );
  INV_X1 U9377 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7606) );
  OR2_X1 U9378 ( .A1(n7604), .A2(n10299), .ZN(n7605) );
  OAI21_X1 U9379 ( .B1(n10301), .B2(n7606), .A(n7605), .ZN(P1_U3472) );
  OAI222_X1 U9380 ( .A1(n6173), .A2(P2_U3152), .B1(n9511), .B2(n7608), .C1(
        n7607), .C2(n9508), .ZN(P2_U3338) );
  AOI21_X1 U9381 ( .B1(n7611), .B2(n7610), .A(n7609), .ZN(n7615) );
  AOI22_X1 U9382 ( .A1(n8903), .A2(n8925), .B1(n8902), .B2(n7914), .ZN(n7612)
         );
  NAND2_X1 U9383 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n9024) );
  OAI211_X1 U9384 ( .C1(n7831), .C2(n8906), .A(n7612), .B(n9024), .ZN(n7613)
         );
  AOI21_X1 U9385 ( .B1(n8908), .B2(n7915), .A(n7613), .ZN(n7614) );
  OAI21_X1 U9386 ( .B1(n7615), .B2(n8910), .A(n7614), .ZN(P2_U3233) );
  XNOR2_X1 U9387 ( .A(n7616), .B(n7617), .ZN(n7866) );
  NAND2_X1 U9388 ( .A1(n7692), .A2(n7618), .ZN(n7619) );
  XNOR2_X1 U9389 ( .A(n7868), .B(n7619), .ZN(n7620) );
  AOI222_X1 U9390 ( .A1(n10313), .A2(n7620), .B1(n8925), .B2(n10316), .C1(
        n8927), .C2(n10317), .ZN(n7857) );
  INV_X1 U9391 ( .A(n7621), .ZN(n7696) );
  AOI21_X1 U9392 ( .B1(n7622), .B2(n7696), .A(n7882), .ZN(n7863) );
  AOI22_X1 U9393 ( .A1(n7863), .A2(n10398), .B1(n7622), .B2(n10396), .ZN(n7623) );
  OAI211_X1 U9394 ( .C1(n9475), .C2(n7866), .A(n7857), .B(n7623), .ZN(n7625)
         );
  NAND2_X1 U9395 ( .A1(n7625), .A2(n10423), .ZN(n7624) );
  OAI21_X1 U9396 ( .B1(n10423), .B2(n8091), .A(n7624), .ZN(P2_U3527) );
  INV_X1 U9397 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7627) );
  NAND2_X1 U9398 ( .A1(n7625), .A2(n10407), .ZN(n7626) );
  OAI21_X1 U9399 ( .B1(n10407), .B2(n7627), .A(n7626), .ZN(P2_U3472) );
  INV_X1 U9400 ( .A(n7628), .ZN(n7629) );
  AOI21_X1 U9401 ( .B1(n7634), .B2(n7630), .A(n7629), .ZN(n7631) );
  OAI222_X1 U9402 ( .A1(n10017), .A2(n7849), .B1(n10014), .B2(n7632), .C1(
        n10045), .C2(n7631), .ZN(n10296) );
  INV_X1 U9403 ( .A(n10296), .ZN(n7645) );
  OAI21_X1 U9404 ( .B1(n7635), .B2(n7634), .A(n7633), .ZN(n10298) );
  INV_X1 U9405 ( .A(n10028), .ZN(n9925) );
  INV_X1 U9406 ( .A(n7636), .ZN(n7638) );
  OAI211_X1 U9407 ( .C1(n7638), .C2(n5026), .A(n10181), .B(n7637), .ZN(n10294)
         );
  AOI22_X1 U9408 ( .A1(n10062), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7639), .B2(
        n10051), .ZN(n7642) );
  NAND2_X1 U9409 ( .A1(n9920), .A2(n7640), .ZN(n7641) );
  OAI211_X1 U9410 ( .C1(n10294), .C2(n9903), .A(n7642), .B(n7641), .ZN(n7643)
         );
  AOI21_X1 U9411 ( .B1(n10298), .B2(n9925), .A(n7643), .ZN(n7644) );
  OAI21_X1 U9412 ( .B1(n7645), .B2(n10062), .A(n7644), .ZN(P1_U3284) );
  XNOR2_X1 U9413 ( .A(n7841), .B(n7843), .ZN(n7647) );
  XNOR2_X1 U9414 ( .A(n7646), .B(n7647), .ZN(n7655) );
  NOR2_X1 U9415 ( .A1(n9654), .A2(n7946), .ZN(n7651) );
  OAI21_X1 U9416 ( .B1(n9657), .B2(n7649), .A(n7648), .ZN(n7650) );
  AOI211_X1 U9417 ( .C1(n7652), .C2(n9660), .A(n7651), .B(n7650), .ZN(n7654)
         );
  NAND2_X1 U9418 ( .A1(n4380), .A2(n10179), .ZN(n7653) );
  OAI211_X1 U9419 ( .C1(n7655), .C2(n9636), .A(n7654), .B(n7653), .ZN(P1_U3219) );
  NOR2_X2 U9420 ( .A1(n7657), .A2(n7656), .ZN(n10332) );
  NOR2_X1 U9421 ( .A1(n9300), .A2(n10332), .ZN(n7756) );
  INV_X1 U9422 ( .A(n7659), .ZN(n10354) );
  AOI22_X1 U9423 ( .A1(n10354), .A2(n10313), .B1(n10316), .B2(n7313), .ZN(
        n10356) );
  OAI22_X1 U9424 ( .A1(n10337), .A2(n10356), .B1(n7658), .B2(n9359), .ZN(n7661) );
  NOR2_X1 U9425 ( .A1(n9366), .A2(n7659), .ZN(n7660) );
  AOI211_X1 U9426 ( .C1(n10337), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7661), .B(
        n7660), .ZN(n7662) );
  OAI21_X1 U9427 ( .B1(n7756), .B2(n7663), .A(n7662), .ZN(P2_U3296) );
  XOR2_X1 U9428 ( .A(n7665), .B(n7664), .Z(n7674) );
  NAND2_X1 U9429 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8303) );
  OAI21_X1 U9430 ( .B1(n9741), .B2(n7666), .A(n8303), .ZN(n7672) );
  OAI211_X1 U9431 ( .C1(n7669), .C2(n7668), .A(n7667), .B(n9695), .ZN(n7670)
         );
  INV_X1 U9432 ( .A(n7670), .ZN(n7671) );
  AOI211_X1 U9433 ( .C1(n9733), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7672), .B(
        n7671), .ZN(n7673) );
  OAI21_X1 U9434 ( .B1(n9745), .B2(n7674), .A(n7673), .ZN(P1_U3254) );
  NAND2_X1 U9435 ( .A1(n7676), .A2(n7675), .ZN(n7677) );
  XOR2_X1 U9436 ( .A(n7681), .B(n7677), .Z(n10375) );
  NAND2_X1 U9437 ( .A1(n7678), .A2(n7679), .ZN(n7680) );
  XOR2_X1 U9438 ( .A(n7681), .B(n7680), .Z(n7682) );
  AOI222_X1 U9439 ( .A1(n10313), .A2(n7682), .B1(n8928), .B2(n10316), .C1(
        n8930), .C2(n10317), .ZN(n10377) );
  MUX2_X1 U9440 ( .A(n7281), .B(n10377), .S(n10335), .Z(n7690) );
  INV_X1 U9441 ( .A(n10332), .ZN(n9194) );
  OR2_X1 U9442 ( .A1(n7683), .A2(n6497), .ZN(n7684) );
  NAND2_X1 U9443 ( .A1(n7723), .A2(n7684), .ZN(n10376) );
  INV_X1 U9444 ( .A(n7685), .ZN(n7686) );
  OAI22_X1 U9445 ( .A1(n9194), .A2(n10376), .B1(n7686), .B2(n9359), .ZN(n7687)
         );
  AOI21_X1 U9446 ( .B1(n9300), .B2(n7688), .A(n7687), .ZN(n7689) );
  OAI211_X1 U9447 ( .C1(n10375), .C2(n9366), .A(n7690), .B(n7689), .ZN(
        P2_U3292) );
  XNOR2_X1 U9448 ( .A(n7691), .B(n7694), .ZN(n10394) );
  INV_X1 U9449 ( .A(n10394), .ZN(n7704) );
  OAI21_X1 U9450 ( .B1(n7694), .B2(n7693), .A(n7692), .ZN(n7695) );
  AOI222_X1 U9451 ( .A1(n10313), .A2(n7695), .B1(n8926), .B2(n10316), .C1(
        n8928), .C2(n10317), .ZN(n10389) );
  MUX2_X1 U9452 ( .A(n7284), .B(n10389), .S(n10335), .Z(n7703) );
  INV_X1 U9453 ( .A(n7724), .ZN(n7697) );
  OAI211_X1 U9454 ( .C1(n10391), .C2(n7697), .A(n7696), .B(n10398), .ZN(n10388) );
  INV_X1 U9455 ( .A(n7698), .ZN(n7699) );
  OAI22_X1 U9456 ( .A1(n10388), .A2(n7714), .B1(n7699), .B2(n9359), .ZN(n7700)
         );
  AOI21_X1 U9457 ( .B1(n9300), .B2(n7701), .A(n7700), .ZN(n7702) );
  OAI211_X1 U9458 ( .C1(n9366), .C2(n7704), .A(n7703), .B(n7702), .ZN(P2_U3290) );
  INV_X1 U9459 ( .A(n7705), .ZN(n7706) );
  AOI21_X1 U9460 ( .B1(n6440), .B2(n7707), .A(n7706), .ZN(n7708) );
  OAI222_X1 U9461 ( .A1(n9312), .A2(n5808), .B1(n6215), .B2(n7709), .C1(n9351), 
        .C2(n7708), .ZN(n10366) );
  NOR2_X1 U9462 ( .A1(n10335), .A2(n7710), .ZN(n7716) );
  NAND2_X1 U9463 ( .A1(n7741), .A2(n10398), .ZN(n7744) );
  INV_X1 U9464 ( .A(n7744), .ZN(n7712) );
  NAND2_X1 U9465 ( .A1(n7720), .A2(n10329), .ZN(n7711) );
  NAND2_X1 U9466 ( .A1(n7712), .A2(n7711), .ZN(n10364) );
  OAI22_X1 U9467 ( .A1(n7714), .A2(n10364), .B1(n7713), .B2(n9359), .ZN(n7715)
         );
  AOI211_X1 U9468 ( .C1(n10366), .C2(n10335), .A(n7716), .B(n7715), .ZN(n7722)
         );
  NAND2_X1 U9469 ( .A1(n7718), .A2(n7717), .ZN(n7719) );
  XNOR2_X1 U9470 ( .A(n6440), .B(n7719), .ZN(n10368) );
  AOI22_X1 U9471 ( .A1(n9196), .A2(n10368), .B1(n9300), .B2(n7720), .ZN(n7721)
         );
  NAND2_X1 U9472 ( .A1(n7722), .A2(n7721), .ZN(P2_U3294) );
  INV_X1 U9473 ( .A(n7723), .ZN(n7725) );
  OAI211_X1 U9474 ( .C1(n7725), .C2(n10383), .A(n10398), .B(n7724), .ZN(n10382) );
  NOR2_X1 U9475 ( .A1(n10382), .A2(n6278), .ZN(n7732) );
  INV_X1 U9476 ( .A(n7727), .ZN(n7728) );
  AOI21_X1 U9477 ( .B1(n7726), .B2(n7737), .A(n7728), .ZN(n7729) );
  OAI222_X1 U9478 ( .A1(n6215), .A2(n7731), .B1(n9312), .B2(n7730), .C1(n9351), 
        .C2(n7729), .ZN(n10384) );
  AOI211_X1 U9479 ( .C1(n10330), .C2(n7733), .A(n7732), .B(n10384), .ZN(n7734)
         );
  MUX2_X1 U9480 ( .A(n7735), .B(n7734), .S(n10335), .Z(n7740) );
  XNOR2_X1 U9481 ( .A(n7736), .B(n7737), .ZN(n10386) );
  AOI22_X1 U9482 ( .A1(n10386), .A2(n9196), .B1(n9300), .B2(n7738), .ZN(n7739)
         );
  NAND2_X1 U9483 ( .A1(n7740), .A2(n7739), .ZN(P2_U3291) );
  OAI21_X1 U9484 ( .B1(n7741), .B2(n6279), .A(n10390), .ZN(n7742) );
  INV_X1 U9485 ( .A(n7742), .ZN(n7743) );
  MUX2_X1 U9486 ( .A(n7744), .B(n7743), .S(n5807), .Z(n10370) );
  NAND3_X1 U9487 ( .A1(n7705), .A2(n4729), .A3(n7746), .ZN(n7747) );
  NAND2_X1 U9488 ( .A1(n7678), .A2(n7747), .ZN(n7748) );
  AOI222_X1 U9489 ( .A1(n10313), .A2(n7748), .B1(n8929), .B2(n10316), .C1(
        n10315), .C2(n10317), .ZN(n10371) );
  MUX2_X1 U9490 ( .A(n7749), .B(n10371), .S(n10335), .Z(n7755) );
  AND2_X1 U9491 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  XNOR2_X1 U9492 ( .A(n7752), .B(n4729), .ZN(n10373) );
  AOI22_X1 U9493 ( .A1(n10373), .A2(n9196), .B1(n10330), .B2(n7753), .ZN(n7754) );
  OAI211_X1 U9494 ( .C1(n7756), .C2(n10370), .A(n7755), .B(n7754), .ZN(
        P2_U3293) );
  AOI22_X1 U9495 ( .A1(n9920), .A2(n7758), .B1(n10051), .B2(n7757), .ZN(n7759)
         );
  OAI21_X1 U9496 ( .B1(n9923), .B2(n7760), .A(n7759), .ZN(n7763) );
  MUX2_X1 U9497 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7761), .S(n9940), .Z(n7762)
         );
  AOI211_X1 U9498 ( .C1(n8406), .C2(n7764), .A(n7763), .B(n7762), .ZN(n7765)
         );
  INV_X1 U9499 ( .A(n7765), .ZN(P1_U3285) );
  INV_X1 U9500 ( .A(n7766), .ZN(n7769) );
  OAI222_X1 U9501 ( .A1(n10232), .A2(n7769), .B1(P1_U3084), .B2(n8561), .C1(
        n7767), .C2(n8444), .ZN(P1_U3332) );
  OAI222_X1 U9502 ( .A1(n9508), .A2(n7770), .B1(n9511), .B2(n7769), .C1(n7768), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  XOR2_X1 U9503 ( .A(n7772), .B(n7771), .Z(n7780) );
  NAND2_X1 U9504 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8426) );
  OAI21_X1 U9505 ( .B1(n9741), .B2(n7773), .A(n8426), .ZN(n7778) );
  XOR2_X1 U9506 ( .A(n7775), .B(n7774), .Z(n7776) );
  NOR2_X1 U9507 ( .A1(n7776), .A2(n9745), .ZN(n7777) );
  AOI211_X1 U9508 ( .C1(n9733), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7778), .B(
        n7777), .ZN(n7779) );
  OAI21_X1 U9509 ( .B1(n9746), .B2(n7780), .A(n7779), .ZN(P1_U3255) );
  OAI211_X1 U9510 ( .C1(n7783), .C2(n7782), .A(n7781), .B(n8888), .ZN(n7788)
         );
  OAI22_X1 U9511 ( .A1(n8906), .A2(n8785), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7784), .ZN(n7786) );
  OAI22_X1 U9512 ( .A1(n8863), .A2(n7877), .B1(n8862), .B2(n8230), .ZN(n7785)
         );
  AOI211_X1 U9513 ( .C1(n8908), .C2(n8229), .A(n7786), .B(n7785), .ZN(n7787)
         );
  NAND2_X1 U9514 ( .A1(n7788), .A2(n7787), .ZN(P2_U3219) );
  NAND2_X1 U9515 ( .A1(n7789), .A2(n8612), .ZN(n7790) );
  XOR2_X1 U9516 ( .A(n7790), .B(n8484), .Z(n7795) );
  INV_X1 U9517 ( .A(n8484), .ZN(n7791) );
  XNOR2_X1 U9518 ( .A(n7792), .B(n7791), .ZN(n10178) );
  AOI22_X1 U9519 ( .A1(n10041), .A2(n9670), .B1(n10043), .B2(n9668), .ZN(n7793) );
  OAI21_X1 U9520 ( .B1(n10178), .B2(n10000), .A(n7793), .ZN(n7794) );
  AOI21_X1 U9521 ( .B1(n7795), .B2(n4705), .A(n7794), .ZN(n10177) );
  AOI21_X1 U9522 ( .B1(n10174), .B2(n7797), .A(n7796), .ZN(n10175) );
  INV_X1 U9523 ( .A(n10174), .ZN(n7799) );
  AOI22_X1 U9524 ( .A1(n10062), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7853), .B2(
        n10051), .ZN(n7798) );
  OAI21_X1 U9525 ( .B1(n7799), .B2(n10054), .A(n7798), .ZN(n7801) );
  NOR2_X1 U9526 ( .A1(n10178), .A2(n10057), .ZN(n7800) );
  AOI211_X1 U9527 ( .C1(n10175), .C2(n10060), .A(n7801), .B(n7800), .ZN(n7802)
         );
  OAI21_X1 U9528 ( .B1(n10177), .B2(n10062), .A(n7802), .ZN(P1_U3282) );
  AOI21_X1 U9529 ( .B1(n9361), .B2(n7804), .A(n7803), .ZN(n7805) );
  INV_X1 U9530 ( .A(n7805), .ZN(n7808) );
  INV_X1 U9531 ( .A(n8254), .ZN(n7806) );
  OAI21_X1 U9532 ( .B1(n7808), .B2(n7807), .A(n7806), .ZN(n7809) );
  NOR2_X1 U9533 ( .A1(n7809), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8253) );
  AOI21_X1 U9534 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7809), .A(n8253), .ZN(
        n7820) );
  INV_X1 U9535 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7810) );
  NAND2_X1 U9536 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8904) );
  OAI21_X1 U9537 ( .B1(n9097), .B2(n7810), .A(n8904), .ZN(n7811) );
  AOI21_X1 U9538 ( .B1(n9077), .B2(n8259), .A(n7811), .ZN(n7819) );
  NOR2_X1 U9539 ( .A1(n7812), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7813) );
  AOI21_X1 U9540 ( .B1(n7815), .B2(n7814), .A(n7813), .ZN(n8260) );
  XOR2_X1 U9541 ( .A(n8259), .B(n8260), .Z(n7817) );
  AND2_X1 U9542 ( .A1(n7817), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8258) );
  INV_X1 U9543 ( .A(n8258), .ZN(n7816) );
  OAI211_X1 U9544 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n7817), .A(n7816), .B(
        n9088), .ZN(n7818) );
  OAI211_X1 U9545 ( .C1(n7820), .C2(n9094), .A(n7819), .B(n7818), .ZN(P2_U3260) );
  INV_X1 U9546 ( .A(n10402), .ZN(n7838) );
  NAND2_X1 U9547 ( .A1(n7823), .A2(n7829), .ZN(n7824) );
  NAND2_X1 U9548 ( .A1(n7822), .A2(n7824), .ZN(n7921) );
  NAND2_X1 U9549 ( .A1(n7826), .A2(n7915), .ZN(n7827) );
  NAND2_X1 U9550 ( .A1(n7934), .A2(n7827), .ZN(n7917) );
  OAI22_X1 U9551 ( .A1(n7917), .A2(n6279), .B1(n7828), .B2(n10390), .ZN(n7837)
         );
  XNOR2_X1 U9552 ( .A(n7830), .B(n5907), .ZN(n7836) );
  INV_X1 U9553 ( .A(n9318), .ZN(n7880) );
  NAND2_X1 U9554 ( .A1(n7921), .A2(n7880), .ZN(n7835) );
  OAI22_X1 U9555 ( .A1(n7832), .A2(n6215), .B1(n7831), .B2(n9312), .ZN(n7833)
         );
  INV_X1 U9556 ( .A(n7833), .ZN(n7834) );
  OAI211_X1 U9557 ( .C1(n9351), .C2(n7836), .A(n7835), .B(n7834), .ZN(n7918)
         );
  AOI211_X1 U9558 ( .C1(n7838), .C2(n7921), .A(n7837), .B(n7918), .ZN(n7890)
         );
  NAND2_X1 U9559 ( .A1(n10405), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7839) );
  OAI21_X1 U9560 ( .B1(n7890), .B2(n10405), .A(n7839), .ZN(P2_U3478) );
  NOR2_X1 U9561 ( .A1(n7646), .A2(n7840), .ZN(n7844) );
  INV_X1 U9562 ( .A(n7646), .ZN(n7842) );
  OAI22_X1 U9563 ( .A1(n7844), .A2(n7843), .B1(n7842), .B2(n7841), .ZN(n7848)
         );
  XNOR2_X1 U9564 ( .A(n7846), .B(n7845), .ZN(n7847) );
  XNOR2_X1 U9565 ( .A(n7848), .B(n7847), .ZN(n7856) );
  NOR2_X1 U9566 ( .A1(n9657), .A2(n7849), .ZN(n7852) );
  OAI21_X1 U9567 ( .B1(n9654), .B2(n8270), .A(n7850), .ZN(n7851) );
  AOI211_X1 U9568 ( .C1(n7853), .C2(n9660), .A(n7852), .B(n7851), .ZN(n7855)
         );
  NAND2_X1 U9569 ( .A1(n10174), .A2(n4380), .ZN(n7854) );
  OAI211_X1 U9570 ( .C1(n7856), .C2(n9636), .A(n7855), .B(n7854), .ZN(P1_U3229) );
  MUX2_X1 U9571 ( .A(n7858), .B(n7857), .S(n10335), .Z(n7865) );
  INV_X1 U9572 ( .A(n7859), .ZN(n7860) );
  OAI22_X1 U9573 ( .A1(n9356), .A2(n7861), .B1(n9359), .B2(n7860), .ZN(n7862)
         );
  AOI21_X1 U9574 ( .B1(n7863), .B2(n10332), .A(n7862), .ZN(n7864) );
  OAI211_X1 U9575 ( .C1(n9366), .C2(n7866), .A(n7865), .B(n7864), .ZN(P2_U3289) );
  OAI21_X1 U9576 ( .B1(n7616), .B2(n7868), .A(n7867), .ZN(n7869) );
  XNOR2_X1 U9577 ( .A(n7869), .B(n7873), .ZN(n7881) );
  INV_X1 U9578 ( .A(n7881), .ZN(n10403) );
  INV_X1 U9579 ( .A(n7870), .ZN(n7871) );
  NAND2_X1 U9580 ( .A1(n10335), .A2(n7871), .ZN(n9327) );
  NAND2_X1 U9581 ( .A1(n7872), .A2(n7873), .ZN(n7874) );
  AOI21_X1 U9582 ( .B1(n7875), .B2(n7874), .A(n9351), .ZN(n7879) );
  OAI22_X1 U9583 ( .A1(n7877), .A2(n9312), .B1(n7876), .B2(n6215), .ZN(n7878)
         );
  AOI211_X1 U9584 ( .C1(n7881), .C2(n7880), .A(n7879), .B(n7878), .ZN(n10401)
         );
  MUX2_X1 U9585 ( .A(n7286), .B(n10401), .S(n10335), .Z(n7889) );
  INV_X1 U9586 ( .A(n7882), .ZN(n7884) );
  INV_X1 U9587 ( .A(n7826), .ZN(n7883) );
  AOI21_X1 U9588 ( .B1(n10397), .B2(n7884), .A(n7883), .ZN(n10399) );
  OAI22_X1 U9589 ( .A1(n9356), .A2(n7886), .B1(n9359), .B2(n7885), .ZN(n7887)
         );
  AOI21_X1 U9590 ( .B1(n10399), .B2(n10332), .A(n7887), .ZN(n7888) );
  OAI211_X1 U9591 ( .C1(n10403), .C2(n9327), .A(n7889), .B(n7888), .ZN(
        P2_U3288) );
  OR2_X1 U9592 ( .A1(n7890), .A2(n10420), .ZN(n7891) );
  OAI21_X1 U9593 ( .B1(n10423), .B2(n7892), .A(n7891), .ZN(P2_U3529) );
  OAI21_X1 U9594 ( .B1(n7893), .B2(P1_REG2_REG_15__SCAN_IN), .A(n9695), .ZN(
        n7901) );
  NAND2_X1 U9595 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9655) );
  OAI21_X1 U9596 ( .B1(n9741), .B2(n4673), .A(n9655), .ZN(n7899) );
  INV_X1 U9597 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7897) );
  INV_X1 U9598 ( .A(n7894), .ZN(n7896) );
  AOI211_X1 U9599 ( .C1(n7897), .C2(n7896), .A(n9745), .B(n7895), .ZN(n7898)
         );
  AOI211_X1 U9600 ( .C1(n9733), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7899), .B(
        n7898), .ZN(n7900) );
  OAI21_X1 U9601 ( .B1(n7902), .B2(n7901), .A(n7900), .ZN(P1_U3256) );
  NAND2_X1 U9602 ( .A1(n7904), .A2(n7903), .ZN(n7905) );
  XOR2_X1 U9603 ( .A(n7906), .B(n7905), .Z(n7913) );
  NAND2_X1 U9604 ( .A1(n9604), .A2(n9668), .ZN(n7908) );
  OAI211_X1 U9605 ( .C1(n7909), .C2(n9654), .A(n7908), .B(n7907), .ZN(n7910)
         );
  AOI21_X1 U9606 ( .B1(n8278), .B2(n9660), .A(n7910), .ZN(n7912) );
  NAND2_X1 U9607 ( .A1(n8411), .A2(n4380), .ZN(n7911) );
  OAI211_X1 U9608 ( .C1(n7913), .C2(n9636), .A(n7912), .B(n7911), .ZN(P1_U3234) );
  INV_X1 U9609 ( .A(n9327), .ZN(n7922) );
  AOI22_X1 U9610 ( .A1(n9300), .A2(n7915), .B1(n10330), .B2(n7914), .ZN(n7916)
         );
  OAI21_X1 U9611 ( .B1(n7917), .B2(n9194), .A(n7916), .ZN(n7920) );
  MUX2_X1 U9612 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7918), .S(n10335), .Z(n7919)
         );
  AOI211_X1 U9613 ( .C1(n7922), .C2(n7921), .A(n7920), .B(n7919), .ZN(n7923)
         );
  INV_X1 U9614 ( .A(n7923), .ZN(P2_U3287) );
  INV_X1 U9615 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7938) );
  NOR2_X1 U9616 ( .A1(n7925), .A2(n7924), .ZN(n8368) );
  AND2_X1 U9617 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  OR2_X1 U9618 ( .A1(n8368), .A2(n7926), .ZN(n8235) );
  OR2_X1 U9619 ( .A1(n8235), .A2(n9318), .ZN(n7933) );
  AOI21_X1 U9620 ( .B1(n7927), .B2(n5930), .A(n9351), .ZN(n7931) );
  NAND2_X1 U9621 ( .A1(n8924), .A2(n10317), .ZN(n7928) );
  OAI21_X1 U9622 ( .B1(n8785), .B2(n9312), .A(n7928), .ZN(n7929) );
  AOI21_X1 U9623 ( .B1(n7931), .B2(n7930), .A(n7929), .ZN(n7932) );
  NAND2_X1 U9624 ( .A1(n7933), .A2(n7932), .ZN(n8227) );
  NAND2_X1 U9625 ( .A1(n7934), .A2(n8229), .ZN(n7935) );
  AND2_X1 U9626 ( .A1(n8375), .A2(n7935), .ZN(n8232) );
  AOI22_X1 U9627 ( .A1(n8232), .A2(n10398), .B1(n8229), .B2(n10396), .ZN(n7936) );
  OAI21_X1 U9628 ( .B1(n8235), .B2(n10402), .A(n7936), .ZN(n7937) );
  NOR2_X1 U9629 ( .A1(n8227), .A2(n7937), .ZN(n7940) );
  MUX2_X1 U9630 ( .A(n7938), .B(n7940), .S(n10407), .Z(n7939) );
  INV_X1 U9631 ( .A(n7939), .ZN(P2_U3481) );
  MUX2_X1 U9632 ( .A(n7941), .B(n7940), .S(n10423), .Z(n7942) );
  INV_X1 U9633 ( .A(n7942), .ZN(P2_U3530) );
  INV_X1 U9634 ( .A(n4380), .ZN(n9663) );
  XNOR2_X1 U9635 ( .A(n7943), .B(n7944), .ZN(n7945) );
  NAND2_X1 U9636 ( .A1(n7945), .A2(n9650), .ZN(n7952) );
  NOR2_X1 U9637 ( .A1(n9657), .A2(n7946), .ZN(n7950) );
  OAI21_X1 U9638 ( .B1(n9654), .B2(n7948), .A(n7947), .ZN(n7949) );
  AOI211_X1 U9639 ( .C1(n8398), .C2(n9660), .A(n7950), .B(n7949), .ZN(n7951)
         );
  OAI211_X1 U9640 ( .C1(n8286), .C2(n9663), .A(n7952), .B(n7951), .ZN(n8226)
         );
  AOI22_X1 U9641 ( .A1(n8439), .A2(keyinput86), .B1(keyinput104), .B2(n8345), 
        .ZN(n7953) );
  OAI221_X1 U9642 ( .B1(n8439), .B2(keyinput86), .C1(n8345), .C2(keyinput104), 
        .A(n7953), .ZN(n7960) );
  INV_X1 U9643 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7955) );
  AOI22_X1 U9644 ( .A1(n7955), .A2(keyinput64), .B1(n9596), .B2(keyinput18), 
        .ZN(n7954) );
  OAI221_X1 U9645 ( .B1(n7955), .B2(keyinput64), .C1(n9596), .C2(keyinput18), 
        .A(n7954), .ZN(n7959) );
  AOI22_X1 U9646 ( .A1(n5106), .A2(keyinput91), .B1(keyinput37), .B2(n7957), 
        .ZN(n7956) );
  OAI221_X1 U9647 ( .B1(n5106), .B2(keyinput91), .C1(n7957), .C2(keyinput37), 
        .A(n7956), .ZN(n7958) );
  NOR3_X1 U9648 ( .A1(n7960), .A2(n7959), .A3(n7958), .ZN(n7984) );
  INV_X1 U9649 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8192) );
  INV_X1 U9650 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8342) );
  AOI22_X1 U9651 ( .A1(n8192), .A2(keyinput119), .B1(keyinput63), .B2(n8342), 
        .ZN(n7961) );
  OAI221_X1 U9652 ( .B1(n8192), .B2(keyinput119), .C1(n8342), .C2(keyinput63), 
        .A(n7961), .ZN(n7967) );
  AOI22_X1 U9653 ( .A1(n7963), .A2(keyinput95), .B1(keyinput38), .B2(n8178), 
        .ZN(n7962) );
  OAI221_X1 U9654 ( .B1(n7963), .B2(keyinput95), .C1(n8178), .C2(keyinput38), 
        .A(n7962), .ZN(n7966) );
  AOI22_X1 U9655 ( .A1(n8189), .A2(keyinput46), .B1(keyinput127), .B2(n8187), 
        .ZN(n7964) );
  OAI221_X1 U9656 ( .B1(n8189), .B2(keyinput46), .C1(n8187), .C2(keyinput127), 
        .A(n7964), .ZN(n7965) );
  NOR3_X1 U9657 ( .A1(n7967), .A2(n7966), .A3(n7965), .ZN(n7983) );
  INV_X1 U9658 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7969) );
  AOI22_X1 U9659 ( .A1(n8179), .A2(keyinput61), .B1(keyinput125), .B2(n7969), 
        .ZN(n7968) );
  OAI221_X1 U9660 ( .B1(n8179), .B2(keyinput61), .C1(n7969), .C2(keyinput125), 
        .A(n7968), .ZN(n7975) );
  AOI22_X1 U9661 ( .A1(n8150), .A2(keyinput0), .B1(keyinput23), .B2(n10200), 
        .ZN(n7970) );
  OAI221_X1 U9662 ( .B1(n8150), .B2(keyinput0), .C1(n10200), .C2(keyinput23), 
        .A(n7970), .ZN(n7974) );
  INV_X1 U9663 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n7972) );
  INV_X1 U9664 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8203) );
  AOI22_X1 U9665 ( .A1(n7972), .A2(keyinput30), .B1(keyinput11), .B2(n8203), 
        .ZN(n7971) );
  OAI221_X1 U9666 ( .B1(n7972), .B2(keyinput30), .C1(n8203), .C2(keyinput11), 
        .A(n7971), .ZN(n7973) );
  NOR3_X1 U9667 ( .A1(n7975), .A2(n7974), .A3(n7973), .ZN(n7982) );
  AOI22_X1 U9668 ( .A1(n8207), .A2(keyinput12), .B1(keyinput10), .B2(n10409), 
        .ZN(n7976) );
  OAI221_X1 U9669 ( .B1(n8207), .B2(keyinput12), .C1(n10409), .C2(keyinput10), 
        .A(n7976), .ZN(n7980) );
  INV_X1 U9670 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7978) );
  AOI22_X1 U9671 ( .A1(n7978), .A2(keyinput126), .B1(n8346), .B2(keyinput16), 
        .ZN(n7977) );
  OAI221_X1 U9672 ( .B1(n7978), .B2(keyinput126), .C1(n8346), .C2(keyinput16), 
        .A(n7977), .ZN(n7979) );
  NOR2_X1 U9673 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  NAND4_X1 U9674 ( .A1(n7984), .A2(n7983), .A3(n7982), .A4(n7981), .ZN(n8043)
         );
  AOI22_X1 U9675 ( .A1(n8191), .A2(keyinput92), .B1(keyinput1), .B2(P2_U3152), 
        .ZN(n7985) );
  OAI221_X1 U9676 ( .B1(n8191), .B2(keyinput92), .C1(P2_U3152), .C2(keyinput1), 
        .A(n7985), .ZN(n7988) );
  INV_X1 U9677 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8148) );
  AOI22_X1 U9678 ( .A1(n8148), .A2(keyinput28), .B1(n8417), .B2(keyinput35), 
        .ZN(n7986) );
  OAI221_X1 U9679 ( .B1(n8148), .B2(keyinput28), .C1(n8417), .C2(keyinput35), 
        .A(n7986), .ZN(n7987) );
  NOR2_X1 U9680 ( .A1(n7988), .A2(n7987), .ZN(n8020) );
  INV_X1 U9681 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10264) );
  XNOR2_X1 U9682 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput68), .ZN(n7990) );
  XNOR2_X1 U9683 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput106), .ZN(n7989) );
  OAI211_X1 U9684 ( .C1(n10264), .C2(keyinput59), .A(n7990), .B(n7989), .ZN(
        n7996) );
  XNOR2_X1 U9685 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput14), .ZN(n7994) );
  XNOR2_X1 U9686 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput39), .ZN(n7993) );
  XNOR2_X1 U9687 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput49), .ZN(n7992) );
  XNOR2_X1 U9688 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput62), .ZN(n7991) );
  NAND4_X1 U9689 ( .A1(n7994), .A2(n7993), .A3(n7992), .A4(n7991), .ZN(n7995)
         );
  NOR2_X1 U9690 ( .A1(n7996), .A2(n7995), .ZN(n8019) );
  XNOR2_X1 U9691 ( .A(P1_REG3_REG_25__SCAN_IN), .B(keyinput101), .ZN(n8000) );
  XNOR2_X1 U9692 ( .A(P1_REG0_REG_11__SCAN_IN), .B(keyinput50), .ZN(n7999) );
  XNOR2_X1 U9693 ( .A(P1_REG3_REG_10__SCAN_IN), .B(keyinput3), .ZN(n7998) );
  XNOR2_X1 U9694 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput100), .ZN(n7997) );
  NAND4_X1 U9695 ( .A1(n8000), .A2(n7999), .A3(n7998), .A4(n7997), .ZN(n8006)
         );
  XNOR2_X1 U9696 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput54), .ZN(n8004) );
  XNOR2_X1 U9697 ( .A(P1_REG3_REG_14__SCAN_IN), .B(keyinput27), .ZN(n8003) );
  XNOR2_X1 U9698 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput123), .ZN(n8002) );
  XNOR2_X1 U9699 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput32), .ZN(n8001) );
  NAND4_X1 U9700 ( .A1(n8004), .A2(n8003), .A3(n8002), .A4(n8001), .ZN(n8005)
         );
  NOR2_X1 U9701 ( .A1(n8006), .A2(n8005), .ZN(n8018) );
  XNOR2_X1 U9702 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput70), .ZN(n8010) );
  XNOR2_X1 U9703 ( .A(P2_REG1_REG_12__SCAN_IN), .B(keyinput80), .ZN(n8009) );
  XNOR2_X1 U9704 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput121), .ZN(n8008) );
  XNOR2_X1 U9705 ( .A(P2_REG1_REG_28__SCAN_IN), .B(keyinput52), .ZN(n8007) );
  NAND4_X1 U9706 ( .A1(n8010), .A2(n8009), .A3(n8008), .A4(n8007), .ZN(n8016)
         );
  XNOR2_X1 U9707 ( .A(P2_REG1_REG_14__SCAN_IN), .B(keyinput114), .ZN(n8014) );
  XNOR2_X1 U9708 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput6), .ZN(n8013) );
  XNOR2_X1 U9709 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput107), .ZN(n8012) );
  XNOR2_X1 U9710 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput124), .ZN(n8011) );
  NAND4_X1 U9711 ( .A1(n8014), .A2(n8013), .A3(n8012), .A4(n8011), .ZN(n8015)
         );
  NOR2_X1 U9712 ( .A1(n8016), .A2(n8015), .ZN(n8017) );
  NAND4_X1 U9713 ( .A1(n8020), .A2(n8019), .A3(n8018), .A4(n8017), .ZN(n8042)
         );
  AOI22_X1 U9714 ( .A1(n9777), .A2(keyinput56), .B1(n9518), .B2(keyinput115), 
        .ZN(n8021) );
  OAI221_X1 U9715 ( .B1(n9777), .B2(keyinput56), .C1(n9518), .C2(keyinput115), 
        .A(n8021), .ZN(n8030) );
  INV_X1 U9716 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10256) );
  INV_X1 U9717 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9070) );
  AOI22_X1 U9718 ( .A1(n10256), .A2(keyinput87), .B1(keyinput26), .B2(n9070), 
        .ZN(n8022) );
  OAI221_X1 U9719 ( .B1(n10256), .B2(keyinput87), .C1(n9070), .C2(keyinput26), 
        .A(n8022), .ZN(n8029) );
  INV_X1 U9720 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10340) );
  AOI22_X1 U9721 ( .A1(n10340), .A2(keyinput2), .B1(n8024), .B2(keyinput25), 
        .ZN(n8023) );
  OAI221_X1 U9722 ( .B1(n10340), .B2(keyinput2), .C1(n8024), .C2(keyinput25), 
        .A(n8023), .ZN(n8028) );
  INV_X1 U9723 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U9724 ( .A1(n10258), .A2(keyinput34), .B1(keyinput71), .B2(n8026), 
        .ZN(n8025) );
  OAI221_X1 U9725 ( .B1(n10258), .B2(keyinput34), .C1(n8026), .C2(keyinput71), 
        .A(n8025), .ZN(n8027) );
  OR4_X1 U9726 ( .A1(n8030), .A2(n8029), .A3(n8028), .A4(n8027), .ZN(n8040) );
  INV_X1 U9727 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8181) );
  AOI22_X1 U9728 ( .A1(n8032), .A2(keyinput47), .B1(keyinput42), .B2(n8181), 
        .ZN(n8031) );
  OAI221_X1 U9729 ( .B1(n8032), .B2(keyinput47), .C1(n8181), .C2(keyinput42), 
        .A(n8031), .ZN(n8039) );
  INV_X1 U9730 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U9731 ( .A1(n8034), .A2(keyinput122), .B1(keyinput93), .B2(n10460), 
        .ZN(n8033) );
  OAI221_X1 U9732 ( .B1(n8034), .B2(keyinput122), .C1(n10460), .C2(keyinput93), 
        .A(n8033), .ZN(n8038) );
  AOI22_X1 U9733 ( .A1(n6916), .A2(keyinput94), .B1(n8036), .B2(keyinput15), 
        .ZN(n8035) );
  OAI221_X1 U9734 ( .B1(n6916), .B2(keyinput94), .C1(n8036), .C2(keyinput15), 
        .A(n8035), .ZN(n8037) );
  OR4_X1 U9735 ( .A1(n8040), .A2(n8039), .A3(n8038), .A4(n8037), .ZN(n8041) );
  NOR3_X1 U9736 ( .A1(n8043), .A2(n8042), .A3(n8041), .ZN(n8123) );
  INV_X1 U9737 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8182) );
  AOI22_X1 U9738 ( .A1(n8182), .A2(keyinput48), .B1(keyinput77), .B2(n10415), 
        .ZN(n8044) );
  OAI221_X1 U9739 ( .B1(n8182), .B2(keyinput48), .C1(n10415), .C2(keyinput77), 
        .A(n8044), .ZN(n8053) );
  AOI22_X1 U9740 ( .A1(n10304), .A2(keyinput4), .B1(keyinput19), .B2(n10343), 
        .ZN(n8045) );
  OAI221_X1 U9741 ( .B1(n10304), .B2(keyinput4), .C1(n10343), .C2(keyinput19), 
        .A(n8045), .ZN(n8052) );
  INV_X1 U9742 ( .A(P1_RD_REG_SCAN_IN), .ZN(n10236) );
  AOI22_X1 U9743 ( .A1(n10236), .A2(keyinput13), .B1(keyinput96), .B2(n8047), 
        .ZN(n8046) );
  OAI221_X1 U9744 ( .B1(n10236), .B2(keyinput13), .C1(n8047), .C2(keyinput96), 
        .A(n8046), .ZN(n8051) );
  AOI22_X1 U9745 ( .A1(n8049), .A2(keyinput112), .B1(n8211), .B2(keyinput7), 
        .ZN(n8048) );
  OAI221_X1 U9746 ( .B1(n8049), .B2(keyinput112), .C1(n8211), .C2(keyinput7), 
        .A(n8048), .ZN(n8050) );
  NOR4_X1 U9747 ( .A1(n8053), .A2(n8052), .A3(n8051), .A4(n8050), .ZN(n8122)
         );
  INV_X1 U9748 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8055) );
  INV_X1 U9749 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U9750 ( .A1(n8055), .A2(keyinput111), .B1(n10250), .B2(keyinput9), 
        .ZN(n8054) );
  OAI221_X1 U9751 ( .B1(n8055), .B2(keyinput111), .C1(n10250), .C2(keyinput9), 
        .A(n8054), .ZN(n8060) );
  INV_X1 U9752 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U9753 ( .A1(n8057), .A2(keyinput102), .B1(n10263), .B2(keyinput44), 
        .ZN(n8056) );
  OAI221_X1 U9754 ( .B1(n8057), .B2(keyinput102), .C1(n10263), .C2(keyinput44), 
        .A(n8056), .ZN(n8059) );
  INV_X1 U9755 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10272) );
  XNOR2_X1 U9756 ( .A(n10272), .B(keyinput105), .ZN(n8058) );
  NOR3_X1 U9757 ( .A1(n8060), .A2(n8059), .A3(n8058), .ZN(n8076) );
  AOI22_X1 U9758 ( .A1(n8188), .A2(keyinput84), .B1(keyinput113), .B2(n6062), 
        .ZN(n8061) );
  OAI221_X1 U9759 ( .B1(n8188), .B2(keyinput84), .C1(n6062), .C2(keyinput113), 
        .A(n8061), .ZN(n8065) );
  AOI22_X1 U9760 ( .A1(n10342), .A2(keyinput20), .B1(n8063), .B2(keyinput89), 
        .ZN(n8062) );
  OAI221_X1 U9761 ( .B1(n10342), .B2(keyinput20), .C1(n8063), .C2(keyinput89), 
        .A(n8062), .ZN(n8064) );
  NOR2_X1 U9762 ( .A1(n8065), .A2(n8064), .ZN(n8075) );
  INV_X1 U9763 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8067) );
  INV_X1 U9764 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U9765 ( .A1(n8067), .A2(keyinput45), .B1(n10260), .B2(keyinput67), 
        .ZN(n8066) );
  OAI221_X1 U9766 ( .B1(n8067), .B2(keyinput45), .C1(n10260), .C2(keyinput67), 
        .A(n8066), .ZN(n8073) );
  AOI22_X1 U9767 ( .A1(n8163), .A2(keyinput117), .B1(n8069), .B2(keyinput43), 
        .ZN(n8068) );
  OAI221_X1 U9768 ( .B1(n8163), .B2(keyinput117), .C1(n8069), .C2(keyinput43), 
        .A(n8068), .ZN(n8072) );
  INV_X1 U9769 ( .A(SI_11_), .ZN(n8160) );
  AOI22_X1 U9770 ( .A1(n8160), .A2(keyinput60), .B1(n8161), .B2(keyinput120), 
        .ZN(n8070) );
  OAI221_X1 U9771 ( .B1(n8160), .B2(keyinput60), .C1(n8161), .C2(keyinput120), 
        .A(n8070), .ZN(n8071) );
  NOR3_X1 U9772 ( .A1(n8073), .A2(n8072), .A3(n8071), .ZN(n8074) );
  NAND3_X1 U9773 ( .A1(n8076), .A2(n8075), .A3(n8074), .ZN(n8120) );
  XNOR2_X1 U9774 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput97), .ZN(n8080) );
  XNOR2_X1 U9775 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput99), .ZN(n8079) );
  XNOR2_X1 U9776 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput90), .ZN(n8078) );
  XNOR2_X1 U9777 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput76), .ZN(n8077) );
  NAND4_X1 U9778 ( .A1(n8080), .A2(n8079), .A3(n8078), .A4(n8077), .ZN(n8086)
         );
  XNOR2_X1 U9779 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput79), .ZN(n8084) );
  XNOR2_X1 U9780 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput73), .ZN(n8083) );
  XNOR2_X1 U9781 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput74), .ZN(n8082) );
  XNOR2_X1 U9782 ( .A(SI_8_), .B(keyinput66), .ZN(n8081) );
  NAND4_X1 U9783 ( .A1(n8084), .A2(n8083), .A3(n8082), .A4(n8081), .ZN(n8085)
         );
  NOR2_X1 U9784 ( .A1(n8086), .A2(n8085), .ZN(n8100) );
  XNOR2_X1 U9785 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput51), .ZN(n8090) );
  XNOR2_X1 U9786 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput57), .ZN(n8089) );
  XNOR2_X1 U9787 ( .A(SI_6_), .B(keyinput8), .ZN(n8088) );
  XNOR2_X1 U9788 ( .A(keyinput83), .B(P2_REG3_REG_2__SCAN_IN), .ZN(n8087) );
  AND4_X1 U9789 ( .A1(n8090), .A2(n8089), .A3(n8088), .A4(n8087), .ZN(n8099)
         );
  XNOR2_X1 U9790 ( .A(keyinput103), .B(n8091), .ZN(n8093) );
  XNOR2_X1 U9791 ( .A(keyinput75), .B(n10334), .ZN(n8092) );
  NOR2_X1 U9792 ( .A1(n8093), .A2(n8092), .ZN(n8098) );
  INV_X1 U9793 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8149) );
  XNOR2_X1 U9794 ( .A(keyinput78), .B(n8149), .ZN(n8096) );
  INV_X1 U9795 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8094) );
  XNOR2_X1 U9796 ( .A(keyinput53), .B(n8094), .ZN(n8095) );
  NOR2_X1 U9797 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  NAND4_X1 U9798 ( .A1(n8100), .A2(n8099), .A3(n8098), .A4(n8097), .ZN(n8119)
         );
  AOI22_X1 U9799 ( .A1(n10421), .A2(keyinput85), .B1(keyinput58), .B2(n8102), 
        .ZN(n8101) );
  OAI221_X1 U9800 ( .B1(n10421), .B2(keyinput85), .C1(n8102), .C2(keyinput58), 
        .A(n8101), .ZN(n8106) );
  AOI22_X1 U9801 ( .A1(n10344), .A2(keyinput69), .B1(n8104), .B2(keyinput65), 
        .ZN(n8103) );
  OAI221_X1 U9802 ( .B1(n10344), .B2(keyinput69), .C1(n8104), .C2(keyinput65), 
        .A(n8103), .ZN(n8105) );
  NOR2_X1 U9803 ( .A1(n8106), .A2(n8105), .ZN(n8117) );
  XNOR2_X1 U9804 ( .A(keyinput33), .B(n4567), .ZN(n8108) );
  INV_X1 U9805 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8355) );
  XNOR2_X1 U9806 ( .A(keyinput41), .B(n8355), .ZN(n8107) );
  NOR2_X1 U9807 ( .A1(n8108), .A2(n8107), .ZN(n8116) );
  XNOR2_X1 U9808 ( .A(keyinput5), .B(n8109), .ZN(n8111) );
  XNOR2_X1 U9809 ( .A(keyinput22), .B(n5176), .ZN(n8110) );
  NOR2_X1 U9810 ( .A1(n8111), .A2(n8110), .ZN(n8115) );
  AOI22_X1 U9811 ( .A1(n10341), .A2(keyinput24), .B1(n8210), .B2(keyinput55), 
        .ZN(n8112) );
  OAI221_X1 U9812 ( .B1(n10341), .B2(keyinput24), .C1(n8210), .C2(keyinput55), 
        .A(n8112), .ZN(n8113) );
  INV_X1 U9813 ( .A(n8113), .ZN(n8114) );
  NAND4_X1 U9814 ( .A1(n8117), .A2(n8116), .A3(n8115), .A4(n8114), .ZN(n8118)
         );
  NOR3_X1 U9815 ( .A1(n8120), .A2(n8119), .A3(n8118), .ZN(n8121) );
  AND3_X1 U9816 ( .A1(n8123), .A2(n8122), .A3(n8121), .ZN(n8224) );
  INV_X1 U9817 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n8340) );
  INV_X1 U9818 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8125) );
  AOI22_X1 U9819 ( .A1(n8340), .A2(keyinput31), .B1(n8125), .B2(keyinput108), 
        .ZN(n8124) );
  OAI221_X1 U9820 ( .B1(n8340), .B2(keyinput31), .C1(n8125), .C2(keyinput108), 
        .A(n8124), .ZN(n8134) );
  INV_X1 U9821 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8128) );
  INV_X1 U9822 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8127) );
  AOI22_X1 U9823 ( .A1(n8128), .A2(keyinput36), .B1(keyinput82), .B2(n8127), 
        .ZN(n8126) );
  OAI221_X1 U9824 ( .B1(n8128), .B2(keyinput36), .C1(n8127), .C2(keyinput82), 
        .A(n8126), .ZN(n8133) );
  AOI22_X1 U9825 ( .A1(n8180), .A2(keyinput118), .B1(keyinput17), .B2(n8354), 
        .ZN(n8129) );
  OAI221_X1 U9826 ( .B1(n8180), .B2(keyinput118), .C1(n8354), .C2(keyinput17), 
        .A(n8129), .ZN(n8132) );
  INV_X1 U9827 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U9828 ( .A1(n10267), .A2(keyinput116), .B1(keyinput88), .B2(n8341), 
        .ZN(n8130) );
  OAI221_X1 U9829 ( .B1(n10267), .B2(keyinput116), .C1(n8341), .C2(keyinput88), 
        .A(n8130), .ZN(n8131) );
  NOR4_X1 U9830 ( .A1(n8134), .A2(n8133), .A3(n8132), .A4(n8131), .ZN(n8223)
         );
  INV_X1 U9831 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8136) );
  AOI22_X1 U9832 ( .A1(n8137), .A2(keyinput109), .B1(keyinput98), .B2(n8136), 
        .ZN(n8135) );
  OAI221_X1 U9833 ( .B1(n8137), .B2(keyinput109), .C1(n8136), .C2(keyinput98), 
        .A(n8135), .ZN(n8146) );
  AOI22_X1 U9834 ( .A1(n9054), .A2(keyinput40), .B1(n6923), .B2(keyinput110), 
        .ZN(n8138) );
  OAI221_X1 U9835 ( .B1(n9054), .B2(keyinput40), .C1(n6923), .C2(keyinput110), 
        .A(n8138), .ZN(n8145) );
  AOI22_X1 U9836 ( .A1(n8140), .A2(keyinput29), .B1(keyinput21), .B2(n7749), 
        .ZN(n8139) );
  OAI221_X1 U9837 ( .B1(n8140), .B2(keyinput29), .C1(n7749), .C2(keyinput21), 
        .A(n8139), .ZN(n8144) );
  INV_X1 U9838 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8142) );
  INV_X1 U9839 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U9840 ( .A1(n8142), .A2(keyinput81), .B1(n10259), .B2(keyinput72), 
        .ZN(n8141) );
  OAI221_X1 U9841 ( .B1(n8142), .B2(keyinput81), .C1(n10259), .C2(keyinput72), 
        .A(n8141), .ZN(n8143) );
  NOR4_X1 U9842 ( .A1(n8146), .A2(n8145), .A3(n8144), .A4(n8143), .ZN(n8222)
         );
  NAND2_X1 U9843 ( .A1(n8341), .A2(n8340), .ZN(n8356) );
  INV_X1 U9844 ( .A(n8356), .ZN(n10470) );
  NOR2_X1 U9845 ( .A1(P2_STATE_REG_SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n8147) );
  NOR4_X1 U9846 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n8354), .A3(n8346), .A4(
        n10460), .ZN(n8155) );
  NOR4_X1 U9847 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .A3(n8149), .A4(n8148), .ZN(n8154) );
  NOR4_X1 U9848 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .A3(P1_REG3_REG_10__SCAN_IN), .A4(n8150), .ZN(n8151) );
  NAND3_X1 U9849 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .A3(
        n8151), .ZN(n8152) );
  NOR3_X1 U9850 ( .A1(n8152), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P1_IR_REG_20__SCAN_IN), .ZN(n8153) );
  NAND3_X1 U9851 ( .A1(n8155), .A2(n8154), .A3(n8153), .ZN(n8156) );
  NOR4_X1 U9852 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        n8157), .A4(n8156), .ZN(n8158) );
  NAND4_X1 U9853 ( .A1(n8159), .A2(P2_DATAO_REG_26__SCAN_IN), .A3(n10470), 
        .A4(n8158), .ZN(n8176) );
  NAND4_X1 U9854 ( .A1(SI_16_), .A2(P1_REG0_REG_21__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_REG1_REG_17__SCAN_IN), .ZN(n8175) );
  NAND4_X1 U9855 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(n8161), .A3(n8160), .A4(
        n6238), .ZN(n8174) );
  NOR4_X1 U9856 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(P2_REG2_REG_3__SCAN_IN), 
        .A3(P2_REG2_REG_30__SCAN_IN), .A4(n9054), .ZN(n8172) );
  NOR4_X1 U9857 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(P1_REG0_REG_23__SCAN_IN), 
        .A3(P1_REG2_REG_13__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8171) );
  NOR4_X1 U9858 ( .A1(n8162), .A2(P2_DATAO_REG_13__SCAN_IN), .A3(
        P1_REG3_REG_27__SCAN_IN), .A4(P2_IR_REG_0__SCAN_IN), .ZN(n8169) );
  NAND4_X1 U9859 ( .A1(SI_19_), .A2(P2_IR_REG_6__SCAN_IN), .A3(
        P2_DATAO_REG_31__SCAN_IN), .A4(n8163), .ZN(n8167) );
  NAND4_X1 U9860 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_REG1_REG_19__SCAN_IN), 
        .A3(n8165), .A4(n8164), .ZN(n8166) );
  NOR4_X1 U9861 ( .A1(P1_REG2_REG_29__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .A3(n8167), .A4(n8166), .ZN(n8168) );
  AND4_X1 U9862 ( .A1(n8169), .A2(P2_D_REG_19__SCAN_IN), .A3(n8168), .A4(n5748), .ZN(n8170) );
  NAND3_X1 U9863 ( .A1(n8172), .A2(n8171), .A3(n8170), .ZN(n8173) );
  NOR4_X1 U9864 ( .A1(n8176), .A2(n8175), .A3(n8174), .A4(n8173), .ZN(n8219)
         );
  NAND4_X1 U9865 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(SI_31_), .A3(n8178), .A4(
        n8177), .ZN(n8186) );
  NAND4_X1 U9866 ( .A1(SI_20_), .A2(P1_REG2_REG_18__SCAN_IN), .A3(n8179), .A4(
        n8255), .ZN(n8185) );
  NAND4_X1 U9867 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P2_REG0_REG_20__SCAN_IN), 
        .A3(P2_REG0_REG_9__SCAN_IN), .A4(n8180), .ZN(n8184) );
  NAND4_X1 U9868 ( .A1(n8182), .A2(n10343), .A3(n8181), .A4(n10415), .ZN(n8183) );
  NOR4_X1 U9869 ( .A1(n8186), .A2(n8185), .A3(n8184), .A4(n8183), .ZN(n8218)
         );
  NAND4_X1 U9870 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(n8189), .A3(n8188), .A4(
        n8187), .ZN(n8190) );
  NOR3_X1 U9871 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_REG1_REG_7__SCAN_IN), 
        .A3(n8190), .ZN(n8217) );
  NAND4_X1 U9872 ( .A1(P1_REG0_REG_20__SCAN_IN), .A2(P2_REG3_REG_2__SCAN_IN), 
        .A3(P2_REG1_REG_1__SCAN_IN), .A4(n8191), .ZN(n8194) );
  NAND4_X1 U9873 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(n10334), .A3(n9070), .A4(
        n8192), .ZN(n8193) );
  NOR3_X1 U9874 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(n8194), .A3(n8193), .ZN(
        n8196) );
  NOR2_X1 U9875 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n8195) );
  AND4_X1 U9876 ( .A1(n8196), .A2(P1_REG0_REG_9__SCAN_IN), .A3(
        P1_REG2_REG_9__SCAN_IN), .A4(n8195), .ZN(n8209) );
  NAND4_X1 U9877 ( .A1(n8199), .A2(n8198), .A3(n8197), .A4(SI_1_), .ZN(n8202)
         );
  NAND4_X1 U9878 ( .A1(n8200), .A2(P2_DATAO_REG_6__SCAN_IN), .A3(SI_6_), .A4(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8201) );
  NOR2_X1 U9879 ( .A1(n8202), .A2(n8201), .ZN(n8208) );
  NAND4_X1 U9880 ( .A1(n8203), .A2(P1_REG3_REG_12__SCAN_IN), .A3(
        P1_REG2_REG_6__SCAN_IN), .A4(P1_REG1_REG_3__SCAN_IN), .ZN(n8205) );
  NAND4_X1 U9881 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P2_DATAO_REG_5__SCAN_IN), 
        .A3(P2_DATAO_REG_4__SCAN_IN), .A4(P2_DATAO_REG_3__SCAN_IN), .ZN(n8204)
         );
  NOR2_X1 U9882 ( .A1(n8205), .A2(n8204), .ZN(n8206) );
  NAND4_X1 U9883 ( .A1(n8209), .A2(n8208), .A3(n8207), .A4(n8206), .ZN(n8215)
         );
  NAND4_X1 U9884 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_REG1_REG_11__SCAN_IN), 
        .A3(P1_REG0_REG_11__SCAN_IN), .A4(n10260), .ZN(n8214) );
  NAND4_X1 U9885 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), 
        .A3(P2_REG0_REG_27__SCAN_IN), .A4(n8210), .ZN(n8213) );
  NAND4_X1 U9886 ( .A1(n8032), .A2(n8211), .A3(P1_REG2_REG_0__SCAN_IN), .A4(
        P1_REG3_REG_1__SCAN_IN), .ZN(n8212) );
  NOR4_X1 U9887 ( .A1(n8215), .A2(n8214), .A3(n8213), .A4(n8212), .ZN(n8216)
         );
  AND4_X1 U9888 ( .A1(n8219), .A2(n8218), .A3(n8217), .A4(n8216), .ZN(n8220)
         );
  OAI21_X1 U9889 ( .B1(n8220), .B2(keyinput59), .A(n10264), .ZN(n8221) );
  NAND4_X1 U9890 ( .A1(n8224), .A2(n8223), .A3(n8222), .A4(n8221), .ZN(n8225)
         );
  XNOR2_X1 U9891 ( .A(n8226), .B(n8225), .ZN(P1_U3215) );
  MUX2_X1 U9892 ( .A(n8227), .B(P2_REG2_REG_10__SCAN_IN), .S(n10337), .Z(n8228) );
  INV_X1 U9893 ( .A(n8228), .ZN(n8234) );
  OAI22_X1 U9894 ( .A1(n9356), .A2(n6172), .B1(n9359), .B2(n8230), .ZN(n8231)
         );
  AOI21_X1 U9895 ( .B1(n8232), .B2(n10332), .A(n8231), .ZN(n8233) );
  OAI211_X1 U9896 ( .C1(n8235), .C2(n9327), .A(n8234), .B(n8233), .ZN(P2_U3286) );
  INV_X1 U9897 ( .A(n8240), .ZN(n8238) );
  OR2_X1 U9898 ( .A1(n8236), .A2(P1_U3084), .ZN(n8729) );
  NAND2_X1 U9899 ( .A1(n10230), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8237) );
  OAI211_X1 U9900 ( .C1(n8238), .C2(n10232), .A(n8729), .B(n8237), .ZN(
        P1_U3330) );
  NAND2_X1 U9901 ( .A1(n8240), .A2(n8239), .ZN(n8242) );
  OAI211_X1 U9902 ( .C1(n8243), .C2(n9508), .A(n8242), .B(n8241), .ZN(P2_U3335) );
  XOR2_X1 U9903 ( .A(n8245), .B(n8244), .Z(n8251) );
  NAND2_X1 U9904 ( .A1(n9604), .A2(n9667), .ZN(n8247) );
  OAI211_X1 U9905 ( .C1(n10015), .C2(n9654), .A(n8247), .B(n8246), .ZN(n8248)
         );
  AOI21_X1 U9906 ( .B1(n8330), .B2(n9660), .A(n8248), .ZN(n8250) );
  NAND2_X1 U9907 ( .A1(n10170), .A2(n4380), .ZN(n8249) );
  OAI211_X1 U9908 ( .C1(n8251), .C2(n9636), .A(n8250), .B(n8249), .ZN(P1_U3222) );
  INV_X1 U9909 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8252) );
  MUX2_X1 U9910 ( .A(n8252), .B(P2_REG2_REG_16__SCAN_IN), .S(n9061), .Z(n9047)
         );
  XOR2_X1 U9911 ( .A(n9047), .B(n9049), .Z(n8266) );
  NOR2_X1 U9912 ( .A1(n8255), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8816) );
  NOR2_X1 U9913 ( .A1(n9090), .A2(n8256), .ZN(n8257) );
  AOI211_X1 U9914 ( .C1(n9056), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8816), .B(
        n8257), .ZN(n8265) );
  XOR2_X1 U9915 ( .A(n9061), .B(P2_REG1_REG_16__SCAN_IN), .Z(n8262) );
  AOI21_X1 U9916 ( .B1(n8260), .B2(n8259), .A(n8258), .ZN(n8261) );
  NAND2_X1 U9917 ( .A1(n8261), .A2(n8262), .ZN(n9060) );
  OAI21_X1 U9918 ( .B1(n8262), .B2(n8261), .A(n9060), .ZN(n8263) );
  NAND2_X1 U9919 ( .A1(n8263), .A2(n9088), .ZN(n8264) );
  OAI211_X1 U9920 ( .C1(n8266), .C2(n9094), .A(n8265), .B(n8264), .ZN(P2_U3261) );
  OR2_X1 U9921 ( .A1(n8267), .A2(n8486), .ZN(n8268) );
  AND2_X1 U9922 ( .A1(n8324), .A2(n8268), .ZN(n8272) );
  INV_X1 U9923 ( .A(n8272), .ZN(n8414) );
  NAND2_X1 U9924 ( .A1(n10043), .A2(n10040), .ZN(n8269) );
  OAI21_X1 U9925 ( .B1(n8270), .B2(n10014), .A(n8269), .ZN(n8271) );
  AOI21_X1 U9926 ( .B1(n8272), .B2(n10048), .A(n8271), .ZN(n8276) );
  INV_X1 U9927 ( .A(n8486), .ZN(n8637) );
  XNOR2_X1 U9928 ( .A(n8273), .B(n8637), .ZN(n8274) );
  NAND2_X1 U9929 ( .A1(n8274), .A2(n4705), .ZN(n8275) );
  NAND2_X1 U9930 ( .A1(n8276), .A2(n8275), .ZN(n8416) );
  NAND2_X1 U9931 ( .A1(n8416), .A2(n9940), .ZN(n8283) );
  NAND2_X1 U9932 ( .A1(n8285), .A2(n8411), .ZN(n8277) );
  AND2_X1 U9933 ( .A1(n5060), .A2(n8277), .ZN(n8412) );
  INV_X1 U9934 ( .A(n8411), .ZN(n8280) );
  AOI22_X1 U9935 ( .A1(n10062), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8278), .B2(
        n10051), .ZN(n8279) );
  OAI21_X1 U9936 ( .B1(n8280), .B2(n10054), .A(n8279), .ZN(n8281) );
  AOI21_X1 U9937 ( .B1(n8412), .B2(n10060), .A(n8281), .ZN(n8282) );
  OAI211_X1 U9938 ( .C1(n8414), .C2(n10057), .A(n8283), .B(n8282), .ZN(
        P1_U3280) );
  XNOR2_X1 U9939 ( .A(n8284), .B(n8472), .ZN(n8405) );
  OAI211_X1 U9940 ( .C1(n8286), .C2(n7796), .A(n8285), .B(n10181), .ZN(n8401)
         );
  OAI21_X1 U9941 ( .B1(n8286), .B2(n10295), .A(n8401), .ZN(n8295) );
  INV_X1 U9942 ( .A(n8636), .ZN(n8290) );
  NAND2_X1 U9943 ( .A1(n8287), .A2(n8613), .ZN(n8288) );
  NAND2_X1 U9944 ( .A1(n8288), .A2(n8472), .ZN(n8289) );
  OAI211_X1 U9945 ( .C1(n8291), .C2(n8290), .A(n8289), .B(n4705), .ZN(n8294)
         );
  AOI22_X1 U9946 ( .A1(n10041), .A2(n9669), .B1(n10043), .B2(n9667), .ZN(n8293) );
  NAND2_X1 U9947 ( .A1(n8405), .A2(n10048), .ZN(n8292) );
  NAND3_X1 U9948 ( .A1(n8294), .A2(n8293), .A3(n8292), .ZN(n8402) );
  AOI211_X1 U9949 ( .C1(n10292), .C2(n8405), .A(n8295), .B(n8402), .ZN(n8298)
         );
  NAND2_X1 U9950 ( .A1(n10299), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8296) );
  OAI21_X1 U9951 ( .B1(n8298), .B2(n10299), .A(n8296), .ZN(P1_U3484) );
  NAND2_X1 U9952 ( .A1(n10306), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8297) );
  OAI21_X1 U9953 ( .B1(n8298), .B2(n10306), .A(n8297), .ZN(P1_U3533) );
  XNOR2_X1 U9954 ( .A(n8300), .B(n8299), .ZN(n8301) );
  XNOR2_X1 U9955 ( .A(n8302), .B(n8301), .ZN(n8308) );
  NAND2_X1 U9956 ( .A1(n9604), .A2(n10040), .ZN(n8304) );
  OAI211_X1 U9957 ( .C1(n9656), .C2(n9654), .A(n8304), .B(n8303), .ZN(n8306)
         );
  NOR2_X1 U9958 ( .A1(n10055), .A2(n9663), .ZN(n8305) );
  AOI211_X1 U9959 ( .C1(n10052), .C2(n9660), .A(n8306), .B(n8305), .ZN(n8307)
         );
  OAI21_X1 U9960 ( .B1(n8308), .B2(n9636), .A(n8307), .ZN(P1_U3232) );
  NAND2_X1 U9961 ( .A1(n8310), .A2(n8309), .ZN(n8311) );
  XNOR2_X1 U9962 ( .A(n8311), .B(n8316), .ZN(n8312) );
  AOI222_X1 U9963 ( .A1(n10313), .A2(n8312), .B1(n8922), .B2(n10317), .C1(
        n8920), .C2(n10316), .ZN(n9468) );
  INV_X1 U9964 ( .A(n8389), .ZN(n8313) );
  AOI21_X1 U9965 ( .B1(n9465), .B2(n4774), .A(n8313), .ZN(n9466) );
  AOI22_X1 U9966 ( .A1(n10337), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8783), .B2(
        n10330), .ZN(n8314) );
  OAI21_X1 U9967 ( .B1(n8790), .B2(n9356), .A(n8314), .ZN(n8318) );
  XNOR2_X1 U9968 ( .A(n8315), .B(n8316), .ZN(n9469) );
  NOR2_X1 U9969 ( .A1(n9469), .A2(n9366), .ZN(n8317) );
  AOI211_X1 U9970 ( .C1(n9466), .C2(n10332), .A(n8318), .B(n8317), .ZN(n8319)
         );
  OAI21_X1 U9971 ( .B1(n9468), .B2(n10337), .A(n8319), .ZN(P2_U3284) );
  NAND2_X1 U9972 ( .A1(n8321), .A2(n8320), .ZN(n8322) );
  XNOR2_X1 U9973 ( .A(n8322), .B(n8489), .ZN(n8329) );
  NAND2_X1 U9974 ( .A1(n8324), .A2(n8323), .ZN(n8326) );
  NAND2_X1 U9975 ( .A1(n8326), .A2(n8325), .ZN(n10034) );
  OAI21_X1 U9976 ( .B1(n8326), .B2(n8325), .A(n10034), .ZN(n10173) );
  AOI22_X1 U9977 ( .A1(n10041), .A2(n9667), .B1(n10043), .B2(n9666), .ZN(n8327) );
  OAI21_X1 U9978 ( .B1(n10173), .B2(n10000), .A(n8327), .ZN(n8328) );
  AOI21_X1 U9979 ( .B1(n8329), .B2(n4705), .A(n8328), .ZN(n10172) );
  AOI211_X1 U9980 ( .C1(n10170), .C2(n5060), .A(n10287), .B(n10049), .ZN(
        n10169) );
  AOI22_X1 U9981 ( .A1(n10062), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8330), .B2(
        n10051), .ZN(n8331) );
  OAI21_X1 U9982 ( .B1(n5029), .B2(n10054), .A(n8331), .ZN(n8333) );
  NOR2_X1 U9983 ( .A1(n10173), .A2(n10057), .ZN(n8332) );
  AOI211_X1 U9984 ( .C1(n10169), .C2(n10031), .A(n8333), .B(n8332), .ZN(n8334)
         );
  OAI21_X1 U9985 ( .B1(n10062), .B2(n10172), .A(n8334), .ZN(P1_U3279) );
  NOR2_X1 U9986 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8335) );
  AOI21_X1 U9987 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n8335), .ZN(n10431) );
  NOR2_X1 U9988 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8336) );
  AOI21_X1 U9989 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n8336), .ZN(n10434) );
  NOR2_X1 U9990 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8337) );
  AOI21_X1 U9991 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n8337), .ZN(n10437) );
  NOR2_X1 U9992 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8338) );
  AOI21_X1 U9993 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n8338), .ZN(n10440) );
  NOR2_X1 U9994 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8339) );
  AOI21_X1 U9995 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n8339), .ZN(n10443) );
  INV_X1 U9996 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8358) );
  INV_X1 U9997 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10467) );
  NOR2_X1 U9998 ( .A1(n8341), .A2(n8340), .ZN(n10469) );
  NOR2_X1 U9999 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8350) );
  AOI22_X1 U10000 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n7277), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(n8342), .ZN(n10478) );
  NAND2_X1 U10001 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n8348) );
  XNOR2_X1 U10002 ( .A(n8343), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U10003 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .B1(n8346), .B2(n8345), .ZN(n10474) );
  AOI21_X1 U10004 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10424) );
  INV_X1 U10005 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10428) );
  NAND3_X1 U10006 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10426) );
  OAI21_X1 U10007 ( .B1(n10424), .B2(n10428), .A(n10426), .ZN(n10473) );
  NAND2_X1 U10008 ( .A1(n10474), .A2(n10473), .ZN(n8344) );
  OAI21_X1 U10009 ( .B1(n8346), .B2(n8345), .A(n8344), .ZN(n10475) );
  NAND2_X1 U10010 ( .A1(n10476), .A2(n10475), .ZN(n8347) );
  NAND2_X1 U10011 ( .A1(n8348), .A2(n8347), .ZN(n10477) );
  NOR2_X1 U10012 ( .A1(n10478), .A2(n10477), .ZN(n8349) );
  NOR2_X1 U10013 ( .A1(n8350), .A2(n8349), .ZN(n8351) );
  NOR2_X1 U10014 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n8351), .ZN(n10456) );
  AND2_X1 U10015 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n8351), .ZN(n10455) );
  NOR2_X1 U10016 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10455), .ZN(n8352) );
  NOR2_X1 U10017 ( .A1(n10456), .A2(n8352), .ZN(n10454) );
  AOI22_X1 U10018 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .B1(n8355), .B2(n8354), .ZN(n10453) );
  NAND2_X1 U10019 ( .A1(n10454), .A2(n10453), .ZN(n8353) );
  NOR2_X1 U10020 ( .A1(n10467), .A2(n10466), .ZN(n8357) );
  NAND2_X1 U10021 ( .A1(n10467), .A2(n10466), .ZN(n10465) );
  OAI21_X1 U10022 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(n8357), .A(n10465), .ZN(
        n8359) );
  NOR2_X1 U10023 ( .A1(n8358), .A2(n8359), .ZN(n8360) );
  INV_X1 U10024 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10464) );
  XOR2_X1 U10025 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n8359), .Z(n10463) );
  NAND2_X1 U10026 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8361) );
  OAI21_X1 U10027 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n8361), .ZN(n10451) );
  NAND2_X1 U10028 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n8362) );
  OAI21_X1 U10029 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8362), .ZN(n10448) );
  AOI21_X1 U10030 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10447), .ZN(n10446) );
  NOR2_X1 U10031 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8363) );
  AOI21_X1 U10032 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n8363), .ZN(n10445) );
  NAND2_X1 U10033 ( .A1(n10446), .A2(n10445), .ZN(n10444) );
  OAI21_X1 U10034 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10444), .ZN(n10442) );
  NAND2_X1 U10035 ( .A1(n10443), .A2(n10442), .ZN(n10441) );
  OAI21_X1 U10036 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10441), .ZN(n10439) );
  NAND2_X1 U10037 ( .A1(n10440), .A2(n10439), .ZN(n10438) );
  OAI21_X1 U10038 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10438), .ZN(n10436) );
  NAND2_X1 U10039 ( .A1(n10437), .A2(n10436), .ZN(n10435) );
  OAI21_X1 U10040 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10435), .ZN(n10433) );
  NAND2_X1 U10041 ( .A1(n10434), .A2(n10433), .ZN(n10432) );
  OAI21_X1 U10042 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10432), .ZN(n10430) );
  NAND2_X1 U10043 ( .A1(n10431), .A2(n10430), .ZN(n10429) );
  OAI21_X1 U10044 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10429), .ZN(n10459) );
  NOR2_X1 U10045 ( .A1(n10460), .A2(n10459), .ZN(n8364) );
  NAND2_X1 U10046 ( .A1(n10460), .A2(n10459), .ZN(n10458) );
  OAI21_X1 U10047 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n8364), .A(n10458), .ZN(
        n8366) );
  XNOR2_X1 U10048 ( .A(n9751), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n8365) );
  XNOR2_X1 U10049 ( .A(n8366), .B(n8365), .ZN(ADD_1071_U4) );
  NOR2_X1 U10050 ( .A1(n8368), .A2(n8367), .ZN(n8370) );
  XNOR2_X1 U10051 ( .A(n8369), .B(n8370), .ZN(n9474) );
  XNOR2_X1 U10052 ( .A(n8372), .B(n8371), .ZN(n8373) );
  AOI222_X1 U10053 ( .A1(n10313), .A2(n8373), .B1(n8921), .B2(n10316), .C1(
        n8923), .C2(n10317), .ZN(n9473) );
  MUX2_X1 U10054 ( .A(n7332), .B(n9473), .S(n10335), .Z(n8380) );
  AOI21_X1 U10055 ( .B1(n9470), .B2(n8375), .A(n8374), .ZN(n9471) );
  INV_X1 U10056 ( .A(n9470), .ZN(n8377) );
  INV_X1 U10057 ( .A(n8873), .ZN(n8376) );
  OAI22_X1 U10058 ( .A1(n9356), .A2(n8377), .B1(n8376), .B2(n9359), .ZN(n8378)
         );
  AOI21_X1 U10059 ( .B1(n9471), .B2(n10332), .A(n8378), .ZN(n8379) );
  OAI211_X1 U10060 ( .C1(n9474), .C2(n9366), .A(n8380), .B(n8379), .ZN(
        P2_U3285) );
  NAND2_X1 U10061 ( .A1(n8381), .A2(n8382), .ZN(n9332) );
  OAI21_X1 U10062 ( .B1(n8382), .B2(n8381), .A(n9332), .ZN(n8388) );
  NAND2_X1 U10063 ( .A1(n8383), .A2(n8382), .ZN(n8384) );
  NAND2_X1 U10064 ( .A1(n8385), .A2(n8384), .ZN(n9464) );
  AOI22_X1 U10065 ( .A1(n8921), .A2(n10317), .B1(n10316), .B2(n9334), .ZN(
        n8386) );
  OAI21_X1 U10066 ( .B1(n9464), .B2(n9318), .A(n8386), .ZN(n8387) );
  AOI21_X1 U10067 ( .B1(n10313), .B2(n8388), .A(n8387), .ZN(n9463) );
  NAND2_X1 U10068 ( .A1(n8389), .A2(n9460), .ZN(n8390) );
  AND2_X1 U10069 ( .A1(n4397), .A2(n8390), .ZN(n9461) );
  AOI22_X1 U10070 ( .A1(n10337), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8847), 
        .B2(n10330), .ZN(n8391) );
  OAI21_X1 U10071 ( .B1(n4772), .B2(n9356), .A(n8391), .ZN(n8393) );
  NOR2_X1 U10072 ( .A1(n9464), .A2(n9327), .ZN(n8392) );
  AOI211_X1 U10073 ( .C1(n9461), .C2(n10332), .A(n8393), .B(n8392), .ZN(n8394)
         );
  OAI21_X1 U10074 ( .B1(n10337), .B2(n9463), .A(n8394), .ZN(P2_U3283) );
  INV_X1 U10075 ( .A(n8395), .ZN(n8409) );
  OAI222_X1 U10076 ( .A1(n10232), .A2(n8409), .B1(P1_U3084), .B2(n8397), .C1(
        n8396), .C2(n8444), .ZN(P1_U3329) );
  AOI22_X1 U10077 ( .A1(n8399), .A2(n9920), .B1(n10051), .B2(n8398), .ZN(n8400) );
  OAI21_X1 U10078 ( .B1(n8401), .B2(n9903), .A(n8400), .ZN(n8404) );
  MUX2_X1 U10079 ( .A(n8402), .B(P1_REG2_REG_10__SCAN_IN), .S(n10062), .Z(
        n8403) );
  AOI211_X1 U10080 ( .C1(n8406), .C2(n8405), .A(n8404), .B(n8403), .ZN(n8407)
         );
  INV_X1 U10081 ( .A(n8407), .ZN(P1_U3281) );
  OAI222_X1 U10082 ( .A1(n8410), .A2(P2_U3152), .B1(n9511), .B2(n8409), .C1(
        n8408), .C2(n9508), .ZN(P2_U3334) );
  AOI22_X1 U10083 ( .A1(n8412), .A2(n10181), .B1(n10180), .B2(n8411), .ZN(
        n8413) );
  OAI21_X1 U10084 ( .B1(n8414), .B2(n10186), .A(n8413), .ZN(n8415) );
  NOR2_X1 U10085 ( .A1(n8416), .A2(n8415), .ZN(n8419) );
  MUX2_X1 U10086 ( .A(n8417), .B(n8419), .S(n10308), .Z(n8418) );
  INV_X1 U10087 ( .A(n8418), .ZN(P1_U3534) );
  INV_X1 U10088 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8420) );
  MUX2_X1 U10089 ( .A(n8420), .B(n8419), .S(n10301), .Z(n8421) );
  INV_X1 U10090 ( .A(n8421), .ZN(P1_U3487) );
  XNOR2_X1 U10091 ( .A(n8423), .B(n8422), .ZN(n8424) );
  XNOR2_X1 U10092 ( .A(n8425), .B(n8424), .ZN(n8431) );
  OAI21_X1 U10093 ( .B1(n9657), .B2(n10015), .A(n8426), .ZN(n8427) );
  AOI21_X1 U10094 ( .B1(n9632), .B2(n9978), .A(n8427), .ZN(n8428) );
  OAI21_X1 U10095 ( .B1(n9629), .B2(n10022), .A(n8428), .ZN(n8429) );
  AOI21_X1 U10096 ( .B1(n10159), .B2(n4380), .A(n8429), .ZN(n8430) );
  OAI21_X1 U10097 ( .B1(n8431), .B2(n9636), .A(n8430), .ZN(P1_U3213) );
  INV_X1 U10098 ( .A(n8432), .ZN(n8436) );
  OAI222_X1 U10099 ( .A1(n8444), .A2(n8434), .B1(n10232), .B2(n8436), .C1(
        n8433), .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U10100 ( .A1(n9508), .A2(n8437), .B1(n9506), .B2(n8436), .C1(n8435), .C2(P2_U3152), .ZN(P2_U3333) );
  INV_X1 U10101 ( .A(n8438), .ZN(n9510) );
  OAI222_X1 U10102 ( .A1(n10232), .A2(n9510), .B1(P1_U3084), .B2(n8440), .C1(
        n8439), .C2(n8444), .ZN(P1_U3327) );
  INV_X1 U10103 ( .A(n8441), .ZN(n8448) );
  OAI222_X1 U10104 ( .A1(n8444), .A2(n8443), .B1(n10232), .B2(n8448), .C1(
        n8442), .C2(P1_U3084), .ZN(P1_U3331) );
  INV_X1 U10105 ( .A(n8465), .ZN(n10225) );
  OAI222_X1 U10106 ( .A1(n9508), .A2(n8446), .B1(n9506), .B2(n10225), .C1(
        n8445), .C2(P2_U3152), .ZN(P2_U3329) );
  OAI222_X1 U10107 ( .A1(n9508), .A2(n8449), .B1(n9511), .B2(n8448), .C1(n8447), .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U10108 ( .A1(n8451), .A2(n8450), .ZN(n9374) );
  NOR2_X1 U10109 ( .A1(n10337), .A2(n9374), .ZN(n9101) );
  AOI21_X1 U10110 ( .B1(n10337), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9101), .ZN(
        n8453) );
  NAND2_X1 U10111 ( .A1(n9369), .A2(n9300), .ZN(n8452) );
  OAI211_X1 U10112 ( .C1(n9371), .C2(n9194), .A(n8453), .B(n8452), .ZN(
        P2_U3265) );
  NAND2_X1 U10113 ( .A1(n7001), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U10114 ( .A1(n8457), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U10115 ( .A1(n7002), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8458) );
  NAND3_X1 U10116 ( .A1(n8460), .A2(n8459), .A3(n8458), .ZN(n9664) );
  NAND2_X1 U10117 ( .A1(n8731), .A2(n8464), .ZN(n8462) );
  NAND2_X1 U10118 ( .A1(n8466), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8461) );
  NOR2_X1 U10119 ( .A1(n10067), .A2(n9769), .ZN(n8503) );
  INV_X1 U10120 ( .A(n8503), .ZN(n8463) );
  NAND2_X1 U10121 ( .A1(n8708), .A2(n8463), .ZN(n8560) );
  INV_X1 U10122 ( .A(n8720), .ZN(n8500) );
  NAND2_X1 U10123 ( .A1(n8465), .A2(n8464), .ZN(n8468) );
  NAND2_X1 U10124 ( .A1(n8466), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10125 ( .A1(n10077), .A2(n8469), .ZN(n8703) );
  INV_X1 U10126 ( .A(n8470), .ZN(n8697) );
  INV_X1 U10127 ( .A(n8678), .ZN(n8471) );
  INV_X1 U10128 ( .A(n9986), .ZN(n9976) );
  INV_X1 U10129 ( .A(n8472), .ZN(n8488) );
  NAND4_X1 U10130 ( .A1(n8476), .A2(n8475), .A3(n8474), .A4(n8473), .ZN(n8480)
         );
  NOR4_X1 U10131 ( .A1(n8480), .A2(n8479), .A3(n8478), .A4(n8477), .ZN(n8481)
         );
  NAND4_X1 U10132 ( .A1(n8484), .A2(n8483), .A3(n8482), .A4(n8481), .ZN(n8485)
         );
  NOR2_X1 U10133 ( .A1(n8486), .A2(n8485), .ZN(n8487) );
  NAND4_X1 U10134 ( .A1(n5705), .A2(n8489), .A3(n8488), .A4(n8487), .ZN(n8490)
         );
  NOR2_X1 U10135 ( .A1(n8490), .A2(n10026), .ZN(n8491) );
  NAND4_X1 U10136 ( .A1(n9969), .A2(n9976), .A3(n9994), .A4(n8491), .ZN(n8492)
         );
  NOR2_X1 U10137 ( .A1(n9956), .A2(n8492), .ZN(n8493) );
  NAND4_X1 U10138 ( .A1(n9891), .A2(n9913), .A3(n9930), .A4(n8493), .ZN(n8494)
         );
  NOR2_X1 U10139 ( .A1(n9884), .A2(n8494), .ZN(n8496) );
  INV_X1 U10140 ( .A(n9847), .ZN(n8495) );
  OR2_X1 U10141 ( .A1(n9846), .A2(n8495), .ZN(n9870) );
  NAND4_X1 U10142 ( .A1(n9842), .A2(n8685), .A3(n8496), .A4(n9870), .ZN(n8497)
         );
  NOR3_X1 U10143 ( .A1(n9798), .A2(n9821), .A3(n8497), .ZN(n8498) );
  NAND2_X1 U10144 ( .A1(n10067), .A2(n9769), .ZN(n8586) );
  AND4_X1 U10145 ( .A1(n10071), .A2(n8697), .A3(n8498), .A4(n8586), .ZN(n8499)
         );
  NAND2_X1 U10146 ( .A1(n8500), .A2(n8499), .ZN(n8501) );
  NOR2_X1 U10147 ( .A1(n8560), .A2(n8501), .ZN(n8559) );
  NOR2_X1 U10148 ( .A1(n4392), .A2(n9857), .ZN(n8716) );
  INV_X1 U10149 ( .A(n9756), .ZN(n10063) );
  NAND2_X1 U10150 ( .A1(n10063), .A2(n8503), .ZN(n8504) );
  AND2_X1 U10151 ( .A1(n8699), .A2(n8704), .ZN(n8553) );
  INV_X1 U10152 ( .A(n8553), .ZN(n8589) );
  NAND2_X1 U10153 ( .A1(n8675), .A2(n8505), .ZN(n8506) );
  AND2_X1 U10154 ( .A1(n8506), .A2(n8673), .ZN(n8507) );
  NAND2_X1 U10155 ( .A1(n8507), .A2(n8678), .ZN(n8667) );
  INV_X1 U10156 ( .A(n9975), .ZN(n8509) );
  NAND2_X1 U10157 ( .A1(n8532), .A2(n10010), .ZN(n8629) );
  NAND4_X1 U10158 ( .A1(n8627), .A2(n8642), .A3(n5063), .A4(n8607), .ZN(n8508)
         );
  OR3_X1 U10159 ( .A1(n8509), .A2(n8629), .A3(n8508), .ZN(n8510) );
  NOR2_X1 U10160 ( .A1(n8537), .A2(n8510), .ZN(n8511) );
  NAND3_X1 U10161 ( .A1(n8657), .A2(n8603), .A3(n8511), .ZN(n8512) );
  NOR2_X1 U10162 ( .A1(n8667), .A2(n8512), .ZN(n8582) );
  INV_X1 U10163 ( .A(n7410), .ZN(n8515) );
  NAND2_X1 U10164 ( .A1(n8514), .A2(n8513), .ZN(n8573) );
  NOR2_X1 U10165 ( .A1(n8515), .A2(n8573), .ZN(n8525) );
  NAND2_X1 U10166 ( .A1(n8609), .A2(n8604), .ZN(n8522) );
  NOR2_X1 U10167 ( .A1(n8578), .A2(n8516), .ZN(n8517) );
  NOR2_X1 U10168 ( .A1(n8522), .A2(n8517), .ZN(n8577) );
  INV_X1 U10169 ( .A(n8518), .ZN(n8520) );
  OR2_X1 U10170 ( .A1(n8520), .A2(n8519), .ZN(n8569) );
  AOI21_X1 U10171 ( .B1(n8569), .B2(n8521), .A(n4690), .ZN(n8523) );
  AOI21_X1 U10172 ( .B1(n8523), .B2(n8606), .A(n8522), .ZN(n8524) );
  AOI21_X1 U10173 ( .B1(n8525), .B2(n8577), .A(n8524), .ZN(n8546) );
  INV_X1 U10174 ( .A(n8603), .ZN(n8539) );
  INV_X1 U10175 ( .A(n8642), .ZN(n8526) );
  OAI21_X1 U10176 ( .B1(n8526), .B2(n8634), .A(n8636), .ZN(n8530) );
  INV_X1 U10177 ( .A(n8527), .ZN(n8528) );
  NAND2_X1 U10178 ( .A1(n8618), .A2(n8528), .ZN(n8529) );
  NAND2_X1 U10179 ( .A1(n8529), .A2(n8638), .ZN(n8624) );
  AOI21_X1 U10180 ( .B1(n8627), .B2(n8530), .A(n8624), .ZN(n8533) );
  NAND2_X1 U10181 ( .A1(n8619), .A2(n8531), .ZN(n8625) );
  NAND2_X1 U10182 ( .A1(n8625), .A2(n8532), .ZN(n8644) );
  OAI21_X1 U10183 ( .B1(n8533), .B2(n8629), .A(n8644), .ZN(n8536) );
  INV_X1 U10184 ( .A(n8640), .ZN(n8535) );
  INV_X1 U10185 ( .A(n8650), .ZN(n8534) );
  AOI211_X1 U10186 ( .C1(n9975), .C2(n8536), .A(n8535), .B(n8534), .ZN(n8538)
         );
  NOR4_X1 U10187 ( .A1(n4990), .A2(n8539), .A3(n8538), .A4(n8537), .ZN(n8543)
         );
  INV_X1 U10188 ( .A(n8675), .ZN(n8669) );
  NAND2_X1 U10189 ( .A1(n8657), .A2(n8540), .ZN(n8659) );
  INV_X1 U10190 ( .A(n8541), .ZN(n8602) );
  NOR2_X1 U10191 ( .A1(n8659), .A2(n8602), .ZN(n8542) );
  NAND2_X1 U10192 ( .A1(n8671), .A2(n8656), .ZN(n8662) );
  NOR4_X1 U10193 ( .A1(n8543), .A2(n8669), .A3(n8542), .A4(n8662), .ZN(n8545)
         );
  INV_X1 U10194 ( .A(n8544), .ZN(n8676) );
  OAI21_X1 U10195 ( .B1(n8545), .B2(n8667), .A(n8676), .ZN(n8580) );
  AOI21_X1 U10196 ( .B1(n8582), .B2(n8546), .A(n8580), .ZN(n8548) );
  OR2_X1 U10197 ( .A1(n8599), .A2(n8682), .ZN(n8584) );
  NAND2_X1 U10198 ( .A1(n8597), .A2(n8595), .ZN(n8683) );
  AOI21_X1 U10199 ( .B1(n5000), .B2(n8683), .A(n8547), .ZN(n8583) );
  OAI211_X1 U10200 ( .C1(n8548), .C2(n8584), .A(n8583), .B(n8694), .ZN(n8555)
         );
  INV_X1 U10201 ( .A(n8694), .ZN(n8550) );
  OAI211_X1 U10202 ( .C1(n8550), .C2(n8549), .A(n9765), .B(n8695), .ZN(n8552)
         );
  INV_X1 U10203 ( .A(n8703), .ZN(n8551) );
  AOI21_X1 U10204 ( .B1(n8553), .B2(n8552), .A(n8551), .ZN(n8587) );
  INV_X1 U10205 ( .A(n9664), .ZN(n9754) );
  NAND2_X1 U10206 ( .A1(n10067), .A2(n9754), .ZN(n8554) );
  AND2_X1 U10207 ( .A1(n8586), .A2(n8554), .ZN(n8707) );
  OAI211_X1 U10208 ( .C1(n8589), .C2(n8555), .A(n8587), .B(n8707), .ZN(n8556)
         );
  AND3_X1 U10209 ( .A1(n8715), .A2(n9857), .A3(n8556), .ZN(n8557) );
  AOI211_X1 U10210 ( .C1(n8720), .C2(n9857), .A(n8719), .B(n8557), .ZN(n8558)
         );
  INV_X1 U10211 ( .A(n8560), .ZN(n8591) );
  AOI21_X1 U10212 ( .B1(n6650), .B2(n10282), .A(n8561), .ZN(n8567) );
  INV_X1 U10213 ( .A(n8562), .ZN(n8566) );
  INV_X1 U10214 ( .A(n8563), .ZN(n8565) );
  AOI211_X1 U10215 ( .C1(n8567), .C2(n8566), .A(n8565), .B(n8564), .ZN(n8572)
         );
  INV_X1 U10216 ( .A(n8568), .ZN(n8571) );
  INV_X1 U10217 ( .A(n8569), .ZN(n8570) );
  OAI211_X1 U10218 ( .C1(n8572), .C2(n8571), .A(n8570), .B(n8575), .ZN(n8579)
         );
  NAND4_X1 U10219 ( .A1(n8606), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n8576)
         );
  OAI211_X1 U10220 ( .C1(n8579), .C2(n8578), .A(n8577), .B(n8576), .ZN(n8581)
         );
  AOI21_X1 U10221 ( .B1(n8582), .B2(n8581), .A(n8580), .ZN(n8585) );
  INV_X1 U10222 ( .A(n9798), .ZN(n9784) );
  OAI211_X1 U10223 ( .C1(n8585), .C2(n8584), .A(n9784), .B(n8583), .ZN(n8588)
         );
  OAI211_X1 U10224 ( .C1(n8589), .C2(n8588), .A(n8587), .B(n8586), .ZN(n8590)
         );
  AOI21_X1 U10225 ( .B1(n8591), .B2(n8590), .A(n8720), .ZN(n8592) );
  XNOR2_X1 U10226 ( .A(n8592), .B(n9857), .ZN(n8593) );
  NAND2_X1 U10227 ( .A1(n8593), .A2(n4392), .ZN(n8723) );
  INV_X1 U10228 ( .A(n8702), .ZN(n8714) );
  INV_X1 U10229 ( .A(n8594), .ZN(n9828) );
  OAI211_X1 U10230 ( .C1(n9828), .C2(n8595), .A(n9804), .B(n8597), .ZN(n8596)
         );
  INV_X1 U10231 ( .A(n8596), .ZN(n8601) );
  AND2_X1 U10232 ( .A1(n8597), .A2(n8682), .ZN(n8598) );
  NOR2_X1 U10233 ( .A1(n8599), .A2(n8598), .ZN(n8600) );
  MUX2_X1 U10234 ( .A(n8601), .B(n8600), .S(n8702), .Z(n8686) );
  MUX2_X1 U10235 ( .A(n8603), .B(n8602), .S(n8714), .Z(n8654) );
  NAND2_X1 U10236 ( .A1(n8605), .A2(n8604), .ZN(n8608) );
  NAND3_X1 U10237 ( .A1(n8608), .A2(n8607), .A3(n8606), .ZN(n8610) );
  NAND2_X1 U10238 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  INV_X1 U10239 ( .A(n8612), .ZN(n8614) );
  NAND3_X1 U10240 ( .A1(n8616), .A2(n8636), .A3(n8615), .ZN(n8621) );
  AND4_X1 U10241 ( .A1(n8637), .A2(n8618), .A3(n8617), .A4(n8714), .ZN(n8620)
         );
  NAND2_X1 U10242 ( .A1(n8629), .A2(n8619), .ZN(n8623) );
  NAND4_X1 U10243 ( .A1(n8621), .A2(n8620), .A3(n9975), .A4(n8623), .ZN(n8648)
         );
  MUX2_X1 U10244 ( .A(n8640), .B(n9975), .S(n8702), .Z(n8633) );
  OAI211_X1 U10245 ( .C1(n8625), .C2(n8624), .A(n8623), .B(n8622), .ZN(n8632)
         );
  INV_X1 U10246 ( .A(n8638), .ZN(n8626) );
  NOR2_X1 U10247 ( .A1(n8627), .A2(n8626), .ZN(n8628) );
  OR2_X1 U10248 ( .A1(n8629), .A2(n8628), .ZN(n8630) );
  NAND4_X1 U10249 ( .A1(n8644), .A2(n8702), .A3(n8630), .A4(n8640), .ZN(n8631)
         );
  NAND2_X1 U10250 ( .A1(n8635), .A2(n8634), .ZN(n8643) );
  AND4_X1 U10251 ( .A1(n8638), .A2(n8637), .A3(n8702), .A4(n8636), .ZN(n8639)
         );
  NAND2_X1 U10252 ( .A1(n8640), .A2(n8639), .ZN(n8641) );
  AOI21_X1 U10253 ( .B1(n8643), .B2(n8642), .A(n8641), .ZN(n8645) );
  NAND2_X1 U10254 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND3_X1 U10255 ( .A1(n8648), .A2(n8647), .A3(n8646), .ZN(n8652) );
  MUX2_X1 U10256 ( .A(n8650), .B(n8649), .S(n8714), .Z(n8651) );
  NAND3_X1 U10257 ( .A1(n8652), .A2(n9969), .A3(n8651), .ZN(n8653) );
  NAND2_X1 U10258 ( .A1(n8654), .A2(n8653), .ZN(n8661) );
  NAND3_X1 U10259 ( .A1(n8661), .A2(n8656), .A3(n8655), .ZN(n8658) );
  NAND3_X1 U10260 ( .A1(n8658), .A2(n5711), .A3(n8657), .ZN(n8666) );
  INV_X1 U10261 ( .A(n8659), .ZN(n8660) );
  NAND2_X1 U10262 ( .A1(n8661), .A2(n8660), .ZN(n8664) );
  INV_X1 U10263 ( .A(n8662), .ZN(n8663) );
  NAND2_X1 U10264 ( .A1(n8664), .A2(n8663), .ZN(n8665) );
  INV_X1 U10265 ( .A(n8667), .ZN(n8668) );
  OAI21_X1 U10266 ( .B1(n8672), .B2(n8669), .A(n8668), .ZN(n8670) );
  NAND2_X1 U10267 ( .A1(n8670), .A2(n8676), .ZN(n8681) );
  NAND2_X1 U10268 ( .A1(n8674), .A2(n8673), .ZN(n8677) );
  NAND3_X1 U10269 ( .A1(n8677), .A2(n8676), .A3(n8675), .ZN(n8679) );
  NAND2_X1 U10270 ( .A1(n8679), .A2(n8678), .ZN(n8680) );
  NOR2_X1 U10271 ( .A1(n8683), .A2(n8682), .ZN(n8684) );
  MUX2_X1 U10272 ( .A(n8687), .B(n9804), .S(n8702), .Z(n8690) );
  MUX2_X1 U10273 ( .A(n9829), .B(n10094), .S(n8702), .Z(n8691) );
  MUX2_X1 U10274 ( .A(n4568), .B(n9519), .S(n8702), .Z(n8688) );
  OAI21_X1 U10275 ( .B1(n8690), .B2(n8689), .A(n8688), .ZN(n8693) );
  INV_X1 U10276 ( .A(n8691), .ZN(n8692) );
  MUX2_X1 U10277 ( .A(n8695), .B(n8694), .S(n8702), .Z(n8696) );
  OAI211_X1 U10278 ( .C1(n8698), .C2(n9798), .A(n8697), .B(n8696), .ZN(n8701)
         );
  MUX2_X1 U10279 ( .A(n8699), .B(n9765), .S(n8702), .Z(n8700) );
  AND2_X1 U10280 ( .A1(n8701), .A2(n8700), .ZN(n8706) );
  MUX2_X1 U10281 ( .A(n8704), .B(n8703), .S(n8702), .Z(n8705) );
  INV_X1 U10282 ( .A(n8707), .ZN(n8709) );
  NAND2_X1 U10283 ( .A1(n8708), .A2(n8714), .ZN(n8710) );
  INV_X1 U10284 ( .A(n8716), .ZN(n8718) );
  NOR3_X1 U10285 ( .A1(n8720), .A2(n8726), .A3(n8719), .ZN(n8721) );
  NOR4_X1 U10286 ( .A1(n8725), .A2(n10213), .A3(n8724), .A4(n4391), .ZN(n8728)
         );
  OAI21_X1 U10287 ( .B1(n8726), .B2(n8729), .A(P1_B_REG_SCAN_IN), .ZN(n8727)
         );
  OAI22_X1 U10288 ( .A1(n8730), .A2(n8729), .B1(n8728), .B2(n8727), .ZN(
        P1_U3240) );
  INV_X1 U10289 ( .A(n8731), .ZN(n10222) );
  OAI222_X1 U10290 ( .A1(n9508), .A2(n8732), .B1(n9506), .B2(n10222), .C1(
        P2_U3152), .C2(n5778), .ZN(P2_U3328) );
  OAI211_X1 U10291 ( .C1(n8735), .C2(n8734), .A(n8733), .B(n8888), .ZN(n8739)
         );
  AOI22_X1 U10292 ( .A1(n8914), .A2(n8874), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8738) );
  AOI22_X1 U10293 ( .A1(n8916), .A2(n8903), .B1(n9124), .B2(n8902), .ZN(n8737)
         );
  NAND2_X1 U10294 ( .A1(n9389), .A2(n8908), .ZN(n8736) );
  NAND4_X1 U10295 ( .A1(n8739), .A2(n8738), .A3(n8737), .A4(n8736), .ZN(
        P2_U3216) );
  OAI21_X1 U10296 ( .B1(n8741), .B2(n8740), .A(n8804), .ZN(n8742) );
  NAND2_X1 U10297 ( .A1(n8742), .A2(n8888), .ZN(n8750) );
  OR2_X1 U10298 ( .A1(n8743), .A2(n6215), .ZN(n8745) );
  OR2_X1 U10299 ( .A1(n9311), .A2(n9312), .ZN(n8744) );
  NAND2_X1 U10300 ( .A1(n8745), .A2(n8744), .ZN(n9353) );
  INV_X1 U10301 ( .A(n9353), .ZN(n8747) );
  OAI21_X1 U10302 ( .B1(n8797), .B2(n8747), .A(n8746), .ZN(n8748) );
  AOI21_X1 U10303 ( .B1(n9358), .B2(n8902), .A(n8748), .ZN(n8749) );
  OAI211_X1 U10304 ( .C1(n9357), .C2(n8897), .A(n8750), .B(n8749), .ZN(
        P2_U3217) );
  XOR2_X1 U10305 ( .A(n8826), .B(n8827), .Z(n8754) );
  AOI22_X1 U10306 ( .A1(n8874), .A2(n9181), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8752) );
  AOI22_X1 U10307 ( .A1(n8903), .A2(n9224), .B1(n8902), .B2(n9188), .ZN(n8751)
         );
  OAI211_X1 U10308 ( .C1(n9409), .C2(n8897), .A(n8752), .B(n8751), .ZN(n8753)
         );
  AOI21_X1 U10309 ( .B1(n8754), .B2(n8888), .A(n8753), .ZN(n8755) );
  INV_X1 U10310 ( .A(n8755), .ZN(P2_U3218) );
  OAI21_X1 U10311 ( .B1(n8758), .B2(n8757), .A(n8756), .ZN(n8759) );
  NAND2_X1 U10312 ( .A1(n8759), .A2(n8888), .ZN(n8762) );
  INV_X1 U10313 ( .A(n8774), .ZN(n9223) );
  AOI22_X1 U10314 ( .A1(n9223), .A2(n10316), .B1(n10317), .B2(n6015), .ZN(
        n9263) );
  NAND2_X1 U10315 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9096) );
  OAI21_X1 U10316 ( .B1(n8797), .B2(n9263), .A(n9096), .ZN(n8760) );
  AOI21_X1 U10317 ( .B1(n9267), .B2(n8902), .A(n8760), .ZN(n8761) );
  OAI211_X1 U10318 ( .C1(n9270), .C2(n8897), .A(n8762), .B(n8761), .ZN(
        P2_U3221) );
  AOI22_X1 U10319 ( .A1(n8903), .A2(n6293), .B1(n8874), .B2(n10315), .ZN(n8769) );
  AOI22_X1 U10320 ( .A1(n8908), .A2(n6488), .B1(n8892), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n8768) );
  OAI21_X1 U10321 ( .B1(n8765), .B2(n8764), .A(n8763), .ZN(n8766) );
  NAND2_X1 U10322 ( .A1(n8766), .A2(n8888), .ZN(n8767) );
  NAND3_X1 U10323 ( .A1(n8769), .A2(n8768), .A3(n8767), .ZN(P2_U3224) );
  XNOR2_X1 U10324 ( .A(n8771), .B(n8770), .ZN(n8778) );
  OAI22_X1 U10325 ( .A1(n8906), .A2(n8773), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8772), .ZN(n8776) );
  OAI22_X1 U10326 ( .A1(n8863), .A2(n8774), .B1(n8862), .B2(n9216), .ZN(n8775)
         );
  AOI211_X1 U10327 ( .C1(n9420), .C2(n8908), .A(n8776), .B(n8775), .ZN(n8777)
         );
  OAI21_X1 U10328 ( .B1(n8778), .B2(n8910), .A(n8777), .ZN(P2_U3225) );
  OAI21_X1 U10329 ( .B1(n8781), .B2(n8780), .A(n8779), .ZN(n8782) );
  NAND2_X1 U10330 ( .A1(n8782), .A2(n8888), .ZN(n8789) );
  INV_X1 U10331 ( .A(n8783), .ZN(n8784) );
  OAI22_X1 U10332 ( .A1(n8863), .A2(n8785), .B1(n8862), .B2(n8784), .ZN(n8786)
         );
  AOI211_X1 U10333 ( .C1(n8874), .C2(n8920), .A(n8787), .B(n8786), .ZN(n8788)
         );
  OAI211_X1 U10334 ( .C1(n8790), .C2(n8897), .A(n8789), .B(n8788), .ZN(
        P2_U3226) );
  XNOR2_X1 U10335 ( .A(n8792), .B(n8791), .ZN(n8793) );
  XNOR2_X1 U10336 ( .A(n8794), .B(n8793), .ZN(n8802) );
  OR2_X1 U10337 ( .A1(n9114), .A2(n9312), .ZN(n8796) );
  NAND2_X1 U10338 ( .A1(n9181), .A2(n10317), .ZN(n8795) );
  NAND2_X1 U10339 ( .A1(n8796), .A2(n8795), .ZN(n9147) );
  INV_X1 U10340 ( .A(n8797), .ZN(n8798) );
  AOI22_X1 U10341 ( .A1(n9147), .A2(n8798), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8799) );
  OAI21_X1 U10342 ( .B1(n9155), .B2(n8862), .A(n8799), .ZN(n8800) );
  AOI21_X1 U10343 ( .B1(n9400), .B2(n8908), .A(n8800), .ZN(n8801) );
  OAI21_X1 U10344 ( .B1(n8802), .B2(n8910), .A(n8801), .ZN(P2_U3227) );
  AND2_X1 U10345 ( .A1(n8804), .A2(n8803), .ZN(n8806) );
  NAND2_X1 U10346 ( .A1(n8806), .A2(n8805), .ZN(n8899) );
  INV_X1 U10347 ( .A(n8806), .ZN(n8808) );
  NAND2_X1 U10348 ( .A1(n8808), .A2(n8807), .ZN(n8898) );
  INV_X1 U10349 ( .A(n8898), .ZN(n8809) );
  AOI211_X1 U10350 ( .C1(n8900), .C2(n8899), .A(n8810), .B(n8809), .ZN(n8813)
         );
  INV_X1 U10351 ( .A(n8811), .ZN(n8812) );
  OAI21_X1 U10352 ( .B1(n8813), .B2(n8812), .A(n8888), .ZN(n8818) );
  INV_X1 U10353 ( .A(n9324), .ZN(n8814) );
  OAI22_X1 U10354 ( .A1(n8863), .A2(n9311), .B1(n8862), .B2(n8814), .ZN(n8815)
         );
  AOI211_X1 U10355 ( .C1(n8874), .C2(n9280), .A(n8816), .B(n8815), .ZN(n8817)
         );
  OAI211_X1 U10356 ( .C1(n9326), .C2(n8897), .A(n8818), .B(n8817), .ZN(
        P2_U3228) );
  XNOR2_X1 U10357 ( .A(n8820), .B(n8819), .ZN(n8825) );
  OAI22_X1 U10358 ( .A1(n8906), .A2(n9289), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9054), .ZN(n8823) );
  INV_X1 U10359 ( .A(n8821), .ZN(n9297) );
  OAI22_X1 U10360 ( .A1(n8863), .A2(n9290), .B1(n8862), .B2(n9297), .ZN(n8822)
         );
  AOI211_X1 U10361 ( .C1(n9442), .C2(n8908), .A(n8823), .B(n8822), .ZN(n8824)
         );
  OAI21_X1 U10362 ( .B1(n8825), .B2(n8910), .A(n8824), .ZN(P2_U3230) );
  AOI21_X1 U10363 ( .B1(n8827), .B2(n8826), .A(n4448), .ZN(n8831) );
  XNOR2_X1 U10364 ( .A(n8829), .B(n8828), .ZN(n8830) );
  XNOR2_X1 U10365 ( .A(n8831), .B(n8830), .ZN(n8836) );
  OAI22_X1 U10366 ( .A1(n8906), .A2(n9131), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8832), .ZN(n8834) );
  OAI22_X1 U10367 ( .A1(n8863), .A2(n9206), .B1(n8862), .B2(n9169), .ZN(n8833)
         );
  AOI211_X1 U10368 ( .C1(n9404), .C2(n8908), .A(n8834), .B(n8833), .ZN(n8835)
         );
  OAI21_X1 U10369 ( .B1(n8836), .B2(n8910), .A(n8835), .ZN(P2_U3231) );
  XNOR2_X1 U10370 ( .A(n8838), .B(n8837), .ZN(n8844) );
  OAI22_X1 U10371 ( .A1(n8906), .A2(n9248), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8839), .ZN(n8842) );
  INV_X1 U10372 ( .A(n9235), .ZN(n8840) );
  OAI22_X1 U10373 ( .A1(n8863), .A2(n9247), .B1(n8862), .B2(n8840), .ZN(n8841)
         );
  AOI211_X1 U10374 ( .C1(n9425), .C2(n8908), .A(n8842), .B(n8841), .ZN(n8843)
         );
  OAI21_X1 U10375 ( .B1(n8844), .B2(n8910), .A(n8843), .ZN(P2_U3235) );
  XNOR2_X1 U10376 ( .A(n8846), .B(n8845), .ZN(n8853) );
  AOI22_X1 U10377 ( .A1(n8903), .A2(n8921), .B1(n8902), .B2(n8847), .ZN(n8849)
         );
  OAI211_X1 U10378 ( .C1(n8850), .C2(n8906), .A(n8849), .B(n8848), .ZN(n8851)
         );
  AOI21_X1 U10379 ( .B1(n8908), .B2(n9460), .A(n8851), .ZN(n8852) );
  OAI21_X1 U10380 ( .B1(n8853), .B2(n8910), .A(n8852), .ZN(P2_U3236) );
  NAND2_X1 U10381 ( .A1(n8855), .A2(n8854), .ZN(n8859) );
  XNOR2_X1 U10382 ( .A(n8857), .B(n8856), .ZN(n8858) );
  XNOR2_X1 U10383 ( .A(n8859), .B(n8858), .ZN(n8867) );
  OAI22_X1 U10384 ( .A1(n8906), .A2(n9206), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8860), .ZN(n8865) );
  INV_X1 U10385 ( .A(n9202), .ZN(n8861) );
  OAI22_X1 U10386 ( .A1(n8863), .A2(n9248), .B1(n8862), .B2(n8861), .ZN(n8864)
         );
  AOI211_X1 U10387 ( .C1(n9415), .C2(n8908), .A(n8865), .B(n8864), .ZN(n8866)
         );
  OAI21_X1 U10388 ( .B1(n8867), .B2(n8910), .A(n8866), .ZN(P2_U3237) );
  NAND2_X1 U10389 ( .A1(n8869), .A2(n8868), .ZN(n8871) );
  XOR2_X1 U10390 ( .A(n8871), .B(n8870), .Z(n8872) );
  NAND2_X1 U10391 ( .A1(n8872), .A2(n8888), .ZN(n8878) );
  AND2_X1 U10392 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9038) );
  AOI21_X1 U10393 ( .B1(n8903), .B2(n8923), .A(n9038), .ZN(n8877) );
  AOI22_X1 U10394 ( .A1(n8874), .A2(n8921), .B1(n8902), .B2(n8873), .ZN(n8876)
         );
  NAND2_X1 U10395 ( .A1(n9470), .A2(n8908), .ZN(n8875) );
  NAND4_X1 U10396 ( .A1(n8878), .A2(n8877), .A3(n8876), .A4(n8875), .ZN(
        P2_U3238) );
  XNOR2_X1 U10397 ( .A(n8880), .B(n8879), .ZN(n8884) );
  AOI22_X1 U10398 ( .A1(n8903), .A2(n9280), .B1(n8902), .B2(n9275), .ZN(n8881)
         );
  NAND2_X1 U10399 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9074) );
  OAI211_X1 U10400 ( .C1(n9247), .C2(n8906), .A(n8881), .B(n9074), .ZN(n8882)
         );
  AOI21_X1 U10401 ( .B1(n9435), .B2(n8908), .A(n8882), .ZN(n8883) );
  OAI21_X1 U10402 ( .B1(n8884), .B2(n8910), .A(n8883), .ZN(P2_U3240) );
  INV_X1 U10403 ( .A(n9394), .ZN(n9141) );
  NAND2_X1 U10404 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  NAND3_X1 U10405 ( .A1(n8889), .A2(n8888), .A3(n8887), .ZN(n8896) );
  NAND2_X1 U10406 ( .A1(n8890), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8891) );
  OAI211_X1 U10407 ( .C1(P2_REG3_REG_26__SCAN_IN), .C2(P2_STATE_REG_SCAN_IN), 
        .A(n8892), .B(n8891), .ZN(n8893) );
  OAI21_X1 U10408 ( .B1(n9132), .B2(n8906), .A(n8893), .ZN(n8894) );
  AOI21_X1 U10409 ( .B1(n8903), .B2(n9165), .A(n8894), .ZN(n8895) );
  OAI211_X1 U10410 ( .C1(n9141), .C2(n8897), .A(n8896), .B(n8895), .ZN(
        P2_U3242) );
  NAND2_X1 U10411 ( .A1(n8899), .A2(n8898), .ZN(n8901) );
  XNOR2_X1 U10412 ( .A(n8901), .B(n8900), .ZN(n8911) );
  AOI22_X1 U10413 ( .A1(n8903), .A2(n9334), .B1(n8902), .B2(n9339), .ZN(n8905)
         );
  OAI211_X1 U10414 ( .C1(n9290), .C2(n8906), .A(n8905), .B(n8904), .ZN(n8907)
         );
  AOI21_X1 U10415 ( .B1(n9450), .B2(n8908), .A(n8907), .ZN(n8909) );
  OAI21_X1 U10416 ( .B1(n8911), .B2(n8910), .A(n8909), .ZN(P2_U3243) );
  MUX2_X1 U10417 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8912), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10418 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8913), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10419 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8914), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10420 ( .A(n8915), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8917), .Z(
        P2_U3579) );
  MUX2_X1 U10421 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8916), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10422 ( .A(n9165), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8917), .Z(
        P2_U3577) );
  MUX2_X1 U10423 ( .A(n9181), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8917), .Z(
        P2_U3576) );
  MUX2_X1 U10424 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9164), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10425 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9224), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10426 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8918), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10427 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9223), .S(P2_U3966), .Z(
        P2_U3572) );
  INV_X1 U10428 ( .A(n9247), .ZN(n9281) );
  MUX2_X1 U10429 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9281), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10430 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n6015), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10431 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9280), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10432 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9335), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10433 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8919), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10434 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9334), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10435 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8920), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10436 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8921), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10437 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8922), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10438 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8923), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10439 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8924), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10440 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8925), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10441 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8926), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10442 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8927), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10443 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8928), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10444 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8929), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10445 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8930), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10446 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n10315), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10447 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n7313), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U10448 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6293), .S(P2_U3966), .Z(
        P2_U3552) );
  AND2_X1 U10449 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n8935) );
  MUX2_X1 U10450 ( .A(n10334), .B(P2_REG2_REG_1__SCAN_IN), .S(n8931), .Z(n8934) );
  INV_X1 U10451 ( .A(n8932), .ZN(n8933) );
  OAI211_X1 U10452 ( .C1(n8935), .C2(n8934), .A(n9051), .B(n8933), .ZN(n8943)
         );
  AOI22_X1 U10453 ( .A1(n9056), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8942) );
  NAND2_X1 U10454 ( .A1(n9077), .A2(n8936), .ZN(n8941) );
  OAI211_X1 U10455 ( .C1(n8939), .C2(n8938), .A(n9088), .B(n8937), .ZN(n8940)
         );
  NAND4_X1 U10456 ( .A1(n8943), .A2(n8942), .A3(n8941), .A4(n8940), .ZN(
        P2_U3246) );
  MUX2_X1 U10457 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7749), .S(n8944), .Z(n8947)
         );
  INV_X1 U10458 ( .A(n8945), .ZN(n8946) );
  NAND2_X1 U10459 ( .A1(n8947), .A2(n8946), .ZN(n8949) );
  OAI211_X1 U10460 ( .C1(n8950), .C2(n8949), .A(n9051), .B(n8948), .ZN(n8958)
         );
  AOI22_X1 U10461 ( .A1(n9056), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n8957) );
  NAND2_X1 U10462 ( .A1(n9077), .A2(n8951), .ZN(n8956) );
  OAI211_X1 U10463 ( .C1(n8954), .C2(n8953), .A(n9088), .B(n8952), .ZN(n8955)
         );
  NAND4_X1 U10464 ( .A1(n8958), .A2(n8957), .A3(n8956), .A4(n8955), .ZN(
        P2_U3248) );
  INV_X1 U10465 ( .A(n8959), .ZN(n8962) );
  MUX2_X1 U10466 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7735), .S(n8960), .Z(n8961)
         );
  NAND3_X1 U10467 ( .A1(n8963), .A2(n8962), .A3(n8961), .ZN(n8964) );
  NAND3_X1 U10468 ( .A1(n9051), .A2(n8976), .A3(n8964), .ZN(n8973) );
  NAND2_X1 U10469 ( .A1(n9077), .A2(n8965), .ZN(n8972) );
  NOR2_X1 U10470 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5860), .ZN(n8966) );
  AOI21_X1 U10471 ( .B1(n9056), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8966), .ZN(
        n8971) );
  OAI211_X1 U10472 ( .C1(n8969), .C2(n8968), .A(n9088), .B(n8967), .ZN(n8970)
         );
  NAND4_X1 U10473 ( .A1(n8973), .A2(n8972), .A3(n8971), .A4(n8970), .ZN(
        P2_U3250) );
  INV_X1 U10474 ( .A(n8991), .ZN(n8978) );
  NAND3_X1 U10475 ( .A1(n8976), .A2(n8975), .A3(n8974), .ZN(n8977) );
  NAND3_X1 U10476 ( .A1(n9051), .A2(n8978), .A3(n8977), .ZN(n8988) );
  NAND2_X1 U10477 ( .A1(n9077), .A2(n8979), .ZN(n8987) );
  INV_X1 U10478 ( .A(n8980), .ZN(n8981) );
  AOI21_X1 U10479 ( .B1(n9056), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8981), .ZN(
        n8986) );
  OAI211_X1 U10480 ( .C1(n8984), .C2(n8983), .A(n9088), .B(n8982), .ZN(n8985)
         );
  NAND4_X1 U10481 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(
        P2_U3251) );
  INV_X1 U10482 ( .A(n9005), .ZN(n8993) );
  NOR3_X1 U10483 ( .A1(n8991), .A2(n8990), .A3(n8989), .ZN(n8992) );
  NOR3_X1 U10484 ( .A1(n8993), .A2(n8992), .A3(n9094), .ZN(n8994) );
  AOI21_X1 U10485 ( .B1(n9077), .B2(n8995), .A(n8994), .ZN(n9002) );
  OAI211_X1 U10486 ( .C1(n8998), .C2(n8997), .A(n9088), .B(n8996), .ZN(n9000)
         );
  NAND2_X1 U10487 ( .A1(n9056), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n8999) );
  NAND4_X1 U10488 ( .A1(n9002), .A2(n9001), .A3(n9000), .A4(n8999), .ZN(
        P2_U3252) );
  INV_X1 U10489 ( .A(n9023), .ZN(n9007) );
  NAND3_X1 U10490 ( .A1(n9005), .A2(n9004), .A3(n9003), .ZN(n9006) );
  NAND3_X1 U10491 ( .A1(n9007), .A2(n9051), .A3(n9006), .ZN(n9017) );
  INV_X1 U10492 ( .A(n9008), .ZN(n9011) );
  NOR2_X1 U10493 ( .A1(n9090), .A2(n9009), .ZN(n9010) );
  AOI211_X1 U10494 ( .C1(n9056), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n9011), .B(
        n9010), .ZN(n9016) );
  OAI211_X1 U10495 ( .C1(n9014), .C2(n9013), .A(n9088), .B(n9012), .ZN(n9015)
         );
  NAND3_X1 U10496 ( .A1(n9017), .A2(n9016), .A3(n9015), .ZN(P2_U3253) );
  INV_X1 U10497 ( .A(n9018), .ZN(n9020) );
  MUX2_X1 U10498 ( .A(n7287), .B(P2_REG2_REG_9__SCAN_IN), .S(n9029), .Z(n9019)
         );
  NAND2_X1 U10499 ( .A1(n9020), .A2(n9019), .ZN(n9022) );
  OAI211_X1 U10500 ( .C1(n9023), .C2(n9022), .A(n9021), .B(n9051), .ZN(n9033)
         );
  INV_X1 U10501 ( .A(n9024), .ZN(n9025) );
  AOI21_X1 U10502 ( .B1(n9056), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n9025), .ZN(
        n9032) );
  OAI211_X1 U10503 ( .C1(n9028), .C2(n9027), .A(n9026), .B(n9088), .ZN(n9031)
         );
  NAND2_X1 U10504 ( .A1(n9077), .A2(n9029), .ZN(n9030) );
  NAND4_X1 U10505 ( .A1(n9033), .A2(n9032), .A3(n9031), .A4(n9030), .ZN(
        P2_U3254) );
  OAI21_X1 U10506 ( .B1(n9036), .B2(n9035), .A(n9034), .ZN(n9037) );
  NAND2_X1 U10507 ( .A1(n9037), .A2(n9051), .ZN(n9046) );
  AOI21_X1 U10508 ( .B1(n9056), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9038), .ZN(
        n9045) );
  OAI211_X1 U10509 ( .C1(n9041), .C2(n9040), .A(n9039), .B(n9088), .ZN(n9044)
         );
  NAND2_X1 U10510 ( .A1(n9077), .A2(n9042), .ZN(n9043) );
  NAND4_X1 U10511 ( .A1(n9046), .A2(n9045), .A3(n9044), .A4(n9043), .ZN(
        P2_U3256) );
  NAND2_X1 U10512 ( .A1(n9061), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9050) );
  INV_X1 U10513 ( .A(n9047), .ZN(n9048) );
  INV_X1 U10514 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9298) );
  XNOR2_X1 U10515 ( .A(n9072), .B(n9298), .ZN(n9052) );
  OAI211_X1 U10516 ( .C1(n9053), .C2(n9052), .A(n9051), .B(n9066), .ZN(n9058)
         );
  NOR2_X1 U10517 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9054), .ZN(n9055) );
  AOI21_X1 U10518 ( .B1(n9056), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9055), .ZN(
        n9057) );
  OAI211_X1 U10519 ( .C1(n9090), .C2(n9059), .A(n9058), .B(n9057), .ZN(n9065)
         );
  OAI21_X1 U10520 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n9061), .A(n9060), .ZN(
        n9063) );
  XNOR2_X1 U10521 ( .A(n9072), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9062) );
  NOR2_X1 U10522 ( .A1(n9062), .A2(n9063), .ZN(n9071) );
  AOI211_X1 U10523 ( .C1(n9063), .C2(n9062), .A(n9071), .B(n9092), .ZN(n9064)
         );
  OR2_X1 U10524 ( .A1(n9065), .A2(n9064), .ZN(P2_U3262) );
  NAND2_X1 U10525 ( .A1(n9072), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U10526 ( .A1(n9067), .A2(n9066), .ZN(n9068) );
  AOI21_X1 U10527 ( .B1(n9069), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9081), .ZN(
        n9079) );
  XNOR2_X1 U10528 ( .A(n9083), .B(n9070), .ZN(n9086) );
  AOI21_X1 U10529 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9072), .A(n9071), .ZN(
        n9085) );
  XNOR2_X1 U10530 ( .A(n9086), .B(n9085), .ZN(n9073) );
  NAND2_X1 U10531 ( .A1(n9088), .A2(n9073), .ZN(n9075) );
  OAI211_X1 U10532 ( .C1(n10460), .C2(n9097), .A(n9075), .B(n9074), .ZN(n9076)
         );
  AOI21_X1 U10533 ( .B1(n9083), .B2(n9077), .A(n9076), .ZN(n9078) );
  OAI21_X1 U10534 ( .B1(n9079), .B2(n9094), .A(n9078), .ZN(P2_U3263) );
  NOR2_X1 U10535 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  XNOR2_X1 U10536 ( .A(n9082), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n9095) );
  INV_X1 U10537 ( .A(n9095), .ZN(n9091) );
  NOR2_X1 U10538 ( .A1(n9083), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9084) );
  AOI21_X1 U10539 ( .B1(n9086), .B2(n9085), .A(n9084), .ZN(n9087) );
  XNOR2_X1 U10540 ( .A(n9087), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U10541 ( .A1(n9088), .A2(n9093), .ZN(n9089) );
  INV_X1 U10542 ( .A(n9099), .ZN(n9373) );
  NAND2_X1 U10543 ( .A1(n4441), .A2(n9100), .ZN(n9372) );
  NAND3_X1 U10544 ( .A1(n9373), .A2(n10332), .A3(n9372), .ZN(n9103) );
  AOI21_X1 U10545 ( .B1(n10337), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9101), .ZN(
        n9102) );
  OAI211_X1 U10546 ( .C1(n4781), .C2(n9356), .A(n9103), .B(n9102), .ZN(
        P2_U3266) );
  NAND2_X1 U10547 ( .A1(n9104), .A2(n10332), .ZN(n9107) );
  AOI22_X1 U10548 ( .A1(n9105), .A2(n10330), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n10337), .ZN(n9106) );
  OAI211_X1 U10549 ( .C1(n9108), .C2(n9356), .A(n9107), .B(n9106), .ZN(n9109)
         );
  AOI21_X1 U10550 ( .B1(n9110), .B2(n9196), .A(n9109), .ZN(n9111) );
  OAI21_X1 U10551 ( .B1(n9112), .B2(n10337), .A(n9111), .ZN(P2_U3268) );
  AOI21_X1 U10552 ( .B1(n9113), .B2(n9120), .A(n9351), .ZN(n9118) );
  OAI22_X1 U10553 ( .A1(n9115), .A2(n9312), .B1(n9114), .B2(n6215), .ZN(n9116)
         );
  AOI21_X1 U10554 ( .B1(n9118), .B2(n9117), .A(n9116), .ZN(n9392) );
  OAI21_X1 U10555 ( .B1(n9121), .B2(n9120), .A(n9119), .ZN(n9388) );
  OR2_X1 U10556 ( .A1(n9127), .A2(n9133), .ZN(n9122) );
  AND2_X1 U10557 ( .A1(n9123), .A2(n9122), .ZN(n9390) );
  NAND2_X1 U10558 ( .A1(n9390), .A2(n10332), .ZN(n9126) );
  AOI22_X1 U10559 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(n10337), .B1(n9124), 
        .B2(n10330), .ZN(n9125) );
  OAI211_X1 U10560 ( .C1(n9127), .C2(n9356), .A(n9126), .B(n9125), .ZN(n9128)
         );
  AOI21_X1 U10561 ( .B1(n9388), .B2(n9196), .A(n9128), .ZN(n9129) );
  OAI21_X1 U10562 ( .B1(n10337), .B2(n9392), .A(n9129), .ZN(P2_U3269) );
  AOI211_X1 U10563 ( .C1(n9394), .C2(n4418), .A(n6279), .B(n9133), .ZN(n9134)
         );
  NOR2_X1 U10564 ( .A1(n9135), .A2(n9134), .ZN(n9396) );
  OAI21_X1 U10565 ( .B1(n9135), .B2(n9154), .A(n10335), .ZN(n9144) );
  OAI21_X1 U10566 ( .B1(n9138), .B2(n9137), .A(n9136), .ZN(n9395) );
  AOI22_X1 U10567 ( .A1(n10337), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n9139), 
        .B2(n10330), .ZN(n9140) );
  OAI21_X1 U10568 ( .B1(n9141), .B2(n9356), .A(n9140), .ZN(n9142) );
  AOI21_X1 U10569 ( .B1(n9395), .B2(n9196), .A(n9142), .ZN(n9143) );
  OAI21_X1 U10570 ( .B1(n9396), .B2(n9144), .A(n9143), .ZN(P2_U3270) );
  INV_X1 U10571 ( .A(n9145), .ZN(n9146) );
  AOI21_X1 U10572 ( .B1(n9146), .B2(n4549), .A(n9351), .ZN(n9149) );
  AOI21_X1 U10573 ( .B1(n9149), .B2(n9148), .A(n9147), .ZN(n9402) );
  OAI21_X1 U10574 ( .B1(n9151), .B2(n4549), .A(n9150), .ZN(n9398) );
  XNOR2_X1 U10575 ( .A(n9168), .B(n9152), .ZN(n9153) );
  NOR2_X1 U10576 ( .A1(n9153), .A2(n6279), .ZN(n9399) );
  AND2_X1 U10577 ( .A1(n10335), .A2(n9154), .ZN(n9304) );
  NAND2_X1 U10578 ( .A1(n9399), .A2(n9304), .ZN(n9159) );
  INV_X1 U10579 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9156) );
  OAI22_X1 U10580 ( .A1(n10335), .A2(n9156), .B1(n9155), .B2(n9359), .ZN(n9157) );
  AOI21_X1 U10581 ( .B1(n9400), .B2(n9300), .A(n9157), .ZN(n9158) );
  NAND2_X1 U10582 ( .A1(n9159), .A2(n9158), .ZN(n9160) );
  AOI21_X1 U10583 ( .B1(n9398), .B2(n9196), .A(n9160), .ZN(n9161) );
  OAI21_X1 U10584 ( .B1(n10337), .B2(n9402), .A(n9161), .ZN(P2_U3271) );
  XNOR2_X1 U10585 ( .A(n9163), .B(n9162), .ZN(n9166) );
  AOI222_X1 U10586 ( .A1(n10313), .A2(n9166), .B1(n9165), .B2(n10316), .C1(
        n9164), .C2(n10317), .ZN(n9407) );
  NOR2_X1 U10587 ( .A1(n9187), .A2(n9172), .ZN(n9167) );
  NOR2_X1 U10588 ( .A1(n9168), .A2(n9167), .ZN(n9405) );
  INV_X1 U10589 ( .A(n9169), .ZN(n9170) );
  AOI22_X1 U10590 ( .A1(n10337), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9170), 
        .B2(n10330), .ZN(n9171) );
  OAI21_X1 U10591 ( .B1(n9172), .B2(n9356), .A(n9171), .ZN(n9176) );
  XNOR2_X1 U10592 ( .A(n9174), .B(n9173), .ZN(n9408) );
  NOR2_X1 U10593 ( .A1(n9408), .A2(n9366), .ZN(n9175) );
  AOI211_X1 U10594 ( .C1(n9405), .C2(n10332), .A(n9176), .B(n9175), .ZN(n9177)
         );
  OAI21_X1 U10595 ( .B1(n10337), .B2(n9407), .A(n9177), .ZN(P2_U3272) );
  OAI21_X1 U10596 ( .B1(n9180), .B2(n9179), .A(n9178), .ZN(n9182) );
  AOI222_X1 U10597 ( .A1(n10313), .A2(n9182), .B1(n9181), .B2(n10316), .C1(
        n9224), .C2(n10317), .ZN(n9413) );
  OAI21_X1 U10598 ( .B1(n9185), .B2(n9184), .A(n9183), .ZN(n9414) );
  INV_X1 U10599 ( .A(n9414), .ZN(n9197) );
  NOR2_X1 U10600 ( .A1(n9201), .A2(n9409), .ZN(n9186) );
  OR2_X1 U10601 ( .A1(n9187), .A2(n9186), .ZN(n9410) );
  INV_X1 U10602 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9190) );
  INV_X1 U10603 ( .A(n9188), .ZN(n9189) );
  OAI22_X1 U10604 ( .A1(n10335), .A2(n9190), .B1(n9189), .B2(n9359), .ZN(n9191) );
  AOI21_X1 U10605 ( .B1(n9192), .B2(n9300), .A(n9191), .ZN(n9193) );
  OAI21_X1 U10606 ( .B1(n9410), .B2(n9194), .A(n9193), .ZN(n9195) );
  AOI21_X1 U10607 ( .B1(n9197), .B2(n9196), .A(n9195), .ZN(n9198) );
  OAI21_X1 U10608 ( .B1(n10337), .B2(n9413), .A(n9198), .ZN(P2_U3273) );
  XNOR2_X1 U10609 ( .A(n9200), .B(n9199), .ZN(n9419) );
  AOI21_X1 U10610 ( .B1(n9415), .B2(n9214), .A(n9201), .ZN(n9416) );
  AOI22_X1 U10611 ( .A1(n10337), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9202), 
        .B2(n10330), .ZN(n9203) );
  OAI21_X1 U10612 ( .B1(n4787), .B2(n9356), .A(n9203), .ZN(n9210) );
  AOI21_X1 U10613 ( .B1(n9204), .B2(n9205), .A(n9351), .ZN(n9208) );
  OAI22_X1 U10614 ( .A1(n9206), .A2(n9312), .B1(n9248), .B2(n6215), .ZN(n9207)
         );
  AOI21_X1 U10615 ( .B1(n9208), .B2(n4806), .A(n9207), .ZN(n9418) );
  NOR2_X1 U10616 ( .A1(n9418), .A2(n10337), .ZN(n9209) );
  AOI211_X1 U10617 ( .C1(n9416), .C2(n10332), .A(n9210), .B(n9209), .ZN(n9211)
         );
  OAI21_X1 U10618 ( .B1(n9419), .B2(n9366), .A(n9211), .ZN(P2_U3274) );
  XNOR2_X1 U10619 ( .A(n9212), .B(n9213), .ZN(n9424) );
  INV_X1 U10620 ( .A(n9214), .ZN(n9215) );
  AOI21_X1 U10621 ( .B1(n9420), .B2(n9232), .A(n9215), .ZN(n9421) );
  INV_X1 U10622 ( .A(n9216), .ZN(n9217) );
  AOI22_X1 U10623 ( .A1(n10337), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9217), 
        .B2(n10330), .ZN(n9218) );
  OAI21_X1 U10624 ( .B1(n9219), .B2(n9356), .A(n9218), .ZN(n9227) );
  OAI21_X1 U10625 ( .B1(n9220), .B2(n9222), .A(n9221), .ZN(n9225) );
  AOI222_X1 U10626 ( .A1(n10313), .A2(n9225), .B1(n9224), .B2(n10316), .C1(
        n9223), .C2(n10317), .ZN(n9423) );
  NOR2_X1 U10627 ( .A1(n9423), .A2(n10337), .ZN(n9226) );
  AOI211_X1 U10628 ( .C1(n9421), .C2(n10332), .A(n9227), .B(n9226), .ZN(n9228)
         );
  OAI21_X1 U10629 ( .B1(n9424), .B2(n9366), .A(n9228), .ZN(P2_U3275) );
  OAI21_X1 U10630 ( .B1(n9231), .B2(n9230), .A(n9229), .ZN(n9429) );
  INV_X1 U10631 ( .A(n9265), .ZN(n9234) );
  INV_X1 U10632 ( .A(n9232), .ZN(n9233) );
  AOI21_X1 U10633 ( .B1(n9425), .B2(n9234), .A(n9233), .ZN(n9426) );
  AOI22_X1 U10634 ( .A1(n10337), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9235), 
        .B2(n10330), .ZN(n9236) );
  OAI21_X1 U10635 ( .B1(n9237), .B2(n9356), .A(n9236), .ZN(n9252) );
  NAND2_X1 U10636 ( .A1(n9239), .A2(n9238), .ZN(n9279) );
  NAND2_X1 U10637 ( .A1(n9279), .A2(n9240), .ZN(n9260) );
  INV_X1 U10638 ( .A(n9255), .ZN(n9258) );
  NAND3_X1 U10639 ( .A1(n9260), .A2(n9258), .A3(n9259), .ZN(n9257) );
  AOI21_X1 U10640 ( .B1(n9257), .B2(n9242), .A(n9241), .ZN(n9246) );
  INV_X1 U10641 ( .A(n9244), .ZN(n9245) );
  NOR3_X1 U10642 ( .A1(n9246), .A2(n9245), .A3(n9351), .ZN(n9250) );
  OAI22_X1 U10643 ( .A1(n9248), .A2(n9312), .B1(n9247), .B2(n6215), .ZN(n9249)
         );
  NOR2_X1 U10644 ( .A1(n9250), .A2(n9249), .ZN(n9428) );
  NOR2_X1 U10645 ( .A1(n9428), .A2(n10337), .ZN(n9251) );
  AOI211_X1 U10646 ( .C1(n9426), .C2(n10332), .A(n9252), .B(n9251), .ZN(n9253)
         );
  OAI21_X1 U10647 ( .B1(n9366), .B2(n9429), .A(n9253), .ZN(P2_U3276) );
  OAI21_X1 U10648 ( .B1(n9256), .B2(n9255), .A(n9254), .ZN(n9434) );
  INV_X1 U10649 ( .A(n9257), .ZN(n9262) );
  AOI21_X1 U10650 ( .B1(n9260), .B2(n9259), .A(n9258), .ZN(n9261) );
  OAI21_X1 U10651 ( .B1(n9262), .B2(n9261), .A(n10313), .ZN(n9264) );
  NAND2_X1 U10652 ( .A1(n9264), .A2(n9263), .ZN(n9430) );
  INV_X1 U10653 ( .A(n9274), .ZN(n9266) );
  AOI211_X1 U10654 ( .C1(n9432), .C2(n9266), .A(n6279), .B(n9265), .ZN(n9431)
         );
  NAND2_X1 U10655 ( .A1(n9431), .A2(n9304), .ZN(n9269) );
  AOI22_X1 U10656 ( .A1(n10337), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9267), 
        .B2(n10330), .ZN(n9268) );
  OAI211_X1 U10657 ( .C1(n9270), .C2(n9356), .A(n9269), .B(n9268), .ZN(n9271)
         );
  AOI21_X1 U10658 ( .B1(n9430), .B2(n10335), .A(n9271), .ZN(n9272) );
  OAI21_X1 U10659 ( .B1(n9434), .B2(n9366), .A(n9272), .ZN(P2_U3277) );
  XOR2_X1 U10660 ( .A(n9278), .B(n9273), .Z(n9439) );
  AOI21_X1 U10661 ( .B1(n9435), .B2(n9302), .A(n9274), .ZN(n9436) );
  AOI22_X1 U10662 ( .A1(n10337), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9275), 
        .B2(n10330), .ZN(n9276) );
  OAI21_X1 U10663 ( .B1(n9277), .B2(n9356), .A(n9276), .ZN(n9284) );
  XNOR2_X1 U10664 ( .A(n9279), .B(n9278), .ZN(n9282) );
  AOI222_X1 U10665 ( .A1(n10313), .A2(n9282), .B1(n9281), .B2(n10316), .C1(
        n9280), .C2(n10317), .ZN(n9438) );
  NOR2_X1 U10666 ( .A1(n9438), .A2(n10337), .ZN(n9283) );
  AOI211_X1 U10667 ( .C1(n9436), .C2(n10332), .A(n9284), .B(n9283), .ZN(n9285)
         );
  OAI21_X1 U10668 ( .B1(n9439), .B2(n9366), .A(n9285), .ZN(P2_U3278) );
  NAND2_X1 U10669 ( .A1(n9309), .A2(n9286), .ZN(n9287) );
  XNOR2_X1 U10670 ( .A(n9287), .B(n9292), .ZN(n9288) );
  OAI222_X1 U10671 ( .A1(n6215), .A2(n9290), .B1(n9312), .B2(n9289), .C1(n9288), .C2(n9351), .ZN(n9440) );
  AOI21_X1 U10672 ( .B1(n9291), .B2(n9293), .A(n9292), .ZN(n9296) );
  INV_X1 U10673 ( .A(n9294), .ZN(n9295) );
  NOR2_X1 U10674 ( .A1(n9296), .A2(n9295), .ZN(n9444) );
  OAI22_X1 U10675 ( .A1(n10335), .A2(n9298), .B1(n9297), .B2(n9359), .ZN(n9299) );
  AOI21_X1 U10676 ( .B1(n9442), .B2(n9300), .A(n9299), .ZN(n9306) );
  AOI21_X1 U10677 ( .B1(n9301), .B2(n9442), .A(n6279), .ZN(n9303) );
  AND2_X1 U10678 ( .A1(n9303), .A2(n9302), .ZN(n9441) );
  NAND2_X1 U10679 ( .A1(n9441), .A2(n9304), .ZN(n9305) );
  OAI211_X1 U10680 ( .C1(n9444), .C2(n9366), .A(n9306), .B(n9305), .ZN(n9307)
         );
  AOI21_X1 U10681 ( .B1(n10335), .B2(n9440), .A(n9307), .ZN(n9308) );
  INV_X1 U10682 ( .A(n9308), .ZN(P2_U3279) );
  OAI21_X1 U10683 ( .B1(n9315), .B2(n9310), .A(n9309), .ZN(n9321) );
  OAI22_X1 U10684 ( .A1(n9313), .A2(n9312), .B1(n9311), .B2(n6215), .ZN(n9320)
         );
  NAND2_X1 U10685 ( .A1(n9343), .A2(n9314), .ZN(n9316) );
  NAND2_X1 U10686 ( .A1(n9316), .A2(n9315), .ZN(n9317) );
  NAND2_X1 U10687 ( .A1(n9291), .A2(n9317), .ZN(n9449) );
  NOR2_X1 U10688 ( .A1(n9449), .A2(n9318), .ZN(n9319) );
  AOI211_X1 U10689 ( .C1(n10313), .C2(n9321), .A(n9320), .B(n9319), .ZN(n9448)
         );
  INV_X1 U10690 ( .A(n9337), .ZN(n9323) );
  INV_X1 U10691 ( .A(n9301), .ZN(n9322) );
  AOI21_X1 U10692 ( .B1(n9445), .B2(n9323), .A(n9322), .ZN(n9446) );
  AOI22_X1 U10693 ( .A1(n10337), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9324), 
        .B2(n10330), .ZN(n9325) );
  OAI21_X1 U10694 ( .B1(n9326), .B2(n9356), .A(n9325), .ZN(n9329) );
  NOR2_X1 U10695 ( .A1(n9449), .A2(n9327), .ZN(n9328) );
  AOI211_X1 U10696 ( .C1(n9446), .C2(n10332), .A(n9329), .B(n9328), .ZN(n9330)
         );
  OAI21_X1 U10697 ( .B1(n9448), .B2(n10337), .A(n9330), .ZN(P2_U3280) );
  NAND2_X1 U10698 ( .A1(n9332), .A2(n9331), .ZN(n9352) );
  NOR2_X1 U10699 ( .A1(n9352), .A2(n9364), .ZN(n9350) );
  AOI21_X1 U10700 ( .B1(n9357), .B2(n9334), .A(n9350), .ZN(n9333) );
  XNOR2_X1 U10701 ( .A(n9333), .B(n9345), .ZN(n9336) );
  AOI222_X1 U10702 ( .A1(n10313), .A2(n9336), .B1(n9335), .B2(n10316), .C1(
        n9334), .C2(n10317), .ZN(n9453) );
  INV_X1 U10703 ( .A(n9355), .ZN(n9338) );
  AOI21_X1 U10704 ( .B1(n9450), .B2(n9338), .A(n9337), .ZN(n9451) );
  AOI22_X1 U10705 ( .A1(n10337), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9339), 
        .B2(n10330), .ZN(n9340) );
  OAI21_X1 U10706 ( .B1(n9341), .B2(n9356), .A(n9340), .ZN(n9348) );
  INV_X1 U10707 ( .A(n9342), .ZN(n9346) );
  INV_X1 U10708 ( .A(n9343), .ZN(n9344) );
  AOI21_X1 U10709 ( .B1(n9346), .B2(n9345), .A(n9344), .ZN(n9454) );
  NOR2_X1 U10710 ( .A1(n9454), .A2(n9366), .ZN(n9347) );
  AOI211_X1 U10711 ( .C1(n9451), .C2(n10332), .A(n9348), .B(n9347), .ZN(n9349)
         );
  OAI21_X1 U10712 ( .B1(n10337), .B2(n9453), .A(n9349), .ZN(P2_U3281) );
  AOI211_X1 U10713 ( .C1(n9364), .C2(n9352), .A(n9351), .B(n9350), .ZN(n9354)
         );
  NOR2_X1 U10714 ( .A1(n9354), .A2(n9353), .ZN(n9458) );
  AOI21_X1 U10715 ( .B1(n9455), .B2(n4397), .A(n9355), .ZN(n9456) );
  NOR2_X1 U10716 ( .A1(n9357), .A2(n9356), .ZN(n9363) );
  INV_X1 U10717 ( .A(n9358), .ZN(n9360) );
  OAI22_X1 U10718 ( .A1(n10335), .A2(n9361), .B1(n9360), .B2(n9359), .ZN(n9362) );
  AOI211_X1 U10719 ( .C1(n9456), .C2(n10332), .A(n9363), .B(n9362), .ZN(n9368)
         );
  XNOR2_X1 U10720 ( .A(n9365), .B(n9364), .ZN(n9459) );
  OR2_X1 U10721 ( .A1(n9459), .A2(n9366), .ZN(n9367) );
  OAI211_X1 U10722 ( .C1(n9458), .C2(n10337), .A(n9368), .B(n9367), .ZN(
        P2_U3282) );
  NAND2_X1 U10723 ( .A1(n9369), .A2(n10396), .ZN(n9370) );
  OAI211_X1 U10724 ( .C1(n9371), .C2(n6279), .A(n9370), .B(n9374), .ZN(n9476)
         );
  MUX2_X1 U10725 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9476), .S(n10423), .Z(
        P2_U3551) );
  NAND3_X1 U10726 ( .A1(n9373), .A2(n10398), .A3(n9372), .ZN(n9375) );
  OAI211_X1 U10727 ( .C1(n4781), .C2(n10390), .A(n9375), .B(n9374), .ZN(n9477)
         );
  MUX2_X1 U10728 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9477), .S(n10423), .Z(
        P2_U3550) );
  NAND3_X1 U10729 ( .A1(n9377), .A2(n9376), .A3(n10393), .ZN(n9381) );
  NAND2_X1 U10730 ( .A1(n9378), .A2(n10396), .ZN(n9379) );
  AND3_X1 U10731 ( .A1(n9381), .A2(n9380), .A3(n9379), .ZN(n9383) );
  INV_X1 U10732 ( .A(n9388), .ZN(n9393) );
  AOI22_X1 U10733 ( .A1(n9390), .A2(n10398), .B1(n9389), .B2(n10396), .ZN(
        n9391) );
  OAI211_X1 U10734 ( .C1(n9393), .C2(n9475), .A(n9392), .B(n9391), .ZN(n9478)
         );
  MUX2_X1 U10735 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9478), .S(n10423), .Z(
        P2_U3547) );
  AOI22_X1 U10736 ( .A1(n9395), .A2(n10393), .B1(n9394), .B2(n10396), .ZN(
        n9397) );
  NAND2_X1 U10737 ( .A1(n9397), .A2(n9396), .ZN(n9479) );
  MUX2_X1 U10738 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9479), .S(n10423), .Z(
        P2_U3546) );
  INV_X1 U10739 ( .A(n9398), .ZN(n9403) );
  AOI21_X1 U10740 ( .B1(n9400), .B2(n10396), .A(n9399), .ZN(n9401) );
  OAI211_X1 U10741 ( .C1(n9403), .C2(n9475), .A(n9402), .B(n9401), .ZN(n9480)
         );
  MUX2_X1 U10742 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9480), .S(n10423), .Z(
        P2_U3545) );
  AOI22_X1 U10743 ( .A1(n9405), .A2(n10398), .B1(n9404), .B2(n10396), .ZN(
        n9406) );
  OAI211_X1 U10744 ( .C1(n9408), .C2(n9475), .A(n9407), .B(n9406), .ZN(n9481)
         );
  MUX2_X1 U10745 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9481), .S(n10423), .Z(
        P2_U3544) );
  OAI22_X1 U10746 ( .A1(n9410), .A2(n6279), .B1(n9409), .B2(n10390), .ZN(n9411) );
  INV_X1 U10747 ( .A(n9411), .ZN(n9412) );
  OAI211_X1 U10748 ( .C1(n9414), .C2(n9475), .A(n9413), .B(n9412), .ZN(n9482)
         );
  MUX2_X1 U10749 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9482), .S(n10423), .Z(
        P2_U3543) );
  AOI22_X1 U10750 ( .A1(n9416), .A2(n10398), .B1(n9415), .B2(n10396), .ZN(
        n9417) );
  OAI211_X1 U10751 ( .C1(n9419), .C2(n9475), .A(n9418), .B(n9417), .ZN(n9483)
         );
  MUX2_X1 U10752 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9483), .S(n10423), .Z(
        P2_U3542) );
  AOI22_X1 U10753 ( .A1(n9421), .A2(n10398), .B1(n9420), .B2(n10396), .ZN(
        n9422) );
  OAI211_X1 U10754 ( .C1(n9424), .C2(n9475), .A(n9423), .B(n9422), .ZN(n9484)
         );
  MUX2_X1 U10755 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9484), .S(n10423), .Z(
        P2_U3541) );
  AOI22_X1 U10756 ( .A1(n9426), .A2(n10398), .B1(n9425), .B2(n10396), .ZN(
        n9427) );
  OAI211_X1 U10757 ( .C1(n9429), .C2(n9475), .A(n9428), .B(n9427), .ZN(n9485)
         );
  MUX2_X1 U10758 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9485), .S(n10423), .Z(
        P2_U3540) );
  AOI211_X1 U10759 ( .C1(n9432), .C2(n10396), .A(n9431), .B(n9430), .ZN(n9433)
         );
  OAI21_X1 U10760 ( .B1(n9475), .B2(n9434), .A(n9433), .ZN(n9486) );
  MUX2_X1 U10761 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9486), .S(n10423), .Z(
        P2_U3539) );
  AOI22_X1 U10762 ( .A1(n9436), .A2(n10398), .B1(n9435), .B2(n10396), .ZN(
        n9437) );
  OAI211_X1 U10763 ( .C1(n9439), .C2(n9475), .A(n9438), .B(n9437), .ZN(n9487)
         );
  MUX2_X1 U10764 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9487), .S(n10423), .Z(
        P2_U3538) );
  AOI211_X1 U10765 ( .C1(n9442), .C2(n10396), .A(n9441), .B(n9440), .ZN(n9443)
         );
  OAI21_X1 U10766 ( .B1(n9475), .B2(n9444), .A(n9443), .ZN(n9488) );
  MUX2_X1 U10767 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9488), .S(n10423), .Z(
        P2_U3537) );
  AOI22_X1 U10768 ( .A1(n9446), .A2(n10398), .B1(n9445), .B2(n10396), .ZN(
        n9447) );
  OAI211_X1 U10769 ( .C1(n10402), .C2(n9449), .A(n9448), .B(n9447), .ZN(n9489)
         );
  MUX2_X1 U10770 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9489), .S(n10423), .Z(
        P2_U3536) );
  AOI22_X1 U10771 ( .A1(n9451), .A2(n10398), .B1(n9450), .B2(n10396), .ZN(
        n9452) );
  OAI211_X1 U10772 ( .C1(n9475), .C2(n9454), .A(n9453), .B(n9452), .ZN(n9490)
         );
  MUX2_X1 U10773 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9490), .S(n10423), .Z(
        P2_U3535) );
  AOI22_X1 U10774 ( .A1(n9456), .A2(n10398), .B1(n9455), .B2(n10396), .ZN(
        n9457) );
  OAI211_X1 U10775 ( .C1(n9475), .C2(n9459), .A(n9458), .B(n9457), .ZN(n9491)
         );
  MUX2_X1 U10776 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9491), .S(n10423), .Z(
        P2_U3534) );
  AOI22_X1 U10777 ( .A1(n9461), .A2(n10398), .B1(n9460), .B2(n10396), .ZN(
        n9462) );
  OAI211_X1 U10778 ( .C1(n10402), .C2(n9464), .A(n9463), .B(n9462), .ZN(n9492)
         );
  MUX2_X1 U10779 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9492), .S(n10423), .Z(
        P2_U3533) );
  AOI22_X1 U10780 ( .A1(n9466), .A2(n10398), .B1(n9465), .B2(n10396), .ZN(
        n9467) );
  OAI211_X1 U10781 ( .C1(n9475), .C2(n9469), .A(n9468), .B(n9467), .ZN(n9493)
         );
  MUX2_X1 U10782 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9493), .S(n10423), .Z(
        P2_U3532) );
  AOI22_X1 U10783 ( .A1(n9471), .A2(n10398), .B1(n9470), .B2(n10396), .ZN(
        n9472) );
  OAI211_X1 U10784 ( .C1(n9475), .C2(n9474), .A(n9473), .B(n9472), .ZN(n9494)
         );
  MUX2_X1 U10785 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9494), .S(n10423), .Z(
        P2_U3531) );
  MUX2_X1 U10786 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9476), .S(n10407), .Z(
        P2_U3519) );
  MUX2_X1 U10787 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9477), .S(n10407), .Z(
        P2_U3518) );
  MUX2_X1 U10788 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9478), .S(n10407), .Z(
        P2_U3515) );
  MUX2_X1 U10789 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9479), .S(n10407), .Z(
        P2_U3514) );
  MUX2_X1 U10790 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9480), .S(n10407), .Z(
        P2_U3513) );
  MUX2_X1 U10791 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9481), .S(n10407), .Z(
        P2_U3512) );
  MUX2_X1 U10792 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9482), .S(n10407), .Z(
        P2_U3511) );
  MUX2_X1 U10793 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9483), .S(n10407), .Z(
        P2_U3510) );
  MUX2_X1 U10794 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9484), .S(n10407), .Z(
        P2_U3509) );
  MUX2_X1 U10795 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9485), .S(n10407), .Z(
        P2_U3508) );
  MUX2_X1 U10796 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9486), .S(n10407), .Z(
        P2_U3507) );
  MUX2_X1 U10797 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9487), .S(n10407), .Z(
        P2_U3505) );
  MUX2_X1 U10798 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9488), .S(n10407), .Z(
        P2_U3502) );
  MUX2_X1 U10799 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9489), .S(n10407), .Z(
        P2_U3499) );
  MUX2_X1 U10800 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9490), .S(n10407), .Z(
        P2_U3496) );
  MUX2_X1 U10801 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9491), .S(n10407), .Z(
        P2_U3493) );
  MUX2_X1 U10802 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9492), .S(n10407), .Z(
        P2_U3490) );
  MUX2_X1 U10803 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9493), .S(n10407), .Z(
        P2_U3487) );
  MUX2_X1 U10804 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9494), .S(n10407), .Z(
        P2_U3484) );
  INV_X1 U10805 ( .A(n9495), .ZN(n10219) );
  NOR4_X1 U10806 ( .A1(n5774), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9497), .A4(
        P2_U3152), .ZN(n9498) );
  AOI21_X1 U10807 ( .B1(n9499), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9498), .ZN(
        n9500) );
  OAI21_X1 U10808 ( .B1(n10219), .B2(n9506), .A(n9500), .ZN(P2_U3327) );
  INV_X1 U10809 ( .A(n9501), .ZN(n10228) );
  OAI222_X1 U10810 ( .A1(n9503), .A2(P2_U3152), .B1(n9511), .B2(n10228), .C1(
        n9502), .C2(n9508), .ZN(P2_U3330) );
  INV_X1 U10811 ( .A(n9504), .ZN(n10233) );
  OAI222_X1 U10812 ( .A1(n9507), .A2(P2_U3152), .B1(n9506), .B2(n10233), .C1(
        n9505), .C2(n9508), .ZN(P2_U3331) );
  OAI222_X1 U10813 ( .A1(n9512), .A2(P2_U3152), .B1(n9511), .B2(n9510), .C1(
        n9509), .C2(n9508), .ZN(P2_U3332) );
  MUX2_X1 U10814 ( .A(n9513), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10815 ( .A(n9515), .B(n9514), .ZN(n9516) );
  XNOR2_X1 U10816 ( .A(n9517), .B(n9516), .ZN(n9524) );
  OAI22_X1 U10817 ( .A1(n9793), .A2(n9629), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9518), .ZN(n9521) );
  NOR2_X1 U10818 ( .A1(n9519), .A2(n9657), .ZN(n9520) );
  AOI211_X1 U10819 ( .C1(n9632), .C2(n9786), .A(n9521), .B(n9520), .ZN(n9523)
         );
  NAND2_X1 U10820 ( .A1(n10089), .A2(n4380), .ZN(n9522) );
  OAI211_X1 U10821 ( .C1(n9524), .C2(n9636), .A(n9523), .B(n9522), .ZN(
        P1_U3212) );
  NAND2_X1 U10822 ( .A1(n9526), .A2(n9525), .ZN(n9527) );
  XOR2_X1 U10823 ( .A(n9528), .B(n9527), .Z(n9534) );
  AOI22_X1 U10824 ( .A1(n9864), .A2(n9632), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9530) );
  NAND2_X1 U10825 ( .A1(n9867), .A2(n9660), .ZN(n9529) );
  OAI211_X1 U10826 ( .C1(n9531), .C2(n9657), .A(n9530), .B(n9529), .ZN(n9532)
         );
  AOI21_X1 U10827 ( .B1(n10109), .B2(n4380), .A(n9532), .ZN(n9533) );
  OAI21_X1 U10828 ( .B1(n9534), .B2(n9636), .A(n9533), .ZN(P1_U3214) );
  OAI21_X1 U10829 ( .B1(n9537), .B2(n9536), .A(n9535), .ZN(n9541) );
  NAND2_X1 U10830 ( .A1(n9538), .A2(n9539), .ZN(n9622) );
  NAND2_X1 U10831 ( .A1(n9622), .A2(n9621), .ZN(n9626) );
  NAND2_X1 U10832 ( .A1(n9626), .A2(n9623), .ZN(n9540) );
  XOR2_X1 U10833 ( .A(n9541), .B(n9540), .Z(n9548) );
  NAND2_X1 U10834 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U10835 ( .A1(n9962), .A2(n9604), .ZN(n9542) );
  OAI211_X1 U10836 ( .C1(n9543), .C2(n9654), .A(n9750), .B(n9542), .ZN(n9544)
         );
  AOI21_X1 U10837 ( .B1(n9935), .B2(n9660), .A(n9544), .ZN(n9547) );
  NAND2_X1 U10838 ( .A1(n10133), .A2(n4380), .ZN(n9546) );
  OAI211_X1 U10839 ( .C1(n9548), .C2(n9636), .A(n9547), .B(n9546), .ZN(
        P1_U3217) );
  NAND2_X1 U10840 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  XOR2_X1 U10841 ( .A(n9552), .B(n9551), .Z(n9557) );
  AOI22_X1 U10842 ( .A1(n9931), .A2(n9604), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9554) );
  NAND2_X1 U10843 ( .A1(n9894), .A2(n9632), .ZN(n9553) );
  OAI211_X1 U10844 ( .C1(n9629), .C2(n9899), .A(n9554), .B(n9553), .ZN(n9555)
         );
  AOI21_X1 U10845 ( .B1(n10118), .B2(n4380), .A(n9555), .ZN(n9556) );
  OAI21_X1 U10846 ( .B1(n9557), .B2(n9636), .A(n9556), .ZN(P1_U3221) );
  XNOR2_X1 U10847 ( .A(n9559), .B(n9558), .ZN(n9560) );
  NAND2_X1 U10848 ( .A1(n9560), .A2(n9650), .ZN(n9566) );
  NOR2_X1 U10849 ( .A1(n9836), .A2(n9629), .ZN(n9564) );
  OAI22_X1 U10850 ( .A1(n9562), .A2(n9657), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9561), .ZN(n9563) );
  AOI211_X1 U10851 ( .C1(n9829), .C2(n9632), .A(n9564), .B(n9563), .ZN(n9565)
         );
  OAI211_X1 U10852 ( .C1(n9839), .C2(n9663), .A(n9566), .B(n9565), .ZN(
        P1_U3223) );
  INV_X1 U10853 ( .A(n10149), .ZN(n9985) );
  NOR2_X1 U10854 ( .A1(n9648), .A2(n9647), .ZN(n9646) );
  NAND2_X1 U10855 ( .A1(n9580), .A2(n9571), .ZN(n9572) );
  NOR3_X1 U10856 ( .A1(n9646), .A2(n9651), .A3(n9572), .ZN(n9583) );
  OAI21_X1 U10857 ( .B1(n9646), .B2(n9651), .A(n9572), .ZN(n9573) );
  INV_X1 U10858 ( .A(n9573), .ZN(n9574) );
  OAI21_X1 U10859 ( .B1(n9583), .B2(n9574), .A(n9650), .ZN(n9579) );
  OAI21_X1 U10860 ( .B1(n9654), .B2(n9628), .A(n9575), .ZN(n9577) );
  NOR2_X1 U10861 ( .A1(n9629), .A2(n9982), .ZN(n9576) );
  AOI211_X1 U10862 ( .C1(n9604), .C2(n9978), .A(n9577), .B(n9576), .ZN(n9578)
         );
  OAI211_X1 U10863 ( .C1(n9985), .C2(n9663), .A(n9579), .B(n9578), .ZN(
        P1_U3224) );
  INV_X1 U10864 ( .A(n9580), .ZN(n9582) );
  NOR3_X1 U10865 ( .A1(n9583), .A2(n9582), .A3(n9581), .ZN(n9586) );
  INV_X1 U10866 ( .A(n9584), .ZN(n9585) );
  OAI21_X1 U10867 ( .B1(n9586), .B2(n9585), .A(n9650), .ZN(n9591) );
  NAND2_X1 U10868 ( .A1(n9604), .A2(n9998), .ZN(n9587) );
  NAND2_X1 U10869 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9714) );
  OAI211_X1 U10870 ( .C1(n9588), .C2(n9654), .A(n9587), .B(n9714), .ZN(n9589)
         );
  AOI21_X1 U10871 ( .B1(n9966), .B2(n9660), .A(n9589), .ZN(n9590) );
  OAI211_X1 U10872 ( .C1(n9968), .C2(n9663), .A(n9591), .B(n9590), .ZN(
        P1_U3226) );
  INV_X1 U10873 ( .A(n9592), .ZN(n9593) );
  AOI21_X1 U10874 ( .B1(n9595), .B2(n9594), .A(n9593), .ZN(n9601) );
  OAI22_X1 U10875 ( .A1(n9852), .A2(n9657), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9596), .ZN(n9597) );
  AOI21_X1 U10876 ( .B1(n9808), .B2(n9632), .A(n9597), .ZN(n9598) );
  OAI21_X1 U10877 ( .B1(n9629), .B2(n9859), .A(n9598), .ZN(n9599) );
  AOI21_X1 U10878 ( .B1(n10106), .B2(n4380), .A(n9599), .ZN(n9600) );
  OAI21_X1 U10879 ( .B1(n9601), .B2(n9636), .A(n9600), .ZN(P1_U3227) );
  XOR2_X1 U10880 ( .A(n9603), .B(n9602), .Z(n9609) );
  AOI22_X1 U10881 ( .A1(n9876), .A2(n9632), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9606) );
  NAND2_X1 U10882 ( .A1(n9947), .A2(n9604), .ZN(n9605) );
  OAI211_X1 U10883 ( .C1(n9629), .C2(n9918), .A(n9606), .B(n9605), .ZN(n9607)
         );
  AOI21_X1 U10884 ( .B1(n10124), .B2(n4380), .A(n9607), .ZN(n9608) );
  OAI21_X1 U10885 ( .B1(n9609), .B2(n9636), .A(n9608), .ZN(P1_U3231) );
  INV_X1 U10886 ( .A(n9613), .ZN(n9610) );
  NOR2_X1 U10887 ( .A1(n9611), .A2(n9610), .ZN(n9616) );
  AOI21_X1 U10888 ( .B1(n9614), .B2(n9613), .A(n9612), .ZN(n9615) );
  OAI21_X1 U10889 ( .B1(n9616), .B2(n9615), .A(n9650), .ZN(n9620) );
  AOI22_X1 U10890 ( .A1(n9877), .A2(n9632), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9617) );
  OAI21_X1 U10891 ( .B1(n9910), .B2(n9657), .A(n9617), .ZN(n9618) );
  AOI21_X1 U10892 ( .B1(n9881), .B2(n9660), .A(n9618), .ZN(n9619) );
  OAI211_X1 U10893 ( .C1(n9883), .C2(n9663), .A(n9620), .B(n9619), .ZN(
        P1_U3233) );
  INV_X1 U10894 ( .A(n9623), .ZN(n9627) );
  AOI21_X1 U10895 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9624) );
  NOR2_X1 U10896 ( .A1(n9624), .A2(n9636), .ZN(n9625) );
  OAI21_X1 U10897 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(n9634) );
  NAND2_X1 U10898 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9725) );
  OAI21_X1 U10899 ( .B1(n9657), .B2(n9628), .A(n9725), .ZN(n9631) );
  NOR2_X1 U10900 ( .A1(n9629), .A2(n9952), .ZN(n9630) );
  AOI211_X1 U10901 ( .C1(n9632), .C2(n9947), .A(n9631), .B(n9630), .ZN(n9633)
         );
  OAI211_X1 U10902 ( .C1(n9955), .C2(n9663), .A(n9634), .B(n9633), .ZN(
        P1_U3236) );
  AOI21_X1 U10903 ( .B1(n9635), .B2(n9637), .A(n9636), .ZN(n9639) );
  NAND2_X1 U10904 ( .A1(n9639), .A2(n9638), .ZN(n9645) );
  OAI22_X1 U10905 ( .A1(n9853), .A2(n9657), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9640), .ZN(n9643) );
  NOR2_X1 U10906 ( .A1(n9641), .A2(n9654), .ZN(n9642) );
  AOI211_X1 U10907 ( .C1(n9814), .C2(n9660), .A(n9643), .B(n9642), .ZN(n9644)
         );
  OAI211_X1 U10908 ( .C1(n4568), .C2(n9663), .A(n9645), .B(n9644), .ZN(
        P1_U3238) );
  INV_X1 U10909 ( .A(n10154), .ZN(n10006) );
  INV_X1 U10910 ( .A(n9646), .ZN(n9652) );
  OAI21_X1 U10911 ( .B1(n9651), .B2(n9648), .A(n9647), .ZN(n9649) );
  OAI211_X1 U10912 ( .C1(n9652), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9662)
         );
  NOR2_X1 U10913 ( .A1(n9654), .A2(n9653), .ZN(n9659) );
  OAI21_X1 U10914 ( .B1(n9657), .B2(n9656), .A(n9655), .ZN(n9658) );
  AOI211_X1 U10915 ( .C1(n10004), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9661)
         );
  OAI211_X1 U10916 ( .C1(n10006), .C2(n9663), .A(n9662), .B(n9661), .ZN(
        P1_U3239) );
  MUX2_X1 U10917 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9664), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10918 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9665), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10919 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9786), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10920 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9807), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10921 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9829), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10922 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9808), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10923 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9864), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10924 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9877), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10925 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9894), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10926 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9876), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10927 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9931), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10928 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9947), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10929 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9962), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10930 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9979), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10931 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9998), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10932 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9978), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10933 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10042), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10934 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9666), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10935 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n10040), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10936 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9667), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10937 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9668), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10938 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9669), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10939 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9670), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10940 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9671), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10941 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9672), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10942 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9673), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10943 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9674), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10944 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9675), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10945 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n7134), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10946 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6650), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10947 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9676), .S(P1_U4006), .Z(
        P1_U3555) );
  NAND2_X1 U10948 ( .A1(n9678), .A2(n9677), .ZN(n9679) );
  AOI21_X1 U10949 ( .B1(n9680), .B2(n9679), .A(n9745), .ZN(n9681) );
  AOI211_X1 U10950 ( .C1(n9733), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9682), .B(
        n9681), .ZN(n9691) );
  NAND2_X1 U10951 ( .A1(n9684), .A2(n9683), .ZN(n9685) );
  AOI21_X1 U10952 ( .B1(n9686), .B2(n9685), .A(n9746), .ZN(n9687) );
  AOI21_X1 U10953 ( .B1(n9696), .B2(n9688), .A(n9687), .ZN(n9690) );
  NAND3_X1 U10954 ( .A1(n9691), .A2(n9690), .A3(n9689), .ZN(P1_U3245) );
  XNOR2_X1 U10955 ( .A(n9693), .B(n9692), .ZN(n9694) );
  AOI22_X1 U10956 ( .A1(n9697), .A2(n9696), .B1(n9695), .B2(n9694), .ZN(n9706)
         );
  OAI211_X1 U10957 ( .C1(n9701), .C2(n9700), .A(n9699), .B(n9698), .ZN(n9705)
         );
  NAND2_X1 U10958 ( .A1(n9733), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n9704) );
  INV_X1 U10959 ( .A(n9702), .ZN(n9703) );
  NAND4_X1 U10960 ( .A1(n9706), .A2(n9705), .A3(n9704), .A4(n9703), .ZN(
        P1_U3246) );
  AOI21_X1 U10961 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9711), .A(n9707), .ZN(
        n9709) );
  XNOR2_X1 U10962 ( .A(n9728), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9708) );
  NOR2_X1 U10963 ( .A1(n9709), .A2(n9708), .ZN(n9727) );
  AOI211_X1 U10964 ( .C1(n9709), .C2(n9708), .A(n9727), .B(n9746), .ZN(n9719)
         );
  XNOR2_X1 U10965 ( .A(n9728), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9712) );
  NOR2_X1 U10966 ( .A1(n9713), .A2(n9712), .ZN(n9721) );
  AOI211_X1 U10967 ( .C1(n9713), .C2(n9712), .A(n9721), .B(n9745), .ZN(n9718)
         );
  NAND2_X1 U10968 ( .A1(n9733), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9715) );
  OAI211_X1 U10969 ( .C1(n9741), .C2(n9716), .A(n9715), .B(n9714), .ZN(n9717)
         );
  OR3_X1 U10970 ( .A1(n9719), .A2(n9718), .A3(n9717), .ZN(P1_U3258) );
  XNOR2_X1 U10971 ( .A(n9739), .B(n9720), .ZN(n9723) );
  AOI21_X1 U10972 ( .B1(n9728), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9721), .ZN(
        n9722) );
  NAND2_X1 U10973 ( .A1(n9723), .A2(n9722), .ZN(n9736) );
  OAI21_X1 U10974 ( .B1(n9723), .B2(n9722), .A(n9736), .ZN(n9724) );
  INV_X1 U10975 ( .A(n9724), .ZN(n9735) );
  INV_X1 U10976 ( .A(n9739), .ZN(n9726) );
  OAI21_X1 U10977 ( .B1(n9726), .B2(n9741), .A(n9725), .ZN(n9732) );
  MUX2_X1 U10978 ( .A(n7969), .B(P1_REG2_REG_18__SCAN_IN), .S(n9739), .Z(n9730) );
  AOI211_X1 U10979 ( .C1(n9730), .C2(n9729), .A(n9738), .B(n9746), .ZN(n9731)
         );
  AOI211_X1 U10980 ( .C1(n9733), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9732), .B(
        n9731), .ZN(n9734) );
  OAI21_X1 U10981 ( .B1(n9735), .B2(n9745), .A(n9734), .ZN(P1_U3259) );
  NAND2_X1 U10982 ( .A1(n9747), .A2(n9740), .ZN(n9742) );
  OAI211_X1 U10983 ( .C1(n9743), .C2(n9745), .A(n9742), .B(n9741), .ZN(n9749)
         );
  INV_X1 U10984 ( .A(n9743), .ZN(n9744) );
  OAI22_X1 U10985 ( .A1(n9747), .A2(n9746), .B1(n9745), .B2(n9744), .ZN(n9748)
         );
  NOR2_X1 U10986 ( .A1(n9775), .A2(n10067), .ZN(n9752) );
  XNOR2_X1 U10987 ( .A(n9756), .B(n9752), .ZN(n10065) );
  NAND2_X1 U10988 ( .A1(n10062), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9755) );
  NAND2_X1 U10989 ( .A1(n10239), .A2(P1_B_REG_SCAN_IN), .ZN(n9753) );
  NAND2_X1 U10990 ( .A1(n10043), .A2(n9753), .ZN(n9770) );
  NOR2_X1 U10991 ( .A1(n9770), .A2(n9754), .ZN(n10066) );
  NAND2_X1 U10992 ( .A1(n10066), .A2(n9940), .ZN(n9759) );
  OAI211_X1 U10993 ( .C1(n9756), .C2(n10054), .A(n9755), .B(n9759), .ZN(n9757)
         );
  INV_X1 U10994 ( .A(n9757), .ZN(n9758) );
  OAI21_X1 U10995 ( .B1(n10065), .B2(n9923), .A(n9758), .ZN(P1_U3261) );
  XNOR2_X1 U10996 ( .A(n9775), .B(n10067), .ZN(n10069) );
  INV_X1 U10997 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9760) );
  OAI21_X1 U10998 ( .B1(n9940), .B2(n9760), .A(n9759), .ZN(n9761) );
  AOI21_X1 U10999 ( .B1(n10067), .B2(n9920), .A(n9761), .ZN(n9762) );
  OAI21_X1 U11000 ( .B1(n10069), .B2(n9923), .A(n9762), .ZN(P1_U3262) );
  NOR2_X1 U11001 ( .A1(n10072), .A2(n10074), .ZN(n9763) );
  XNOR2_X1 U11002 ( .A(n9763), .B(n10071), .ZN(n9783) );
  AOI21_X2 U11003 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9767) );
  XNOR2_X1 U11004 ( .A(n9767), .B(n10076), .ZN(n9773) );
  OAI21_X1 U11005 ( .B1(n9773), .B2(n10045), .A(n9772), .ZN(n10070) );
  AOI21_X1 U11006 ( .B1(n10077), .B2(n9774), .A(n10287), .ZN(n9776) );
  OAI22_X1 U11007 ( .A1(n9778), .A2(n9898), .B1(n9777), .B2(n9940), .ZN(n9779)
         );
  AOI21_X1 U11008 ( .B1(n10077), .B2(n9920), .A(n9779), .ZN(n9780) );
  OAI21_X1 U11009 ( .B1(n10081), .B2(n9903), .A(n9780), .ZN(n9781) );
  AOI21_X1 U11010 ( .B1(n10070), .B2(n9940), .A(n9781), .ZN(n9782) );
  OAI21_X1 U11011 ( .B1(n9783), .B2(n10028), .A(n9782), .ZN(P1_U3355) );
  INV_X1 U11012 ( .A(n9813), .ZN(n9792) );
  INV_X1 U11013 ( .A(n9790), .ZN(n9791) );
  AOI21_X1 U11014 ( .B1(n10089), .B2(n9792), .A(n9791), .ZN(n10090) );
  INV_X1 U11015 ( .A(n9793), .ZN(n9794) );
  AOI22_X1 U11016 ( .A1(n9794), .A2(n10051), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10062), .ZN(n9795) );
  OAI21_X1 U11017 ( .B1(n9796), .B2(n10054), .A(n9795), .ZN(n9802) );
  OAI21_X1 U11018 ( .B1(n9799), .B2(n9798), .A(n9797), .ZN(n9800) );
  INV_X1 U11019 ( .A(n9800), .ZN(n10093) );
  NOR2_X1 U11020 ( .A1(n10093), .A2(n10028), .ZN(n9801) );
  AOI211_X1 U11021 ( .C1(n10090), .C2(n10060), .A(n9802), .B(n9801), .ZN(n9803) );
  OAI21_X1 U11022 ( .B1(n10092), .B2(n10062), .A(n9803), .ZN(P1_U3264) );
  INV_X1 U11023 ( .A(n9804), .ZN(n9805) );
  AOI21_X1 U11024 ( .B1(n10094), .B2(n9833), .A(n9813), .ZN(n10095) );
  AOI22_X1 U11025 ( .A1(n9814), .A2(n10051), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10062), .ZN(n9815) );
  OAI21_X1 U11026 ( .B1(n4568), .B2(n10054), .A(n9815), .ZN(n9825) );
  NAND2_X1 U11027 ( .A1(n9816), .A2(n9817), .ZN(n9819) );
  NAND2_X1 U11028 ( .A1(n9819), .A2(n9818), .ZN(n9822) );
  OAI21_X1 U11029 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9823) );
  INV_X1 U11030 ( .A(n9823), .ZN(n10098) );
  NOR2_X1 U11031 ( .A1(n10098), .A2(n10028), .ZN(n9824) );
  AOI211_X1 U11032 ( .C1(n10095), .C2(n10060), .A(n9825), .B(n9824), .ZN(n9826) );
  OAI21_X1 U11033 ( .B1(n10097), .B2(n10062), .A(n9826), .ZN(P1_U3265) );
  AOI21_X2 U11034 ( .B1(n9832), .B2(n4705), .A(n9831), .ZN(n10102) );
  INV_X1 U11035 ( .A(n9855), .ZN(n9835) );
  INV_X1 U11036 ( .A(n9833), .ZN(n9834) );
  AOI21_X1 U11037 ( .B1(n10099), .B2(n9835), .A(n9834), .ZN(n10100) );
  INV_X1 U11038 ( .A(n9836), .ZN(n9837) );
  AOI22_X1 U11039 ( .A1(n9837), .A2(n10051), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10062), .ZN(n9838) );
  OAI21_X1 U11040 ( .B1(n9839), .B2(n10054), .A(n9838), .ZN(n9844) );
  NAND2_X1 U11041 ( .A1(n9816), .A2(n9840), .ZN(n9841) );
  XOR2_X1 U11042 ( .A(n9842), .B(n9841), .Z(n10103) );
  NOR2_X1 U11043 ( .A1(n10103), .A2(n10028), .ZN(n9843) );
  AOI211_X1 U11044 ( .C1(n10100), .C2(n10060), .A(n9844), .B(n9843), .ZN(n9845) );
  OAI21_X1 U11045 ( .B1(n10102), .B2(n10062), .A(n9845), .ZN(P1_U3266) );
  OR2_X1 U11046 ( .A1(n9871), .A2(n9846), .ZN(n9848) );
  NAND2_X1 U11047 ( .A1(n9848), .A2(n9847), .ZN(n9849) );
  XNOR2_X1 U11048 ( .A(n9849), .B(n9851), .ZN(n10107) );
  OAI21_X1 U11049 ( .B1(n9854), .B2(n9866), .A(n10181), .ZN(n9856) );
  NOR2_X1 U11050 ( .A1(n9856), .A2(n9855), .ZN(n10105) );
  NAND2_X1 U11051 ( .A1(n10105), .A2(n9857), .ZN(n9858) );
  OAI21_X1 U11052 ( .B1(n9898), .B2(n9859), .A(n9858), .ZN(n9860) );
  OAI21_X1 U11053 ( .B1(n10104), .B2(n9860), .A(n9940), .ZN(n9862) );
  AOI22_X1 U11054 ( .A1(n10106), .A2(n9920), .B1(n10062), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9861) );
  OAI211_X1 U11055 ( .C1(n10107), .C2(n10028), .A(n9862), .B(n9861), .ZN(
        P1_U3267) );
  XNOR2_X1 U11056 ( .A(n9863), .B(n9870), .ZN(n9865) );
  AOI222_X1 U11057 ( .A1(n4705), .A2(n9865), .B1(n9864), .B2(n10043), .C1(
        n9894), .C2(n10041), .ZN(n10111) );
  AOI211_X1 U11058 ( .C1(n10109), .C2(n9879), .A(n10287), .B(n9866), .ZN(
        n10108) );
  AOI22_X1 U11059 ( .A1(n9867), .A2(n10051), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10062), .ZN(n9868) );
  OAI21_X1 U11060 ( .B1(n9869), .B2(n10054), .A(n9868), .ZN(n9873) );
  XNOR2_X1 U11061 ( .A(n9871), .B(n9870), .ZN(n10112) );
  NOR2_X1 U11062 ( .A1(n10112), .A2(n10028), .ZN(n9872) );
  AOI211_X1 U11063 ( .C1(n10108), .C2(n10031), .A(n9873), .B(n9872), .ZN(n9874) );
  OAI21_X1 U11064 ( .B1(n10111), .B2(n10062), .A(n9874), .ZN(P1_U3268) );
  XNOR2_X1 U11065 ( .A(n9875), .B(n9884), .ZN(n9878) );
  AOI222_X1 U11066 ( .A1(n4705), .A2(n9878), .B1(n9877), .B2(n10043), .C1(
        n9876), .C2(n10041), .ZN(n10116) );
  INV_X1 U11067 ( .A(n9901), .ZN(n9880) );
  AOI21_X1 U11068 ( .B1(n10113), .B2(n9880), .A(n5035), .ZN(n10114) );
  AOI22_X1 U11069 ( .A1(n9881), .A2(n10051), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10062), .ZN(n9882) );
  OAI21_X1 U11070 ( .B1(n9883), .B2(n10054), .A(n9882), .ZN(n9887) );
  XNOR2_X1 U11071 ( .A(n9885), .B(n9884), .ZN(n10117) );
  NOR2_X1 U11072 ( .A1(n10117), .A2(n10028), .ZN(n9886) );
  AOI211_X1 U11073 ( .C1(n10114), .C2(n10060), .A(n9887), .B(n9886), .ZN(n9888) );
  OAI21_X1 U11074 ( .B1(n10116), .B2(n10062), .A(n9888), .ZN(P1_U3269) );
  XNOR2_X1 U11075 ( .A(n9890), .B(n9889), .ZN(n10121) );
  XNOR2_X1 U11076 ( .A(n9892), .B(n9891), .ZN(n9893) );
  NAND2_X1 U11077 ( .A1(n9893), .A2(n4705), .ZN(n9896) );
  AOI22_X1 U11078 ( .A1(n9894), .A2(n10043), .B1(n9931), .B2(n10041), .ZN(
        n9895) );
  NAND2_X1 U11079 ( .A1(n9896), .A2(n9895), .ZN(n10123) );
  NAND2_X1 U11080 ( .A1(n10123), .A2(n9940), .ZN(n9907) );
  INV_X1 U11081 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9897) );
  OAI22_X1 U11082 ( .A1(n9899), .A2(n9898), .B1(n9897), .B2(n9940), .ZN(n9905)
         );
  NAND2_X1 U11083 ( .A1(n10118), .A2(n9917), .ZN(n9900) );
  NAND2_X1 U11084 ( .A1(n9900), .A2(n10181), .ZN(n9902) );
  OR2_X1 U11085 ( .A1(n9902), .A2(n9901), .ZN(n10119) );
  NOR2_X1 U11086 ( .A1(n10119), .A2(n9903), .ZN(n9904) );
  AOI211_X1 U11087 ( .C1(n9920), .C2(n10118), .A(n9905), .B(n9904), .ZN(n9906)
         );
  OAI211_X1 U11088 ( .C1(n10121), .C2(n10028), .A(n9907), .B(n9906), .ZN(
        P1_U3270) );
  XNOR2_X1 U11089 ( .A(n9908), .B(n9913), .ZN(n9912) );
  OAI22_X1 U11090 ( .A1(n9910), .A2(n10017), .B1(n9909), .B2(n10014), .ZN(
        n9911) );
  AOI21_X1 U11091 ( .B1(n9912), .B2(n4705), .A(n9911), .ZN(n10130) );
  INV_X1 U11092 ( .A(n9913), .ZN(n9914) );
  XNOR2_X1 U11093 ( .A(n9915), .B(n9914), .ZN(n10128) );
  NAND2_X1 U11094 ( .A1(n10124), .A2(n9934), .ZN(n9916) );
  NAND2_X1 U11095 ( .A1(n9917), .A2(n9916), .ZN(n10126) );
  INV_X1 U11096 ( .A(n9918), .ZN(n9919) );
  AOI22_X1 U11097 ( .A1(n9919), .A2(n10051), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n10062), .ZN(n9922) );
  NAND2_X1 U11098 ( .A1(n10124), .A2(n9920), .ZN(n9921) );
  OAI211_X1 U11099 ( .C1(n10126), .C2(n9923), .A(n9922), .B(n9921), .ZN(n9924)
         );
  AOI21_X1 U11100 ( .B1(n10128), .B2(n9925), .A(n9924), .ZN(n9926) );
  OAI21_X1 U11101 ( .B1(n10130), .B2(n10062), .A(n9926), .ZN(P1_U3271) );
  XOR2_X1 U11102 ( .A(n9927), .B(n9930), .Z(n10137) );
  OAI21_X1 U11103 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(n9932) );
  AOI222_X1 U11104 ( .A1(n4705), .A2(n9932), .B1(n9931), .B2(n10043), .C1(
        n9962), .C2(n10041), .ZN(n10136) );
  INV_X1 U11105 ( .A(n10136), .ZN(n9941) );
  INV_X1 U11106 ( .A(n10133), .ZN(n9938) );
  NAND2_X1 U11107 ( .A1(n9949), .A2(n10133), .ZN(n9933) );
  AND2_X1 U11108 ( .A1(n9934), .A2(n9933), .ZN(n10134) );
  NAND2_X1 U11109 ( .A1(n10134), .A2(n10060), .ZN(n9937) );
  AOI22_X1 U11110 ( .A1(n9935), .A2(n10051), .B1(n10062), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9936) );
  OAI211_X1 U11111 ( .C1(n9938), .C2(n10054), .A(n9937), .B(n9936), .ZN(n9939)
         );
  AOI21_X1 U11112 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n9942) );
  OAI21_X1 U11113 ( .B1(n10028), .B2(n10137), .A(n9942), .ZN(P1_U3272) );
  INV_X1 U11114 ( .A(n9943), .ZN(n9944) );
  AOI21_X1 U11115 ( .B1(n9961), .B2(n9945), .A(n9944), .ZN(n9946) );
  XOR2_X1 U11116 ( .A(n9956), .B(n9946), .Z(n9948) );
  AOI222_X1 U11117 ( .A1(n4705), .A2(n9948), .B1(n9947), .B2(n10043), .C1(
        n9979), .C2(n10041), .ZN(n10141) );
  INV_X1 U11118 ( .A(n9964), .ZN(n9951) );
  INV_X1 U11119 ( .A(n9949), .ZN(n9950) );
  AOI21_X1 U11120 ( .B1(n10138), .B2(n9951), .A(n9950), .ZN(n10139) );
  INV_X1 U11121 ( .A(n9952), .ZN(n9953) );
  AOI22_X1 U11122 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n10062), .B1(n9953), 
        .B2(n10051), .ZN(n9954) );
  OAI21_X1 U11123 ( .B1(n9955), .B2(n10054), .A(n9954), .ZN(n9959) );
  XNOR2_X1 U11124 ( .A(n9957), .B(n9956), .ZN(n10142) );
  NOR2_X1 U11125 ( .A1(n10142), .A2(n10028), .ZN(n9958) );
  AOI211_X1 U11126 ( .C1(n10139), .C2(n10060), .A(n9959), .B(n9958), .ZN(n9960) );
  OAI21_X1 U11127 ( .B1(n10141), .B2(n10062), .A(n9960), .ZN(P1_U3273) );
  XOR2_X1 U11128 ( .A(n9961), .B(n9969), .Z(n9963) );
  AOI222_X1 U11129 ( .A1(n4705), .A2(n9963), .B1(n9962), .B2(n10043), .C1(
        n9998), .C2(n10041), .ZN(n10146) );
  INV_X1 U11130 ( .A(n9981), .ZN(n9965) );
  AOI211_X1 U11131 ( .C1(n10144), .C2(n9965), .A(n10287), .B(n9964), .ZN(
        n10143) );
  AOI22_X1 U11132 ( .A1(n10062), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9966), 
        .B2(n10051), .ZN(n9967) );
  OAI21_X1 U11133 ( .B1(n9968), .B2(n10054), .A(n9967), .ZN(n9972) );
  XOR2_X1 U11134 ( .A(n9970), .B(n9969), .Z(n10147) );
  NOR2_X1 U11135 ( .A1(n10147), .A2(n10028), .ZN(n9971) );
  AOI211_X1 U11136 ( .C1(n10143), .C2(n10031), .A(n9972), .B(n9971), .ZN(n9973) );
  OAI21_X1 U11137 ( .B1(n10146), .B2(n10062), .A(n9973), .ZN(P1_U3274) );
  NAND2_X1 U11138 ( .A1(n9974), .A2(n9975), .ZN(n9977) );
  XNOR2_X1 U11139 ( .A(n9977), .B(n9976), .ZN(n9980) );
  AOI222_X1 U11140 ( .A1(n4705), .A2(n9980), .B1(n9979), .B2(n10043), .C1(
        n9978), .C2(n10041), .ZN(n10151) );
  AOI211_X1 U11141 ( .C1(n10149), .C2(n10003), .A(n10287), .B(n9981), .ZN(
        n10148) );
  INV_X1 U11142 ( .A(n9982), .ZN(n9983) );
  AOI22_X1 U11143 ( .A1(n10062), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9983), 
        .B2(n10051), .ZN(n9984) );
  OAI21_X1 U11144 ( .B1(n9985), .B2(n10054), .A(n9984), .ZN(n9991) );
  OR2_X1 U11145 ( .A1(n9987), .A2(n9986), .ZN(n9988) );
  NAND2_X1 U11146 ( .A1(n9989), .A2(n9988), .ZN(n10152) );
  NOR2_X1 U11147 ( .A1(n10152), .A2(n10028), .ZN(n9990) );
  AOI211_X1 U11148 ( .C1(n10148), .C2(n10031), .A(n9991), .B(n9990), .ZN(n9992) );
  OAI21_X1 U11149 ( .B1(n10151), .B2(n10062), .A(n9992), .ZN(P1_U3275) );
  OAI21_X1 U11150 ( .B1(n9994), .B2(n9993), .A(n9974), .ZN(n10002) );
  NAND2_X1 U11151 ( .A1(n9995), .A2(n9994), .ZN(n9996) );
  NAND2_X1 U11152 ( .A1(n9997), .A2(n9996), .ZN(n10157) );
  AOI22_X1 U11153 ( .A1(n9998), .A2(n10043), .B1(n10041), .B2(n10042), .ZN(
        n9999) );
  OAI21_X1 U11154 ( .B1(n10157), .B2(n10000), .A(n9999), .ZN(n10001) );
  AOI21_X1 U11155 ( .B1(n10002), .B2(n4705), .A(n10001), .ZN(n10156) );
  AOI211_X1 U11156 ( .C1(n10154), .C2(n10020), .A(n10287), .B(n5045), .ZN(
        n10153) );
  AOI22_X1 U11157 ( .A1(n10062), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10004), 
        .B2(n10051), .ZN(n10005) );
  OAI21_X1 U11158 ( .B1(n10006), .B2(n10054), .A(n10005), .ZN(n10008) );
  NOR2_X1 U11159 ( .A1(n10157), .A2(n10057), .ZN(n10007) );
  AOI211_X1 U11160 ( .C1(n10153), .C2(n10031), .A(n10008), .B(n10007), .ZN(
        n10009) );
  OAI21_X1 U11161 ( .B1(n10062), .B2(n10156), .A(n10009), .ZN(P1_U3276) );
  NAND2_X1 U11162 ( .A1(n10036), .A2(n10010), .ZN(n10013) );
  INV_X1 U11163 ( .A(n10011), .ZN(n10012) );
  AOI211_X1 U11164 ( .C1(n10026), .C2(n10013), .A(n10045), .B(n10012), .ZN(
        n10019) );
  OAI22_X1 U11165 ( .A1(n10017), .A2(n10016), .B1(n10015), .B2(n10014), .ZN(
        n10018) );
  NOR2_X1 U11166 ( .A1(n10019), .A2(n10018), .ZN(n10161) );
  INV_X1 U11167 ( .A(n10050), .ZN(n10021) );
  AOI211_X1 U11168 ( .C1(n10159), .C2(n10021), .A(n10287), .B(n5042), .ZN(
        n10158) );
  INV_X1 U11169 ( .A(n10022), .ZN(n10023) );
  AOI22_X1 U11170 ( .A1(n10062), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n10023), 
        .B2(n10051), .ZN(n10024) );
  OAI21_X1 U11171 ( .B1(n10025), .B2(n10054), .A(n10024), .ZN(n10030) );
  XNOR2_X1 U11172 ( .A(n10027), .B(n10026), .ZN(n10162) );
  NOR2_X1 U11173 ( .A1(n10162), .A2(n10028), .ZN(n10029) );
  AOI211_X1 U11174 ( .C1(n10158), .C2(n10031), .A(n10030), .B(n10029), .ZN(
        n10032) );
  OAI21_X1 U11175 ( .B1(n10161), .B2(n10062), .A(n10032), .ZN(P1_U3277) );
  NAND2_X1 U11176 ( .A1(n10034), .A2(n10033), .ZN(n10035) );
  XNOR2_X1 U11177 ( .A(n10035), .B(n5705), .ZN(n10056) );
  INV_X1 U11178 ( .A(n10036), .ZN(n10037) );
  AOI21_X1 U11179 ( .B1(n10039), .B2(n10038), .A(n10037), .ZN(n10046) );
  AOI22_X1 U11180 ( .A1(n10043), .A2(n10042), .B1(n10041), .B2(n10040), .ZN(
        n10044) );
  OAI21_X1 U11181 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(n10047) );
  AOI21_X1 U11182 ( .B1(n10048), .B2(n10056), .A(n10047), .ZN(n10167) );
  AOI21_X1 U11183 ( .B1(n10164), .B2(n5031), .A(n10050), .ZN(n10165) );
  AOI22_X1 U11184 ( .A1(n10062), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10052), 
        .B2(n10051), .ZN(n10053) );
  OAI21_X1 U11185 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(n10059) );
  INV_X1 U11186 ( .A(n10056), .ZN(n10168) );
  NOR2_X1 U11187 ( .A1(n10168), .A2(n10057), .ZN(n10058) );
  AOI211_X1 U11188 ( .C1(n10165), .C2(n10060), .A(n10059), .B(n10058), .ZN(
        n10061) );
  OAI21_X1 U11189 ( .B1(n10167), .B2(n10062), .A(n10061), .ZN(P1_U3278) );
  AOI21_X1 U11190 ( .B1(n10063), .B2(n10180), .A(n10066), .ZN(n10064) );
  OAI21_X1 U11191 ( .B1(n10065), .B2(n10287), .A(n10064), .ZN(n10188) );
  MUX2_X1 U11192 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10188), .S(n10308), .Z(
        P1_U3554) );
  AOI21_X1 U11193 ( .B1(n10067), .B2(n10180), .A(n10066), .ZN(n10068) );
  OAI21_X1 U11194 ( .B1(n10069), .B2(n10287), .A(n10068), .ZN(n10189) );
  MUX2_X1 U11195 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10189), .S(n10308), .Z(
        P1_U3553) );
  INV_X1 U11196 ( .A(n10070), .ZN(n10083) );
  INV_X1 U11197 ( .A(n10074), .ZN(n10075) );
  INV_X1 U11198 ( .A(n10077), .ZN(n10078) );
  MUX2_X1 U11199 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10190), .S(n10308), .Z(
        P1_U3552) );
  AOI21_X1 U11200 ( .B1(n10180), .B2(n10085), .A(n10084), .ZN(n10086) );
  OAI211_X1 U11201 ( .C1(n10163), .C2(n10088), .A(n10087), .B(n10086), .ZN(
        n10191) );
  MUX2_X1 U11202 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10191), .S(n10308), .Z(
        P1_U3551) );
  AOI22_X1 U11203 ( .A1(n10090), .A2(n10181), .B1(n10180), .B2(n10089), .ZN(
        n10091) );
  OAI211_X1 U11204 ( .C1(n10163), .C2(n10093), .A(n10092), .B(n10091), .ZN(
        n10192) );
  MUX2_X1 U11205 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10192), .S(n10308), .Z(
        P1_U3550) );
  AOI22_X1 U11206 ( .A1(n10095), .A2(n10181), .B1(n10180), .B2(n10094), .ZN(
        n10096) );
  MUX2_X1 U11207 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10193), .S(n10308), .Z(
        P1_U3549) );
  AOI22_X1 U11208 ( .A1(n10100), .A2(n10181), .B1(n10180), .B2(n10099), .ZN(
        n10101) );
  OAI211_X1 U11209 ( .C1(n10163), .C2(n10103), .A(n10102), .B(n10101), .ZN(
        n10194) );
  MUX2_X1 U11210 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10194), .S(n10308), .Z(
        P1_U3548) );
  MUX2_X1 U11211 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10195), .S(n10308), .Z(
        P1_U3547) );
  AOI21_X1 U11212 ( .B1(n10180), .B2(n10109), .A(n10108), .ZN(n10110) );
  OAI211_X1 U11213 ( .C1(n10163), .C2(n10112), .A(n10111), .B(n10110), .ZN(
        n10196) );
  MUX2_X1 U11214 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10196), .S(n10308), .Z(
        P1_U3546) );
  AOI22_X1 U11215 ( .A1(n10114), .A2(n10181), .B1(n10180), .B2(n10113), .ZN(
        n10115) );
  OAI211_X1 U11216 ( .C1(n10163), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        n10197) );
  MUX2_X1 U11217 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10197), .S(n10308), .Z(
        P1_U3545) );
  NAND2_X1 U11218 ( .A1(n10118), .A2(n10180), .ZN(n10120) );
  OAI211_X1 U11219 ( .C1(n10121), .C2(n10163), .A(n10120), .B(n10119), .ZN(
        n10122) );
  MUX2_X1 U11220 ( .A(n10198), .B(P1_REG1_REG_21__SCAN_IN), .S(n10306), .Z(
        P1_U3544) );
  INV_X1 U11221 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10131) );
  INV_X1 U11222 ( .A(n10124), .ZN(n10125) );
  OAI22_X1 U11223 ( .A1(n10126), .A2(n10287), .B1(n10125), .B2(n10295), .ZN(
        n10127) );
  AOI21_X1 U11224 ( .B1(n10128), .B2(n4976), .A(n10127), .ZN(n10129) );
  AND2_X1 U11225 ( .A1(n10130), .A2(n10129), .ZN(n10199) );
  MUX2_X1 U11226 ( .A(n10131), .B(n10199), .S(n10308), .Z(n10132) );
  INV_X1 U11227 ( .A(n10132), .ZN(P1_U3543) );
  AOI22_X1 U11228 ( .A1(n10134), .A2(n10181), .B1(n10180), .B2(n10133), .ZN(
        n10135) );
  OAI211_X1 U11229 ( .C1(n10163), .C2(n10137), .A(n10136), .B(n10135), .ZN(
        n10202) );
  MUX2_X1 U11230 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10202), .S(n10308), .Z(
        P1_U3542) );
  AOI22_X1 U11231 ( .A1(n10139), .A2(n10181), .B1(n10180), .B2(n10138), .ZN(
        n10140) );
  OAI211_X1 U11232 ( .C1(n10163), .C2(n10142), .A(n10141), .B(n10140), .ZN(
        n10203) );
  MUX2_X1 U11233 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10203), .S(n10308), .Z(
        P1_U3541) );
  AOI21_X1 U11234 ( .B1(n10180), .B2(n10144), .A(n10143), .ZN(n10145) );
  OAI211_X1 U11235 ( .C1(n10163), .C2(n10147), .A(n10146), .B(n10145), .ZN(
        n10204) );
  MUX2_X1 U11236 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10204), .S(n10308), .Z(
        P1_U3540) );
  AOI21_X1 U11237 ( .B1(n10180), .B2(n10149), .A(n10148), .ZN(n10150) );
  OAI211_X1 U11238 ( .C1(n10163), .C2(n10152), .A(n10151), .B(n10150), .ZN(
        n10205) );
  MUX2_X1 U11239 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10205), .S(n10308), .Z(
        P1_U3539) );
  AOI21_X1 U11240 ( .B1(n10180), .B2(n10154), .A(n10153), .ZN(n10155) );
  OAI211_X1 U11241 ( .C1(n10186), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        n10206) );
  MUX2_X1 U11242 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10206), .S(n10308), .Z(
        P1_U3538) );
  AOI21_X1 U11243 ( .B1(n10180), .B2(n10159), .A(n10158), .ZN(n10160) );
  OAI211_X1 U11244 ( .C1(n10163), .C2(n10162), .A(n10161), .B(n10160), .ZN(
        n10207) );
  MUX2_X1 U11245 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10207), .S(n10308), .Z(
        P1_U3537) );
  AOI22_X1 U11246 ( .A1(n10165), .A2(n10181), .B1(n10180), .B2(n10164), .ZN(
        n10166) );
  OAI211_X1 U11247 ( .C1(n10186), .C2(n10168), .A(n10167), .B(n10166), .ZN(
        n10208) );
  MUX2_X1 U11248 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10208), .S(n10308), .Z(
        P1_U3536) );
  AOI21_X1 U11249 ( .B1(n10180), .B2(n10170), .A(n10169), .ZN(n10171) );
  OAI211_X1 U11250 ( .C1(n10186), .C2(n10173), .A(n10172), .B(n10171), .ZN(
        n10209) );
  MUX2_X1 U11251 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10209), .S(n10308), .Z(
        P1_U3535) );
  AOI22_X1 U11252 ( .A1(n10175), .A2(n10181), .B1(n10180), .B2(n10174), .ZN(
        n10176) );
  OAI211_X1 U11253 ( .C1(n10186), .C2(n10178), .A(n10177), .B(n10176), .ZN(
        n10210) );
  MUX2_X1 U11254 ( .A(n10210), .B(P1_REG1_REG_9__SCAN_IN), .S(n10306), .Z(
        P1_U3532) );
  AOI22_X1 U11255 ( .A1(n10182), .A2(n10181), .B1(n10180), .B2(n10179), .ZN(
        n10183) );
  OAI211_X1 U11256 ( .C1(n10186), .C2(n10185), .A(n10184), .B(n10183), .ZN(
        n10211) );
  MUX2_X1 U11257 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10211), .S(n10308), .Z(
        P1_U3531) );
  MUX2_X1 U11258 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10187), .S(n10308), .Z(
        P1_U3523) );
  MUX2_X1 U11259 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10188), .S(n10301), .Z(
        P1_U3522) );
  MUX2_X1 U11260 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10189), .S(n10301), .Z(
        P1_U3521) );
  MUX2_X1 U11261 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10190), .S(n10301), .Z(
        P1_U3520) );
  MUX2_X1 U11262 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10191), .S(n10301), .Z(
        P1_U3519) );
  MUX2_X1 U11263 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10192), .S(n10301), .Z(
        P1_U3518) );
  MUX2_X1 U11264 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10193), .S(n10301), .Z(
        P1_U3517) );
  MUX2_X1 U11265 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10194), .S(n10301), .Z(
        P1_U3516) );
  MUX2_X1 U11266 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10195), .S(n10301), .Z(
        P1_U3515) );
  MUX2_X1 U11267 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10196), .S(n10301), .Z(
        P1_U3514) );
  MUX2_X1 U11268 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10197), .S(n10301), .Z(
        P1_U3513) );
  MUX2_X1 U11269 ( .A(n10198), .B(P1_REG0_REG_21__SCAN_IN), .S(n10299), .Z(
        P1_U3512) );
  MUX2_X1 U11270 ( .A(n10200), .B(n10199), .S(n10301), .Z(n10201) );
  INV_X1 U11271 ( .A(n10201), .ZN(P1_U3511) );
  MUX2_X1 U11272 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10202), .S(n10301), .Z(
        P1_U3510) );
  MUX2_X1 U11273 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10203), .S(n10301), .Z(
        P1_U3508) );
  MUX2_X1 U11274 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10204), .S(n10301), .Z(
        P1_U3505) );
  MUX2_X1 U11275 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10205), .S(n10301), .Z(
        P1_U3502) );
  MUX2_X1 U11276 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10206), .S(n10301), .Z(
        P1_U3499) );
  MUX2_X1 U11277 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10207), .S(n10301), .Z(
        P1_U3496) );
  MUX2_X1 U11278 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10208), .S(n10301), .Z(
        P1_U3493) );
  MUX2_X1 U11279 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10209), .S(n10301), .Z(
        P1_U3490) );
  MUX2_X1 U11280 ( .A(n10210), .B(P1_REG0_REG_9__SCAN_IN), .S(n10299), .Z(
        P1_U3481) );
  MUX2_X1 U11281 ( .A(P1_REG0_REG_8__SCAN_IN), .B(n10211), .S(n10301), .Z(
        P1_U3478) );
  MUX2_X1 U11282 ( .A(P1_D_REG_0__SCAN_IN), .B(n10214), .S(n10279), .Z(
        P1_U3440) );
  NOR4_X1 U11283 ( .A1(n10216), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n10215), .ZN(n10217) );
  AOI21_X1 U11284 ( .B1(n10230), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10217), 
        .ZN(n10218) );
  OAI21_X1 U11285 ( .B1(n10219), .B2(n10232), .A(n10218), .ZN(P1_U3322) );
  AOI22_X1 U11286 ( .A1(n10220), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10230), .ZN(n10221) );
  OAI21_X1 U11287 ( .B1(n10222), .B2(n10232), .A(n10221), .ZN(P1_U3323) );
  AOI22_X1 U11288 ( .A1(n10223), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10230), .ZN(n10224) );
  OAI21_X1 U11289 ( .B1(n10225), .B2(n10232), .A(n10224), .ZN(P1_U3324) );
  AOI22_X1 U11290 ( .A1(n10226), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10230), .ZN(n10227) );
  OAI21_X1 U11291 ( .B1(n10228), .B2(n10232), .A(n10227), .ZN(P1_U3325) );
  AOI21_X1 U11292 ( .B1(n10230), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n10229), 
        .ZN(n10231) );
  OAI21_X1 U11293 ( .B1(n10233), .B2(n10232), .A(n10231), .ZN(P1_U3326) );
  INV_X1 U11294 ( .A(n10234), .ZN(n10235) );
  MUX2_X1 U11295 ( .A(n10235), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  XNOR2_X1 U11296 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U11297 ( .A(n10236), .B(P2_RD_REG_SCAN_IN), .Z(U126) );
  INV_X1 U11298 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10244) );
  INV_X1 U11299 ( .A(n10237), .ZN(n10238) );
  OAI21_X1 U11300 ( .B1(n10239), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10238), .ZN(
        n10241) );
  XNOR2_X1 U11301 ( .A(n10241), .B(n10240), .ZN(n10242) );
  OAI22_X1 U11302 ( .A1(n10245), .A2(n10244), .B1(n10243), .B2(n10242), .ZN(
        n10246) );
  INV_X1 U11303 ( .A(n10246), .ZN(n10247) );
  OAI21_X1 U11304 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n8211), .A(n10247), .ZN(
        P1_U3241) );
  INV_X1 U11305 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10248) );
  NOR2_X1 U11306 ( .A1(n10265), .A2(n10248), .ZN(P1_U3292) );
  INV_X1 U11307 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10249) );
  NOR2_X1 U11308 ( .A1(n10265), .A2(n10249), .ZN(P1_U3293) );
  NOR2_X1 U11309 ( .A1(n10279), .A2(n10250), .ZN(P1_U3294) );
  INV_X1 U11310 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10251) );
  NOR2_X1 U11311 ( .A1(n10279), .A2(n10251), .ZN(P1_U3295) );
  INV_X1 U11312 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10252) );
  NOR2_X1 U11313 ( .A1(n10279), .A2(n10252), .ZN(P1_U3296) );
  INV_X1 U11314 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10253) );
  NOR2_X1 U11315 ( .A1(n10279), .A2(n10253), .ZN(P1_U3297) );
  INV_X1 U11316 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10254) );
  NOR2_X1 U11317 ( .A1(n10279), .A2(n10254), .ZN(P1_U3298) );
  INV_X1 U11318 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10255) );
  NOR2_X1 U11319 ( .A1(n10279), .A2(n10255), .ZN(P1_U3299) );
  NOR2_X1 U11320 ( .A1(n10279), .A2(n10256), .ZN(P1_U3300) );
  INV_X1 U11321 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10257) );
  NOR2_X1 U11322 ( .A1(n10265), .A2(n10257), .ZN(P1_U3301) );
  NOR2_X1 U11323 ( .A1(n10265), .A2(n10258), .ZN(P1_U3302) );
  NOR2_X1 U11324 ( .A1(n10265), .A2(n10259), .ZN(P1_U3303) );
  NOR2_X1 U11325 ( .A1(n10265), .A2(n10260), .ZN(P1_U3304) );
  INV_X1 U11326 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10261) );
  NOR2_X1 U11327 ( .A1(n10265), .A2(n10261), .ZN(P1_U3305) );
  INV_X1 U11328 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10262) );
  NOR2_X1 U11329 ( .A1(n10265), .A2(n10262), .ZN(P1_U3306) );
  NOR2_X1 U11330 ( .A1(n10265), .A2(n10263), .ZN(P1_U3307) );
  NOR2_X1 U11331 ( .A1(n10265), .A2(n10264), .ZN(P1_U3308) );
  INV_X1 U11332 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10266) );
  NOR2_X1 U11333 ( .A1(n10279), .A2(n10266), .ZN(P1_U3309) );
  NOR2_X1 U11334 ( .A1(n10279), .A2(n10267), .ZN(P1_U3310) );
  INV_X1 U11335 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10268) );
  NOR2_X1 U11336 ( .A1(n10279), .A2(n10268), .ZN(P1_U3311) );
  INV_X1 U11337 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10269) );
  NOR2_X1 U11338 ( .A1(n10279), .A2(n10269), .ZN(P1_U3312) );
  INV_X1 U11339 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10270) );
  NOR2_X1 U11340 ( .A1(n10279), .A2(n10270), .ZN(P1_U3313) );
  INV_X1 U11341 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10271) );
  NOR2_X1 U11342 ( .A1(n10279), .A2(n10271), .ZN(P1_U3314) );
  NOR2_X1 U11343 ( .A1(n10279), .A2(n10272), .ZN(P1_U3315) );
  INV_X1 U11344 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10273) );
  NOR2_X1 U11345 ( .A1(n10279), .A2(n10273), .ZN(P1_U3316) );
  INV_X1 U11346 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U11347 ( .A1(n10279), .A2(n10274), .ZN(P1_U3317) );
  INV_X1 U11348 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10275) );
  NOR2_X1 U11349 ( .A1(n10279), .A2(n10275), .ZN(P1_U3318) );
  INV_X1 U11350 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10276) );
  NOR2_X1 U11351 ( .A1(n10279), .A2(n10276), .ZN(P1_U3319) );
  INV_X1 U11352 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10277) );
  NOR2_X1 U11353 ( .A1(n10279), .A2(n10277), .ZN(P1_U3320) );
  INV_X1 U11354 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10278) );
  NOR2_X1 U11355 ( .A1(n10279), .A2(n10278), .ZN(P1_U3321) );
  INV_X1 U11356 ( .A(n10280), .ZN(n10285) );
  OAI21_X1 U11357 ( .B1(n10282), .B2(n10295), .A(n10281), .ZN(n10284) );
  AOI211_X1 U11358 ( .C1(n10292), .C2(n10285), .A(n10284), .B(n10283), .ZN(
        n10303) );
  AOI22_X1 U11359 ( .A1(n10301), .A2(n10303), .B1(n5082), .B2(n10299), .ZN(
        P1_U3457) );
  OAI22_X1 U11360 ( .A1(n10288), .A2(n10287), .B1(n10286), .B2(n10295), .ZN(
        n10290) );
  AOI211_X1 U11361 ( .C1(n10292), .C2(n10291), .A(n10290), .B(n10289), .ZN(
        n10305) );
  INV_X1 U11362 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U11363 ( .A1(n10301), .A2(n10305), .B1(n10293), .B2(n10299), .ZN(
        P1_U3463) );
  OAI21_X1 U11364 ( .B1(n5026), .B2(n10295), .A(n10294), .ZN(n10297) );
  AOI211_X1 U11365 ( .C1(n4976), .C2(n10298), .A(n10297), .B(n10296), .ZN(
        n10307) );
  INV_X1 U11366 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U11367 ( .A1(n10301), .A2(n10307), .B1(n10300), .B2(n10299), .ZN(
        P1_U3475) );
  INV_X1 U11368 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U11369 ( .A1(n10308), .A2(n10303), .B1(n10302), .B2(n10306), .ZN(
        P1_U3524) );
  AOI22_X1 U11370 ( .A1(n10308), .A2(n10305), .B1(n10304), .B2(n10306), .ZN(
        P1_U3526) );
  AOI22_X1 U11371 ( .A1(n10308), .A2(n10307), .B1(n6945), .B2(n10306), .ZN(
        P1_U3530) );
  INV_X1 U11372 ( .A(n10309), .ZN(n10310) );
  OR2_X1 U11373 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  OAI211_X1 U11374 ( .C1(n10321), .C2(n10314), .A(n10313), .B(n10312), .ZN(
        n10319) );
  AOI22_X1 U11375 ( .A1(n6293), .A2(n10317), .B1(n10316), .B2(n10315), .ZN(
        n10318) );
  NAND2_X1 U11376 ( .A1(n10319), .A2(n10318), .ZN(n10360) );
  INV_X1 U11377 ( .A(n10360), .ZN(n10324) );
  XNOR2_X1 U11378 ( .A(n10321), .B(n10320), .ZN(n10362) );
  NAND2_X1 U11379 ( .A1(n10362), .A2(n10322), .ZN(n10323) );
  OAI211_X1 U11380 ( .C1(n10326), .C2(n10325), .A(n10324), .B(n10323), .ZN(
        n10327) );
  INV_X1 U11381 ( .A(n10327), .ZN(n10336) );
  NAND2_X1 U11382 ( .A1(n6488), .A2(n10353), .ZN(n10328) );
  NAND2_X1 U11383 ( .A1(n10329), .A2(n10328), .ZN(n10359) );
  INV_X1 U11384 ( .A(n10359), .ZN(n10331) );
  AOI22_X1 U11385 ( .A1(n10332), .A2(n10331), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n10330), .ZN(n10333) );
  OAI221_X1 U11386 ( .B1(n10337), .B2(n10336), .C1(n10335), .C2(n10334), .A(
        n10333), .ZN(P2_U3295) );
  AND2_X1 U11387 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10346), .ZN(P2_U3297) );
  AND2_X1 U11388 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10346), .ZN(P2_U3298) );
  AND2_X1 U11389 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10346), .ZN(P2_U3299) );
  AND2_X1 U11390 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10346), .ZN(P2_U3300) );
  AND2_X1 U11391 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10346), .ZN(P2_U3301) );
  AND2_X1 U11392 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10346), .ZN(P2_U3302) );
  AND2_X1 U11393 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10346), .ZN(P2_U3303) );
  AND2_X1 U11394 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10346), .ZN(P2_U3304) );
  AND2_X1 U11395 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10346), .ZN(P2_U3305) );
  AND2_X1 U11396 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10346), .ZN(P2_U3306) );
  AND2_X1 U11397 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10346), .ZN(P2_U3307) );
  AND2_X1 U11398 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10346), .ZN(P2_U3308) );
  INV_X1 U11399 ( .A(n10346), .ZN(n10349) );
  NOR2_X1 U11400 ( .A1(n10349), .A2(n10340), .ZN(P2_U3309) );
  AND2_X1 U11401 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10346), .ZN(P2_U3310) );
  AND2_X1 U11402 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10346), .ZN(P2_U3311) );
  AND2_X1 U11403 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10346), .ZN(P2_U3312) );
  AND2_X1 U11404 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10346), .ZN(P2_U3313) );
  AND2_X1 U11405 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10346), .ZN(P2_U3314) );
  AND2_X1 U11406 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10346), .ZN(P2_U3315) );
  AND2_X1 U11407 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10346), .ZN(P2_U3316) );
  AND2_X1 U11408 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10346), .ZN(P2_U3317) );
  NOR2_X1 U11409 ( .A1(n10349), .A2(n10341), .ZN(P2_U3318) );
  NOR2_X1 U11410 ( .A1(n10349), .A2(n10342), .ZN(P2_U3319) );
  AND2_X1 U11411 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10346), .ZN(P2_U3320) );
  AND2_X1 U11412 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10346), .ZN(P2_U3321) );
  NOR2_X1 U11413 ( .A1(n10349), .A2(n10343), .ZN(P2_U3322) );
  NOR2_X1 U11414 ( .A1(n10349), .A2(n10344), .ZN(P2_U3323) );
  AND2_X1 U11415 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10346), .ZN(P2_U3324) );
  AND2_X1 U11416 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10346), .ZN(P2_U3325) );
  AND2_X1 U11417 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10346), .ZN(P2_U3326) );
  NAND2_X1 U11418 ( .A1(n10345), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10350) );
  INV_X1 U11419 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U11420 ( .A1(n10348), .A2(n6148), .B1(n10347), .B2(n10346), .ZN(
        P2_U3437) );
  OAI22_X1 U11421 ( .A1(n10351), .A2(n10350), .B1(P2_D_REG_1__SCAN_IN), .B2(
        n10349), .ZN(n10352) );
  INV_X1 U11422 ( .A(n10352), .ZN(P2_U3438) );
  AOI22_X1 U11423 ( .A1(n10354), .A2(n10393), .B1(n10353), .B2(n6229), .ZN(
        n10355) );
  AND2_X1 U11424 ( .A1(n10356), .A2(n10355), .ZN(n10408) );
  INV_X1 U11425 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U11426 ( .A1(n10407), .A2(n10408), .B1(n10357), .B2(n10405), .ZN(
        P2_U3451) );
  NAND2_X1 U11427 ( .A1(n10396), .A2(n6488), .ZN(n10358) );
  OAI21_X1 U11428 ( .B1(n10359), .B2(n6279), .A(n10358), .ZN(n10361) );
  AOI211_X1 U11429 ( .C1(n10393), .C2(n10362), .A(n10361), .B(n10360), .ZN(
        n10410) );
  INV_X1 U11430 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U11431 ( .A1(n10407), .A2(n10410), .B1(n10363), .B2(n10405), .ZN(
        P2_U3454) );
  OAI21_X1 U11432 ( .B1(n10365), .B2(n10390), .A(n10364), .ZN(n10367) );
  AOI211_X1 U11433 ( .C1(n10393), .C2(n10368), .A(n10367), .B(n10366), .ZN(
        n10412) );
  INV_X1 U11434 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U11435 ( .A1(n10407), .A2(n10412), .B1(n10369), .B2(n10405), .ZN(
        P2_U3457) );
  NAND2_X1 U11436 ( .A1(n10371), .A2(n10370), .ZN(n10372) );
  AOI21_X1 U11437 ( .B1(n10393), .B2(n10373), .A(n10372), .ZN(n10414) );
  INV_X1 U11438 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U11439 ( .A1(n10407), .A2(n10414), .B1(n10374), .B2(n10405), .ZN(
        P2_U3460) );
  INV_X1 U11440 ( .A(n10375), .ZN(n10380) );
  OAI22_X1 U11441 ( .A1(n10376), .A2(n6279), .B1(n6497), .B2(n10390), .ZN(
        n10379) );
  INV_X1 U11442 ( .A(n10377), .ZN(n10378) );
  AOI211_X1 U11443 ( .C1(n10393), .C2(n10380), .A(n10379), .B(n10378), .ZN(
        n10416) );
  INV_X1 U11444 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U11445 ( .A1(n10407), .A2(n10416), .B1(n10381), .B2(n10405), .ZN(
        P2_U3463) );
  OAI21_X1 U11446 ( .B1(n10383), .B2(n10390), .A(n10382), .ZN(n10385) );
  AOI211_X1 U11447 ( .C1(n10393), .C2(n10386), .A(n10385), .B(n10384), .ZN(
        n10418) );
  INV_X1 U11448 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U11449 ( .A1(n10407), .A2(n10418), .B1(n10387), .B2(n10405), .ZN(
        P2_U3466) );
  OAI211_X1 U11450 ( .C1(n10391), .C2(n10390), .A(n10389), .B(n10388), .ZN(
        n10392) );
  AOI21_X1 U11451 ( .B1(n10394), .B2(n10393), .A(n10392), .ZN(n10419) );
  INV_X1 U11452 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U11453 ( .A1(n10407), .A2(n10419), .B1(n10395), .B2(n10405), .ZN(
        P2_U3469) );
  AOI22_X1 U11454 ( .A1(n10399), .A2(n10398), .B1(n10397), .B2(n10396), .ZN(
        n10400) );
  OAI211_X1 U11455 ( .C1(n10403), .C2(n10402), .A(n10401), .B(n10400), .ZN(
        n10404) );
  INV_X1 U11456 ( .A(n10404), .ZN(n10422) );
  INV_X1 U11457 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U11458 ( .A1(n10407), .A2(n10422), .B1(n10406), .B2(n10405), .ZN(
        P2_U3475) );
  AOI22_X1 U11459 ( .A1(n10423), .A2(n10408), .B1(n7386), .B2(n10420), .ZN(
        P2_U3520) );
  AOI22_X1 U11460 ( .A1(n10423), .A2(n10410), .B1(n10409), .B2(n10420), .ZN(
        P2_U3521) );
  INV_X1 U11461 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U11462 ( .A1(n10423), .A2(n10412), .B1(n10411), .B2(n10420), .ZN(
        P2_U3522) );
  INV_X1 U11463 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U11464 ( .A1(n10423), .A2(n10414), .B1(n10413), .B2(n10420), .ZN(
        P2_U3523) );
  AOI22_X1 U11465 ( .A1(n10423), .A2(n10416), .B1(n10415), .B2(n10420), .ZN(
        P2_U3524) );
  INV_X1 U11466 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U11467 ( .A1(n10423), .A2(n10418), .B1(n10417), .B2(n10420), .ZN(
        P2_U3525) );
  AOI22_X1 U11468 ( .A1(n10423), .A2(n10419), .B1(n7300), .B2(n10420), .ZN(
        P2_U3526) );
  AOI22_X1 U11469 ( .A1(n10423), .A2(n10422), .B1(n10421), .B2(n10420), .ZN(
        P2_U3528) );
  INV_X1 U11470 ( .A(n10424), .ZN(n10425) );
  NAND2_X1 U11471 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  XOR2_X1 U11472 ( .A(n10428), .B(n10427), .Z(ADD_1071_U5) );
  XOR2_X1 U11473 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11474 ( .B1(n10431), .B2(n10430), .A(n10429), .ZN(ADD_1071_U56) );
  OAI21_X1 U11475 ( .B1(n10434), .B2(n10433), .A(n10432), .ZN(ADD_1071_U57) );
  OAI21_X1 U11476 ( .B1(n10437), .B2(n10436), .A(n10435), .ZN(ADD_1071_U58) );
  OAI21_X1 U11477 ( .B1(n10440), .B2(n10439), .A(n10438), .ZN(ADD_1071_U59) );
  OAI21_X1 U11478 ( .B1(n10443), .B2(n10442), .A(n10441), .ZN(ADD_1071_U60) );
  OAI21_X1 U11479 ( .B1(n10446), .B2(n10445), .A(n10444), .ZN(ADD_1071_U61) );
  AOI21_X1 U11480 ( .B1(n10449), .B2(n10448), .A(n10447), .ZN(ADD_1071_U62) );
  AOI21_X1 U11481 ( .B1(n10452), .B2(n10451), .A(n10450), .ZN(ADD_1071_U63) );
  XOR2_X1 U11482 ( .A(n10454), .B(n10453), .Z(ADD_1071_U50) );
  NOR2_X1 U11483 ( .A1(n10456), .A2(n10455), .ZN(n10457) );
  XOR2_X1 U11484 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10457), .Z(ADD_1071_U51) );
  OAI21_X1 U11485 ( .B1(n10460), .B2(n10459), .A(n10458), .ZN(n10461) );
  XNOR2_X1 U11486 ( .A(n10461), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11487 ( .B1(n10464), .B2(n10463), .A(n10462), .ZN(ADD_1071_U47) );
  OAI21_X1 U11488 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(n10468) );
  XNOR2_X1 U11489 ( .A(n10468), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(ADD_1071_U48)
         );
  NOR2_X1 U11490 ( .A1(n10470), .A2(n10469), .ZN(n10471) );
  XOR2_X1 U11491 ( .A(n10472), .B(n10471), .Z(ADD_1071_U49) );
  XOR2_X1 U11492 ( .A(n10474), .B(n10473), .Z(ADD_1071_U54) );
  XOR2_X1 U11493 ( .A(n10476), .B(n10475), .Z(ADD_1071_U53) );
  XNOR2_X1 U11494 ( .A(n10478), .B(n10477), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4921 ( .A(n5080), .Z(n10216) );
  CLKBUF_X1 U4937 ( .A(n5720), .Z(n4391) );
  CLKBUF_X1 U4961 ( .A(n10265), .Z(n10279) );
  CLKBUF_X1 U5072 ( .A(n5699), .Z(n4392) );
endmodule

