

module b15_C_AntiSAT_k_128_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3012, n3013, n3014, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824;

  INV_X2 U34600 ( .A(n6106), .ZN(n4374) );
  INV_X1 U34610 ( .A(n6614), .ZN(n6075) );
  OR2_X1 U34620 ( .A1(n4578), .A2(n3499), .ZN(n3506) );
  AND2_X1 U34630 ( .A1(n3945), .A2(n3944), .ZN(n4465) );
  CLKBUF_X2 U34640 ( .A(n3962), .Z(n4054) );
  CLKBUF_X1 U34650 ( .A(n4031), .Z(n5312) );
  CLKBUF_X2 U3466 ( .A(n3313), .Z(n3229) );
  BUF_X1 U3467 ( .A(n3241), .Z(n3696) );
  CLKBUF_X1 U34680 ( .A(n3864), .Z(n3666) );
  CLKBUF_X1 U34690 ( .A(n3759), .Z(n3855) );
  CLKBUF_X2 U34700 ( .A(n3209), .Z(n3718) );
  CLKBUF_X2 U34710 ( .A(n3760), .Z(n3854) );
  INV_X1 U34740 ( .A(n3018), .ZN(n3166) );
  NOR2_X1 U3475 ( .A1(n4235), .A2(n3162), .ZN(n4094) );
  INV_X1 U3476 ( .A(n4235), .ZN(n3154) );
  NAND2_X2 U3477 ( .A1(n3086), .A2(n3085), .ZN(n5325) );
  AND4_X1 U3478 ( .A1(n3084), .A2(n3083), .A3(n3082), .A4(n3081), .ZN(n3085)
         );
  CLKBUF_X2 U3479 ( .A(n3140), .Z(n3829) );
  AND4_X1 U3480 ( .A1(n3071), .A2(n3070), .A3(n3069), .A4(n3068), .ZN(n3072)
         );
  AND4_X1 U3481 ( .A1(n3059), .A2(n3058), .A3(n3057), .A4(n3056), .ZN(n3075)
         );
  NAND2_X2 U3482 ( .A1(n3055), .A2(n3026), .ZN(n4419) );
  AOI22_X1 U3483 ( .A1(n3241), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3084) );
  AND4_X1 U3484 ( .A1(n3046), .A2(n3045), .A3(n3044), .A4(n3043), .ZN(n3025)
         );
  AND2_X4 U3485 ( .A1(n5409), .A2(n4478), .ZN(n3241) );
  AND2_X2 U3486 ( .A1(n5409), .A2(n3042), .ZN(n3313) );
  NOR2_X1 U3487 ( .A1(n4185), .A2(n4031), .ZN(n4467) );
  NAND2_X1 U3488 ( .A1(n3032), .A2(n3025), .ZN(n3127) );
  AND2_X1 U3489 ( .A1(n3953), .A2(n3952), .ZN(n3954) );
  NAND2_X1 U3490 ( .A1(n5325), .A2(n4419), .ZN(n5324) );
  AND2_X1 U3493 ( .A1(n5448), .A2(n5447), .ZN(n5623) );
  AOI211_X1 U3494 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5443), .A(n5442), .B(n5441), .ZN(n5444) );
  INV_X1 U3495 ( .A(n6615), .ZN(n6060) );
  OR2_X4 U3496 ( .A1(n5689), .A2(n5688), .ZN(n5691) );
  AND4_X4 U3497 ( .A1(n3075), .A2(n3074), .A3(n3073), .A4(n3072), .ZN(n3018)
         );
  AOI21_X2 U3498 ( .B1(n4355), .B2(n4354), .A(n4100), .ZN(n6188) );
  INV_X2 U3499 ( .A(n4916), .ZN(n3555) );
  AND2_X4 U3500 ( .A1(n3500), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3042)
         );
  AND4_X2 U3501 ( .A1(n4184), .A2(n3167), .A3(n3173), .A4(n4290), .ZN(n3168)
         );
  CLKBUF_X3 U3502 ( .A(n4078), .Z(n4721) );
  OAI21_X2 U3504 ( .B1(n4526), .B2(STATE2_REG_0__SCAN_IN), .A(n3280), .ZN(
        n3465) );
  OAI21_X2 U3505 ( .B1(n4077), .B2(n4147), .A(n4076), .ZN(n4106) );
  OAI22_X2 U3506 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n5661), .B1(n5671), .B2(n5419), .ZN(n5420) );
  NOR2_X1 U3507 ( .A1(n5626), .A2(n5652), .ZN(n4180) );
  BUF_X2 U3509 ( .A(n3829), .Z(n3853) );
  AND2_X1 U3510 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U3511 ( .A1(n4178), .A2(n4177), .ZN(n5626) );
  OR2_X1 U3512 ( .A1(n5695), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5696)
         );
  NAND2_X1 U3513 ( .A1(n5414), .A2(n4173), .ZN(n5695) );
  NAND2_X1 U3514 ( .A1(n5708), .A2(n4171), .ZN(n5414) );
  CLKBUF_X1 U3515 ( .A(n5353), .Z(n3021) );
  AOI21_X1 U3516 ( .B1(n4982), .B2(n4161), .A(n3027), .ZN(n5291) );
  XNOR2_X1 U3517 ( .A(n4053), .B(n4052), .ZN(n5367) );
  NAND2_X1 U3518 ( .A1(n6178), .A2(n6177), .ZN(n6180) );
  NAND2_X1 U3519 ( .A1(n3497), .A2(n3496), .ZN(n4443) );
  BUF_X1 U3520 ( .A(n4077), .Z(n4578) );
  AND2_X1 U3521 ( .A1(n3283), .A2(n3490), .ZN(n3016) );
  NAND2_X2 U3522 ( .A1(n5586), .A2(n4425), .ZN(n5931) );
  NAND2_X1 U3523 ( .A1(n3287), .A2(n3286), .ZN(n4348) );
  NAND2_X1 U3524 ( .A1(n3258), .A2(n4148), .ZN(n3464) );
  NOR2_X2 U3525 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4529), .ZN(n5072) );
  CLKBUF_X1 U3526 ( .A(n3172), .Z(n3183) );
  INV_X1 U3527 ( .A(n3191), .ZN(n4245) );
  CLKBUF_X1 U3528 ( .A(n4094), .Z(n4236) );
  NAND2_X1 U3529 ( .A1(n4448), .A2(n5312), .ZN(n4034) );
  NOR2_X1 U3530 ( .A1(n4468), .A2(n5324), .ZN(n4221) );
  INV_X1 U3532 ( .A(n4931), .ZN(n4553) );
  OR2_X1 U3533 ( .A1(n3240), .A2(n3239), .ZN(n4151) );
  AND4_X1 U3534 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .ZN(n3126)
         );
  AND4_X1 U3535 ( .A1(n3063), .A2(n3062), .A3(n3061), .A4(n3060), .ZN(n3074)
         );
  AND4_X1 U3536 ( .A1(n3067), .A2(n3066), .A3(n3065), .A4(n3064), .ZN(n3073)
         );
  AND4_X1 U3537 ( .A1(n3114), .A2(n3113), .A3(n3112), .A4(n3111), .ZN(n3125)
         );
  AND4_X1 U3538 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3104)
         );
  AND4_X1 U3539 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .ZN(n3106)
         );
  AND4_X1 U3540 ( .A1(n3122), .A2(n3121), .A3(n3120), .A4(n3119), .ZN(n3123)
         );
  AND4_X1 U3541 ( .A1(n3040), .A2(n3039), .A3(n3038), .A4(n3037), .ZN(n3032)
         );
  AND4_X1 U3542 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3105)
         );
  BUF_X2 U3543 ( .A(n3228), .Z(n3857) );
  BUF_X2 U3544 ( .A(n3260), .Z(n3836) );
  BUF_X2 U3545 ( .A(n3234), .Z(n3856) );
  CLKBUF_X1 U3546 ( .A(n3500), .Z(n4481) );
  NOR2_X2 U3547 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3019) );
  NOR2_X2 U3548 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4509) );
  INV_X1 U3549 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3500) );
  OR2_X2 U3551 ( .A1(n6051), .A2(n6050), .ZN(n6053) );
  OAI21_X1 U3552 ( .B1(n5716), .B2(n4169), .A(n4168), .ZN(n4170) );
  AND2_X1 U3553 ( .A1(n5646), .A2(n3013), .ZN(n5616) );
  AND2_X1 U3554 ( .A1(n5644), .A2(n4253), .ZN(n3013) );
  NOR2_X1 U3555 ( .A1(n4180), .A2(n4179), .ZN(n3014) );
  INV_X1 U3556 ( .A(n3127), .ZN(n3164) );
  NOR2_X1 U3557 ( .A1(n4180), .A2(n4179), .ZN(n5646) );
  NAND2_X1 U3559 ( .A1(n3283), .A2(n3490), .ZN(n3017) );
  NAND2_X1 U3560 ( .A1(n3014), .A2(n5644), .ZN(n5638) );
  INV_X2 U3561 ( .A(n4577), .ZN(n3308) );
  NAND2_X1 U3562 ( .A1(n4542), .A2(n3185), .ZN(n3165) );
  AND2_X4 U3563 ( .A1(n3034), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5409)
         );
  AND2_X2 U3564 ( .A1(n5508), .A2(n5422), .ZN(n5421) );
  OR2_X2 U3565 ( .A1(n4960), .A2(n4961), .ZN(n5170) );
  NOR2_X4 U3566 ( .A1(n5582), .A2(n4020), .ZN(n5508) );
  NAND2_X2 U3567 ( .A1(n3506), .A2(n3505), .ZN(n4442) );
  AND4_X2 U3568 ( .A1(n3054), .A2(n3053), .A3(n3052), .A4(n3051), .ZN(n3026)
         );
  NAND2_X1 U3569 ( .A1(n3508), .A2(n3498), .ZN(n4077) );
  AND2_X4 U3570 ( .A1(n5406), .A2(n3042), .ZN(n3133) );
  AND2_X2 U3571 ( .A1(n3307), .A2(n3306), .ZN(n4577) );
  INV_X1 U3572 ( .A(n3203), .ZN(n3020) );
  XNOR2_X1 U3573 ( .A(n3466), .B(n3465), .ZN(n4519) );
  XNOR2_X2 U3574 ( .A(n3958), .B(n4361), .ZN(n5034) );
  OAI21_X2 U3575 ( .B1(n4027), .B2(EBX_REG_1__SCAN_IN), .A(n3954), .ZN(n3958)
         );
  XNOR2_X1 U3576 ( .A(n4200), .B(n4266), .ZN(n4277) );
  AND2_X1 U3577 ( .A1(n4105), .A2(n4104), .ZN(n6177) );
  OAI21_X2 U3578 ( .B1(n3024), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5418), 
        .ZN(n5671) );
  NAND2_X1 U3579 ( .A1(n4984), .A2(n4983), .ZN(n4982) );
  OAI21_X1 U3580 ( .B1(n4198), .B2(n4266), .A(n4181), .ZN(n4182) );
  AND2_X1 U3581 ( .A1(n5409), .A2(n3042), .ZN(n3023) );
  NOR2_X1 U3582 ( .A1(n4465), .A2(n5994), .ZN(n4370) );
  AOI22_X1 U3583 ( .A1(n3241), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3132) );
  AND2_X1 U3584 ( .A1(n5390), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3843) );
  OAI21_X1 U3585 ( .B1(n3943), .B2(n3942), .A(n3941), .ZN(n3944) );
  INV_X1 U3586 ( .A(n6490), .ZN(n5994) );
  OR2_X1 U3587 ( .A1(n5681), .A2(n5578), .ZN(n3685) );
  INV_X1 U3588 ( .A(n3843), .ZN(n3881) );
  CLKBUF_X1 U3589 ( .A(n3946), .Z(n3753) );
  INV_X1 U3590 ( .A(n3946), .ZN(n3878) );
  NAND2_X1 U3591 ( .A1(n3915), .A2(n3166), .ZN(n3935) );
  AND2_X1 U3592 ( .A1(n3175), .A2(n3558), .ZN(n5390) );
  OR2_X2 U3593 ( .A1(n3139), .A2(n3138), .ZN(n4080) );
  OR3_X1 U3594 ( .A1(n6598), .A2(n6279), .A3(n3947), .ZN(n4966) );
  AND2_X1 U3595 ( .A1(n4676), .A2(n4675), .ZN(n4678) );
  INV_X1 U3596 ( .A(n3962), .ZN(n4448) );
  AND2_X1 U3597 ( .A1(n6475), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3885) );
  OR2_X1 U3598 ( .A1(n3777), .A2(n3776), .ZN(n3821) );
  INV_X1 U3599 ( .A(n3732), .ZN(n3731) );
  NOR2_X1 U3600 ( .A1(n3557), .A2(n6801), .ZN(n3601) );
  NOR2_X1 U3601 ( .A1(n4224), .A2(n4050), .ZN(n4053) );
  INV_X1 U3602 ( .A(n4031), .ZN(n5800) );
  AND2_X1 U3603 ( .A1(n4250), .A2(n4249), .ZN(n4477) );
  NOR2_X2 U3604 ( .A1(n5178), .A2(n4454), .ZN(n4676) );
  NAND2_X1 U3605 ( .A1(n4215), .A2(n4214), .ZN(n4255) );
  OR2_X1 U3607 ( .A1(n4623), .A2(n3022), .ZN(n4842) );
  INV_X1 U3608 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6480) );
  INV_X1 U3609 ( .A(n5586), .ZN(n6098) );
  AND2_X1 U3610 ( .A1(n5586), .A2(n4426), .ZN(n5173) );
  INV_X1 U3611 ( .A(n6197), .ZN(n5946) );
  INV_X1 U3612 ( .A(n6165), .ZN(n6193) );
  NAND2_X1 U3613 ( .A1(n4186), .A2(n4370), .ZN(n6165) );
  NOR2_X1 U3614 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  INV_X1 U3615 ( .A(n5367), .ZN(n5380) );
  INV_X1 U3616 ( .A(n6262), .ZN(n6277) );
  INV_X1 U3617 ( .A(n6255), .ZN(n6273) );
  NAND2_X1 U3618 ( .A1(n3321), .A2(n3507), .ZN(n3528) );
  INV_X1 U3619 ( .A(n3508), .ZN(n3321) );
  OR2_X1 U3620 ( .A1(n3319), .A2(n3318), .ZN(n4124) );
  INV_X1 U3621 ( .A(n4080), .ZN(n3162) );
  AND2_X1 U3622 ( .A1(n4931), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3915) );
  NAND2_X1 U3623 ( .A1(n4417), .A2(n3294), .ZN(n3920) );
  OR2_X1 U3624 ( .A1(n3304), .A2(n3303), .ZN(n4109) );
  NAND2_X1 U3625 ( .A1(n3866), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3065) );
  OR2_X1 U3626 ( .A1(n3166), .A2(n6596), .ZN(n4417) );
  NOR2_X1 U3627 ( .A1(n3602), .A2(n5262), .ZN(n3603) );
  INV_X1 U3628 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3518) );
  NAND2_X1 U3629 ( .A1(n3171), .A2(n3170), .ZN(n3227) );
  OR2_X1 U3630 ( .A1(n4931), .A2(n6596), .ZN(n3294) );
  OR2_X1 U3631 ( .A1(n3271), .A2(n3270), .ZN(n4092) );
  NAND2_X1 U3632 ( .A1(n3282), .A2(n3281), .ZN(n3490) );
  INV_X1 U3633 ( .A(n3920), .ZN(n3943) );
  AND2_X1 U3634 ( .A1(n3904), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3906)
         );
  NOR2_X1 U3635 ( .A1(n3935), .A2(n4147), .ZN(n3936) );
  AND2_X1 U3636 ( .A1(n3289), .A2(n4567), .ZN(n4798) );
  AOI21_X1 U3637 ( .B1(n6595), .B2(n6493), .A(n5408), .ZN(n4529) );
  INV_X1 U3638 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6460) );
  INV_X1 U3639 ( .A(n4210), .ZN(n4470) );
  NAND2_X1 U3640 ( .A1(n5006), .A2(n4058), .ZN(n6608) );
  INV_X1 U3641 ( .A(n3285), .ZN(n3287) );
  CLKBUF_X1 U3642 ( .A(n3284), .Z(n3285) );
  INV_X1 U3643 ( .A(n6608), .ZN(n6025) );
  AND2_X1 U3644 ( .A1(n3973), .A2(n3972), .ZN(n4675) );
  OR2_X1 U3645 ( .A1(n5621), .A2(n3878), .ZN(n3851) );
  NAND2_X1 U3646 ( .A1(n3820), .A2(n3819), .ZN(n3849) );
  INV_X1 U3647 ( .A(n3821), .ZN(n3820) );
  CLKBUF_X1 U3648 ( .A(n5445), .Z(n5458) );
  OR2_X1 U3650 ( .A1(n3775), .A2(n5653), .ZN(n3777) );
  OR2_X1 U3651 ( .A1(n3780), .A2(n3779), .ZN(n5469) );
  AND2_X1 U3652 ( .A1(n5657), .A2(n3753), .ZN(n3754) );
  NAND2_X1 U3653 ( .A1(n3710), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3732)
         );
  AND2_X1 U3654 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3678), .ZN(n3679)
         );
  OR2_X1 U3655 ( .A1(n5897), .A2(n3878), .ZN(n3683) );
  AND2_X1 U3656 ( .A1(n3641), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3643)
         );
  NAND2_X1 U3657 ( .A1(n3643), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3677)
         );
  AND2_X1 U3659 ( .A1(n3572), .A2(n3571), .ZN(n5019) );
  BUF_X1 U3660 ( .A(n5021), .Z(n5244) );
  NOR2_X1 U3661 ( .A1(n6620), .A2(n3538), .ZN(n3556) );
  NAND2_X1 U3662 ( .A1(n3380), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3538)
         );
  NAND2_X1 U3663 ( .A1(n3408), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3382)
         );
  INV_X1 U3664 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3381) );
  NOR2_X1 U3665 ( .A1(n3382), .A2(n3381), .ZN(n3380) );
  NAND2_X1 U3666 ( .A1(n3445), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3428)
         );
  INV_X1 U3667 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3427) );
  NOR2_X1 U3668 ( .A1(n3529), .A2(n3518), .ZN(n3346) );
  NAND2_X1 U3669 ( .A1(n3346), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3352)
         );
  AND2_X2 U3670 ( .A1(n4613), .A2(n3537), .ZN(n4903) );
  AND2_X1 U3671 ( .A1(n4557), .A2(n4614), .ZN(n3537) );
  NAND2_X1 U3672 ( .A1(n3530), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3529)
         );
  INV_X1 U3673 ( .A(n3484), .ZN(n3501) );
  NAND2_X1 U3674 ( .A1(n3501), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3513)
         );
  NAND2_X1 U3675 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3484) );
  AND2_X1 U3676 ( .A1(n5818), .A2(n5627), .ZN(n4179) );
  NAND2_X1 U3677 ( .A1(n5659), .A2(n5417), .ZN(n5677) );
  NOR2_X2 U3678 ( .A1(n5677), .A2(n5678), .ZN(n5676) );
  OR2_X1 U3679 ( .A1(n5818), .A2(n4172), .ZN(n4173) );
  CLKBUF_X1 U3680 ( .A(n5708), .Z(n5709) );
  OR2_X1 U3681 ( .A1(n5625), .A2(n5980), .ZN(n5360) );
  AND2_X1 U3682 ( .A1(n3983), .A2(n3982), .ZN(n4911) );
  NOR2_X2 U3683 ( .A1(n6053), .A2(n4911), .ZN(n4979) );
  CLKBUF_X1 U3684 ( .A(n4982), .Z(n5269) );
  INV_X1 U3685 ( .A(n5175), .ZN(n3966) );
  AND2_X1 U3686 ( .A1(n4036), .A2(n4031), .ZN(n4360) );
  OAI211_X1 U3687 ( .C1(n3203), .C2(n5413), .A(n3201), .B(n3200), .ZN(n3276)
         );
  INV_X1 U3688 ( .A(n5390), .ZN(n5399) );
  AND2_X2 U3689 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4479) );
  AND2_X1 U3690 ( .A1(n4346), .A2(n4446), .ZN(n6452) );
  OR2_X1 U3691 ( .A1(n5016), .A2(n5403), .ZN(n5125) );
  AND2_X1 U3692 ( .A1(n4760), .A2(n5192), .ZN(n5844) );
  INV_X1 U3693 ( .A(n4841), .ZN(n4869) );
  NOR2_X1 U3694 ( .A1(n4578), .A2(n4721), .ZN(n6381) );
  INV_X1 U3695 ( .A(n4419), .ZN(n4542) );
  INV_X1 U3696 ( .A(n6337), .ZN(n6387) );
  OR2_X1 U3697 ( .A1(n4842), .A2(n4869), .ZN(n4805) );
  OR2_X1 U3698 ( .A1(n5896), .A2(n4069), .ZN(n5437) );
  AND2_X1 U3699 ( .A1(n4966), .A2(n4936), .ZN(n6614) );
  INV_X1 U3700 ( .A(n6611), .ZN(n6035) );
  AND2_X1 U3701 ( .A1(n4966), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6054) );
  CLKBUF_X1 U3702 ( .A(n3475), .Z(n6385) );
  AND2_X1 U3703 ( .A1(n6060), .A2(n5004), .ZN(n6065) );
  OR2_X1 U3704 ( .A1(n4446), .A2(n5994), .ZN(n4453) );
  INV_X1 U3705 ( .A(n5325), .ZN(n5585) );
  INV_X1 U3706 ( .A(n5623), .ZN(n5596) );
  NAND2_X1 U3707 ( .A1(n4424), .A2(n4423), .ZN(n5586) );
  AND2_X1 U3708 ( .A1(n4422), .A2(n4421), .ZN(n4423) );
  INV_X1 U3709 ( .A(n5173), .ZN(n5255) );
  AND2_X1 U3710 ( .A1(n4373), .A2(n4372), .ZN(n6116) );
  INV_X1 U3711 ( .A(n6159), .ZN(n6153) );
  XNOR2_X1 U3712 ( .A(n3949), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4935)
         );
  OR2_X1 U3713 ( .A1(n3948), .A2(n4279), .ZN(n3949) );
  NOR2_X1 U3714 ( .A1(n5817), .A2(n4271), .ZN(n5790) );
  OR2_X1 U3715 ( .A1(n5951), .A2(n4270), .ZN(n5817) );
  NOR2_X1 U3716 ( .A1(n5980), .A2(n5981), .ZN(n5959) );
  AND2_X1 U3717 ( .A1(n4986), .A2(n4985), .ZN(n6214) );
  INV_X1 U3718 ( .A(n6254), .ZN(n6279) );
  INV_X1 U3719 ( .A(n5974), .ZN(n4366) );
  INV_X1 U3720 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6447) );
  XNOR2_X1 U3721 ( .A(n3464), .B(n3463), .ZN(n3466) );
  CLKBUF_X1 U3722 ( .A(n4492), .Z(n5016) );
  INV_X1 U3724 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5413) );
  INV_X1 U3725 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3034) );
  INV_X1 U3726 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3036) );
  INV_X1 U3727 ( .A(n5158), .ZN(n6368) );
  OR2_X1 U3728 ( .A1(n6288), .A2(n5116), .ZN(n5158) );
  INV_X1 U3729 ( .A(n5063), .ZN(n5099) );
  AND2_X1 U3730 ( .A1(n6477), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6490) );
  INV_X1 U3731 ( .A(n4283), .ZN(n4284) );
  OAI21_X1 U3732 ( .B1(n5593), .B2(n5352), .A(n4282), .ZN(n4283) );
  INV_X1 U3733 ( .A(n5376), .ZN(n5377) );
  OAI21_X1 U3734 ( .B1(n5380), .B2(n6255), .A(n5375), .ZN(n5376) );
  AOI211_X1 U3735 ( .C1(n5374), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5373), .B(n5372), .ZN(n5375) );
  AND2_X1 U3736 ( .A1(n4274), .A2(n3029), .ZN(n4275) );
  AND2_X2 U3737 ( .A1(n4150), .A2(n4149), .ZN(n3024) );
  OAI21_X1 U3738 ( .B1(n3203), .B2(n3204), .A(n3208), .ZN(n3286) );
  NAND2_X1 U3739 ( .A1(n5276), .A2(n4160), .ZN(n3027) );
  NAND2_X1 U3740 ( .A1(n5818), .A2(n6792), .ZN(n3028) );
  INV_X1 U3741 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U3742 ( .A1(n6081), .A2(n5585), .ZN(n6077) );
  AND2_X1 U3743 ( .A1(n4979), .A2(n4978), .ZN(n4977) );
  INV_X1 U3744 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3512) );
  INV_X1 U3745 ( .A(n6388), .ZN(n6382) );
  OR2_X1 U3746 ( .A1(n5371), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3029)
         );
  INV_X1 U3747 ( .A(n4917), .ZN(n3554) );
  OR2_X1 U3748 ( .A1(n4956), .A2(n4955), .ZN(n4975) );
  AND2_X1 U3749 ( .A1(n4902), .A2(n3462), .ZN(n3030) );
  OR2_X1 U3750 ( .A1(n4070), .A2(n4193), .ZN(n3031) );
  AND2_X1 U3751 ( .A1(n6159), .A2(n4309), .ZN(n6156) );
  NAND2_X1 U3752 ( .A1(n3030), .A2(n4903), .ZN(n4916) );
  AND2_X1 U3753 ( .A1(n6081), .A2(n5325), .ZN(n6085) );
  INV_X1 U3754 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3204) );
  OR2_X1 U3755 ( .A1(n3014), .A2(n5617), .ZN(n3033) );
  INV_X4 U3756 ( .A(n3024), .ZN(n5818) );
  AND2_X1 U3757 ( .A1(n6382), .A2(n4188), .ZN(n6192) );
  INV_X1 U3758 ( .A(n3951), .ZN(n4036) );
  NAND2_X1 U3759 ( .A1(n4447), .A2(n3161), .ZN(n4239) );
  NOR2_X1 U3760 ( .A1(n5003), .A2(n3910), .ZN(n3928) );
  AND2_X1 U3761 ( .A1(n6447), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3913)
         );
  OR2_X1 U3762 ( .A1(n3331), .A2(n3330), .ZN(n4123) );
  NAND2_X1 U3763 ( .A1(n3893), .A2(n3892), .ZN(n3897) );
  INV_X1 U3764 ( .A(n5324), .ZN(n4234) );
  OR2_X1 U3765 ( .A1(n3220), .A2(n3219), .ZN(n3223) );
  AOI21_X1 U3766 ( .B1(n3897), .B2(n3895), .A(n3894), .ZN(n3903) );
  AND2_X1 U3767 ( .A1(n3938), .A2(n3929), .ZN(n3909) );
  INV_X1 U3768 ( .A(n3963), .ZN(n3951) );
  INV_X1 U3769 ( .A(n3677), .ZN(n3678) );
  BUF_X1 U3771 ( .A(n3261), .Z(n3831) );
  AND2_X1 U3772 ( .A1(n3920), .A2(n4140), .ZN(n3520) );
  OR2_X1 U3773 ( .A1(n3343), .A2(n3342), .ZN(n4140) );
  INV_X1 U3774 ( .A(n3223), .ZN(n4079) );
  AND2_X1 U3775 ( .A1(n3903), .A2(n4353), .ZN(n3905) );
  NAND2_X1 U3776 ( .A1(n3164), .A2(n4419), .ZN(n3159) );
  XNOR2_X1 U3777 ( .A(n4150), .B(n3345), .ZN(n4138) );
  INV_X1 U3778 ( .A(n3849), .ZN(n3848) );
  INV_X1 U3779 ( .A(n3711), .ZN(n3710) );
  INV_X1 U3780 ( .A(n3601), .ZN(n3602) );
  OR2_X1 U3781 ( .A1(n5325), .A2(n6475), .ZN(n3584) );
  NAND2_X1 U3782 ( .A1(n3524), .A2(n3523), .ZN(n4122) );
  NAND2_X1 U3783 ( .A1(n3519), .A2(n3520), .ZN(n4150) );
  OR2_X1 U3784 ( .A1(n3906), .A2(n3905), .ZN(n3942) );
  OR2_X1 U3785 ( .A1(n3251), .A2(n3250), .ZN(n4093) );
  AND2_X1 U3786 ( .A1(n6025), .A2(n4064), .ZN(n5259) );
  AND2_X1 U3787 ( .A1(n3971), .A2(n3970), .ZN(n4454) );
  BUF_X1 U3788 ( .A(n3159), .Z(n4447) );
  NAND2_X1 U3789 ( .A1(n3848), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3948)
         );
  NAND2_X1 U3790 ( .A1(n3679), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3711)
         );
  NAND2_X1 U3791 ( .A1(n3556), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3557)
         );
  AND2_X1 U3792 ( .A1(n3412), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3408)
         );
  AND2_X1 U3793 ( .A1(n5818), .A2(n5980), .ZN(n5361) );
  INV_X1 U3794 ( .A(n3024), .ZN(n5625) );
  NAND2_X1 U3795 ( .A1(n4129), .A2(n4128), .ZN(n4135) );
  NOR2_X1 U3797 ( .A1(n3254), .A2(n6596), .ZN(n3257) );
  INV_X1 U3798 ( .A(n4205), .ZN(n3193) );
  INV_X1 U3799 ( .A(n6054), .ZN(n6619) );
  NOR2_X1 U3800 ( .A1(n3428), .A2(n3427), .ZN(n3412) );
  AND2_X1 U3801 ( .A1(n4935), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3950) );
  XNOR2_X1 U3802 ( .A(n4348), .B(n6294), .ZN(n4466) );
  AND2_X1 U3803 ( .A1(n4966), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U3804 ( .A1(n3351), .A2(n3350), .ZN(n4902) );
  NAND2_X1 U3805 ( .A1(n3731), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3775)
         );
  AND2_X1 U3806 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n3603), .ZN(n3641)
         );
  NOR2_X1 U3807 ( .A1(n4956), .A2(n4955), .ZN(n5105) );
  INV_X1 U3808 ( .A(n3352), .ZN(n3445) );
  INV_X1 U3809 ( .A(n6187), .ZN(n5702) );
  AND2_X1 U3810 ( .A1(n5787), .A2(n4262), .ZN(n5767) );
  AND2_X1 U3811 ( .A1(n5824), .A2(n4261), .ZN(n5787) );
  NAND2_X1 U3812 ( .A1(n4477), .A2(n4255), .ZN(n6250) );
  OR2_X1 U3813 ( .A1(n5997), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6254) );
  INV_X1 U3814 ( .A(n3889), .ZN(n4252) );
  INV_X1 U3816 ( .A(n3022), .ZN(n4860) );
  OR2_X1 U3817 ( .A1(n4692), .A2(n4841), .ZN(n6293) );
  INV_X1 U3818 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6456) );
  INV_X1 U3819 ( .A(n6338), .ZN(n6388) );
  INV_X1 U3820 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U3821 ( .A1(n3293), .A2(n3292), .ZN(n6294) );
  OR2_X1 U3822 ( .A1(n6570), .A2(n4529), .ZN(n4566) );
  AOI21_X1 U3823 ( .B1(n6447), .B2(STATE2_REG_3__SCAN_IN), .A(n4799), .ZN(
        n6337) );
  AND2_X1 U3824 ( .A1(n5006), .A2(n4934), .ZN(n6611) );
  AND2_X1 U3825 ( .A1(n4056), .A2(n4055), .ZN(n6058) );
  AND2_X1 U3826 ( .A1(n4966), .A2(n3950), .ZN(n6615) );
  NOR2_X2 U3827 ( .A1(n5562), .A2(n5561), .ZN(n5564) );
  INV_X1 U3828 ( .A(n6077), .ZN(n6084) );
  AND2_X1 U3829 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  AND2_X1 U3830 ( .A1(n5586), .A2(n5326), .ZN(n6099) );
  OR2_X1 U3831 ( .A1(n4309), .A2(n4538), .ZN(n4422) );
  INV_X1 U3832 ( .A(n4422), .ZN(n6157) );
  AND2_X1 U3833 ( .A1(n5580), .A2(n5579), .ZN(n5902) );
  NAND2_X1 U3834 ( .A1(n3555), .A2(n3554), .ZN(n5020) );
  OR2_X1 U3835 ( .A1(n4975), .A2(n4974), .ZN(n5236) );
  NOR2_X1 U3836 ( .A1(n3513), .A2(n3512), .ZN(n3530) );
  AND2_X1 U3837 ( .A1(n6165), .A2(n4190), .ZN(n6187) );
  NOR2_X1 U3838 ( .A1(n5758), .A2(n4273), .ZN(n5746) );
  AND2_X1 U3839 ( .A1(n5790), .A2(n5660), .ZN(n5770) );
  AND2_X1 U3840 ( .A1(n5333), .A2(n5332), .ZN(n6020) );
  OR2_X1 U3841 ( .A1(n4257), .A2(n4987), .ZN(n5969) );
  NOR2_X1 U3842 ( .A1(n6250), .A2(n6230), .ZN(n6238) );
  OR2_X1 U3843 ( .A1(n5976), .A2(n4366), .ZN(n6280) );
  OR2_X1 U3844 ( .A1(n5972), .A2(n4366), .ZN(n6227) );
  NOR2_X1 U3845 ( .A1(n6571), .A2(n4465), .ZN(n5408) );
  INV_X1 U3846 ( .A(n4768), .ZN(n4794) );
  AND3_X1 U3847 ( .A1(n4725), .A2(n5189), .A3(n4578), .ZN(n5882) );
  INV_X1 U3848 ( .A(n4753), .ZN(n4610) );
  INV_X1 U3849 ( .A(n4691), .ZN(n4717) );
  INV_X1 U3850 ( .A(n6293), .ZN(n6322) );
  INV_X1 U3851 ( .A(n6326), .ZN(n6370) );
  INV_X1 U3852 ( .A(n5188), .ZN(n5231) );
  INV_X1 U3853 ( .A(n6445), .ZN(n6430) );
  INV_X1 U3854 ( .A(n4805), .ZN(n4899) );
  OAI211_X1 U3855 ( .C1(n6571), .C2(n5075), .A(n5074), .B(n5073), .ZN(n5100)
         );
  INV_X1 U3856 ( .A(n5352), .ZN(n6181) );
  AND2_X1 U3857 ( .A1(n6480), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U3858 ( .A1(n4301), .A2(n4299), .ZN(n6598) );
  AND2_X1 U3859 ( .A1(n4071), .A2(n3031), .ZN(n4072) );
  INV_X1 U3860 ( .A(n6058), .ZN(n6624) );
  INV_X2 U3861 ( .A(n6118), .ZN(n6132) );
  OR2_X1 U3862 ( .A1(n6116), .A2(n4374), .ZN(n6118) );
  INV_X1 U3863 ( .A(n6116), .ZN(n6135) );
  INV_X1 U3864 ( .A(n6156), .ZN(n6143) );
  NAND2_X1 U3865 ( .A1(n4370), .A2(n4306), .ZN(n6159) );
  OR2_X1 U3866 ( .A1(n6187), .A2(n4435), .ZN(n6197) );
  NAND2_X1 U3867 ( .A1(n4255), .A2(n4219), .ZN(n6262) );
  INV_X1 U3868 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5395) );
  INV_X1 U3869 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4353) );
  AND2_X1 U3870 ( .A1(n4636), .A2(n4635), .ZN(n4674) );
  OR2_X1 U3871 ( .A1(n4769), .A2(n4841), .ZN(n5884) );
  INV_X1 U3872 ( .A(n4724), .ZN(n4759) );
  OR2_X1 U3873 ( .A1(n4692), .A2(n4869), .ZN(n4691) );
  OR2_X1 U3874 ( .A1(n6288), .A2(n6287), .ZN(n6326) );
  NAND2_X1 U3875 ( .A1(n4861), .A2(n4869), .ZN(n5188) );
  NAND2_X1 U3876 ( .A1(n6381), .A2(n4800), .ZN(n6434) );
  NAND2_X1 U3877 ( .A1(n6381), .A2(n5189), .ZN(n6445) );
  NOR2_X1 U3878 ( .A1(n4804), .A2(n4803), .ZN(n4840) );
  OR2_X1 U3879 ( .A1(n4842), .A2(n4841), .ZN(n5103) );
  OR2_X1 U3880 ( .A1(n4623), .A2(n6287), .ZN(n5063) );
  NOR2_X4 U3881 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4478) );
  INV_X1 U3882 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3035) );
  AND2_X2 U3883 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n3035), .ZN(n3041)
         );
  AND2_X4 U3884 ( .A1(n3041), .A2(n3019), .ZN(n3759) );
  AOI22_X1 U3885 ( .A1(n3241), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3040) );
  AND2_X2 U3886 ( .A1(n3036), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5406)
         );
  AND2_X2 U3887 ( .A1(n5406), .A2(n4479), .ZN(n3076) );
  AOI22_X1 U3888 ( .A1(n3076), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3039) );
  AND2_X4 U3889 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5398) );
  AND2_X2 U3890 ( .A1(n3041), .A2(n5398), .ZN(n3128) );
  AND2_X2 U3891 ( .A1(n3019), .A2(n4479), .ZN(n3234) );
  AOI22_X1 U3892 ( .A1(n3128), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3234), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3038) );
  AND2_X2 U3893 ( .A1(n5409), .A2(n3041), .ZN(n3140) );
  AOI22_X1 U3895 ( .A1(n3140), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3037) );
  AND2_X4 U3896 ( .A1(n5409), .A2(n4479), .ZN(n3261) );
  AOI22_X1 U3897 ( .A1(n3133), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3046) );
  AND2_X2 U3898 ( .A1(n5406), .A2(n4478), .ZN(n3260) );
  AND2_X2 U3899 ( .A1(n3042), .A2(n4509), .ZN(n3760) );
  AOI22_X1 U3900 ( .A1(n3260), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3760), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3045) );
  AND2_X2 U3901 ( .A1(n3041), .A2(n5406), .ZN(n3228) );
  AND2_X2 U3902 ( .A1(n4478), .A2(n5398), .ZN(n3209) );
  AOI22_X1 U3903 ( .A1(n3228), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3044) );
  AND2_X4 U3904 ( .A1(n3042), .A2(n5398), .ZN(n3866) );
  AND2_X4 U3905 ( .A1(n4509), .A2(n4478), .ZN(n3214) );
  AOI22_X1 U3906 ( .A1(n3866), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3043) );
  AOI22_X1 U3907 ( .A1(n3241), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3128), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3050) );
  AOI22_X1 U3908 ( .A1(n3228), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3049) );
  AOI22_X1 U3909 ( .A1(n3140), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3760), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3048) );
  AOI22_X1 U3910 ( .A1(n3234), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3047) );
  AND4_X2 U3911 ( .A1(n3050), .A2(n3049), .A3(n3048), .A4(n3047), .ZN(n3055)
         );
  AOI22_X1 U3912 ( .A1(n3076), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3023), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3054) );
  AOI22_X1 U3913 ( .A1(n3133), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U3914 ( .A1(n3866), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3052) );
  AOI22_X1 U3915 ( .A1(n3261), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3916 ( .A1(n3133), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3059) );
  NAND2_X1 U3917 ( .A1(n3260), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3058) );
  NAND2_X1 U3918 ( .A1(n3261), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3057)
         );
  NAND2_X1 U3919 ( .A1(n3145), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3056)
         );
  NAND2_X1 U3920 ( .A1(n3228), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3063) );
  NAND2_X1 U3921 ( .A1(n3140), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3062)
         );
  NAND2_X1 U3922 ( .A1(n3759), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3061) );
  NAND2_X1 U3923 ( .A1(n3760), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3060) );
  BUF_X2 U3924 ( .A(n3076), .Z(n3830) );
  NAND2_X1 U3925 ( .A1(n3830), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3067)
         );
  NAND2_X1 U3926 ( .A1(n3313), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3066) );
  NAND2_X1 U3927 ( .A1(n3214), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3064) );
  NAND2_X1 U3928 ( .A1(n3241), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3071) );
  NAND2_X1 U3930 ( .A1(n3128), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3070)
         );
  NAND2_X1 U3931 ( .A1(n3234), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3069)
         );
  NAND2_X1 U3932 ( .A1(n3209), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3068) );
  NAND2_X1 U3933 ( .A1(n3159), .A2(n3018), .ZN(n3152) );
  AOI22_X1 U3934 ( .A1(n3133), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3080) );
  AOI22_X1 U3935 ( .A1(n3864), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3079) );
  AOI22_X1 U3936 ( .A1(n3261), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3078) );
  AOI22_X1 U3937 ( .A1(n3866), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3077) );
  AOI22_X1 U3939 ( .A1(n3234), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3083) );
  AOI22_X1 U3940 ( .A1(n3140), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3760), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3082) );
  AOI22_X1 U3941 ( .A1(n3228), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3081) );
  OR2_X2 U3942 ( .A1(n3152), .A2(n5585), .ZN(n4203) );
  NAND2_X1 U3943 ( .A1(n3228), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3944 ( .A1(n3140), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3089)
         );
  NAND2_X1 U3945 ( .A1(n3759), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3946 ( .A1(n3760), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U3947 ( .A1(n3133), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U3948 ( .A1(n3260), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3093) );
  NAND2_X1 U3949 ( .A1(n3261), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3092)
         );
  NAND2_X1 U3950 ( .A1(n3145), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3091)
         );
  NAND2_X1 U3951 ( .A1(n3830), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3098)
         );
  NAND2_X1 U3952 ( .A1(n3313), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3953 ( .A1(n3866), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U3954 ( .A1(n3214), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3095) );
  NAND2_X1 U3955 ( .A1(n3241), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3102) );
  NAND2_X1 U3956 ( .A1(n3128), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3101)
         );
  NAND2_X1 U3957 ( .A1(n3234), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3100)
         );
  NAND2_X1 U3958 ( .A1(n3209), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3099) );
  NAND4_X4 U3960 ( .A1(n3106), .A2(n3105), .A3(n3104), .A4(n3103), .ZN(n4205)
         );
  NAND2_X1 U3961 ( .A1(n3829), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3110)
         );
  NAND2_X1 U3962 ( .A1(n3759), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3109) );
  NAND2_X1 U3963 ( .A1(n3133), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U3964 ( .A1(n3214), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3965 ( .A1(n3241), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3114) );
  NAND2_X1 U3966 ( .A1(n3261), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3113)
         );
  NAND2_X1 U3967 ( .A1(n3260), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3112) );
  NAND2_X1 U3968 ( .A1(n3760), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3111) );
  NAND2_X1 U3969 ( .A1(n3830), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3118)
         );
  NAND2_X1 U3970 ( .A1(n3313), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3117) );
  NAND2_X1 U3971 ( .A1(n3866), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3116) );
  NAND2_X1 U3972 ( .A1(n3145), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3115)
         );
  NAND2_X1 U3974 ( .A1(n3228), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3122) );
  NAND2_X1 U3975 ( .A1(n3128), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3121)
         );
  NAND2_X1 U3976 ( .A1(n3234), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3120)
         );
  NAND2_X1 U3977 ( .A1(n3209), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3119) );
  NAND4_X4 U3978 ( .A1(n3126), .A2(n3125), .A3(n3124), .A4(n3123), .ZN(n4931)
         );
  AND2_X2 U3979 ( .A1(n3193), .A2(n4931), .ZN(n6594) );
  BUF_X4 U3980 ( .A(n3127), .Z(n3185) );
  NAND2_X2 U3981 ( .A1(n3018), .A2(n3185), .ZN(n3178) );
  AOI22_X1 U3982 ( .A1(n3228), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U3983 ( .A1(n3140), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3760), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U3984 ( .A1(n3234), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3129) );
  NAND4_X1 U3985 ( .A1(n3132), .A2(n3131), .A3(n3130), .A4(n3129), .ZN(n3139)
         );
  AOI22_X1 U3986 ( .A1(n3133), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U3987 ( .A1(n3864), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3136) );
  AOI22_X1 U3988 ( .A1(n3261), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U3989 ( .A1(n3866), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3134) );
  NAND4_X1 U3990 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3138)
         );
  NAND2_X2 U3991 ( .A1(n4080), .A2(n4205), .ZN(n4031) );
  AOI21_X1 U3992 ( .B1(n4203), .B2(n6594), .A(n4467), .ZN(n3158) );
  AND2_X2 U3993 ( .A1(n4542), .A2(n5325), .ZN(n3175) );
  AOI22_X1 U3994 ( .A1(n3140), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3760), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U3995 ( .A1(n3864), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U3996 ( .A1(n3261), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U3997 ( .A1(n3228), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3234), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3141) );
  NAND4_X1 U3998 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n3151)
         );
  AOI22_X1 U3999 ( .A1(n3241), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4000 ( .A1(n3133), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4001 ( .A1(n3128), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4002 ( .A1(n3214), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3146) );
  NAND4_X1 U4003 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3150)
         );
  OAI21_X1 U4004 ( .B1(n3152), .B2(n3175), .A(n4235), .ZN(n3157) );
  OAI21_X1 U4005 ( .B1(n3018), .B2(n4419), .A(n3159), .ZN(n3153) );
  INV_X1 U4006 ( .A(n3153), .ZN(n3155) );
  NAND2_X1 U4007 ( .A1(n3155), .A2(n3154), .ZN(n3156) );
  NAND2_X1 U4008 ( .A1(n3165), .A2(n4080), .ZN(n3177) );
  NAND4_X1 U4009 ( .A1(n3157), .A2(n3156), .A3(n5325), .A4(n3177), .ZN(n3190)
         );
  NOR2_X2 U4010 ( .A1(n4931), .A2(n4205), .ZN(n5003) );
  NAND2_X1 U4011 ( .A1(n3190), .A2(n5003), .ZN(n4243) );
  NAND2_X1 U4012 ( .A1(n3158), .A2(n4243), .ZN(n3172) );
  INV_X1 U4013 ( .A(n3172), .ZN(n3169) );
  NAND2_X1 U4014 ( .A1(n3178), .A2(n5325), .ZN(n3160) );
  NAND2_X1 U4015 ( .A1(n3160), .A2(n5324), .ZN(n3161) );
  INV_X1 U4016 ( .A(n4094), .ZN(n3186) );
  NOR2_X2 U4017 ( .A1(n4239), .A2(n3186), .ZN(n4184) );
  INV_X1 U4018 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6505) );
  XNOR2_X1 U4019 ( .A(n6505), .B(STATE_REG_2__SCAN_IN), .ZN(n4057) );
  INV_X1 U4020 ( .A(n4057), .ZN(n3163) );
  NAND2_X1 U4021 ( .A1(n3193), .A2(n3163), .ZN(n3189) );
  NAND2_X1 U4022 ( .A1(n3189), .A2(n3012), .ZN(n3167) );
  NAND2_X1 U4023 ( .A1(n3165), .A2(n3166), .ZN(n3173) );
  NAND2_X1 U4024 ( .A1(n4553), .A2(n4205), .ZN(n4290) );
  AOI21_X2 U4025 ( .B1(n3169), .B2(n3168), .A(n6596), .ZN(n3288) );
  NAND2_X1 U4026 ( .A1(n3288), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3171) );
  NOR2_X1 U4027 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6489) );
  NAND2_X1 U4028 ( .A1(n6489), .A2(n6596), .ZN(n4189) );
  MUX2_X1 U4029 ( .A(n4189), .B(n6477), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3170) );
  NAND2_X1 U4030 ( .A1(n3173), .A2(n4080), .ZN(n3174) );
  OAI21_X1 U4031 ( .B1(n4239), .B2(n3174), .A(n4205), .ZN(n3181) );
  NOR2_X1 U4032 ( .A1(n4235), .A2(n4080), .ZN(n4449) );
  AND2_X1 U4033 ( .A1(n4449), .A2(n4553), .ZN(n4244) );
  NAND2_X1 U4034 ( .A1(n6489), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3176) );
  AOI21_X1 U4035 ( .B1(n4244), .B2(n3175), .A(n3176), .ZN(n3180) );
  NAND2_X1 U4036 ( .A1(n3177), .A2(n6594), .ZN(n3179) );
  OR2_X1 U4037 ( .A1(n3178), .A2(n4931), .ZN(n3191) );
  INV_X1 U4038 ( .A(n5003), .ZN(n4287) );
  OAI211_X1 U4039 ( .C1(n4553), .C2(n4235), .A(n3191), .B(n4287), .ZN(n4233)
         );
  NAND4_X1 U4040 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n4233), .ZN(n3182)
         );
  NOR2_X2 U4041 ( .A1(n3183), .A2(n3182), .ZN(n3226) );
  INV_X1 U4042 ( .A(n3226), .ZN(n3184) );
  NAND2_X2 U4043 ( .A1(n3227), .A2(n3184), .ZN(n3275) );
  NAND3_X1 U4044 ( .A1(n4449), .A2(n5003), .A3(n3012), .ZN(n4468) );
  INV_X1 U4045 ( .A(n4221), .ZN(n3195) );
  NOR2_X1 U4046 ( .A1(n3186), .A2(n3185), .ZN(n3188) );
  INV_X1 U4047 ( .A(n4203), .ZN(n3187) );
  AND2_X2 U4048 ( .A1(n3188), .A2(n3187), .ZN(n4210) );
  AND2_X2 U4049 ( .A1(n4210), .A2(n4931), .ZN(n4307) );
  NAND2_X1 U4050 ( .A1(n4307), .A2(n3189), .ZN(n3194) );
  INV_X1 U4051 ( .A(n3190), .ZN(n3192) );
  AND2_X2 U4052 ( .A1(n3192), .A2(n4245), .ZN(n3889) );
  NAND2_X2 U4053 ( .A1(n3889), .A2(n4538), .ZN(n4473) );
  NAND3_X1 U4054 ( .A1(n3195), .A2(n3194), .A3(n4473), .ZN(n3196) );
  NAND2_X1 U4055 ( .A1(n3196), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3200) );
  INV_X1 U4056 ( .A(n3200), .ZN(n3199) );
  INV_X1 U4057 ( .A(n4189), .ZN(n3291) );
  XNOR2_X1 U4058 ( .A(n6447), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6289)
         );
  INV_X1 U4059 ( .A(n6477), .ZN(n3290) );
  AND2_X1 U4060 ( .A1(n3290), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3197)
         );
  AOI21_X1 U4061 ( .B1(n3291), .B2(n6289), .A(n3197), .ZN(n3201) );
  NAND2_X1 U4062 ( .A1(n3201), .A2(n5413), .ZN(n3198) );
  NAND2_X1 U4063 ( .A1(n3199), .A2(n3198), .ZN(n3277) );
  NAND2_X1 U4064 ( .A1(n3275), .A2(n3277), .ZN(n3202) );
  INV_X1 U4065 ( .A(n3288), .ZN(n3203) );
  NAND2_X1 U4066 ( .A1(n3202), .A2(n3276), .ZN(n3284) );
  AND2_X1 U4067 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4068 ( .A1(n3205), .A2(n6460), .ZN(n6378) );
  INV_X1 U4069 ( .A(n3205), .ZN(n3206) );
  NAND2_X1 U4070 ( .A1(n3206), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U4071 ( .A1(n6378), .A2(n3207), .ZN(n4582) );
  AOI22_X1 U4072 ( .A1(n3291), .A2(n4582), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3290), .ZN(n3208) );
  XNOR2_X1 U4073 ( .A(n3284), .B(n3286), .ZN(n4492) );
  NAND2_X1 U4074 ( .A1(n4492), .A2(n6596), .ZN(n3222) );
  INV_X1 U4075 ( .A(n4417), .ZN(n3279) );
  AOI22_X1 U4076 ( .A1(n3696), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4077 ( .A1(n3857), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4078 ( .A1(n3853), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4079 ( .A1(n3856), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3210) );
  NAND4_X1 U4080 ( .A1(n3213), .A2(n3212), .A3(n3211), .A4(n3210), .ZN(n3220)
         );
  AOI22_X1 U4081 ( .A1(n3784), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4082 ( .A1(n3666), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U4083 ( .A1(n3831), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4084 ( .A1(n3866), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3215) );
  NAND4_X1 U4085 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n3219)
         );
  NAND2_X1 U4086 ( .A1(n3279), .A2(n3223), .ZN(n3221) );
  NAND2_X1 U4087 ( .A1(n3222), .A2(n3221), .ZN(n3225) );
  INV_X1 U4088 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4662) );
  OAI22_X1 U4089 ( .A1(n3935), .A2(n4662), .B1(n4079), .B2(n3294), .ZN(n3224)
         );
  XNOR2_X1 U4090 ( .A(n3225), .B(n3224), .ZN(n3491) );
  INV_X1 U4091 ( .A(n3491), .ZN(n3283) );
  XNOR2_X1 U4092 ( .A(n3227), .B(n3226), .ZN(n3475) );
  NAND2_X1 U4093 ( .A1(n3475), .A2(n6596), .ZN(n3471) );
  AOI22_X1 U4094 ( .A1(n3857), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4095 ( .A1(n3853), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U4096 ( .A1(n3784), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3231) );
  AOI22_X1 U4097 ( .A1(n3666), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3023), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3230) );
  NAND4_X1 U4098 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n3240)
         );
  AOI22_X1 U4099 ( .A1(n3696), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4100 ( .A1(n3856), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4101 ( .A1(n3866), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4102 ( .A1(n3854), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3235) );
  NAND4_X1 U4103 ( .A1(n3238), .A2(n3237), .A3(n3236), .A4(n3235), .ZN(n3239)
         );
  NOR2_X1 U4104 ( .A1(n4417), .A2(n4151), .ZN(n3259) );
  NAND2_X1 U4105 ( .A1(n3018), .A2(n4151), .ZN(n3254) );
  AOI22_X1 U4106 ( .A1(n3857), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3696), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4107 ( .A1(n3784), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4108 ( .A1(n3313), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4109 ( .A1(n3856), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3242) );
  NAND4_X1 U4110 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3251)
         );
  AOI22_X1 U4111 ( .A1(n3128), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4112 ( .A1(n3853), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4113 ( .A1(n3261), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4114 ( .A1(n3666), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3246) );
  NAND4_X1 U4115 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3250)
         );
  INV_X1 U4116 ( .A(n4093), .ZN(n3252) );
  MUX2_X1 U4117 ( .A(n3259), .B(n3257), .S(n3252), .Z(n3472) );
  INV_X1 U4118 ( .A(n3472), .ZN(n3253) );
  NAND2_X1 U4119 ( .A1(n3471), .A2(n3253), .ZN(n3256) );
  INV_X1 U4120 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4666) );
  AOI21_X1 U4121 ( .B1(n4553), .B2(n4093), .A(n6596), .ZN(n3255) );
  OAI211_X1 U4122 ( .C1(n3935), .C2(n4666), .A(n3255), .B(n3254), .ZN(n3473)
         );
  NAND2_X1 U4123 ( .A1(n3256), .A2(n3473), .ZN(n3258) );
  INV_X1 U4124 ( .A(n3257), .ZN(n4148) );
  INV_X1 U4125 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4642) );
  INV_X1 U4126 ( .A(n3259), .ZN(n3274) );
  INV_X1 U4127 ( .A(n3294), .ZN(n3272) );
  AOI22_X1 U4128 ( .A1(n3853), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4129 ( .A1(n3133), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4130 ( .A1(n3831), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4131 ( .A1(n3128), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3262) );
  NAND4_X1 U4132 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3271)
         );
  AOI22_X1 U4133 ( .A1(n3864), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4134 ( .A1(n3855), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4135 ( .A1(n3857), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4136 ( .A1(n3863), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3266) );
  NAND4_X1 U4137 ( .A1(n3269), .A2(n3268), .A3(n3267), .A4(n3266), .ZN(n3270)
         );
  NAND2_X1 U4138 ( .A1(n3272), .A2(n4092), .ZN(n3273) );
  OAI211_X1 U4139 ( .C1(n3935), .C2(n4642), .A(n3274), .B(n3273), .ZN(n3463)
         );
  NAND2_X1 U4140 ( .A1(n3277), .A2(n3276), .ZN(n3278) );
  XNOR2_X2 U4141 ( .A(n3275), .B(n3278), .ZN(n4526) );
  NAND2_X1 U4142 ( .A1(n3279), .A2(n4092), .ZN(n3280) );
  OAI21_X1 U4143 ( .B1(n3464), .B2(n3463), .A(n3465), .ZN(n3282) );
  NAND2_X1 U4144 ( .A1(n3464), .A2(n3463), .ZN(n3281) );
  NAND2_X1 U4145 ( .A1(n3020), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3293) );
  NOR3_X1 U4146 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6460), .A3(n6456), 
        .ZN(n6339) );
  NAND2_X1 U4147 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6339), .ZN(n6333) );
  NAND2_X1 U4148 ( .A1(n6377), .A2(n6333), .ZN(n3289) );
  NOR3_X1 U4149 ( .A1(n6377), .A2(n6460), .A3(n6456), .ZN(n5067) );
  NAND2_X1 U4150 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5067), .ZN(n4567) );
  AOI22_X1 U4151 ( .A1(n3291), .A2(n4798), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3290), .ZN(n3292) );
  NAND2_X1 U4152 ( .A1(n4466), .A2(n6596), .ZN(n3307) );
  INV_X1 U4153 ( .A(n3935), .ZN(n3305) );
  AOI22_X1 U4154 ( .A1(n3696), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4155 ( .A1(n3857), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4156 ( .A1(n3853), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4157 ( .A1(n3856), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3295) );
  NAND4_X1 U4158 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3304)
         );
  AOI22_X1 U4159 ( .A1(n3784), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4160 ( .A1(n3666), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4161 ( .A1(n3831), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4162 ( .A1(n4483), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3299) );
  NAND4_X1 U4163 ( .A1(n3302), .A2(n3301), .A3(n3300), .A4(n3299), .ZN(n3303)
         );
  AOI22_X1 U4164 ( .A1(n3305), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3920), 
        .B2(n4109), .ZN(n3306) );
  NAND2_X2 U4165 ( .A1(n3016), .A2(n3308), .ZN(n3508) );
  INV_X1 U4166 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U4167 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3789), .B1(n3241), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4168 ( .A1(n3857), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4169 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3853), .B1(n3854), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4170 ( .A1(n3856), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3309) );
  NAND4_X1 U4171 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3319)
         );
  AOI22_X1 U4172 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3836), .B1(n3784), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4173 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3666), .B1(n3229), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4174 ( .A1(n3831), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4175 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4483), .B1(n3863), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3314) );
  NAND4_X1 U4176 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3318)
         );
  NAND2_X1 U4177 ( .A1(n3920), .A2(n4124), .ZN(n3320) );
  OAI21_X1 U4178 ( .B1(n3935), .B2(n4658), .A(n3320), .ZN(n3507) );
  INV_X1 U4179 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4646) );
  AOI22_X1 U4180 ( .A1(n3696), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4181 ( .A1(n3857), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4182 ( .A1(n3853), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4183 ( .A1(n3856), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3322) );
  NAND4_X1 U4184 ( .A1(n3325), .A2(n3324), .A3(n3323), .A4(n3322), .ZN(n3331)
         );
  AOI22_X1 U4185 ( .A1(n3784), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4186 ( .A1(n3666), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4187 ( .A1(n3831), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4188 ( .A1(n4483), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3326) );
  NAND4_X1 U4189 ( .A1(n3329), .A2(n3328), .A3(n3327), .A4(n3326), .ZN(n3330)
         );
  NAND2_X1 U4190 ( .A1(n3920), .A2(n4123), .ZN(n3332) );
  OAI21_X1 U4191 ( .B1(n3935), .B2(n4646), .A(n3332), .ZN(n3527) );
  INV_X1 U4192 ( .A(n3527), .ZN(n3333) );
  NOR2_X2 U4193 ( .A1(n3528), .A2(n3333), .ZN(n3519) );
  AOI22_X1 U4194 ( .A1(n3696), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4195 ( .A1(n3857), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4196 ( .A1(n3853), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4197 ( .A1(n3856), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3334) );
  NAND4_X1 U4198 ( .A1(n3337), .A2(n3336), .A3(n3335), .A4(n3334), .ZN(n3343)
         );
  AOI22_X1 U4199 ( .A1(n3784), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4200 ( .A1(n3666), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4201 ( .A1(n3831), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4202 ( .A1(n4483), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3338) );
  NAND4_X1 U4203 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3342)
         );
  INV_X1 U4204 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U4205 ( .A1(n3920), .A2(n4151), .ZN(n3344) );
  OAI21_X1 U4206 ( .B1(n3935), .B2(n4673), .A(n3344), .ZN(n3345) );
  INV_X2 U4207 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6475) );
  NOR2_X2 U4208 ( .A1(n4419), .A2(n6475), .ZN(n3547) );
  NAND2_X1 U4209 ( .A1(n4138), .A2(n3547), .ZN(n3351) );
  INV_X2 U4210 ( .A(n3584), .ZN(n3886) );
  AOI22_X1 U4211 ( .A1(n3886), .A2(EAX_REG_7__SCAN_IN), .B1(n3885), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3349) );
  OR2_X1 U4212 ( .A1(n3346), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3347) );
  NAND2_X1 U4213 ( .A1(n3347), .A2(n3352), .ZN(n6169) );
  NOR2_X1 U4214 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3946) );
  NAND2_X1 U4215 ( .A1(n6169), .A2(n3753), .ZN(n3348) );
  AND2_X1 U4216 ( .A1(n3349), .A2(n3348), .ZN(n3350) );
  INV_X1 U4217 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6620) );
  XOR2_X1 U4218 ( .A(n6620), .B(n3538), .Z(n6613) );
  AOI22_X1 U4219 ( .A1(n3857), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3356) );
  CLKBUF_X2 U4220 ( .A(n3133), .Z(n3784) );
  AOI22_X1 U4221 ( .A1(n3784), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3831), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4222 ( .A1(n3696), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4223 ( .A1(n4483), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3353) );
  NAND4_X1 U4224 ( .A1(n3356), .A2(n3355), .A3(n3354), .A4(n3353), .ZN(n3362)
         );
  AOI22_X1 U4225 ( .A1(n3666), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4226 ( .A1(n3855), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4227 ( .A1(n3789), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4228 ( .A1(n3836), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3357) );
  NAND4_X1 U4229 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3361)
         );
  OR2_X1 U4230 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  AOI22_X1 U4231 ( .A1(n3547), .A2(n3363), .B1(n3885), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U4232 ( .A1(n3886), .A2(EAX_REG_14__SCAN_IN), .ZN(n3364) );
  OAI211_X1 U4233 ( .C1(n6613), .C2(n3878), .A(n3365), .B(n3364), .ZN(n4906)
         );
  XNOR2_X1 U4234 ( .A(n3380), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5521)
         );
  AOI22_X1 U4235 ( .A1(n3857), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4236 ( .A1(n3666), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4237 ( .A1(n3831), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4238 ( .A1(n3696), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3366) );
  NAND4_X1 U4239 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3375)
         );
  AOI22_X1 U4240 ( .A1(n3784), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4241 ( .A1(n3853), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4242 ( .A1(n3789), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4243 ( .A1(n3214), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3370) );
  NAND4_X1 U4244 ( .A1(n3373), .A2(n3372), .A3(n3371), .A4(n3370), .ZN(n3374)
         );
  OAI21_X1 U4245 ( .B1(n3375), .B2(n3374), .A(n3547), .ZN(n3378) );
  NAND2_X1 U4246 ( .A1(n3886), .A2(EAX_REG_13__SCAN_IN), .ZN(n3377) );
  NAND2_X1 U4247 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3376)
         );
  NAND3_X1 U4248 ( .A1(n3378), .A2(n3377), .A3(n3376), .ZN(n3379) );
  AOI21_X1 U4249 ( .B1(n5521), .B2(n3753), .A(n3379), .ZN(n5107) );
  INV_X1 U4250 ( .A(n5107), .ZN(n3444) );
  AOI21_X1 U4251 ( .B1(n3382), .B2(n3381), .A(n3380), .ZN(n6029) );
  OR2_X1 U4252 ( .A1(n6029), .A2(n3878), .ZN(n3397) );
  AOI22_X1 U4253 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3857), .B1(n3696), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4254 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3229), .B1(n3830), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4255 ( .A1(n3784), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4256 ( .A1(n3831), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3383) );
  NAND4_X1 U4257 ( .A1(n3386), .A2(n3385), .A3(n3384), .A4(n3383), .ZN(n3392)
         );
  AOI22_X1 U4258 ( .A1(n3789), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4259 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3853), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4260 ( .A1(n3856), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4261 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4483), .B1(n3863), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3387) );
  NAND4_X1 U4262 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3391)
         );
  OAI21_X1 U4263 ( .B1(n3392), .B2(n3391), .A(n3547), .ZN(n3395) );
  NAND2_X1 U4264 ( .A1(n3886), .A2(EAX_REG_12__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4265 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3393)
         );
  AND3_X1 U4266 ( .A1(n3395), .A2(n3394), .A3(n3393), .ZN(n3396) );
  AND2_X1 U4267 ( .A1(n3397), .A2(n3396), .ZN(n5167) );
  INV_X1 U4268 ( .A(n5167), .ZN(n3443) );
  AOI22_X1 U4269 ( .A1(n3857), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4270 ( .A1(n3853), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3831), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4271 ( .A1(n3789), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4272 ( .A1(n3229), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3398) );
  NAND4_X1 U4273 ( .A1(n3401), .A2(n3400), .A3(n3399), .A4(n3398), .ZN(n3407)
         );
  AOI22_X1 U4274 ( .A1(n3836), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4275 ( .A1(n3784), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4276 ( .A1(n3696), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4277 ( .A1(n3666), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3402) );
  NAND4_X1 U4278 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3406)
         );
  NOR2_X1 U4279 ( .A1(n3407), .A2(n3406), .ZN(n3411) );
  INV_X1 U4280 ( .A(n3547), .ZN(n3499) );
  XNOR2_X1 U4281 ( .A(n3408), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5347)
         );
  NAND2_X1 U4282 ( .A1(n5347), .A2(n3753), .ZN(n3410) );
  AOI22_X1 U4283 ( .A1(n3886), .A2(EAX_REG_11__SCAN_IN), .B1(n3885), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3409) );
  OAI211_X1 U4284 ( .C1(n3411), .C2(n3499), .A(n3410), .B(n3409), .ZN(n4959)
         );
  XOR2_X1 U4285 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3412), .Z(n6041) );
  INV_X1 U4286 ( .A(n6041), .ZN(n5282) );
  AOI22_X1 U4287 ( .A1(n3857), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4288 ( .A1(n3784), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4289 ( .A1(n3831), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4290 ( .A1(n3229), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3413) );
  NAND4_X1 U4291 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3422)
         );
  AOI22_X1 U4292 ( .A1(n3696), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4293 ( .A1(n3853), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4294 ( .A1(n3856), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4295 ( .A1(n3666), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3417) );
  NAND4_X1 U4296 ( .A1(n3420), .A2(n3419), .A3(n3418), .A4(n3417), .ZN(n3421)
         );
  OAI21_X1 U4297 ( .B1(n3422), .B2(n3421), .A(n3547), .ZN(n3425) );
  NAND2_X1 U4298 ( .A1(n3886), .A2(EAX_REG_10__SCAN_IN), .ZN(n3424) );
  NAND2_X1 U4299 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3423)
         );
  NAND3_X1 U4300 ( .A1(n3425), .A2(n3424), .A3(n3423), .ZN(n3426) );
  AOI21_X1 U4301 ( .B1(n5282), .B2(n3753), .A(n3426), .ZN(n5237) );
  XNOR2_X1 U4302 ( .A(n3428), .B(n3427), .ZN(n5271) );
  AOI22_X1 U4303 ( .A1(n3759), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4304 ( .A1(n3831), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4305 ( .A1(n3857), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4306 ( .A1(n3229), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3429) );
  NAND4_X1 U4307 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3438)
         );
  AOI22_X1 U4308 ( .A1(n3853), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3784), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4309 ( .A1(n3696), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4310 ( .A1(n3789), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4311 ( .A1(n3666), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3433) );
  NAND4_X1 U4312 ( .A1(n3436), .A2(n3435), .A3(n3434), .A4(n3433), .ZN(n3437)
         );
  OAI21_X1 U4313 ( .B1(n3438), .B2(n3437), .A(n3547), .ZN(n3441) );
  NAND2_X1 U4314 ( .A1(n3886), .A2(EAX_REG_9__SCAN_IN), .ZN(n3440) );
  NAND2_X1 U4315 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3439)
         );
  NAND3_X1 U4316 ( .A1(n3441), .A2(n3440), .A3(n3439), .ZN(n3442) );
  AOI21_X1 U4317 ( .B1(n5271), .B2(n3753), .A(n3442), .ZN(n4974) );
  NOR2_X1 U4318 ( .A1(n5237), .A2(n4974), .ZN(n4957) );
  AND2_X1 U4319 ( .A1(n4959), .A2(n4957), .ZN(n4958) );
  AND2_X1 U4320 ( .A1(n3443), .A2(n4958), .ZN(n5104) );
  NAND2_X1 U4321 ( .A1(n3444), .A2(n5104), .ZN(n3461) );
  XOR2_X1 U4322 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3445), .Z(n4998) );
  INV_X1 U4323 ( .A(n4998), .ZN(n3460) );
  AOI22_X1 U4324 ( .A1(n3853), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4325 ( .A1(n3784), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3831), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4326 ( .A1(n3854), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4327 ( .A1(n3666), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3446) );
  NAND4_X1 U4328 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(n3455)
         );
  AOI22_X1 U4329 ( .A1(n3857), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4330 ( .A1(n3759), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4331 ( .A1(n3789), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4332 ( .A1(n3229), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3450) );
  NAND4_X1 U4333 ( .A1(n3453), .A2(n3452), .A3(n3451), .A4(n3450), .ZN(n3454)
         );
  OAI21_X1 U4334 ( .B1(n3455), .B2(n3454), .A(n3547), .ZN(n3458) );
  NAND2_X1 U4335 ( .A1(n3886), .A2(EAX_REG_8__SCAN_IN), .ZN(n3457) );
  NAND2_X1 U4336 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3456)
         );
  NAND3_X1 U4337 ( .A1(n3458), .A2(n3457), .A3(n3456), .ZN(n3459) );
  AOI21_X1 U4338 ( .B1(n3460), .B2(n3946), .A(n3459), .ZN(n4955) );
  NOR2_X1 U4339 ( .A1(n3461), .A2(n4955), .ZN(n4904) );
  AND2_X1 U4340 ( .A1(n4906), .A2(n4904), .ZN(n3462) );
  NAND2_X1 U4341 ( .A1(n4519), .A2(n3547), .ZN(n3470) );
  AOI22_X1 U4342 ( .A1(n3886), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6475), .ZN(n3468) );
  AND2_X1 U4343 ( .A1(n4234), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3483) );
  NAND2_X1 U4344 ( .A1(n3483), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3467) );
  AND2_X1 U4345 ( .A1(n3468), .A2(n3467), .ZN(n3469) );
  NAND2_X1 U4346 ( .A1(n3470), .A2(n3469), .ZN(n4413) );
  NAND2_X1 U4347 ( .A1(n3471), .A2(n3473), .ZN(n3474) );
  MUX2_X2 U4348 ( .A(n3474), .B(n3473), .S(n3472), .Z(n4841) );
  AOI21_X1 U4349 ( .B1(n4841), .B2(n3175), .A(n6475), .ZN(n4434) );
  NAND2_X1 U4350 ( .A1(n6385), .A2(n3547), .ZN(n3480) );
  INV_X1 U4351 ( .A(n3483), .ZN(n3511) );
  NAND2_X1 U4352 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6475), .ZN(n3477)
         );
  NAND2_X1 U4353 ( .A1(n3886), .A2(EAX_REG_0__SCAN_IN), .ZN(n3476) );
  OAI211_X1 U4354 ( .C1(n3511), .C2(n5395), .A(n3477), .B(n3476), .ZN(n3478)
         );
  INV_X1 U4355 ( .A(n3478), .ZN(n3479) );
  NAND2_X1 U4356 ( .A1(n3480), .A2(n3479), .ZN(n4433) );
  NAND2_X1 U4357 ( .A1(n4434), .A2(n4433), .ZN(n4432) );
  INV_X1 U4358 ( .A(n4433), .ZN(n3481) );
  NAND2_X1 U4359 ( .A1(n3481), .A2(n3946), .ZN(n3482) );
  NAND2_X1 U4360 ( .A1(n4432), .A2(n3482), .ZN(n4415) );
  NAND2_X1 U4361 ( .A1(n4413), .A2(n4415), .ZN(n4414) );
  NAND2_X1 U4362 ( .A1(n3483), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3489) );
  OAI21_X1 U4363 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3484), .ZN(n6196) );
  NAND2_X1 U4364 ( .A1(n6196), .A2(n3946), .ZN(n3486) );
  NAND2_X1 U4365 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3485)
         );
  NAND2_X1 U4366 ( .A1(n3486), .A2(n3485), .ZN(n3487) );
  AOI21_X1 U4367 ( .B1(n3886), .B2(EAX_REG_2__SCAN_IN), .A(n3487), .ZN(n3488)
         );
  AND2_X1 U4368 ( .A1(n3489), .A2(n3488), .ZN(n3493) );
  NAND2_X1 U4369 ( .A1(n4414), .A2(n3493), .ZN(n4428) );
  XNOR2_X1 U4370 ( .A(n3491), .B(n3490), .ZN(n4078) );
  NAND2_X1 U4371 ( .A1(n4721), .A2(n3547), .ZN(n3492) );
  INV_X1 U4372 ( .A(n3885), .ZN(n3735) );
  NAND2_X1 U4373 ( .A1(n3492), .A2(n3735), .ZN(n4427) );
  NAND2_X1 U4374 ( .A1(n4428), .A2(n4427), .ZN(n3497) );
  INV_X1 U4375 ( .A(n4414), .ZN(n3495) );
  INV_X1 U4376 ( .A(n3493), .ZN(n3494) );
  NAND2_X1 U4377 ( .A1(n3495), .A2(n3494), .ZN(n3496) );
  NAND2_X1 U4378 ( .A1(n3017), .A2(n4577), .ZN(n3498) );
  OAI21_X1 U4379 ( .B1(n3501), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3513), 
        .ZN(n6186) );
  AOI22_X1 U4380 ( .A1(n6186), .A2(n3753), .B1(n3885), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3503) );
  NAND2_X1 U4381 ( .A1(n3886), .A2(EAX_REG_3__SCAN_IN), .ZN(n3502) );
  OAI211_X1 U4382 ( .C1(n3511), .C2(n4481), .A(n3503), .B(n3502), .ZN(n3504)
         );
  INV_X1 U4383 ( .A(n3504), .ZN(n3505) );
  XNOR2_X1 U4384 ( .A(n3508), .B(n3507), .ZN(n4108) );
  NAND2_X1 U4385 ( .A1(n4108), .A2(n3547), .ZN(n3517) );
  NAND2_X1 U4386 ( .A1(n6475), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3510)
         );
  NAND2_X1 U4387 ( .A1(n3886), .A2(EAX_REG_4__SCAN_IN), .ZN(n3509) );
  OAI211_X1 U4388 ( .C1(n3511), .C2(n4353), .A(n3510), .B(n3509), .ZN(n3515)
         );
  AOI21_X1 U4389 ( .B1(n3513), .B2(n3512), .A(n3530), .ZN(n5529) );
  NOR2_X1 U4390 ( .A1(n5529), .A2(n3878), .ZN(n3514) );
  AOI21_X1 U4391 ( .B1(n3515), .B2(n3878), .A(n3514), .ZN(n3516) );
  NAND2_X1 U4392 ( .A1(n3517), .A2(n3516), .ZN(n4441) );
  AND3_X2 U4393 ( .A1(n4443), .A2(n4442), .A3(n4441), .ZN(n4613) );
  XOR2_X1 U4394 ( .A(n3518), .B(n3529), .Z(n4951) );
  INV_X1 U4395 ( .A(n3519), .ZN(n3524) );
  INV_X1 U4396 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4650) );
  INV_X1 U4397 ( .A(n3520), .ZN(n3521) );
  OAI21_X1 U4398 ( .B1(n3935), .B2(n4650), .A(n3521), .ZN(n3522) );
  INV_X1 U4399 ( .A(n3522), .ZN(n3523) );
  NAND2_X1 U4400 ( .A1(n4122), .A2(n3547), .ZN(n3526) );
  AOI22_X1 U4401 ( .A1(n3886), .A2(EAX_REG_6__SCAN_IN), .B1(n3885), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3525) );
  OAI211_X1 U4402 ( .C1(n4951), .C2(n3878), .A(n3526), .B(n3525), .ZN(n4557)
         );
  XNOR2_X1 U4403 ( .A(n3528), .B(n3527), .ZN(n4116) );
  NAND2_X1 U4404 ( .A1(n4116), .A2(n3547), .ZN(n3536) );
  INV_X1 U4405 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3533) );
  OAI21_X1 U4406 ( .B1(n3530), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3529), 
        .ZN(n6176) );
  NAND2_X1 U4407 ( .A1(n6176), .A2(n3753), .ZN(n3532) );
  NAND2_X1 U4408 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3531)
         );
  OAI211_X1 U4409 ( .C1(n3584), .C2(n3533), .A(n3532), .B(n3531), .ZN(n3534)
         );
  INV_X1 U4410 ( .A(n3534), .ZN(n3535) );
  NAND2_X1 U4411 ( .A1(n3536), .A2(n3535), .ZN(n4614) );
  XNOR2_X1 U4412 ( .A(n3556), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5719)
         );
  AOI22_X1 U4413 ( .A1(n3853), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3784), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4414 ( .A1(n3855), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4415 ( .A1(n3857), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4416 ( .A1(n3831), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4417 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3549)
         );
  AOI22_X1 U4418 ( .A1(n3696), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4419 ( .A1(n3666), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4420 ( .A1(n3789), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4421 ( .A1(n4483), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3543) );
  NAND4_X1 U4422 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3548)
         );
  OAI21_X1 U4423 ( .B1(n3549), .B2(n3548), .A(n3547), .ZN(n3552) );
  NAND2_X1 U4424 ( .A1(n3886), .A2(EAX_REG_15__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U4425 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3550)
         );
  NAND3_X1 U4426 ( .A1(n3552), .A2(n3551), .A3(n3550), .ZN(n3553) );
  AOI21_X1 U4427 ( .B1(n5719), .B2(n3753), .A(n3553), .ZN(n4917) );
  INV_X1 U4428 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6801) );
  AOI21_X1 U4429 ( .B1(n3557), .B2(n6801), .A(n3601), .ZN(n5711) );
  OR2_X1 U4430 ( .A1(n5711), .A2(n3878), .ZN(n3572) );
  AND2_X1 U4431 ( .A1(n3185), .A2(n3166), .ZN(n3558) );
  AOI22_X1 U4432 ( .A1(n3857), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3696), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4433 ( .A1(n3853), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3831), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4434 ( .A1(n3855), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4435 ( .A1(n3789), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4436 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3568)
         );
  AOI22_X1 U4437 ( .A1(n3666), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4438 ( .A1(n3836), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4439 ( .A1(n4483), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4440 ( .A1(n3784), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4441 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3567)
         );
  OR2_X1 U4442 ( .A1(n3568), .A2(n3567), .ZN(n3570) );
  INV_X1 U4443 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4321) );
  OAI22_X1 U4444 ( .A1(n3584), .A2(n4321), .B1(n3735), .B2(n6801), .ZN(n3569)
         );
  AOI21_X1 U4445 ( .B1(n3843), .B2(n3570), .A(n3569), .ZN(n3571) );
  NOR2_X2 U4446 ( .A1(n5020), .A2(n5019), .ZN(n5021) );
  INV_X1 U4447 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5262) );
  XNOR2_X1 U4448 ( .A(n3601), .B(n5262), .ZN(n5947) );
  AOI22_X1 U4449 ( .A1(n3696), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4450 ( .A1(n3857), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4451 ( .A1(n3853), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4452 ( .A1(n3856), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4453 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3582)
         );
  AOI22_X1 U4454 ( .A1(n3784), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4455 ( .A1(n3666), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4456 ( .A1(n3831), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4457 ( .A1(n4483), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3577) );
  NAND4_X1 U4458 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3581)
         );
  OR2_X1 U4459 ( .A1(n3582), .A2(n3581), .ZN(n3586) );
  INV_X1 U4460 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4398) );
  INV_X1 U4461 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6593) );
  OAI21_X1 U4462 ( .B1(n6593), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n6475), 
        .ZN(n3583) );
  OAI21_X1 U4463 ( .B1(n3584), .B2(n4398), .A(n3583), .ZN(n3585) );
  AOI21_X1 U4464 ( .B1(n3843), .B2(n3586), .A(n3585), .ZN(n3587) );
  AOI21_X1 U4465 ( .B1(n5947), .B2(n3753), .A(n3587), .ZN(n5243) );
  AND2_X2 U4466 ( .A1(n5021), .A2(n5243), .ZN(n5242) );
  AOI22_X1 U4467 ( .A1(n3857), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4468 ( .A1(n3855), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3784), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4469 ( .A1(n3831), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4470 ( .A1(n3856), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3588) );
  NAND4_X1 U4471 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3597)
         );
  AOI22_X1 U4472 ( .A1(n3853), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4473 ( .A1(n3696), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4474 ( .A1(n3866), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4475 ( .A1(n3229), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3592) );
  NAND4_X1 U4476 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3596)
         );
  NOR2_X1 U4477 ( .A1(n3597), .A2(n3596), .ZN(n3598) );
  OR2_X1 U4478 ( .A1(n3881), .A2(n3598), .ZN(n3610) );
  OAI21_X1 U4479 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6593), .A(n6475), 
        .ZN(n3599) );
  INV_X1 U4480 ( .A(n3599), .ZN(n3600) );
  AOI21_X1 U4481 ( .B1(n3886), .B2(EAX_REG_18__SCAN_IN), .A(n3600), .ZN(n3609)
         );
  INV_X1 U4482 ( .A(n3641), .ZN(n3607) );
  INV_X1 U4483 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3605) );
  INV_X1 U4484 ( .A(n3603), .ZN(n3604) );
  NAND2_X1 U4485 ( .A1(n3605), .A2(n3604), .ZN(n3606) );
  NAND2_X1 U4486 ( .A1(n3607), .A2(n3606), .ZN(n6023) );
  NOR2_X1 U4487 ( .A1(n6023), .A2(n3878), .ZN(n3608) );
  AOI21_X1 U4488 ( .B1(n3610), .B2(n3609), .A(n3608), .ZN(n5334) );
  NAND2_X1 U4489 ( .A1(n5242), .A2(n5334), .ZN(n5306) );
  AOI22_X1 U4490 ( .A1(n3855), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4491 ( .A1(n3666), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4492 ( .A1(n3789), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4493 ( .A1(n3784), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3611) );
  NAND4_X1 U4494 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(n3620)
         );
  AOI22_X1 U4495 ( .A1(n3853), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3831), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4496 ( .A1(n3857), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4497 ( .A1(n3696), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4498 ( .A1(n4483), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3615) );
  NAND4_X1 U4499 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3619)
         );
  NOR2_X1 U4500 ( .A1(n3620), .A2(n3619), .ZN(n3624) );
  NAND2_X1 U4501 ( .A1(n6475), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3621)
         );
  NAND2_X1 U4502 ( .A1(n3878), .A2(n3621), .ZN(n3622) );
  AOI21_X1 U4503 ( .B1(n3886), .B2(EAX_REG_19__SCAN_IN), .A(n3622), .ZN(n3623)
         );
  OAI21_X1 U4504 ( .B1(n3881), .B2(n3624), .A(n3623), .ZN(n3626) );
  INV_X1 U4505 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5701) );
  XNOR2_X1 U4506 ( .A(n3641), .B(n5701), .ZN(n5704) );
  NAND2_X1 U4507 ( .A1(n5704), .A2(n3753), .ZN(n3625) );
  NAND2_X1 U4508 ( .A1(n3626), .A2(n3625), .ZN(n5307) );
  OR2_X2 U4509 ( .A1(n5306), .A2(n5307), .ZN(n5689) );
  AOI22_X1 U4510 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3857), .B1(n3759), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4511 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3836), .B1(n3261), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4512 ( .A1(n3853), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4513 ( .A1(n3666), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4514 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3636)
         );
  AOI22_X1 U4515 ( .A1(n3696), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4516 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3784), .B1(n4483), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4517 ( .A1(n3856), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4518 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3229), .B1(n3863), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3631) );
  NAND4_X1 U4519 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n3635)
         );
  NOR2_X1 U4520 ( .A1(n3636), .A2(n3635), .ZN(n3640) );
  OAI21_X1 U4521 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6593), .A(n6475), 
        .ZN(n3637) );
  INV_X1 U4522 ( .A(n3637), .ZN(n3638) );
  AOI21_X1 U4523 ( .B1(n3886), .B2(EAX_REG_20__SCAN_IN), .A(n3638), .ZN(n3639)
         );
  OAI21_X1 U4524 ( .B1(n3881), .B2(n3640), .A(n3639), .ZN(n3646) );
  INV_X1 U4525 ( .A(n3643), .ZN(n3642) );
  INV_X1 U4526 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U4527 ( .A1(n3642), .A2(n5687), .ZN(n3644) );
  AND2_X1 U4528 ( .A1(n3644), .A2(n3677), .ZN(n5919) );
  NAND2_X1 U4529 ( .A1(n5919), .A2(n3946), .ZN(n3645) );
  NAND2_X1 U4530 ( .A1(n3646), .A2(n3645), .ZN(n5688) );
  AOI22_X1 U4531 ( .A1(n3696), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4532 ( .A1(n3784), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4533 ( .A1(n3836), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4534 ( .A1(n4483), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3647) );
  NAND4_X1 U4535 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(n3656)
         );
  AOI22_X1 U4536 ( .A1(n3857), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4537 ( .A1(n3666), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4538 ( .A1(n3856), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4539 ( .A1(n3853), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3651) );
  NAND4_X1 U4540 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3655)
         );
  NOR2_X1 U4541 ( .A1(n3656), .A2(n3655), .ZN(n3659) );
  INV_X1 U4542 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5910) );
  OAI21_X1 U4543 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5910), .A(n3878), .ZN(
        n3657) );
  AOI21_X1 U4544 ( .B1(n3886), .B2(EAX_REG_21__SCAN_IN), .A(n3657), .ZN(n3658)
         );
  OAI21_X1 U4545 ( .B1(n3881), .B2(n3659), .A(n3658), .ZN(n3661) );
  XNOR2_X1 U4546 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3677), .ZN(n5912)
         );
  NAND2_X1 U4547 ( .A1(n5912), .A2(n3946), .ZN(n3660) );
  NAND2_X1 U4548 ( .A1(n3661), .A2(n3660), .ZN(n5681) );
  AOI22_X1 U4549 ( .A1(n3853), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4550 ( .A1(n3784), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3831), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4551 ( .A1(n3229), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4552 ( .A1(n3759), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4553 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3672)
         );
  AOI22_X1 U4554 ( .A1(n3857), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3696), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4555 ( .A1(n3128), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4556 ( .A1(n3666), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4557 ( .A1(n3836), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3667) );
  NAND4_X1 U4558 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), .ZN(n3671)
         );
  NOR2_X1 U4559 ( .A1(n3672), .A2(n3671), .ZN(n3676) );
  NAND2_X1 U4560 ( .A1(n6475), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3673)
         );
  NAND2_X1 U4561 ( .A1(n3878), .A2(n3673), .ZN(n3674) );
  AOI21_X1 U4562 ( .B1(n3886), .B2(EAX_REG_22__SCAN_IN), .A(n3674), .ZN(n3675)
         );
  OAI21_X1 U4563 ( .B1(n3881), .B2(n3676), .A(n3675), .ZN(n3684) );
  INV_X1 U4564 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3681) );
  INV_X1 U4565 ( .A(n3679), .ZN(n3680) );
  NAND2_X1 U4566 ( .A1(n3681), .A2(n3680), .ZN(n3682) );
  NAND2_X1 U4567 ( .A1(n3711), .A2(n3682), .ZN(n5897) );
  NAND2_X1 U4568 ( .A1(n3684), .A2(n3683), .ZN(n5578) );
  NOR2_X2 U4569 ( .A1(n5691), .A2(n3685), .ZN(n5505) );
  AOI22_X1 U4570 ( .A1(n3857), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4571 ( .A1(n3831), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4572 ( .A1(n3856), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4573 ( .A1(n3830), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3686) );
  NAND4_X1 U4574 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n3695)
         );
  AOI22_X1 U4575 ( .A1(n3696), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4576 ( .A1(n3853), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4577 ( .A1(n3133), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4578 ( .A1(n3229), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3690) );
  NAND4_X1 U4579 ( .A1(n3693), .A2(n3692), .A3(n3691), .A4(n3690), .ZN(n3694)
         );
  NOR2_X1 U4580 ( .A1(n3695), .A2(n3694), .ZN(n3716) );
  AOI22_X1 U4581 ( .A1(n3696), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4582 ( .A1(n3857), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4583 ( .A1(n3829), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4584 ( .A1(n3856), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3697) );
  NAND4_X1 U4585 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3707)
         );
  AOI22_X1 U4586 ( .A1(n3784), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4587 ( .A1(n3229), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4588 ( .A1(n3831), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4589 ( .A1(n4483), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3702) );
  NAND4_X1 U4590 ( .A1(n3705), .A2(n3704), .A3(n3703), .A4(n3702), .ZN(n3706)
         );
  NOR2_X1 U4591 ( .A1(n3707), .A2(n3706), .ZN(n3717) );
  XOR2_X1 U4592 ( .A(n3716), .B(n3717), .Z(n3708) );
  NAND2_X1 U4593 ( .A1(n3708), .A2(n3843), .ZN(n3715) );
  INV_X1 U4594 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5510) );
  OAI21_X1 U4595 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5510), .A(n3878), .ZN(
        n3709) );
  AOI21_X1 U4596 ( .B1(n3886), .B2(EAX_REG_23__SCAN_IN), .A(n3709), .ZN(n3714)
         );
  NAND2_X1 U4597 ( .A1(n3711), .A2(n5510), .ZN(n3712) );
  NAND2_X1 U4598 ( .A1(n3732), .A2(n3712), .ZN(n5665) );
  NOR2_X1 U4599 ( .A1(n5665), .A2(n3878), .ZN(n3713) );
  AOI21_X1 U4600 ( .B1(n3715), .B2(n3714), .A(n3713), .ZN(n5504) );
  AND2_X2 U4601 ( .A1(n5505), .A2(n5504), .ZN(n5429) );
  NOR2_X1 U4602 ( .A1(n3717), .A2(n3716), .ZN(n3740) );
  AOI22_X1 U4603 ( .A1(n3241), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4604 ( .A1(n3857), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4605 ( .A1(n3829), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4606 ( .A1(n3856), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4607 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3728)
         );
  AOI22_X1 U4608 ( .A1(n3784), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4609 ( .A1(n3864), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4610 ( .A1(n3261), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4611 ( .A1(n3866), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3723) );
  NAND4_X1 U4612 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3727)
         );
  OR2_X1 U4613 ( .A1(n3728), .A2(n3727), .ZN(n3739) );
  INV_X1 U4614 ( .A(n3739), .ZN(n3729) );
  XNOR2_X1 U4615 ( .A(n3740), .B(n3729), .ZN(n3730) );
  NAND2_X1 U4616 ( .A1(n3730), .A2(n3843), .ZN(n3738) );
  INV_X1 U4617 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U4618 ( .A1(n3732), .A2(n6806), .ZN(n3733) );
  NAND2_X1 U4619 ( .A1(n3775), .A2(n3733), .ZN(n5495) );
  NAND2_X1 U4620 ( .A1(n5495), .A2(n3753), .ZN(n3734) );
  OAI21_X1 U4621 ( .B1(n6806), .B2(n3735), .A(n3734), .ZN(n3736) );
  AOI21_X1 U4622 ( .B1(n3886), .B2(EAX_REG_24__SCAN_IN), .A(n3736), .ZN(n3737)
         );
  NAND2_X1 U4623 ( .A1(n3738), .A2(n3737), .ZN(n5428) );
  AND2_X2 U4624 ( .A1(n5429), .A2(n5428), .ZN(n5484) );
  NAND2_X1 U4625 ( .A1(n3740), .A2(n3739), .ZN(n3757) );
  AOI22_X1 U4626 ( .A1(n3784), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4627 ( .A1(n3229), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4628 ( .A1(n3855), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4629 ( .A1(n3866), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3741) );
  NAND4_X1 U4630 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3750)
         );
  AOI22_X1 U4631 ( .A1(n3857), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4632 ( .A1(n3241), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4633 ( .A1(n3856), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4634 ( .A1(n3261), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4635 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3749)
         );
  NOR2_X1 U4636 ( .A1(n3750), .A2(n3749), .ZN(n3758) );
  XOR2_X1 U4637 ( .A(n3757), .B(n3758), .Z(n3751) );
  NAND2_X1 U4638 ( .A1(n3751), .A2(n3843), .ZN(n3756) );
  INV_X1 U4639 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5653) );
  AOI21_X1 U4640 ( .B1(n5653), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3752) );
  AOI21_X1 U4641 ( .B1(n3886), .B2(EAX_REG_25__SCAN_IN), .A(n3752), .ZN(n3755)
         );
  XNOR2_X1 U4642 ( .A(n3775), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5657)
         );
  AOI21_X1 U4643 ( .B1(n3756), .B2(n3755), .A(n3754), .ZN(n5483) );
  NAND2_X2 U4644 ( .A1(n5484), .A2(n5483), .ZN(n5482) );
  NOR2_X1 U4645 ( .A1(n3758), .A2(n3757), .ZN(n3783) );
  AOI22_X1 U4646 ( .A1(n3241), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4647 ( .A1(n3857), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3759), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4648 ( .A1(n3829), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4649 ( .A1(n3856), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3761) );
  NAND4_X1 U4650 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3770)
         );
  AOI22_X1 U4651 ( .A1(n3784), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4652 ( .A1(n3864), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4653 ( .A1(n3831), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4654 ( .A1(n3866), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4655 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3769)
         );
  OR2_X1 U4656 ( .A1(n3770), .A2(n3769), .ZN(n3782) );
  INV_X1 U4657 ( .A(n3782), .ZN(n3771) );
  XNOR2_X1 U4658 ( .A(n3783), .B(n3771), .ZN(n3774) );
  INV_X1 U4659 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3776) );
  NAND2_X1 U4660 ( .A1(n3886), .A2(EAX_REG_26__SCAN_IN), .ZN(n3772) );
  OAI211_X1 U4661 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n3776), .A(n3772), .B(
        n3878), .ZN(n3773) );
  AOI21_X1 U4662 ( .B1(n3774), .B2(n3843), .A(n3773), .ZN(n3780) );
  NAND2_X1 U4663 ( .A1(n3777), .A2(n3776), .ZN(n3778) );
  NAND2_X1 U4664 ( .A1(n3821), .A2(n3778), .ZN(n5647) );
  NOR2_X1 U4665 ( .A1(n5647), .A2(n3878), .ZN(n3779) );
  NOR2_X2 U4666 ( .A1(n5482), .A2(n5469), .ZN(n3781) );
  INV_X1 U4667 ( .A(n3781), .ZN(n5559) );
  NAND2_X1 U4668 ( .A1(n3783), .A2(n3782), .ZN(n3803) );
  AOI22_X1 U4669 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3784), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4670 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3831), .B1(n3830), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4671 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3855), .B1(n3854), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4672 ( .A1(n3856), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4673 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3795)
         );
  AOI22_X1 U4674 ( .A1(n3857), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4675 ( .A1(n3696), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4676 ( .A1(n3866), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4677 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3229), .B1(n3863), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4678 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3794)
         );
  NOR2_X1 U4679 ( .A1(n3795), .A2(n3794), .ZN(n3804) );
  XOR2_X1 U4680 ( .A(n3803), .B(n3804), .Z(n3796) );
  NAND2_X1 U4681 ( .A1(n3796), .A2(n3843), .ZN(n3800) );
  INV_X1 U4682 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5887) );
  NOR2_X1 U4683 ( .A1(n5887), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3797) );
  OR2_X1 U4684 ( .A1(n3797), .A2(n3946), .ZN(n3798) );
  AOI21_X1 U4685 ( .B1(n3886), .B2(EAX_REG_27__SCAN_IN), .A(n3798), .ZN(n3799)
         );
  NAND2_X1 U4686 ( .A1(n3800), .A2(n3799), .ZN(n3802) );
  XNOR2_X1 U4687 ( .A(n3821), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5885)
         );
  NAND2_X1 U4688 ( .A1(n5885), .A2(n3946), .ZN(n3801) );
  NAND2_X1 U4689 ( .A1(n3802), .A2(n3801), .ZN(n5560) );
  NOR2_X2 U4690 ( .A1(n5559), .A2(n5560), .ZN(n5455) );
  NOR2_X1 U4691 ( .A1(n3804), .A2(n3803), .ZN(n3827) );
  AOI22_X1 U4692 ( .A1(n3241), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4693 ( .A1(n3857), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4694 ( .A1(n3829), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4695 ( .A1(n3856), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4696 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3814)
         );
  AOI22_X1 U4697 ( .A1(n3133), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4698 ( .A1(n3864), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4699 ( .A1(n3261), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4700 ( .A1(n3866), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4701 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3813)
         );
  OR2_X1 U4702 ( .A1(n3814), .A2(n3813), .ZN(n3826) );
  INV_X1 U4703 ( .A(n3826), .ZN(n3815) );
  XNOR2_X1 U4704 ( .A(n3827), .B(n3815), .ZN(n3816) );
  NAND2_X1 U4705 ( .A1(n3816), .A2(n3843), .ZN(n3825) );
  NAND2_X1 U4706 ( .A1(n6475), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3817)
         );
  NAND2_X1 U4707 ( .A1(n3878), .A2(n3817), .ZN(n3818) );
  AOI21_X1 U4708 ( .B1(n3886), .B2(EAX_REG_28__SCAN_IN), .A(n3818), .ZN(n3824)
         );
  AND2_X1 U4709 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3819) );
  INV_X1 U4710 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5461) );
  OAI21_X1 U4711 ( .B1(n3821), .B2(n5887), .A(n5461), .ZN(n3822) );
  NAND2_X1 U4712 ( .A1(n3849), .A2(n3822), .ZN(n5633) );
  NOR2_X1 U4713 ( .A1(n5633), .A2(n3878), .ZN(n3823) );
  AOI21_X1 U4714 ( .B1(n3825), .B2(n3824), .A(n3823), .ZN(n5456) );
  NAND2_X1 U4715 ( .A1(n5455), .A2(n5456), .ZN(n5445) );
  NAND2_X1 U4716 ( .A1(n3827), .A2(n3826), .ZN(n3873) );
  AOI22_X1 U4717 ( .A1(n3241), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3789), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4718 ( .A1(n3857), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3829), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4719 ( .A1(n3229), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3830), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4720 ( .A1(n3831), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4483), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3832) );
  NAND4_X1 U4721 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3842)
         );
  AOI22_X1 U4722 ( .A1(n3133), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4723 ( .A1(n3855), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4724 ( .A1(n3856), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4725 ( .A1(n3214), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4726 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3841)
         );
  NOR2_X1 U4727 ( .A1(n3842), .A2(n3841), .ZN(n3874) );
  XOR2_X1 U4728 ( .A(n3873), .B(n3874), .Z(n3844) );
  NAND2_X1 U4729 ( .A1(n3844), .A2(n3843), .ZN(n3847) );
  INV_X1 U4730 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6654) );
  AOI21_X1 U4731 ( .B1(n6654), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3845) );
  AOI21_X1 U4732 ( .B1(n3886), .B2(EAX_REG_29__SCAN_IN), .A(n3845), .ZN(n3846)
         );
  NAND2_X1 U4733 ( .A1(n3847), .A2(n3846), .ZN(n3852) );
  NAND2_X1 U4734 ( .A1(n3849), .A2(n6654), .ZN(n3850) );
  NAND2_X1 U4735 ( .A1(n3948), .A2(n3850), .ZN(n5621) );
  NAND2_X1 U4736 ( .A1(n3852), .A2(n3851), .ZN(n5446) );
  OR2_X2 U4737 ( .A1(n5445), .A2(n5446), .ZN(n5448) );
  AOI22_X1 U4738 ( .A1(n3853), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4739 ( .A1(n3133), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4740 ( .A1(n3855), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4741 ( .A1(n3857), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3856), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4742 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3872)
         );
  AOI22_X1 U4743 ( .A1(n3696), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4744 ( .A1(n3128), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3718), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4745 ( .A1(n3864), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4746 ( .A1(n3866), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4747 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3871)
         );
  NOR2_X1 U4748 ( .A1(n3872), .A2(n3871), .ZN(n3876) );
  NOR2_X1 U4749 ( .A1(n3874), .A2(n3873), .ZN(n3875) );
  XOR2_X1 U4750 ( .A(n3876), .B(n3875), .Z(n3882) );
  NAND2_X1 U4751 ( .A1(n6475), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3877)
         );
  NAND2_X1 U4752 ( .A1(n3878), .A2(n3877), .ZN(n3879) );
  AOI21_X1 U4753 ( .B1(n3886), .B2(EAX_REG_30__SCAN_IN), .A(n3879), .ZN(n3880)
         );
  OAI21_X1 U4754 ( .B1(n3882), .B2(n3881), .A(n3880), .ZN(n3884) );
  XNOR2_X1 U4755 ( .A(n3948), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5438)
         );
  NAND2_X1 U4756 ( .A1(n5438), .A2(n3946), .ZN(n3883) );
  NAND2_X1 U4757 ( .A1(n3884), .A2(n3883), .ZN(n4278) );
  NOR2_X2 U4758 ( .A1(n5448), .A2(n4278), .ZN(n3888) );
  AOI22_X1 U4759 ( .A1(n3886), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n3885), .ZN(n3887) );
  XNOR2_X1 U4760 ( .A(n3888), .B(n3887), .ZN(n5588) );
  XNOR2_X1 U4761 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3901) );
  NAND2_X1 U4762 ( .A1(n3913), .A2(n3901), .ZN(n3891) );
  NAND2_X1 U4763 ( .A1(n6456), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4764 ( .A1(n3891), .A2(n3890), .ZN(n3900) );
  XNOR2_X1 U4765 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3898) );
  NAND2_X1 U4766 ( .A1(n3900), .A2(n3898), .ZN(n3893) );
  NAND2_X1 U4767 ( .A1(n6460), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3892) );
  XNOR2_X1 U4768 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3895) );
  NOR2_X1 U4769 ( .A1(n4481), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3894)
         );
  NAND2_X1 U4770 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3905), .ZN(n3938) );
  INV_X1 U4771 ( .A(n3895), .ZN(n3896) );
  XNOR2_X1 U4772 ( .A(n3897), .B(n3896), .ZN(n3929) );
  INV_X1 U4773 ( .A(n3898), .ZN(n3899) );
  XNOR2_X1 U4774 ( .A(n3900), .B(n3899), .ZN(n3911) );
  XOR2_X1 U4775 ( .A(n3913), .B(n3901), .Z(n3912) );
  AND2_X1 U4776 ( .A1(n3911), .A2(n3912), .ZN(n3902) );
  NAND2_X1 U4777 ( .A1(n3909), .A2(n3902), .ZN(n3907) );
  OR2_X1 U4778 ( .A1(n3903), .A2(n4353), .ZN(n3904) );
  NAND2_X1 U4779 ( .A1(n3907), .A2(n3942), .ZN(n4293) );
  NOR2_X1 U4780 ( .A1(n4252), .A2(n4293), .ZN(n4286) );
  NAND2_X1 U4781 ( .A1(n4286), .A2(n6490), .ZN(n4301) );
  NAND2_X1 U4782 ( .A1(n3185), .A2(n4205), .ZN(n4147) );
  INV_X1 U4783 ( .A(n3942), .ZN(n3908) );
  NAND2_X1 U4784 ( .A1(n3936), .A2(n3908), .ZN(n3945) );
  INV_X1 U4785 ( .A(n3909), .ZN(n3934) );
  AND2_X1 U4786 ( .A1(n4538), .A2(n3185), .ZN(n3910) );
  NAND2_X1 U4787 ( .A1(n3920), .A2(n3911), .ZN(n3927) );
  OAI211_X1 U4788 ( .C1(n3911), .C2(n3935), .A(n3928), .B(n3927), .ZN(n3932)
         );
  AOI21_X1 U4789 ( .B1(n3920), .B2(n4205), .A(n3012), .ZN(n3926) );
  NAND2_X1 U4790 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3912), .ZN(n3925) );
  INV_X1 U4791 ( .A(n3912), .ZN(n3918) );
  INV_X1 U4792 ( .A(n4185), .ZN(n3916) );
  INV_X1 U4793 ( .A(n3913), .ZN(n3914) );
  OAI21_X1 U4794 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6447), .A(n3914), 
        .ZN(n3919) );
  OAI21_X1 U4795 ( .B1(n3916), .B2(n3919), .A(n3915), .ZN(n3917) );
  AOI22_X1 U4796 ( .A1(n3928), .A2(n3917), .B1(n3926), .B2(n3925), .ZN(n3921)
         );
  OAI21_X1 U4797 ( .B1(n3918), .B2(n3921), .A(n3936), .ZN(n3924) );
  INV_X1 U4798 ( .A(n3919), .ZN(n3922) );
  NAND3_X1 U4799 ( .A1(n3922), .A2(n3921), .A3(n3920), .ZN(n3923) );
  OAI211_X1 U4800 ( .C1(n3926), .C2(n3925), .A(n3924), .B(n3923), .ZN(n3931)
         );
  OAI22_X1 U4801 ( .A1(n3929), .A2(n4147), .B1(n3928), .B2(n3927), .ZN(n3930)
         );
  AOI21_X1 U4802 ( .B1(n3932), .B2(n3931), .A(n3930), .ZN(n3933) );
  AOI21_X1 U4803 ( .B1(n3935), .B2(n3934), .A(n3933), .ZN(n3940) );
  INV_X1 U4804 ( .A(n3936), .ZN(n3937) );
  OAI22_X1 U4805 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4353), .B1(n3938), .B2(
        n3937), .ZN(n3939) );
  NOR2_X1 U4806 ( .A1(n3940), .A2(n3939), .ZN(n3941) );
  NAND2_X1 U4807 ( .A1(n4370), .A2(n4307), .ZN(n4299) );
  NOR2_X1 U4808 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6338) );
  NAND2_X1 U4809 ( .A1(n6382), .A2(n6480), .ZN(n5997) );
  NAND2_X1 U4810 ( .A1(n6596), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6603) );
  INV_X1 U4811 ( .A(n6603), .ZN(n4187) );
  AND2_X1 U4812 ( .A1(n3946), .A2(n4187), .ZN(n6487) );
  INV_X1 U4813 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U4814 ( .A1(n6480), .A2(n6475), .ZN(n6595) );
  NOR3_X1 U4815 ( .A1(n6596), .A2(n6571), .A3(n6595), .ZN(n6482) );
  OR2_X1 U4816 ( .A1(n6487), .A2(n6482), .ZN(n3947) );
  INV_X1 U4817 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4279) );
  NAND2_X1 U4818 ( .A1(n5588), .A2(n6615), .ZN(n4073) );
  BUF_X4 U4819 ( .A(n4031), .Z(n4027) );
  NAND2_X1 U4820 ( .A1(n4931), .A2(n4205), .ZN(n3962) );
  NAND2_X1 U4821 ( .A1(n3962), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3953)
         );
  INV_X1 U4822 ( .A(n4080), .ZN(n4549) );
  NAND2_X1 U4823 ( .A1(n4549), .A2(n4931), .ZN(n3963) );
  NAND2_X1 U4824 ( .A1(n3951), .A2(EBX_REG_1__SCAN_IN), .ZN(n3952) );
  NAND2_X1 U4825 ( .A1(n3963), .A2(EBX_REG_0__SCAN_IN), .ZN(n3956) );
  INV_X1 U4826 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U4827 ( .A1(n4031), .A2(n4524), .ZN(n3955) );
  NAND2_X1 U4828 ( .A1(n3956), .A2(n3955), .ZN(n4361) );
  INV_X1 U4829 ( .A(n4361), .ZN(n3957) );
  NOR2_X1 U4830 ( .A1(n3958), .A2(n3957), .ZN(n3959) );
  AOI21_X2 U4831 ( .B1(n5034), .B2(n4448), .A(n3959), .ZN(n4574) );
  MUX2_X1 U4832 ( .A(n4031), .B(n4036), .S(EBX_REG_2__SCAN_IN), .Z(n3961) );
  NAND2_X1 U4833 ( .A1(n4054), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3960)
         );
  NAND2_X1 U4834 ( .A1(n3961), .A2(n3960), .ZN(n4573) );
  NAND2_X1 U4835 ( .A1(n4574), .A2(n4573), .ZN(n5176) );
  INV_X1 U4836 ( .A(n5176), .ZN(n3967) );
  NAND2_X1 U4837 ( .A1(n5312), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3964)
         );
  OAI211_X1 U4838 ( .C1(n4054), .C2(EBX_REG_3__SCAN_IN), .A(n4036), .B(n3964), 
        .ZN(n3965) );
  OAI21_X1 U4839 ( .B1(n4034), .B2(EBX_REG_3__SCAN_IN), .A(n3965), .ZN(n5175)
         );
  NAND2_X1 U4840 ( .A1(n3967), .A2(n3966), .ZN(n5178) );
  INV_X1 U4841 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U4842 ( .A1(n4036), .A2(n6800), .ZN(n3969) );
  INV_X1 U4843 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4456) );
  NAND2_X1 U4844 ( .A1(n4448), .A2(n4456), .ZN(n3968) );
  NAND3_X1 U4845 ( .A1(n3969), .A2(n4027), .A3(n3968), .ZN(n3971) );
  NAND2_X1 U4846 ( .A1(n5800), .A2(n4456), .ZN(n3970) );
  MUX2_X1 U4847 ( .A(n4034), .B(n4027), .S(EBX_REG_5__SCAN_IN), .Z(n3973) );
  INV_X1 U4848 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U4849 ( .A1(n4360), .A2(n6231), .ZN(n3972) );
  INV_X1 U4850 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U4851 ( .A1(n4036), .A2(n6237), .ZN(n3975) );
  INV_X1 U4852 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U4853 ( .A1(n4448), .A2(n5048), .ZN(n3974) );
  NAND3_X1 U4854 ( .A1(n3975), .A2(n4027), .A3(n3974), .ZN(n3977) );
  NAND2_X1 U4855 ( .A1(n5800), .A2(n5048), .ZN(n3976) );
  NAND2_X1 U4856 ( .A1(n3977), .A2(n3976), .ZN(n4559) );
  NAND2_X1 U4857 ( .A1(n4678), .A2(n4559), .ZN(n6051) );
  NAND2_X1 U4858 ( .A1(n5312), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3978)
         );
  OAI211_X1 U4859 ( .C1(n4054), .C2(EBX_REG_7__SCAN_IN), .A(n4036), .B(n3978), 
        .ZN(n3979) );
  OAI21_X1 U4860 ( .B1(n4034), .B2(EBX_REG_7__SCAN_IN), .A(n3979), .ZN(n6050)
         );
  INV_X1 U4861 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U4862 ( .A1(n4036), .A2(n4990), .ZN(n3981) );
  INV_X1 U4863 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U4864 ( .A1(n4448), .A2(n4940), .ZN(n3980) );
  NAND3_X1 U4865 ( .A1(n3981), .A2(n4027), .A3(n3980), .ZN(n3983) );
  NAND2_X1 U4866 ( .A1(n5800), .A2(n4940), .ZN(n3982) );
  MUX2_X1 U4867 ( .A(n4034), .B(n4027), .S(EBX_REG_9__SCAN_IN), .Z(n3985) );
  INV_X1 U4868 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U4869 ( .A1(n4360), .A2(n5286), .ZN(n3984) );
  AND2_X1 U4870 ( .A1(n3985), .A2(n3984), .ZN(n4978) );
  INV_X1 U4871 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4159) );
  NAND2_X1 U4872 ( .A1(n4036), .A2(n4159), .ZN(n3987) );
  INV_X1 U4873 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U4874 ( .A1(n4448), .A2(n6036), .ZN(n3986) );
  NAND3_X1 U4875 ( .A1(n3987), .A2(n4027), .A3(n3986), .ZN(n3989) );
  NAND2_X1 U4876 ( .A1(n5800), .A2(n6036), .ZN(n3988) );
  NAND2_X1 U4877 ( .A1(n3989), .A2(n3988), .ZN(n5238) );
  NAND2_X1 U4878 ( .A1(n4977), .A2(n5238), .ZN(n4960) );
  MUX2_X1 U4879 ( .A(n4034), .B(n4027), .S(EBX_REG_11__SCAN_IN), .Z(n3991) );
  INV_X1 U4880 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6792) );
  NAND2_X1 U4881 ( .A1(n4360), .A2(n6792), .ZN(n3990) );
  NAND2_X1 U4882 ( .A1(n3991), .A2(n3990), .ZN(n4961) );
  INV_X1 U4883 ( .A(n4034), .ZN(n4047) );
  INV_X1 U4884 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U4885 ( .A1(n4047), .A2(n6645), .ZN(n3994) );
  NAND2_X1 U4886 ( .A1(n4031), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3992) );
  OAI211_X1 U4887 ( .C1(n4054), .C2(EBX_REG_13__SCAN_IN), .A(n4036), .B(n3992), 
        .ZN(n3993) );
  AND2_X1 U4888 ( .A1(n3994), .A2(n3993), .ZN(n5108) );
  MUX2_X1 U4889 ( .A(n4027), .B(n4036), .S(EBX_REG_12__SCAN_IN), .Z(n3996) );
  NAND2_X1 U4890 ( .A1(n4054), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3995) );
  NAND2_X1 U4891 ( .A1(n3996), .A2(n3995), .ZN(n5169) );
  NAND2_X1 U4892 ( .A1(n5108), .A2(n5169), .ZN(n3997) );
  NOR2_X2 U4893 ( .A1(n5170), .A2(n3997), .ZN(n5110) );
  MUX2_X1 U4894 ( .A(n4027), .B(n4036), .S(EBX_REG_14__SCAN_IN), .Z(n3999) );
  NAND2_X1 U4895 ( .A1(n4054), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3998) );
  NAND2_X1 U4896 ( .A1(n3999), .A2(n3998), .ZN(n4907) );
  NAND2_X1 U4897 ( .A1(n5110), .A2(n4907), .ZN(n4919) );
  NAND2_X1 U4898 ( .A1(n5312), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4000) );
  OAI211_X1 U4899 ( .C1(n4054), .C2(EBX_REG_15__SCAN_IN), .A(n4036), .B(n4000), 
        .ZN(n4001) );
  OAI21_X1 U4900 ( .B1(n4034), .B2(EBX_REG_15__SCAN_IN), .A(n4001), .ZN(n4920)
         );
  OR2_X2 U4901 ( .A1(n4919), .A2(n4920), .ZN(n5024) );
  MUX2_X1 U4902 ( .A(n4031), .B(n4036), .S(EBX_REG_16__SCAN_IN), .Z(n4003) );
  NAND2_X1 U4903 ( .A1(n4054), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4002) );
  AND2_X1 U4904 ( .A1(n4003), .A2(n4002), .ZN(n5025) );
  OR2_X2 U4905 ( .A1(n5024), .A2(n5025), .ZN(n5246) );
  MUX2_X1 U4906 ( .A(n4034), .B(n4027), .S(EBX_REG_17__SCAN_IN), .Z(n4005) );
  INV_X1 U4907 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U4908 ( .A1(n4360), .A2(n5952), .ZN(n4004) );
  NAND2_X1 U4909 ( .A1(n4005), .A2(n4004), .ZN(n5247) );
  NOR2_X4 U4910 ( .A1(n5246), .A2(n5247), .ZN(n5331) );
  MUX2_X1 U4911 ( .A(n4027), .B(n4036), .S(EBX_REG_19__SCAN_IN), .Z(n4007) );
  NAND2_X1 U4912 ( .A1(n4054), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4006) );
  NAND2_X1 U4913 ( .A1(n4007), .A2(n4006), .ZN(n5314) );
  AND2_X2 U4914 ( .A1(n5331), .A2(n5314), .ZN(n5798) );
  INV_X1 U4915 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5416) );
  NOR2_X1 U4916 ( .A1(n4054), .A2(EBX_REG_20__SCAN_IN), .ZN(n4008) );
  AOI21_X1 U4917 ( .B1(n4360), .B2(n5416), .A(n4008), .ZN(n5801) );
  INV_X1 U4918 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U4919 ( .A1(n4360), .A2(n5957), .ZN(n4009) );
  INV_X1 U4920 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U4921 ( .A1(n4448), .A2(n5338), .ZN(n5310) );
  NAND2_X1 U4922 ( .A1(n4009), .A2(n5310), .ZN(n5311) );
  NAND2_X1 U4923 ( .A1(n5800), .A2(EBX_REG_20__SCAN_IN), .ZN(n4011) );
  NAND2_X1 U4924 ( .A1(n5311), .A2(n5312), .ZN(n4010) );
  OAI211_X1 U4925 ( .C1(n5801), .C2(n5311), .A(n4011), .B(n4010), .ZN(n4012)
         );
  INV_X1 U4926 ( .A(n4012), .ZN(n4013) );
  NAND2_X1 U4927 ( .A1(n5798), .A2(n4013), .ZN(n5784) );
  NAND2_X1 U4928 ( .A1(n5312), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4014) );
  OAI211_X1 U4929 ( .C1(n4054), .C2(EBX_REG_21__SCAN_IN), .A(n4036), .B(n4014), 
        .ZN(n4015) );
  OAI21_X1 U4930 ( .B1(n4034), .B2(EBX_REG_21__SCAN_IN), .A(n4015), .ZN(n5783)
         );
  OR2_X2 U4931 ( .A1(n5784), .A2(n5783), .ZN(n5582) );
  MUX2_X1 U4932 ( .A(n4034), .B(n4027), .S(EBX_REG_23__SCAN_IN), .Z(n4017) );
  INV_X1 U4933 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U4934 ( .A1(n4360), .A2(n5769), .ZN(n4016) );
  AND2_X1 U4935 ( .A1(n4017), .A2(n4016), .ZN(n5507) );
  MUX2_X1 U4936 ( .A(n4027), .B(n4036), .S(EBX_REG_22__SCAN_IN), .Z(n4019) );
  NAND2_X1 U4937 ( .A1(n4054), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4018) );
  NAND2_X1 U4938 ( .A1(n4019), .A2(n4018), .ZN(n5581) );
  NAND2_X1 U4939 ( .A1(n5507), .A2(n5581), .ZN(n4020) );
  MUX2_X1 U4940 ( .A(n4031), .B(n4036), .S(EBX_REG_24__SCAN_IN), .Z(n4022) );
  NAND2_X1 U4941 ( .A1(n4054), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4021) );
  NAND2_X1 U4942 ( .A1(n4022), .A2(n4021), .ZN(n5422) );
  INV_X1 U4943 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U4944 ( .A1(n4047), .A2(n5571), .ZN(n4025) );
  NAND2_X1 U4945 ( .A1(n5312), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4023) );
  OAI211_X1 U4946 ( .C1(n4054), .C2(EBX_REG_25__SCAN_IN), .A(n4036), .B(n4023), 
        .ZN(n4024) );
  AND2_X1 U4947 ( .A1(n4025), .A2(n4024), .ZN(n5479) );
  NAND2_X1 U4948 ( .A1(n5421), .A2(n5479), .ZN(n5481) );
  INV_X1 U4949 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U4950 ( .A1(n4036), .A2(n5629), .ZN(n4028) );
  INV_X1 U4951 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U4952 ( .A1(n4448), .A2(n5568), .ZN(n4026) );
  NAND3_X1 U4953 ( .A1(n4028), .A2(n4027), .A3(n4026), .ZN(n4030) );
  NAND2_X1 U4954 ( .A1(n5800), .A2(n5568), .ZN(n4029) );
  AND2_X1 U4955 ( .A1(n4030), .A2(n4029), .ZN(n5472) );
  OR2_X2 U4956 ( .A1(n5481), .A2(n5472), .ZN(n5562) );
  NAND2_X1 U4957 ( .A1(n4031), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4032) );
  OAI211_X1 U4958 ( .C1(n4054), .C2(EBX_REG_27__SCAN_IN), .A(n4036), .B(n4032), 
        .ZN(n4033) );
  OAI21_X1 U4959 ( .B1(n4034), .B2(EBX_REG_27__SCAN_IN), .A(n4033), .ZN(n5561)
         );
  INV_X1 U4960 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U4961 ( .A1(n4036), .A2(n4035), .ZN(n4037) );
  OAI211_X1 U4962 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4054), .A(n4037), .B(n5312), 
        .ZN(n4039) );
  INV_X1 U4963 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U4964 ( .A1(n5800), .A2(n5557), .ZN(n4038) );
  NAND2_X1 U4965 ( .A1(n4039), .A2(n4038), .ZN(n5460) );
  NAND2_X1 U4966 ( .A1(n5564), .A2(n5460), .ZN(n4041) );
  INV_X1 U4967 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5728) );
  AND2_X1 U4968 ( .A1(n4360), .A2(n5728), .ZN(n4044) );
  NOR2_X1 U4969 ( .A1(n4054), .A2(EBX_REG_29__SCAN_IN), .ZN(n4040) );
  OR3_X2 U4970 ( .A1(n4041), .A2(n4044), .A3(n4040), .ZN(n4228) );
  AND2_X2 U4971 ( .A1(n4228), .A2(n5312), .ZN(n4224) );
  INV_X1 U4972 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5554) );
  OR2_X1 U4973 ( .A1(n4360), .A2(n5554), .ZN(n4043) );
  NAND2_X1 U4974 ( .A1(n4054), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4042) );
  NAND2_X1 U4975 ( .A1(n4043), .A2(n4042), .ZN(n4227) );
  INV_X1 U4976 ( .A(n4044), .ZN(n4046) );
  INV_X1 U4977 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4045) );
  MUX2_X1 U4978 ( .A(n4046), .B(n4045), .S(n5800), .Z(n4049) );
  NAND2_X1 U4979 ( .A1(n4047), .A2(n4045), .ZN(n4048) );
  NAND2_X1 U4980 ( .A1(n4049), .A2(n4048), .ZN(n5449) );
  NOR3_X1 U4981 ( .A1(n5459), .A2(n4227), .A3(n5449), .ZN(n4050) );
  INV_X1 U4982 ( .A(n4360), .ZN(n4051) );
  OAI22_X1 U4983 ( .A1(n4051), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4054), .ZN(n4052) );
  NAND2_X1 U4984 ( .A1(n5006), .A2(EBX_REG_31__SCAN_IN), .ZN(n4060) );
  INV_X1 U4985 ( .A(n4060), .ZN(n4056) );
  NOR2_X1 U4986 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4929) );
  NOR2_X1 U4987 ( .A1(n4054), .A2(n4929), .ZN(n4055) );
  NAND3_X1 U4988 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4066) );
  NAND2_X1 U4989 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5317) );
  INV_X1 U4990 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U4991 ( .A1(n4057), .A2(n6509), .ZN(n6504) );
  NAND2_X1 U4992 ( .A1(n4538), .A2(n6504), .ZN(n4211) );
  AND3_X1 U4993 ( .A1(n4211), .A2(n4929), .A3(n4931), .ZN(n4058) );
  INV_X1 U4994 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6623) );
  INV_X1 U4995 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6520) );
  INV_X1 U4996 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6522) );
  NOR2_X1 U4997 ( .A1(n6520), .A2(n6522), .ZN(n5045) );
  NAND4_X1 U4998 ( .A1(n5045), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_8__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n4925) );
  NAND3_X1 U4999 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n4927) );
  NOR2_X1 U5000 ( .A1(n4925), .A2(n4927), .ZN(n5055) );
  NAND2_X1 U5001 ( .A1(n5055), .A2(REIP_REG_9__SCAN_IN), .ZN(n6039) );
  INV_X1 U5002 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6532) );
  NOR2_X1 U5003 ( .A1(n6039), .A2(n6532), .ZN(n4967) );
  NAND2_X1 U5004 ( .A1(n4967), .A2(REIP_REG_11__SCAN_IN), .ZN(n4965) );
  INV_X1 U5005 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6534) );
  NOR2_X1 U5006 ( .A1(n4965), .A2(n6534), .ZN(n5517) );
  NAND2_X1 U5007 ( .A1(n5517), .A2(REIP_REG_13__SCAN_IN), .ZN(n6607) );
  NOR2_X1 U5008 ( .A1(n6623), .A2(n6607), .ZN(n4064) );
  NAND4_X1 U5009 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5259), .ZN(n6018) );
  NOR2_X1 U5010 ( .A1(n5317), .A2(n6018), .ZN(n5918) );
  NAND2_X1 U5011 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5918), .ZN(n5915) );
  NOR2_X1 U5012 ( .A1(n4066), .A2(n5915), .ZN(n5486) );
  AND3_X1 U5013 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4068) );
  NAND2_X1 U5014 ( .A1(n5486), .A2(n4068), .ZN(n5896) );
  NAND2_X1 U5015 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4069) );
  INV_X1 U5016 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6564) );
  INV_X1 U5017 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6557) );
  NOR4_X1 U5018 ( .A1(n5437), .A2(REIP_REG_31__SCAN_IN), .A3(n6564), .A4(n6557), .ZN(n4062) );
  INV_X1 U5019 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6773) );
  INV_X1 U5020 ( .A(n4929), .ZN(n4059) );
  OR2_X1 U5021 ( .A1(n6504), .A2(n4059), .ZN(n6478) );
  NAND2_X1 U5022 ( .A1(n6594), .A2(n6478), .ZN(n4933) );
  OAI22_X1 U5023 ( .A1(n6773), .A2(n6619), .B1(n4060), .B2(n4933), .ZN(n4061)
         );
  AOI211_X1 U5024 ( .C1(n5367), .C2(n6058), .A(n4062), .B(n4061), .ZN(n4071)
         );
  INV_X1 U5025 ( .A(n5437), .ZN(n4063) );
  NAND2_X1 U5026 ( .A1(n4063), .A2(n6557), .ZN(n5453) );
  NAND2_X1 U5027 ( .A1(n6608), .A2(n4966), .ZN(n5899) );
  INV_X1 U5028 ( .A(n5899), .ZN(n5547) );
  NAND2_X1 U5029 ( .A1(n4064), .A2(n4966), .ZN(n5028) );
  NAND3_X1 U5030 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4065) );
  NOR2_X1 U5031 ( .A1(n5028), .A2(n4065), .ZN(n5261) );
  NAND4_X1 U5032 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        n5261), .A4(REIP_REG_18__SCAN_IN), .ZN(n5898) );
  NOR2_X1 U5033 ( .A1(n5898), .A2(n4066), .ZN(n4067) );
  OR2_X1 U5034 ( .A1(n4067), .A2(n5547), .ZN(n5499) );
  OAI21_X1 U5035 ( .B1(n5547), .B2(n4068), .A(n5499), .ZN(n5889) );
  AOI21_X1 U5036 ( .B1(n6025), .B2(n4069), .A(n5889), .ZN(n5464) );
  NAND2_X1 U5037 ( .A1(n5453), .A2(n5464), .ZN(n5443) );
  AOI21_X1 U5038 ( .B1(n6025), .B2(n6564), .A(n5443), .ZN(n4070) );
  INV_X1 U5039 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4193) );
  NAND2_X1 U5040 ( .A1(n4073), .A2(n4072), .ZN(U2796) );
  NAND2_X1 U5041 ( .A1(n4092), .A2(n4093), .ZN(n4091) );
  NAND2_X1 U5042 ( .A1(n4091), .A2(n4079), .ZN(n4110) );
  INV_X1 U5043 ( .A(n4109), .ZN(n4074) );
  XNOR2_X1 U5044 ( .A(n4110), .B(n4074), .ZN(n4075) );
  NAND2_X1 U5045 ( .A1(n4075), .A2(n6594), .ZN(n4076) );
  INV_X1 U5046 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6268) );
  XNOR2_X1 U5047 ( .A(n4106), .B(n6268), .ZN(n6178) );
  INV_X1 U5048 ( .A(n4147), .ZN(n4137) );
  NAND2_X1 U5049 ( .A1(n4078), .A2(n4137), .ZN(n4084) );
  XNOR2_X1 U5050 ( .A(n4091), .B(n4079), .ZN(n4082) );
  NAND2_X1 U5051 ( .A1(n4553), .A2(n4080), .ZN(n4085) );
  INV_X1 U5052 ( .A(n4085), .ZN(n4081) );
  AOI21_X1 U5053 ( .B1(n4082), .B2(n6594), .A(n4081), .ZN(n4083) );
  NAND2_X1 U5054 ( .A1(n4084), .A2(n4083), .ZN(n6189) );
  NAND2_X1 U5055 ( .A1(n6189), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4101)
         );
  INV_X1 U5056 ( .A(n6594), .ZN(n4220) );
  OAI21_X1 U5057 ( .B1(n4220), .B2(n4093), .A(n4085), .ZN(n4086) );
  INV_X1 U5058 ( .A(n4086), .ZN(n4087) );
  OAI21_X2 U5059 ( .B1(n4841), .B2(n4147), .A(n4087), .ZN(n4359) );
  NAND2_X1 U5060 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4088)
         );
  INV_X1 U5061 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U5062 ( .A1(n4088), .A2(n5382), .ZN(n4090) );
  AND2_X1 U5063 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4089) );
  NAND2_X1 U5064 ( .A1(n4359), .A2(n4089), .ZN(n4099) );
  AND2_X1 U5065 ( .A1(n4090), .A2(n4099), .ZN(n4355) );
  NAND2_X1 U5066 ( .A1(n4519), .A2(n4137), .ZN(n4098) );
  OAI21_X1 U5067 ( .B1(n4093), .B2(n4092), .A(n4091), .ZN(n4095) );
  OAI211_X1 U5068 ( .C1(n4095), .C2(n4220), .A(n4236), .B(n3185), .ZN(n4096)
         );
  INV_X1 U5069 ( .A(n4096), .ZN(n4097) );
  NAND2_X1 U5070 ( .A1(n4098), .A2(n4097), .ZN(n4354) );
  INV_X1 U5071 ( .A(n4099), .ZN(n4100) );
  NAND2_X1 U5072 ( .A1(n4101), .A2(n6188), .ZN(n4105) );
  INV_X1 U5073 ( .A(n6189), .ZN(n4103) );
  INV_X1 U5074 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4102) );
  NAND2_X1 U5075 ( .A1(n4103), .A2(n4102), .ZN(n4104) );
  NAND2_X1 U5076 ( .A1(n4106), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4107)
         );
  NAND2_X1 U5077 ( .A1(n6180), .A2(n4107), .ZN(n4618) );
  NAND2_X1 U5078 ( .A1(n4108), .A2(n4137), .ZN(n4113) );
  NAND2_X1 U5079 ( .A1(n4110), .A2(n4109), .ZN(n4126) );
  XNOR2_X1 U5080 ( .A(n4126), .B(n4124), .ZN(n4111) );
  NAND2_X1 U5081 ( .A1(n4111), .A2(n6594), .ZN(n4112) );
  NAND2_X1 U5082 ( .A1(n4113), .A2(n4112), .ZN(n4114) );
  XNOR2_X1 U5083 ( .A(n4114), .B(n6800), .ZN(n4617) );
  NAND2_X1 U5084 ( .A1(n4618), .A2(n4617), .ZN(n4616) );
  NAND2_X1 U5085 ( .A1(n4114), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4115)
         );
  NAND2_X1 U5086 ( .A1(n4616), .A2(n4115), .ZN(n6170) );
  NAND2_X1 U5087 ( .A1(n4116), .A2(n4137), .ZN(n4121) );
  INV_X1 U5088 ( .A(n4124), .ZN(n4117) );
  OR2_X1 U5089 ( .A1(n4126), .A2(n4117), .ZN(n4118) );
  XNOR2_X1 U5090 ( .A(n4118), .B(n4123), .ZN(n4119) );
  NAND2_X1 U5091 ( .A1(n4119), .A2(n6594), .ZN(n4120) );
  NAND2_X1 U5092 ( .A1(n4121), .A2(n4120), .ZN(n4130) );
  XNOR2_X1 U5093 ( .A(n4130), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6171)
         );
  NOR2_X1 U5094 ( .A1(n6170), .A2(n6171), .ZN(n4945) );
  INV_X1 U5095 ( .A(n4945), .ZN(n4134) );
  NAND3_X1 U5096 ( .A1(n4122), .A2(n4150), .A3(n4137), .ZN(n4129) );
  NAND2_X1 U5097 ( .A1(n4124), .A2(n4123), .ZN(n4125) );
  OR2_X1 U5098 ( .A1(n4126), .A2(n4125), .ZN(n4139) );
  XNOR2_X1 U5099 ( .A(n4139), .B(n4140), .ZN(n4127) );
  NAND2_X1 U5100 ( .A1(n4127), .A2(n6594), .ZN(n4128) );
  XNOR2_X1 U5101 ( .A(n4135), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4950)
         );
  INV_X1 U5102 ( .A(n4130), .ZN(n4131) );
  NAND2_X1 U5103 ( .A1(n4131), .A2(n6231), .ZN(n4946) );
  INV_X1 U5104 ( .A(n4946), .ZN(n4132) );
  NOR2_X1 U5105 ( .A1(n4950), .A2(n4132), .ZN(n4133) );
  NAND2_X1 U5106 ( .A1(n4134), .A2(n4133), .ZN(n4947) );
  NAND2_X1 U5107 ( .A1(n4135), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4136)
         );
  NAND2_X1 U5108 ( .A1(n4947), .A2(n4136), .ZN(n6163) );
  NAND2_X1 U5109 ( .A1(n4138), .A2(n4137), .ZN(n4144) );
  INV_X1 U5110 ( .A(n4139), .ZN(n4141) );
  NAND2_X1 U5111 ( .A1(n4141), .A2(n4140), .ZN(n4153) );
  XNOR2_X1 U5112 ( .A(n4153), .B(n4151), .ZN(n4142) );
  NAND2_X1 U5113 ( .A1(n4142), .A2(n6594), .ZN(n4143) );
  NAND2_X1 U5114 ( .A1(n4144), .A2(n4143), .ZN(n4145) );
  INV_X1 U5115 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6220) );
  XNOR2_X1 U5116 ( .A(n4145), .B(n6220), .ZN(n6162) );
  NAND2_X1 U5117 ( .A1(n6163), .A2(n6162), .ZN(n6161) );
  NAND2_X1 U5118 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4146)
         );
  NAND2_X1 U5119 ( .A1(n6161), .A2(n4146), .ZN(n4984) );
  NOR2_X1 U5120 ( .A1(n4148), .A2(n4147), .ZN(n4149) );
  INV_X1 U5121 ( .A(n4151), .ZN(n4152) );
  OR3_X1 U5122 ( .A1(n4153), .A2(n4152), .A3(n4220), .ZN(n4154) );
  NAND2_X1 U5123 ( .A1(n5818), .A2(n4154), .ZN(n4155) );
  XNOR2_X1 U5124 ( .A(n4155), .B(n4990), .ZN(n4983) );
  NAND2_X1 U5125 ( .A1(n4155), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5268)
         );
  OR2_X1 U5126 ( .A1(n5625), .A2(n5286), .ZN(n5278) );
  OR2_X1 U5127 ( .A1(n5625), .A2(n4159), .ZN(n5342) );
  OR2_X1 U5128 ( .A1(n5625), .A2(n6792), .ZN(n4156) );
  AND2_X1 U5129 ( .A1(n5342), .A2(n4156), .ZN(n4157) );
  AND2_X1 U5130 ( .A1(n5278), .A2(n4157), .ZN(n4158) );
  AND2_X1 U5131 ( .A1(n5268), .A2(n4158), .ZN(n4161) );
  NAND2_X1 U5132 ( .A1(n5818), .A2(n5286), .ZN(n5276) );
  NAND2_X1 U5133 ( .A1(n5818), .A2(n4159), .ZN(n5340) );
  AND2_X1 U5134 ( .A1(n5340), .A2(n3028), .ZN(n4160) );
  INV_X1 U5135 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4258) );
  NOR2_X1 U5136 ( .A1(n5818), .A2(n4258), .ZN(n5294) );
  NAND2_X1 U5137 ( .A1(n5818), .A2(n4258), .ZN(n5292) );
  OAI21_X1 U5138 ( .B1(n5291), .B2(n5294), .A(n5292), .ZN(n5353) );
  XNOR2_X1 U5139 ( .A(n5818), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5354)
         );
  NAND2_X1 U5140 ( .A1(n5353), .A2(n5354), .ZN(n4164) );
  INV_X1 U5141 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4162) );
  NAND2_X1 U5142 ( .A1(n5818), .A2(n4162), .ZN(n4163) );
  NAND2_X1 U5143 ( .A1(n4164), .A2(n4163), .ZN(n5359) );
  INV_X1 U5144 ( .A(n5359), .ZN(n4166) );
  INV_X1 U5145 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5980) );
  INV_X1 U5146 ( .A(n5361), .ZN(n4165) );
  NAND2_X1 U5147 ( .A1(n4166), .A2(n4165), .ZN(n4167) );
  NAND2_X1 U5148 ( .A1(n4167), .A2(n5360), .ZN(n5716) );
  INV_X1 U5149 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5717) );
  NOR2_X1 U5150 ( .A1(n5818), .A2(n5717), .ZN(n4169) );
  NAND2_X1 U5151 ( .A1(n5818), .A2(n5717), .ZN(n4168) );
  INV_X1 U5152 ( .A(n4170), .ZN(n5708) );
  INV_X1 U5153 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U5154 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4270) );
  OAI21_X1 U5155 ( .B1(n5831), .B2(n4270), .A(n5818), .ZN(n4171) );
  AND3_X1 U5156 ( .A1(n5831), .A2(n5952), .A3(n5957), .ZN(n4172) );
  AND2_X1 U5157 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5805) );
  AND2_X1 U5158 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5660) );
  AND2_X1 U5159 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4272) );
  NAND3_X1 U5160 ( .A1(n5805), .A2(n5660), .A3(n4272), .ZN(n4174) );
  NAND2_X1 U5161 ( .A1(n5818), .A2(n4174), .ZN(n4175) );
  NAND2_X1 U5162 ( .A1(n5695), .A2(n4175), .ZN(n4178) );
  NOR2_X1 U5163 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5804) );
  NOR2_X1 U5164 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5776) );
  INV_X1 U5165 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6671) );
  NAND4_X1 U5166 ( .A1(n5804), .A2(n5776), .A3(n6671), .A4(n5769), .ZN(n4176)
         );
  NAND2_X1 U5167 ( .A1(n3024), .A2(n4176), .ZN(n4177) );
  INV_X1 U5168 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5627) );
  XNOR2_X1 U5169 ( .A(n5818), .B(n5627), .ZN(n5652) );
  NOR2_X1 U5170 ( .A1(n3024), .A2(n5629), .ZN(n5644) );
  NAND2_X1 U5171 ( .A1(n5616), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4198) );
  INV_X1 U5172 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4266) );
  NOR2_X1 U5173 ( .A1(n5818), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5643)
         );
  NOR2_X1 U5174 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U5175 ( .A1(n5643), .A2(n5734), .ZN(n5617) );
  NOR2_X1 U5176 ( .A1(n5617), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4197)
         );
  NAND3_X1 U5177 ( .A1(n4180), .A2(n4197), .A3(n4266), .ZN(n4181) );
  XNOR2_X1 U5178 ( .A(n4182), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5378)
         );
  NAND2_X1 U5179 ( .A1(n5399), .A2(n4553), .ZN(n4183) );
  NAND2_X1 U5180 ( .A1(n4184), .A2(n4183), .ZN(n4216) );
  OR2_X1 U5181 ( .A1(n4216), .A2(n4185), .ZN(n6467) );
  INV_X1 U5182 ( .A(n6467), .ZN(n4186) );
  NAND2_X1 U5183 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4187), .ZN(n6497) );
  INV_X1 U5184 ( .A(n6497), .ZN(n4188) );
  NAND2_X1 U5185 ( .A1(n5588), .A2(n6181), .ZN(n4196) );
  NAND2_X1 U5186 ( .A1(n6388), .A2(n4189), .ZN(n6599) );
  NAND2_X1 U5187 ( .A1(n6599), .A2(n6596), .ZN(n4190) );
  NAND2_X1 U5188 ( .A1(n6596), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4192) );
  NAND2_X1 U5189 ( .A1(n6593), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4191) );
  AND2_X1 U5190 ( .A1(n4192), .A2(n4191), .ZN(n4435) );
  NOR2_X1 U5191 ( .A1(n6254), .A2(n4193), .ZN(n5373) );
  NOR2_X1 U5192 ( .A1(n5702), .A2(n6773), .ZN(n4194) );
  AOI211_X1 U5193 ( .C1(n5946), .C2(n4935), .A(n5373), .B(n4194), .ZN(n4195)
         );
  OAI211_X1 U5194 ( .C1(n5378), .C2(n6165), .A(n4196), .B(n4195), .ZN(U2955)
         );
  INV_X1 U5195 ( .A(n4197), .ZN(n4199) );
  OAI21_X1 U5196 ( .B1(n3014), .B2(n4199), .A(n4198), .ZN(n4200) );
  NAND2_X1 U5197 ( .A1(n4252), .A2(n4216), .ZN(n4204) );
  INV_X1 U5198 ( .A(n3165), .ZN(n4202) );
  AND2_X1 U5199 ( .A1(n3165), .A2(n4931), .ZN(n4201) );
  OAI22_X1 U5200 ( .A1(n4203), .A2(n4202), .B1(n4201), .B2(n6594), .ZN(n4241)
         );
  NAND2_X1 U5201 ( .A1(n4204), .A2(n4241), .ZN(n4339) );
  NOR2_X1 U5202 ( .A1(n5399), .A2(n4538), .ZN(n4249) );
  NAND2_X1 U5203 ( .A1(n4465), .A2(n4249), .ZN(n4208) );
  NAND2_X1 U5204 ( .A1(n4205), .A2(n6504), .ZN(n4206) );
  NOR2_X1 U5205 ( .A1(READY_N), .A2(n4293), .ZN(n4343) );
  NAND3_X1 U5206 ( .A1(n4206), .A2(n4343), .A3(n4235), .ZN(n4207) );
  NAND2_X1 U5207 ( .A1(n4208), .A2(n4207), .ZN(n4209) );
  OAI21_X1 U5208 ( .B1(n4339), .B2(n4209), .A(n6490), .ZN(n4215) );
  INV_X1 U5209 ( .A(READY_N), .ZN(n6590) );
  NAND2_X1 U5210 ( .A1(n4211), .A2(n6590), .ZN(n4212) );
  OAI211_X1 U5211 ( .C1(n4470), .C2(n4212), .A(n4931), .B(n5324), .ZN(n4213)
         );
  NAND3_X1 U5212 ( .A1(n4370), .A2(n3154), .A3(n4213), .ZN(n4214) );
  OR2_X1 U5213 ( .A1(n4216), .A2(n4287), .ZN(n4475) );
  AND2_X1 U5214 ( .A1(n6467), .A2(n4475), .ZN(n4218) );
  INV_X1 U5215 ( .A(n4307), .ZN(n4292) );
  OR2_X1 U5216 ( .A1(n4292), .A2(n4538), .ZN(n4337) );
  NAND2_X1 U5217 ( .A1(n4221), .A2(n3166), .ZN(n4217) );
  NAND4_X1 U5218 ( .A1(n4473), .A2(n4218), .A3(n4337), .A4(n4217), .ZN(n4219)
         );
  NAND2_X1 U5219 ( .A1(n4277), .A2(n6277), .ZN(n4276) );
  OR2_X1 U5220 ( .A1(n4470), .A2(n4220), .ZN(n6479) );
  NAND2_X1 U5221 ( .A1(n4221), .A2(n3018), .ZN(n4222) );
  NAND2_X1 U5222 ( .A1(n6479), .A2(n4222), .ZN(n4223) );
  NAND2_X1 U5223 ( .A1(n4255), .A2(n4223), .ZN(n6255) );
  INV_X1 U5224 ( .A(n4224), .ZN(n4232) );
  INV_X1 U5225 ( .A(n5459), .ZN(n4226) );
  INV_X1 U5226 ( .A(n4227), .ZN(n4225) );
  AOI21_X1 U5227 ( .B1(n4228), .B2(n4226), .A(n4225), .ZN(n4231) );
  AOI21_X1 U5228 ( .B1(n5459), .B2(n5800), .A(n4227), .ZN(n4229) );
  AND2_X1 U5229 ( .A1(n4229), .A2(n4228), .ZN(n4230) );
  AOI21_X1 U5230 ( .B1(n4232), .B2(n4231), .A(n4230), .ZN(n5552) );
  NOR2_X1 U5231 ( .A1(n6254), .A2(n6564), .ZN(n4281) );
  OAI21_X1 U5232 ( .B1(n3154), .B2(n4234), .A(n4233), .ZN(n4238) );
  OR2_X1 U5233 ( .A1(n4290), .A2(n4235), .ZN(n4340) );
  AOI21_X1 U5234 ( .B1(n4360), .B2(n4340), .A(n4236), .ZN(n4237) );
  NOR2_X1 U5235 ( .A1(n4238), .A2(n4237), .ZN(n4242) );
  NAND2_X1 U5236 ( .A1(n4239), .A2(n5800), .ZN(n4240) );
  NAND4_X1 U5237 ( .A1(n4243), .A2(n4242), .A3(n4241), .A4(n4240), .ZN(n4472)
         );
  INV_X1 U5238 ( .A(n3175), .ZN(n4247) );
  NAND2_X1 U5239 ( .A1(n5390), .A2(n4244), .ZN(n4495) );
  NAND2_X1 U5240 ( .A1(n4245), .A2(n5800), .ZN(n4246) );
  OAI211_X1 U5241 ( .C1(n4468), .C2(n4247), .A(n4495), .B(n4246), .ZN(n4248)
         );
  NOR2_X1 U5242 ( .A1(n4472), .A2(n4248), .ZN(n4250) );
  INV_X1 U5243 ( .A(n4250), .ZN(n4251) );
  NAND2_X1 U5244 ( .A1(n4255), .A2(n4251), .ZN(n4263) );
  NAND2_X1 U5245 ( .A1(n6250), .A2(n4263), .ZN(n5972) );
  NOR2_X1 U5246 ( .A1(n4252), .A2(n4538), .ZN(n6448) );
  NAND2_X1 U5247 ( .A1(n4255), .A2(n6448), .ZN(n5974) );
  INV_X1 U5248 ( .A(n6227), .ZN(n5369) );
  NAND2_X1 U5249 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4273) );
  NAND2_X1 U5250 ( .A1(n4263), .A2(n5974), .ZN(n6224) );
  NOR2_X1 U5251 ( .A1(n6800), .A2(n6268), .ZN(n6252) );
  INV_X1 U5252 ( .A(n6252), .ZN(n6242) );
  NAND2_X1 U5253 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4254) );
  NOR2_X1 U5254 ( .A1(n6242), .A2(n4254), .ZN(n4986) );
  NAND3_X1 U5255 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4986), .ZN(n4989) );
  NOR2_X1 U5256 ( .A1(n4990), .A2(n6220), .ZN(n5285) );
  NAND3_X1 U5257 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n5285), .ZN(n4257) );
  NOR2_X1 U5258 ( .A1(n4989), .A2(n4257), .ZN(n4268) );
  INV_X1 U5259 ( .A(n4268), .ZN(n5968) );
  INV_X1 U5260 ( .A(n6250), .ZN(n6275) );
  INV_X1 U5261 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U5262 ( .A1(n5384), .A2(n5972), .ZN(n4363) );
  INV_X1 U5263 ( .A(n4255), .ZN(n4256) );
  NAND2_X1 U5264 ( .A1(n4256), .A2(n6254), .ZN(n4365) );
  NAND2_X1 U5265 ( .A1(n4363), .A2(n4365), .ZN(n6222) );
  NOR2_X1 U5266 ( .A1(n6275), .A2(n6222), .ZN(n5794) );
  INV_X1 U5267 ( .A(n5794), .ZN(n4988) );
  NAND2_X1 U5268 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U5269 ( .A1(n4102), .A2(n6271), .ZN(n6270) );
  NAND2_X1 U5270 ( .A1(n6252), .A2(n6270), .ZN(n6230) );
  NAND3_X1 U5271 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6238), .ZN(n4987) );
  AOI22_X1 U5272 ( .A1(n6224), .A2(n5968), .B1(n4988), .B2(n5969), .ZN(n6204)
         );
  INV_X1 U5273 ( .A(n6204), .ZN(n5970) );
  NAND2_X1 U5274 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5828) );
  NOR2_X1 U5275 ( .A1(n4258), .A2(n6792), .ZN(n5297) );
  INV_X1 U5276 ( .A(n5297), .ZN(n5971) );
  NOR2_X1 U5277 ( .A1(n4162), .A2(n5971), .ZN(n5975) );
  NAND2_X1 U5278 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5975), .ZN(n5830) );
  OAI21_X1 U5279 ( .B1(n5828), .B2(n5830), .A(n6227), .ZN(n4259) );
  INV_X1 U5280 ( .A(n4259), .ZN(n4260) );
  NOR2_X1 U5281 ( .A1(n5970), .A2(n4260), .ZN(n5824) );
  INV_X1 U5282 ( .A(n5805), .ZN(n4271) );
  OAI21_X1 U5283 ( .B1(n4271), .B2(n4270), .A(n6227), .ZN(n4261) );
  INV_X1 U5284 ( .A(n5660), .ZN(n5778) );
  NAND2_X1 U5285 ( .A1(n6227), .A2(n5778), .ZN(n4262) );
  NOR2_X1 U5286 ( .A1(n4263), .A2(n5384), .ZN(n5976) );
  INV_X1 U5287 ( .A(n4272), .ZN(n4264) );
  OAI21_X1 U5288 ( .B1(n6280), .B2(n6275), .A(n4264), .ZN(n4265) );
  NAND2_X1 U5289 ( .A1(n5767), .A2(n4265), .ZN(n5761) );
  AOI21_X1 U5290 ( .B1(n6227), .B2(n4273), .A(n5761), .ZN(n5742) );
  OAI21_X1 U5291 ( .B1(n4253), .B2(n5369), .A(n5742), .ZN(n5727) );
  AOI21_X1 U5292 ( .B1(n5728), .B2(n6227), .A(n5727), .ZN(n5368) );
  NOR2_X1 U5293 ( .A1(n5368), .A2(n4266), .ZN(n4267) );
  AOI211_X1 U5294 ( .C1(n6273), .C2(n5552), .A(n4281), .B(n4267), .ZN(n4274)
         );
  NAND2_X1 U5295 ( .A1(n4268), .A2(n6280), .ZN(n5793) );
  NAND2_X1 U5296 ( .A1(n5969), .A2(n5793), .ZN(n6200) );
  NAND2_X1 U5297 ( .A1(n5975), .A2(n6200), .ZN(n5981) );
  AND2_X1 U5298 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4269) );
  NAND2_X1 U5299 ( .A1(n5959), .A2(n4269), .ZN(n5951) );
  NAND2_X1 U5300 ( .A1(n5770), .A2(n4272), .ZN(n5758) );
  NAND3_X1 U5301 ( .A1(n5746), .A2(n4253), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U5302 ( .A1(n4276), .A2(n4275), .ZN(U2988) );
  NAND2_X1 U5303 ( .A1(n4277), .A2(n6193), .ZN(n4285) );
  XNOR2_X2 U5304 ( .A(n5448), .B(n4278), .ZN(n5593) );
  NOR2_X1 U5305 ( .A1(n5702), .A2(n4279), .ZN(n4280) );
  AOI211_X1 U5306 ( .C1(n5946), .C2(n5438), .A(n4281), .B(n4280), .ZN(n4282)
         );
  NAND2_X1 U5307 ( .A1(n4285), .A2(n4284), .ZN(U2956) );
  OR2_X1 U5308 ( .A1(n4286), .A2(n4307), .ZN(n4289) );
  NAND2_X1 U5309 ( .A1(n4465), .A2(n4287), .ZN(n4288) );
  AND2_X1 U5310 ( .A1(n4289), .A2(n4288), .ZN(n5993) );
  INV_X1 U5311 ( .A(n4290), .ZN(n5005) );
  OR2_X1 U5312 ( .A1(n5005), .A2(n6594), .ZN(n4305) );
  NAND2_X1 U5313 ( .A1(n4305), .A2(n6504), .ZN(n6591) );
  NAND2_X1 U5314 ( .A1(n6591), .A2(n6590), .ZN(n4291) );
  NAND2_X1 U5315 ( .A1(n5993), .A2(n4291), .ZN(n6469) );
  AND2_X1 U5316 ( .A1(n6469), .A2(n6490), .ZN(n6002) );
  INV_X1 U5317 ( .A(MORE_REG_SCAN_IN), .ZN(n4298) );
  INV_X1 U5318 ( .A(n4477), .ZN(n4296) );
  NAND3_X1 U5319 ( .A1(n4292), .A2(n6467), .A3(n4475), .ZN(n4294) );
  AOI22_X1 U5320 ( .A1(n4294), .A2(n4465), .B1(n3889), .B2(n4293), .ZN(n4295)
         );
  OAI21_X1 U5321 ( .B1(n4296), .B2(n4465), .A(n4295), .ZN(n6471) );
  NAND2_X1 U5322 ( .A1(n6471), .A2(n6002), .ZN(n4297) );
  OAI21_X1 U5323 ( .B1(n6002), .B2(n4298), .A(n4297), .ZN(U3471) );
  NAND2_X1 U5324 ( .A1(n4299), .A2(n5997), .ZN(n4302) );
  AOI21_X1 U5325 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n4301), .A(n4302), .ZN(
        n4300) );
  INV_X1 U5326 ( .A(n4300), .ZN(U2788) );
  INV_X1 U5327 ( .A(n4301), .ZN(n4303) );
  NOR3_X1 U5328 ( .A1(n4303), .A2(READREQUEST_REG_SCAN_IN), .A3(n4302), .ZN(
        n4304) );
  AOI21_X1 U5329 ( .B1(n6598), .B2(n4305), .A(n4304), .ZN(U3474) );
  INV_X1 U5330 ( .A(n6479), .ZN(n4306) );
  INV_X1 U5331 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4311) );
  AND2_X1 U5332 ( .A1(n4307), .A2(n6590), .ZN(n4308) );
  NAND2_X1 U5333 ( .A1(n4370), .A2(n4308), .ZN(n4309) );
  NAND2_X1 U5334 ( .A1(n6157), .A2(DATAI_9_), .ZN(n4395) );
  NAND2_X1 U5335 ( .A1(n6156), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4310) );
  OAI211_X1 U5336 ( .C1(n6159), .C2(n4311), .A(n4395), .B(n4310), .ZN(U2933)
         );
  INV_X1 U5337 ( .A(EAX_REG_10__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U5338 ( .A1(n6157), .A2(DATAI_10_), .ZN(n4406) );
  NAND2_X1 U5339 ( .A1(n6156), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4312) );
  OAI211_X1 U5340 ( .C1(n6159), .C2(n4313), .A(n4406), .B(n4312), .ZN(U2949)
         );
  INV_X1 U5341 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4315) );
  INV_X1 U5342 ( .A(DATAI_2_), .ZN(n4430) );
  OR2_X1 U5343 ( .A1(n4422), .A2(n4430), .ZN(n4408) );
  NAND2_X1 U5344 ( .A1(n6156), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4314) );
  OAI211_X1 U5345 ( .C1(n6159), .C2(n4315), .A(n4408), .B(n4314), .ZN(U2941)
         );
  INV_X1 U5346 ( .A(DATAI_0_), .ZN(n4518) );
  OR2_X1 U5347 ( .A1(n4422), .A2(n4518), .ZN(n4320) );
  NAND2_X1 U5348 ( .A1(n6156), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4316) );
  OAI211_X1 U5349 ( .C1(n6159), .C2(n6136), .A(n4320), .B(n4316), .ZN(U2939)
         );
  INV_X1 U5350 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U5351 ( .A1(n6157), .A2(DATAI_6_), .ZN(n4411) );
  NAND2_X1 U5352 ( .A1(n6156), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4317) );
  OAI211_X1 U5353 ( .C1(n6159), .C2(n4318), .A(n4411), .B(n4317), .ZN(U2930)
         );
  NAND2_X1 U5354 ( .A1(n6156), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4319) );
  OAI211_X1 U5355 ( .C1(n6159), .C2(n4321), .A(n4320), .B(n4319), .ZN(U2924)
         );
  INV_X1 U5356 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n4323) );
  INV_X1 U5357 ( .A(DATAI_5_), .ZN(n4615) );
  NOR2_X1 U5358 ( .A1(n4422), .A2(n4615), .ZN(n4326) );
  AOI21_X1 U5359 ( .B1(n6153), .B2(EAX_REG_5__SCAN_IN), .A(n4326), .ZN(n4322)
         );
  OAI21_X1 U5360 ( .B1(n6143), .B2(n4323), .A(n4322), .ZN(U2944) );
  INV_X1 U5361 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n4325) );
  INV_X1 U5362 ( .A(DATAI_7_), .ZN(n4682) );
  NOR2_X1 U5363 ( .A1(n4422), .A2(n4682), .ZN(n4329) );
  AOI21_X1 U5364 ( .B1(n6153), .B2(EAX_REG_7__SCAN_IN), .A(n4329), .ZN(n4324)
         );
  OAI21_X1 U5365 ( .B1(n6143), .B2(n4325), .A(n4324), .ZN(U2946) );
  INV_X1 U5366 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4328) );
  AOI21_X1 U5367 ( .B1(n6153), .B2(EAX_REG_21__SCAN_IN), .A(n4326), .ZN(n4327)
         );
  OAI21_X1 U5368 ( .B1(n6143), .B2(n4328), .A(n4327), .ZN(U2929) );
  INV_X1 U5369 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4331) );
  AOI21_X1 U5370 ( .B1(n6153), .B2(EAX_REG_23__SCAN_IN), .A(n4329), .ZN(n4330)
         );
  OAI21_X1 U5371 ( .B1(n6143), .B2(n4331), .A(n4330), .ZN(U2931) );
  INV_X1 U5372 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4333) );
  INV_X1 U5373 ( .A(DATAI_3_), .ZN(n4431) );
  NOR2_X1 U5374 ( .A1(n4422), .A2(n4431), .ZN(n4334) );
  AOI21_X1 U5375 ( .B1(n6153), .B2(EAX_REG_3__SCAN_IN), .A(n4334), .ZN(n4332)
         );
  OAI21_X1 U5376 ( .B1(n6143), .B2(n4333), .A(n4332), .ZN(U2942) );
  INV_X1 U5377 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4336) );
  AOI21_X1 U5378 ( .B1(n6153), .B2(EAX_REG_19__SCAN_IN), .A(n4334), .ZN(n4335)
         );
  OAI21_X1 U5379 ( .B1(n6143), .B2(n4336), .A(n4335), .ZN(U2927) );
  NOR2_X1 U5380 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6571), .ZN(n4528) );
  AOI211_X1 U5381 ( .C1(n4337), .C2(n6504), .A(READY_N), .B(n4465), .ZN(n4338)
         );
  OAI21_X1 U5382 ( .B1(n6448), .B2(n4210), .A(n4338), .ZN(n4342) );
  INV_X1 U5383 ( .A(n4339), .ZN(n4341) );
  NAND3_X1 U5384 ( .A1(n4342), .A2(n4341), .A3(n4340), .ZN(n4345) );
  INV_X1 U5385 ( .A(n4343), .ZN(n4344) );
  OAI22_X1 U5386 ( .A1(n4473), .A2(n4344), .B1(n4465), .B2(n4475), .ZN(n4416)
         );
  NOR2_X1 U5387 ( .A1(n4345), .A2(n4416), .ZN(n4346) );
  NAND2_X1 U5388 ( .A1(n4477), .A2(n4465), .ZN(n4446) );
  INV_X1 U5389 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6001) );
  NOR2_X1 U5390 ( .A1(n6480), .A2(n6475), .ZN(n4513) );
  NAND2_X1 U5391 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4513), .ZN(n6569) );
  OAI22_X1 U5392 ( .A1(n6452), .A2(n5994), .B1(n6001), .B2(n6569), .ZN(n4351)
         );
  NOR2_X1 U5393 ( .A1(n4528), .A2(n4351), .ZN(n6578) );
  INV_X1 U5394 ( .A(n6578), .ZN(n5412) );
  INV_X1 U5395 ( .A(n6294), .ZN(n4347) );
  OR2_X1 U5396 ( .A1(n4348), .A2(n4347), .ZN(n4349) );
  XNOR2_X1 U5397 ( .A(n4349), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5538)
         );
  INV_X1 U5398 ( .A(n4473), .ZN(n4350) );
  NAND2_X1 U5399 ( .A1(n5538), .A2(n4350), .ZN(n4503) );
  NAND2_X1 U5400 ( .A1(n6489), .A2(n4351), .ZN(n4352) );
  OAI22_X1 U5401 ( .A1(n5412), .A2(n4353), .B1(n4503), .B2(n4352), .ZN(U3455)
         );
  XNOR2_X1 U5402 ( .A(n4355), .B(n4354), .ZN(n4464) );
  INV_X1 U5403 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6804) );
  NOR2_X1 U5404 ( .A1(n6254), .A2(n6804), .ZN(n4459) );
  XNOR2_X1 U5405 ( .A(n5034), .B(n4054), .ZN(n4523) );
  NOR2_X1 U5406 ( .A1(n6255), .A2(n4523), .ZN(n4356) );
  AOI211_X1 U5407 ( .C1(n6222), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4459), 
        .B(n4356), .ZN(n4358) );
  OAI211_X1 U5408 ( .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n4366), .A(n6227), 
        .B(n5382), .ZN(n4357) );
  OAI211_X1 U5409 ( .C1(n4464), .C2(n6262), .A(n4358), .B(n4357), .ZN(U3017)
         );
  XNOR2_X1 U5410 ( .A(n4359), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4440)
         );
  NAND2_X1 U5411 ( .A1(n4360), .A2(n5384), .ZN(n4362) );
  AND2_X1 U5412 ( .A1(n4362), .A2(n4361), .ZN(n5543) );
  INV_X1 U5413 ( .A(REIP_REG_0__SCAN_IN), .ZN(n5546) );
  NOR2_X1 U5414 ( .A1(n6254), .A2(n5546), .ZN(n4437) );
  INV_X1 U5415 ( .A(n4363), .ZN(n4364) );
  AOI211_X1 U5416 ( .C1(n6273), .C2(n5543), .A(n4437), .B(n4364), .ZN(n4369)
         );
  INV_X1 U5417 ( .A(n4365), .ZN(n4367) );
  OAI21_X1 U5418 ( .B1(n4367), .B2(n4366), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4368) );
  OAI211_X1 U5419 ( .C1(n4440), .C2(n6262), .A(n4369), .B(n4368), .ZN(U3018)
         );
  INV_X1 U5420 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4376) );
  NAND2_X1 U5421 ( .A1(n6448), .A2(n4370), .ZN(n4371) );
  NAND2_X1 U5422 ( .A1(n4371), .A2(n6159), .ZN(n4373) );
  INV_X1 U5423 ( .A(n6504), .ZN(n4372) );
  NAND2_X1 U5424 ( .A1(n6116), .A2(n4931), .ZN(n6102) );
  NAND2_X1 U5425 ( .A1(n6596), .A2(n4513), .ZN(n6106) );
  AOI22_X1 U5426 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4375) );
  OAI21_X1 U5427 ( .B1(n4376), .B2(n6102), .A(n4375), .ZN(U2893) );
  INV_X1 U5428 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U5429 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4377) );
  OAI21_X1 U5430 ( .B1(n4378), .B2(n6102), .A(n4377), .ZN(U2899) );
  AOI22_X1 U5431 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4379) );
  OAI21_X1 U5432 ( .B1(n4398), .B2(n6102), .A(n4379), .ZN(U2906) );
  INV_X1 U5433 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U5434 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4380) );
  OAI21_X1 U5435 ( .B1(n4409), .B2(n6102), .A(n4380), .ZN(U2905) );
  INV_X1 U5436 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U5437 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4381) );
  OAI21_X1 U5438 ( .B1(n4382), .B2(n6102), .A(n4381), .ZN(U2904) );
  INV_X1 U5439 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4401) );
  AOI22_X1 U5440 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4383) );
  OAI21_X1 U5441 ( .B1(n4401), .B2(n6102), .A(n4383), .ZN(U2903) );
  AOI22_X1 U5442 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4384) );
  OAI21_X1 U5443 ( .B1(n4318), .B2(n6102), .A(n4384), .ZN(U2901) );
  INV_X1 U5444 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U5445 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4385) );
  OAI21_X1 U5446 ( .B1(n4386), .B2(n6102), .A(n4385), .ZN(U2900) );
  AOI22_X1 U5447 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4387) );
  OAI21_X1 U5448 ( .B1(n4311), .B2(n6102), .A(n4387), .ZN(U2898) );
  INV_X1 U5449 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4389) );
  AOI22_X1 U5450 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4388) );
  OAI21_X1 U5451 ( .B1(n4389), .B2(n6102), .A(n4388), .ZN(U2897) );
  INV_X1 U5452 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U5453 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4390) );
  OAI21_X1 U5454 ( .B1(n4391), .B2(n6102), .A(n4390), .ZN(U2895) );
  INV_X1 U5455 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4393) );
  INV_X1 U5456 ( .A(DATAI_4_), .ZN(n4445) );
  OR2_X1 U5457 ( .A1(n4422), .A2(n4445), .ZN(n4400) );
  NAND2_X1 U5458 ( .A1(n6156), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4392) );
  OAI211_X1 U5459 ( .C1(n6159), .C2(n4393), .A(n4400), .B(n4392), .ZN(U2943)
         );
  INV_X1 U5460 ( .A(EAX_REG_9__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U5461 ( .A1(n6156), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4394) );
  OAI211_X1 U5462 ( .C1(n6159), .C2(n4396), .A(n4395), .B(n4394), .ZN(U2948)
         );
  NAND2_X1 U5463 ( .A1(n6157), .A2(DATAI_1_), .ZN(n4403) );
  NAND2_X1 U5464 ( .A1(n6156), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4397) );
  OAI211_X1 U5465 ( .C1(n6159), .C2(n4398), .A(n4403), .B(n4397), .ZN(U2925)
         );
  NAND2_X1 U5466 ( .A1(n6156), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4399) );
  OAI211_X1 U5467 ( .C1(n6159), .C2(n4401), .A(n4400), .B(n4399), .ZN(U2928)
         );
  INV_X1 U5468 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U5469 ( .A1(n6156), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4402) );
  OAI211_X1 U5470 ( .C1(n6159), .C2(n4404), .A(n4403), .B(n4402), .ZN(U2940)
         );
  NAND2_X1 U5471 ( .A1(n6156), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4405) );
  OAI211_X1 U5472 ( .C1(n6159), .C2(n4389), .A(n4406), .B(n4405), .ZN(U2934)
         );
  NAND2_X1 U5473 ( .A1(n6156), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4407) );
  OAI211_X1 U5474 ( .C1(n6159), .C2(n4409), .A(n4408), .B(n4407), .ZN(U2926)
         );
  INV_X1 U5475 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U5476 ( .A1(n6156), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4410) );
  OAI211_X1 U5477 ( .C1(n6159), .C2(n4412), .A(n4411), .B(n4410), .ZN(U2945)
         );
  OAI21_X1 U5478 ( .B1(n4413), .B2(n4415), .A(n4414), .ZN(n5044) );
  NAND2_X1 U5479 ( .A1(n4416), .A2(n6490), .ZN(n4424) );
  INV_X1 U5480 ( .A(n4468), .ZN(n4420) );
  NOR2_X1 U5481 ( .A1(n4417), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4418) );
  AND2_X1 U5482 ( .A1(n4418), .A2(n3886), .ZN(n4451) );
  NAND3_X1 U5483 ( .A1(n4420), .A2(n4451), .A3(n4419), .ZN(n4421) );
  NAND2_X1 U5484 ( .A1(n3165), .A2(n5325), .ZN(n4425) );
  INV_X1 U5485 ( .A(n4425), .ZN(n4426) );
  INV_X1 U5486 ( .A(DATAI_1_), .ZN(n6651) );
  OAI222_X1 U5487 ( .A1(n5044), .A2(n5931), .B1(n5255), .B2(n6651), .C1(n5586), 
        .C2(n4404), .ZN(U2890) );
  NOR2_X1 U5488 ( .A1(n4428), .A2(n4427), .ZN(n4429) );
  NOR2_X1 U5489 ( .A1(n4443), .A2(n4429), .ZN(n6191) );
  INV_X1 U5490 ( .A(n6191), .ZN(n5018) );
  OAI222_X1 U5491 ( .A1(n5018), .A2(n5931), .B1(n5255), .B2(n4430), .C1(n5586), 
        .C2(n4315), .ZN(U2889) );
  XNOR2_X1 U5492 ( .A(n4443), .B(n4442), .ZN(n6083) );
  INV_X1 U5493 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6129) );
  OAI222_X1 U5494 ( .A1(n6083), .A2(n5931), .B1(n5255), .B2(n4431), .C1(n5586), 
        .C2(n6129), .ZN(U2888) );
  OAI21_X1 U5495 ( .B1(n4434), .B2(n4433), .A(n4432), .ZN(n5551) );
  INV_X1 U5496 ( .A(n5551), .ZN(n4438) );
  INV_X1 U5497 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5541) );
  AOI21_X1 U5498 ( .B1(n5702), .B2(n4435), .A(n5541), .ZN(n4436) );
  AOI211_X1 U5499 ( .C1(n4438), .C2(n6181), .A(n4437), .B(n4436), .ZN(n4439)
         );
  OAI21_X1 U5500 ( .B1(n4440), .B2(n6165), .A(n4439), .ZN(U2986) );
  AOI21_X1 U5501 ( .B1(n4443), .B2(n4442), .A(n4441), .ZN(n4444) );
  OR2_X1 U5502 ( .A1(n4613), .A2(n4444), .ZN(n5540) );
  OAI222_X1 U5503 ( .A1(n5540), .A2(n5931), .B1(n5255), .B2(n4445), .C1(n5586), 
        .C2(n4393), .ZN(U2887) );
  INV_X1 U5504 ( .A(n4447), .ZN(n4450) );
  NAND4_X1 U5505 ( .A1(n4451), .A2(n4450), .A3(n4449), .A4(n4448), .ZN(n4452)
         );
  NAND2_X2 U5506 ( .A1(n4453), .A2(n4452), .ZN(n6081) );
  INV_X2 U5507 ( .A(n6085), .ZN(n6078) );
  AND2_X1 U5508 ( .A1(n5178), .A2(n4454), .ZN(n4455) );
  OR2_X1 U5509 ( .A1(n4455), .A2(n4676), .ZN(n6256) );
  OAI22_X1 U5510 ( .A1(n6077), .A2(n6256), .B1(n4456), .B2(n6081), .ZN(n4457)
         );
  INV_X1 U5511 ( .A(n4457), .ZN(n4458) );
  OAI21_X1 U5512 ( .B1(n5540), .B2(n6078), .A(n4458), .ZN(U2855) );
  INV_X1 U5513 ( .A(n5044), .ZN(n4462) );
  AOI21_X1 U5514 ( .B1(n6187), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4459), 
        .ZN(n4460) );
  OAI21_X1 U5515 ( .B1(n6197), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4460), 
        .ZN(n4461) );
  AOI21_X1 U5516 ( .B1(n4462), .B2(n6181), .A(n4461), .ZN(n4463) );
  OAI21_X1 U5517 ( .B1(n4464), .B2(n6165), .A(n4463), .ZN(U2985) );
  INV_X1 U5518 ( .A(n4513), .ZN(n6493) );
  NAND2_X1 U5519 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6001), .ZN(n4508) );
  INV_X1 U5520 ( .A(n4479), .ZN(n4507) );
  INV_X1 U5521 ( .A(n4467), .ZN(n4469) );
  NAND3_X1 U5522 ( .A1(n4470), .A2(n4469), .A3(n4468), .ZN(n4471) );
  NOR2_X1 U5523 ( .A1(n4472), .A2(n4471), .ZN(n4474) );
  NAND2_X1 U5524 ( .A1(n4474), .A2(n4473), .ZN(n5402) );
  NAND2_X1 U5525 ( .A1(n5191), .A2(n5402), .ZN(n4491) );
  INV_X1 U5526 ( .A(n4475), .ZN(n4476) );
  OR2_X1 U5527 ( .A1(n4477), .A2(n4476), .ZN(n4498) );
  MUX2_X1 U5528 ( .A(n4478), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5398), 
        .Z(n4480) );
  NOR2_X1 U5529 ( .A1(n4480), .A2(n4479), .ZN(n4489) );
  AOI21_X1 U5530 ( .B1(n5398), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4481), 
        .ZN(n4482) );
  NOR2_X1 U5531 ( .A1(n4483), .A2(n4482), .ZN(n6575) );
  AND2_X1 U5532 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4485) );
  INV_X1 U5533 ( .A(n4485), .ZN(n4484) );
  MUX2_X1 U5534 ( .A(n4485), .B(n4484), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4486) );
  NAND2_X1 U5535 ( .A1(n6448), .A2(n4486), .ZN(n4487) );
  OAI21_X1 U5536 ( .B1(n6575), .B2(n4495), .A(n4487), .ZN(n4488) );
  AOI21_X1 U5537 ( .B1(n4498), .B2(n4489), .A(n4488), .ZN(n4490) );
  NAND2_X1 U5538 ( .A1(n4491), .A2(n4490), .ZN(n6573) );
  INV_X1 U5539 ( .A(n6452), .ZN(n4501) );
  MUX2_X1 U5540 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6573), .S(n4501), 
        .Z(n6465) );
  NAND2_X1 U5541 ( .A1(n5016), .A2(n5402), .ZN(n4500) );
  XNOR2_X1 U5542 ( .A(n5398), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4497)
         );
  XNOR2_X1 U5543 ( .A(n3204), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4493)
         );
  NAND2_X1 U5544 ( .A1(n6448), .A2(n4493), .ZN(n4494) );
  OAI21_X1 U5545 ( .B1(n4497), .B2(n4495), .A(n4494), .ZN(n4496) );
  AOI21_X1 U5546 ( .B1(n4498), .B2(n4497), .A(n4496), .ZN(n4499) );
  NAND2_X1 U5547 ( .A1(n4500), .A2(n4499), .ZN(n5385) );
  MUX2_X1 U5548 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5385), .S(n4501), 
        .Z(n6461) );
  NAND3_X1 U5549 ( .A1(n6465), .A2(n6461), .A3(n6480), .ZN(n4506) );
  NAND2_X1 U5550 ( .A1(n6452), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4502) );
  NAND2_X1 U5551 ( .A1(n4503), .A2(n4502), .ZN(n4505) );
  NOR2_X1 U5552 ( .A1(n4353), .A2(n4508), .ZN(n4504) );
  AOI21_X1 U5553 ( .B1(n4505), .B2(n6480), .A(n4504), .ZN(n4510) );
  OAI211_X1 U5554 ( .C1(n4508), .C2(n4507), .A(n4506), .B(n4510), .ZN(n6472)
         );
  NAND2_X1 U5555 ( .A1(n4510), .A2(n3019), .ZN(n4511) );
  NAND2_X1 U5556 ( .A1(n6472), .A2(n4511), .ZN(n4514) );
  AOI21_X1 U5557 ( .B1(n4514), .B2(n6001), .A(n6569), .ZN(n4512) );
  OR2_X1 U5558 ( .A1(n5072), .A2(n4512), .ZN(n6285) );
  NAND2_X1 U5559 ( .A1(n4514), .A2(n4513), .ZN(n6485) );
  INV_X1 U5560 ( .A(n6485), .ZN(n4516) );
  INV_X1 U5561 ( .A(n6385), .ZN(n6329) );
  NAND2_X1 U5562 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6571), .ZN(n4627) );
  INV_X1 U5563 ( .A(n4627), .ZN(n5838) );
  OAI22_X1 U5564 ( .A1(n4841), .A2(n6388), .B1(n6329), .B2(n5838), .ZN(n4515)
         );
  OAI21_X1 U5565 ( .B1(n4516), .B2(n4515), .A(n6285), .ZN(n4517) );
  OAI21_X1 U5566 ( .B1(n6285), .B2(n6447), .A(n4517), .ZN(U3465) );
  INV_X1 U5567 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6136) );
  OAI222_X1 U5568 ( .A1(n5551), .A2(n5931), .B1(n5255), .B2(n4518), .C1(n5586), 
        .C2(n6136), .ZN(U2891) );
  INV_X1 U5569 ( .A(n6285), .ZN(n4626) );
  NAND2_X1 U5570 ( .A1(n3022), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6383) );
  XNOR2_X1 U5571 ( .A(n4721), .B(n6383), .ZN(n4520) );
  AOI22_X1 U5572 ( .A1(n4520), .A2(n6338), .B1(n4627), .B2(n5016), .ZN(n4522)
         );
  NAND2_X1 U5573 ( .A1(n4626), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4521) );
  OAI21_X1 U5574 ( .B1(n4626), .B2(n4522), .A(n4521), .ZN(U3463) );
  INV_X1 U5575 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6632) );
  OAI222_X1 U5576 ( .A1(n4523), .A2(n6077), .B1(n6081), .B2(n6632), .C1(n6078), 
        .C2(n5044), .ZN(U2858) );
  INV_X1 U5577 ( .A(n5543), .ZN(n4525) );
  OAI222_X1 U5578 ( .A1(n4525), .A2(n6077), .B1(n6081), .B2(n4524), .C1(n5551), 
        .C2(n6078), .ZN(U2859) );
  NAND2_X1 U5579 ( .A1(n4721), .A2(n3308), .ZN(n4623) );
  NAND2_X1 U5580 ( .A1(n3022), .A2(n4841), .ZN(n6287) );
  AND2_X1 U5581 ( .A1(n6192), .A2(DATAI_31_), .ZN(n6371) );
  INV_X1 U5582 ( .A(n6371), .ZN(n6446) );
  NAND2_X1 U5583 ( .A1(n6192), .A2(DATAI_23_), .ZN(n6327) );
  INV_X1 U5584 ( .A(n6327), .ZN(n6438) );
  NAND2_X1 U5585 ( .A1(n3022), .A2(n4869), .ZN(n5116) );
  NOR2_X2 U5586 ( .A1(n4623), .A2(n5116), .ZN(n4671) );
  NAND2_X1 U5587 ( .A1(DATAI_7_), .A2(n5072), .ZN(n6375) );
  NAND2_X1 U5588 ( .A1(n5191), .A2(n6385), .ZN(n4862) );
  INV_X1 U5589 ( .A(n4526), .ZN(n5403) );
  NAND2_X1 U5590 ( .A1(n5016), .A2(n5403), .ZN(n6295) );
  OR2_X1 U5591 ( .A1(n4862), .A2(n6295), .ZN(n4527) );
  NAND2_X1 U5592 ( .A1(n4527), .A2(n4567), .ZN(n4532) );
  AOI22_X1 U5593 ( .A1(n4532), .A2(n6382), .B1(n5067), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4568) );
  INV_X1 U5594 ( .A(n4528), .ZN(n6570) );
  NOR2_X1 U5595 ( .A1(n4566), .A2(n5585), .ZN(n6437) );
  INV_X1 U5596 ( .A(n6437), .ZN(n5219) );
  OAI22_X1 U5597 ( .A1(n6375), .A2(n4568), .B1(n4567), .B2(n5219), .ZN(n4530)
         );
  AOI21_X1 U5598 ( .B1(n6438), .B2(n4671), .A(n4530), .ZN(n4537) );
  INV_X1 U5599 ( .A(n5072), .ZN(n4799) );
  INV_X1 U5600 ( .A(n4623), .ZN(n4531) );
  AOI21_X1 U5601 ( .B1(n4531), .B2(n3022), .A(n5352), .ZN(n4534) );
  NAND2_X1 U5602 ( .A1(n6382), .A2(n6593), .ZN(n5845) );
  INV_X1 U5603 ( .A(n5845), .ZN(n6296) );
  INV_X1 U5604 ( .A(n4532), .ZN(n4533) );
  OAI21_X1 U5605 ( .B1(n4534), .B2(n6296), .A(n4533), .ZN(n4535) );
  OAI211_X1 U5606 ( .C1(n5067), .C2(n6338), .A(n6337), .B(n4535), .ZN(n4570)
         );
  NAND2_X1 U5607 ( .A1(n4570), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4536)
         );
  OAI211_X1 U5608 ( .C1(n5063), .C2(n6446), .A(n4537), .B(n4536), .ZN(U3147)
         );
  NAND2_X1 U5609 ( .A1(n6181), .A2(DATAI_25_), .ZN(n6403) );
  AND2_X1 U5610 ( .A1(n6192), .A2(DATAI_17_), .ZN(n6399) );
  NAND2_X1 U5611 ( .A1(DATAI_1_), .A2(n5072), .ZN(n6347) );
  NOR2_X1 U5612 ( .A1(n4566), .A2(n4538), .ZN(n6398) );
  INV_X1 U5613 ( .A(n6398), .ZN(n5207) );
  OAI22_X1 U5614 ( .A1(n6347), .A2(n4568), .B1(n4567), .B2(n5207), .ZN(n4539)
         );
  AOI21_X1 U5615 ( .B1(n6399), .B2(n4671), .A(n4539), .ZN(n4541) );
  NAND2_X1 U5616 ( .A1(n4570), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4540)
         );
  OAI211_X1 U5617 ( .C1(n5063), .C2(n6403), .A(n4541), .B(n4540), .ZN(U3141)
         );
  AND2_X1 U5618 ( .A1(n6192), .A2(DATAI_30_), .ZN(n6429) );
  INV_X1 U5619 ( .A(n6429), .ZN(n5876) );
  AND2_X1 U5620 ( .A1(n6192), .A2(DATAI_22_), .ZN(n6364) );
  NAND2_X1 U5621 ( .A1(DATAI_6_), .A2(n5072), .ZN(n6367) );
  NOR2_X1 U5622 ( .A1(n4566), .A2(n4542), .ZN(n6428) );
  INV_X1 U5623 ( .A(n6428), .ZN(n5199) );
  OAI22_X1 U5624 ( .A1(n6367), .A2(n4568), .B1(n4567), .B2(n5199), .ZN(n4543)
         );
  AOI21_X1 U5625 ( .B1(n6364), .B2(n4671), .A(n4543), .ZN(n4545) );
  NAND2_X1 U5626 ( .A1(n4570), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4544)
         );
  OAI211_X1 U5627 ( .C1(n5063), .C2(n5876), .A(n4545), .B(n4544), .ZN(U3146)
         );
  NAND2_X1 U5628 ( .A1(n6192), .A2(DATAI_26_), .ZN(n6409) );
  AND2_X1 U5629 ( .A1(n6192), .A2(DATAI_18_), .ZN(n6405) );
  NAND2_X1 U5630 ( .A1(DATAI_2_), .A2(n5072), .ZN(n6351) );
  NOR2_X1 U5631 ( .A1(n4566), .A2(n3154), .ZN(n6404) );
  INV_X1 U5632 ( .A(n6404), .ZN(n5223) );
  OAI22_X1 U5633 ( .A1(n6351), .A2(n4568), .B1(n4567), .B2(n5223), .ZN(n4546)
         );
  AOI21_X1 U5634 ( .B1(n6405), .B2(n4671), .A(n4546), .ZN(n4548) );
  NAND2_X1 U5635 ( .A1(n4570), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4547)
         );
  OAI211_X1 U5636 ( .C1(n5063), .C2(n6409), .A(n4548), .B(n4547), .ZN(U3142)
         );
  AND2_X1 U5637 ( .A1(n6192), .A2(DATAI_27_), .ZN(n6411) );
  INV_X1 U5638 ( .A(n6411), .ZN(n5864) );
  NAND2_X1 U5639 ( .A1(n6181), .A2(DATAI_19_), .ZN(n6415) );
  INV_X1 U5640 ( .A(n6415), .ZN(n6352) );
  NAND2_X1 U5641 ( .A1(DATAI_3_), .A2(n5072), .ZN(n6355) );
  NOR2_X1 U5642 ( .A1(n4566), .A2(n4549), .ZN(n6410) );
  INV_X1 U5643 ( .A(n6410), .ZN(n5215) );
  OAI22_X1 U5644 ( .A1(n6355), .A2(n4568), .B1(n4567), .B2(n5215), .ZN(n4550)
         );
  AOI21_X1 U5645 ( .B1(n6352), .B2(n4671), .A(n4550), .ZN(n4552) );
  NAND2_X1 U5646 ( .A1(n4570), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4551)
         );
  OAI211_X1 U5647 ( .C1(n5063), .C2(n5864), .A(n4552), .B(n4551), .ZN(U3143)
         );
  AND2_X1 U5648 ( .A1(n6192), .A2(DATAI_24_), .ZN(n6380) );
  INV_X1 U5649 ( .A(n6380), .ZN(n5854) );
  AND2_X1 U5650 ( .A1(n6192), .A2(DATAI_16_), .ZN(n6340) );
  NAND2_X1 U5651 ( .A1(DATAI_0_), .A2(n5072), .ZN(n6343) );
  NOR2_X1 U5652 ( .A1(n4566), .A2(n4553), .ZN(n6379) );
  INV_X1 U5653 ( .A(n6379), .ZN(n5203) );
  OAI22_X1 U5654 ( .A1(n6343), .A2(n4568), .B1(n4567), .B2(n5203), .ZN(n4554)
         );
  AOI21_X1 U5655 ( .B1(n6340), .B2(n4671), .A(n4554), .ZN(n4556) );
  NAND2_X1 U5656 ( .A1(n4570), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4555)
         );
  OAI211_X1 U5657 ( .C1(n5063), .C2(n5854), .A(n4556), .B(n4555), .ZN(U3140)
         );
  AOI21_X1 U5658 ( .B1(n4613), .B2(n4614), .A(n4557), .ZN(n4558) );
  OR2_X1 U5659 ( .A1(n4903), .A2(n4558), .ZN(n5054) );
  OR2_X1 U5660 ( .A1(n4678), .A2(n4559), .ZN(n4560) );
  NAND2_X1 U5661 ( .A1(n6051), .A2(n4560), .ZN(n5046) );
  OAI22_X1 U5662 ( .A1(n5046), .A2(n6077), .B1(n5048), .B2(n6081), .ZN(n4561)
         );
  INV_X1 U5663 ( .A(n4561), .ZN(n4562) );
  OAI21_X1 U5664 ( .B1(n5054), .B2(n6078), .A(n4562), .ZN(U2853) );
  AND2_X1 U5665 ( .A1(n6192), .A2(DATAI_29_), .ZN(n6423) );
  INV_X1 U5666 ( .A(n6423), .ZN(n5872) );
  NAND2_X1 U5667 ( .A1(n6192), .A2(DATAI_21_), .ZN(n6427) );
  INV_X1 U5668 ( .A(n6427), .ZN(n6360) );
  NAND2_X1 U5669 ( .A1(DATAI_5_), .A2(n5072), .ZN(n6363) );
  NOR2_X1 U5670 ( .A1(n4566), .A2(n3012), .ZN(n6422) );
  INV_X1 U5671 ( .A(n6422), .ZN(n5211) );
  OAI22_X1 U5672 ( .A1(n6363), .A2(n4568), .B1(n4567), .B2(n5211), .ZN(n4563)
         );
  AOI21_X1 U5673 ( .B1(n6360), .B2(n4671), .A(n4563), .ZN(n4565) );
  NAND2_X1 U5674 ( .A1(n4570), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4564)
         );
  OAI211_X1 U5675 ( .C1(n5063), .C2(n5872), .A(n4565), .B(n4564), .ZN(U3145)
         );
  AND2_X1 U5676 ( .A1(n6192), .A2(DATAI_28_), .ZN(n6417) );
  INV_X1 U5677 ( .A(n6417), .ZN(n5868) );
  NAND2_X1 U5678 ( .A1(n6181), .A2(DATAI_20_), .ZN(n6421) );
  INV_X1 U5679 ( .A(n6421), .ZN(n6356) );
  NAND2_X1 U5680 ( .A1(DATAI_4_), .A2(n5072), .ZN(n6359) );
  NOR2_X1 U5681 ( .A1(n4566), .A2(n3018), .ZN(n6416) );
  INV_X1 U5682 ( .A(n6416), .ZN(n5229) );
  OAI22_X1 U5683 ( .A1(n6359), .A2(n4568), .B1(n4567), .B2(n5229), .ZN(n4569)
         );
  AOI21_X1 U5684 ( .B1(n6356), .B2(n4671), .A(n4569), .ZN(n4572) );
  NAND2_X1 U5685 ( .A1(n4570), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4571)
         );
  OAI211_X1 U5686 ( .C1(n5063), .C2(n5868), .A(n4572), .B(n4571), .ZN(U3144)
         );
  INV_X1 U5687 ( .A(DATAI_6_), .ZN(n6776) );
  OAI222_X1 U5688 ( .A1(n5054), .A2(n5931), .B1(n5255), .B2(n6776), .C1(n5586), 
        .C2(n4412), .ZN(U2885) );
  OR2_X1 U5689 ( .A1(n4574), .A2(n4573), .ZN(n4575) );
  AND2_X1 U5690 ( .A1(n5176), .A2(n4575), .ZN(n6272) );
  INV_X1 U5691 ( .A(n6081), .ZN(n5583) );
  AOI22_X1 U5692 ( .A1(n6084), .A2(n6272), .B1(n5583), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4576) );
  OAI21_X1 U5693 ( .B1(n5018), .B2(n6078), .A(n4576), .ZN(U2857) );
  NAND2_X1 U5694 ( .A1(n4721), .A2(n4577), .ZN(n6288) );
  OR2_X1 U5695 ( .A1(n6288), .A2(n3022), .ZN(n4692) );
  NAND3_X1 U5696 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6377), .A3(n6456), .ZN(n4687) );
  OR2_X1 U5697 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4687), .ZN(n4607)
         );
  NOR2_X1 U5698 ( .A1(n4582), .A2(n6475), .ZN(n6299) );
  OR2_X1 U5699 ( .A1(n4798), .A2(n6289), .ZN(n4637) );
  INV_X1 U5700 ( .A(n4637), .ZN(n4583) );
  OAI21_X1 U5701 ( .B1(n4583), .B2(n6475), .A(n5072), .ZN(n4632) );
  AOI211_X1 U5702 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4607), .A(n6299), .B(
        n4632), .ZN(n4581) );
  INV_X1 U5703 ( .A(n4721), .ZN(n4725) );
  INV_X1 U5704 ( .A(n5116), .ZN(n4800) );
  NAND3_X1 U5705 ( .A1(n4725), .A2(n4800), .A3(n4578), .ZN(n4753) );
  NOR3_X1 U5706 ( .A1(n6288), .A2(n3022), .A3(n6593), .ZN(n4579) );
  NOR2_X1 U5707 ( .A1(n4579), .A2(n6388), .ZN(n4686) );
  NAND2_X1 U5708 ( .A1(n5016), .A2(n4526), .ZN(n4843) );
  OR2_X1 U5709 ( .A1(n4843), .A2(n6294), .ZN(n4683) );
  OAI211_X1 U5710 ( .C1(n6296), .C2(n4753), .A(n4686), .B(n4683), .ZN(n4580)
         );
  NAND2_X1 U5711 ( .A1(n4581), .A2(n4580), .ZN(n4606) );
  NAND2_X1 U5712 ( .A1(n4606), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4587) );
  INV_X1 U5713 ( .A(n5191), .ZN(n4760) );
  NAND2_X1 U5714 ( .A1(n4760), .A2(n6382), .ZN(n6292) );
  INV_X1 U5715 ( .A(n6292), .ZN(n4584) );
  INV_X1 U5716 ( .A(n4843), .ZN(n4801) );
  AND2_X1 U5717 ( .A1(n4582), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6290) );
  AOI22_X1 U5718 ( .A1(n4584), .A2(n4801), .B1(n6290), .B2(n4583), .ZN(n4608)
         );
  OAI22_X1 U5719 ( .A1(n6359), .A2(n4608), .B1(n5229), .B2(n4607), .ZN(n4585)
         );
  AOI21_X1 U5720 ( .B1(n6417), .B2(n4610), .A(n4585), .ZN(n4586) );
  OAI211_X1 U5721 ( .C1(n4691), .C2(n6421), .A(n4587), .B(n4586), .ZN(U3056)
         );
  INV_X1 U5722 ( .A(n6364), .ZN(n6435) );
  NAND2_X1 U5723 ( .A1(n4606), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4590) );
  OAI22_X1 U5724 ( .A1(n6367), .A2(n4608), .B1(n5199), .B2(n4607), .ZN(n4588)
         );
  AOI21_X1 U5725 ( .B1(n6429), .B2(n4610), .A(n4588), .ZN(n4589) );
  OAI211_X1 U5726 ( .C1(n4691), .C2(n6435), .A(n4590), .B(n4589), .ZN(U3058)
         );
  NAND2_X1 U5727 ( .A1(n4606), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4593) );
  OAI22_X1 U5728 ( .A1(n6355), .A2(n4608), .B1(n5215), .B2(n4607), .ZN(n4591)
         );
  AOI21_X1 U5729 ( .B1(n6411), .B2(n4610), .A(n4591), .ZN(n4592) );
  OAI211_X1 U5730 ( .C1(n4691), .C2(n6415), .A(n4593), .B(n4592), .ZN(U3055)
         );
  INV_X1 U5731 ( .A(n6399), .ZN(n6308) );
  NAND2_X1 U5732 ( .A1(n4606), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4596) );
  INV_X1 U5733 ( .A(n6403), .ZN(n6344) );
  OAI22_X1 U5734 ( .A1(n6347), .A2(n4608), .B1(n5207), .B2(n4607), .ZN(n4594)
         );
  AOI21_X1 U5735 ( .B1(n6344), .B2(n4610), .A(n4594), .ZN(n4595) );
  OAI211_X1 U5736 ( .C1(n4691), .C2(n6308), .A(n4596), .B(n4595), .ZN(U3053)
         );
  NAND2_X1 U5737 ( .A1(n4606), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4599) );
  OAI22_X1 U5738 ( .A1(n6363), .A2(n4608), .B1(n5211), .B2(n4607), .ZN(n4597)
         );
  AOI21_X1 U5739 ( .B1(n6423), .B2(n4610), .A(n4597), .ZN(n4598) );
  OAI211_X1 U5740 ( .C1(n4691), .C2(n6427), .A(n4599), .B(n4598), .ZN(U3057)
         );
  INV_X1 U5741 ( .A(n6340), .ZN(n6397) );
  NAND2_X1 U5742 ( .A1(n4606), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4602) );
  OAI22_X1 U5743 ( .A1(n6343), .A2(n4608), .B1(n5203), .B2(n4607), .ZN(n4600)
         );
  AOI21_X1 U5744 ( .B1(n6380), .B2(n4610), .A(n4600), .ZN(n4601) );
  OAI211_X1 U5745 ( .C1(n4691), .C2(n6397), .A(n4602), .B(n4601), .ZN(U3052)
         );
  INV_X1 U5746 ( .A(n6405), .ZN(n6311) );
  NAND2_X1 U5747 ( .A1(n4606), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4605) );
  INV_X1 U5748 ( .A(n6409), .ZN(n6348) );
  OAI22_X1 U5749 ( .A1(n6351), .A2(n4608), .B1(n5223), .B2(n4607), .ZN(n4603)
         );
  AOI21_X1 U5750 ( .B1(n6348), .B2(n4610), .A(n4603), .ZN(n4604) );
  OAI211_X1 U5751 ( .C1(n4691), .C2(n6311), .A(n4605), .B(n4604), .ZN(U3054)
         );
  NAND2_X1 U5752 ( .A1(n4606), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4612) );
  OAI22_X1 U5753 ( .A1(n6375), .A2(n4608), .B1(n5219), .B2(n4607), .ZN(n4609)
         );
  AOI21_X1 U5754 ( .B1(n6371), .B2(n4610), .A(n4609), .ZN(n4611) );
  OAI211_X1 U5755 ( .C1(n4691), .C2(n6327), .A(n4612), .B(n4611), .ZN(U3059)
         );
  XOR2_X1 U5756 ( .A(n4614), .B(n4613), .Z(n6173) );
  INV_X1 U5757 ( .A(n6173), .ZN(n4680) );
  OAI222_X1 U5758 ( .A1(n5931), .A2(n4680), .B1(n5255), .B2(n4615), .C1(n5586), 
        .C2(n3533), .ZN(U2886) );
  OR2_X1 U5759 ( .A1(n4618), .A2(n4617), .ZN(n4619) );
  NAND2_X1 U5760 ( .A1(n4616), .A2(n4619), .ZN(n6253) );
  OAI22_X1 U5761 ( .A1(n5702), .A2(n3512), .B1(n6254), .B2(n6520), .ZN(n4621)
         );
  NOR2_X1 U5762 ( .A1(n5540), .A2(n5352), .ZN(n4620) );
  AOI211_X1 U5763 ( .C1(n5946), .C2(n5529), .A(n4621), .B(n4620), .ZN(n4622)
         );
  OAI21_X1 U5764 ( .B1(n6165), .B2(n6253), .A(n4622), .ZN(U2982) );
  NOR2_X1 U5765 ( .A1(n6288), .A2(n6383), .ZN(n6328) );
  NOR2_X1 U5766 ( .A1(n6328), .A2(n6381), .ZN(n4625) );
  INV_X1 U5767 ( .A(n4842), .ZN(n4624) );
  NAND2_X1 U5768 ( .A1(n4624), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4846) );
  AOI21_X1 U5769 ( .B1(n4625), .B2(n4846), .A(n6388), .ZN(n4722) );
  NOR2_X1 U5770 ( .A1(n4626), .A2(n4722), .ZN(n4629) );
  NAND2_X1 U5771 ( .A1(n5191), .A2(n4627), .ZN(n4628) );
  OAI211_X1 U5772 ( .C1(n4578), .C2(n5845), .A(n4629), .B(n4628), .ZN(n4630)
         );
  OAI21_X1 U5773 ( .B1(n6285), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n4630), 
        .ZN(n4631) );
  INV_X1 U5774 ( .A(n4631), .ZN(U3462) );
  NOR3_X1 U5775 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4767) );
  NAND2_X1 U5776 ( .A1(n6447), .A2(n4767), .ZN(n4638) );
  AOI211_X1 U5777 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4638), .A(n6290), .B(
        n4632), .ZN(n4636) );
  NAND3_X1 U5778 ( .A1(n4725), .A2(n4860), .A3(n4578), .ZN(n4769) );
  INV_X1 U5779 ( .A(n4769), .ZN(n4633) );
  OAI21_X1 U5780 ( .B1(n4633), .B2(n6388), .A(n5845), .ZN(n4765) );
  NAND2_X1 U5781 ( .A1(n4671), .A2(n5845), .ZN(n4634) );
  OAI211_X1 U5782 ( .C1(n5191), .C2(n5125), .A(n4765), .B(n4634), .ZN(n4635)
         );
  OR2_X1 U5783 ( .A1(n4769), .A2(n4869), .ZN(n4768) );
  INV_X1 U5784 ( .A(n6347), .ZN(n6400) );
  INV_X1 U5785 ( .A(n6299), .ZN(n5841) );
  OAI22_X1 U5786 ( .A1(n6292), .A2(n5125), .B1(n5841), .B2(n4637), .ZN(n4668)
         );
  INV_X1 U5787 ( .A(n4638), .ZN(n4667) );
  AOI22_X1 U5788 ( .A1(n6400), .A2(n4668), .B1(n6398), .B2(n4667), .ZN(n4639)
         );
  OAI21_X1 U5789 ( .B1(n6308), .B2(n4768), .A(n4639), .ZN(n4640) );
  AOI21_X1 U5790 ( .B1(n6344), .B2(n4671), .A(n4640), .ZN(n4641) );
  OAI21_X1 U5791 ( .B1(n4674), .B2(n4642), .A(n4641), .ZN(U3021) );
  INV_X1 U5792 ( .A(n6363), .ZN(n6424) );
  AOI22_X1 U5793 ( .A1(n6424), .A2(n4668), .B1(n6422), .B2(n4667), .ZN(n4643)
         );
  OAI21_X1 U5794 ( .B1(n6427), .B2(n4768), .A(n4643), .ZN(n4644) );
  AOI21_X1 U5795 ( .B1(n6423), .B2(n4671), .A(n4644), .ZN(n4645) );
  OAI21_X1 U5796 ( .B1(n4674), .B2(n4646), .A(n4645), .ZN(U3025) );
  INV_X1 U5797 ( .A(n6367), .ZN(n6431) );
  AOI22_X1 U5798 ( .A1(n6431), .A2(n4668), .B1(n6428), .B2(n4667), .ZN(n4647)
         );
  OAI21_X1 U5799 ( .B1(n6435), .B2(n4768), .A(n4647), .ZN(n4648) );
  AOI21_X1 U5800 ( .B1(n6429), .B2(n4671), .A(n4648), .ZN(n4649) );
  OAI21_X1 U5801 ( .B1(n4674), .B2(n4650), .A(n4649), .ZN(U3026) );
  INV_X1 U5802 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4654) );
  INV_X1 U5803 ( .A(n6355), .ZN(n6412) );
  AOI22_X1 U5804 ( .A1(n6412), .A2(n4668), .B1(n6410), .B2(n4667), .ZN(n4651)
         );
  OAI21_X1 U5805 ( .B1(n6415), .B2(n4768), .A(n4651), .ZN(n4652) );
  AOI21_X1 U5806 ( .B1(n6411), .B2(n4671), .A(n4652), .ZN(n4653) );
  OAI21_X1 U5807 ( .B1(n4674), .B2(n4654), .A(n4653), .ZN(U3023) );
  INV_X1 U5808 ( .A(n6359), .ZN(n6418) );
  AOI22_X1 U5809 ( .A1(n6418), .A2(n4668), .B1(n6416), .B2(n4667), .ZN(n4655)
         );
  OAI21_X1 U5810 ( .B1(n6421), .B2(n4768), .A(n4655), .ZN(n4656) );
  AOI21_X1 U5811 ( .B1(n6417), .B2(n4671), .A(n4656), .ZN(n4657) );
  OAI21_X1 U5812 ( .B1(n4674), .B2(n4658), .A(n4657), .ZN(U3024) );
  INV_X1 U5813 ( .A(n6351), .ZN(n6406) );
  AOI22_X1 U5814 ( .A1(n6406), .A2(n4668), .B1(n6404), .B2(n4667), .ZN(n4659)
         );
  OAI21_X1 U5815 ( .B1(n6311), .B2(n4768), .A(n4659), .ZN(n4660) );
  AOI21_X1 U5816 ( .B1(n6348), .B2(n4671), .A(n4660), .ZN(n4661) );
  OAI21_X1 U5817 ( .B1(n4674), .B2(n4662), .A(n4661), .ZN(U3022) );
  INV_X1 U5818 ( .A(n6343), .ZN(n6394) );
  AOI22_X1 U5819 ( .A1(n6394), .A2(n4668), .B1(n6379), .B2(n4667), .ZN(n4663)
         );
  OAI21_X1 U5820 ( .B1(n6397), .B2(n4768), .A(n4663), .ZN(n4664) );
  AOI21_X1 U5821 ( .B1(n6380), .B2(n4671), .A(n4664), .ZN(n4665) );
  OAI21_X1 U5822 ( .B1(n4674), .B2(n4666), .A(n4665), .ZN(U3020) );
  INV_X1 U5823 ( .A(n6375), .ZN(n6441) );
  AOI22_X1 U5824 ( .A1(n6441), .A2(n4668), .B1(n6437), .B2(n4667), .ZN(n4669)
         );
  OAI21_X1 U5825 ( .B1(n6327), .B2(n4768), .A(n4669), .ZN(n4670) );
  AOI21_X1 U5826 ( .B1(n6371), .B2(n4671), .A(n4670), .ZN(n4672) );
  OAI21_X1 U5827 ( .B1(n4674), .B2(n4673), .A(n4672), .ZN(U3027) );
  NOR2_X1 U5828 ( .A1(n4676), .A2(n4675), .ZN(n4677) );
  OR2_X1 U5829 ( .A1(n4678), .A2(n4677), .ZN(n6239) );
  INV_X1 U5830 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4679) );
  OAI222_X1 U5831 ( .A1(n6239), .A2(n6077), .B1(n6078), .B2(n4680), .C1(n6081), 
        .C2(n4679), .ZN(U2854) );
  NAND2_X1 U5832 ( .A1(n4903), .A2(n4902), .ZN(n4956) );
  OR2_X1 U5833 ( .A1(n4903), .A2(n4902), .ZN(n4681) );
  NAND2_X1 U5834 ( .A1(n4956), .A2(n4681), .ZN(n6164) );
  INV_X1 U5835 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6124) );
  OAI222_X1 U5836 ( .A1(n6164), .A2(n5931), .B1(n5255), .B2(n4682), .C1(n5586), 
        .C2(n6124), .ZN(U2884) );
  OR2_X1 U5837 ( .A1(n4683), .A2(n6329), .ZN(n4684) );
  OR2_X1 U5838 ( .A1(n6447), .A2(n4687), .ZN(n4715) );
  NAND2_X1 U5839 ( .A1(n4684), .A2(n4715), .ZN(n4689) );
  INV_X1 U5840 ( .A(n4687), .ZN(n4685) );
  AOI22_X1 U5841 ( .A1(n4686), .A2(n4689), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4685), .ZN(n4720) );
  INV_X1 U5842 ( .A(n4686), .ZN(n4690) );
  AOI21_X1 U5843 ( .B1(n6388), .B2(n4687), .A(n6387), .ZN(n4688) );
  OAI21_X1 U5844 ( .B1(n4690), .B2(n4689), .A(n4688), .ZN(n4714) );
  NAND2_X1 U5845 ( .A1(n4714), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4695) );
  OAI22_X1 U5846 ( .A1(n5229), .A2(n4715), .B1(n6421), .B2(n6293), .ZN(n4693)
         );
  AOI21_X1 U5847 ( .B1(n6417), .B2(n4717), .A(n4693), .ZN(n4694) );
  OAI211_X1 U5848 ( .C1(n4720), .C2(n6359), .A(n4695), .B(n4694), .ZN(U3064)
         );
  NAND2_X1 U5849 ( .A1(n4714), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4698) );
  OAI22_X1 U5850 ( .A1(n5223), .A2(n4715), .B1(n6311), .B2(n6293), .ZN(n4696)
         );
  AOI21_X1 U5851 ( .B1(n6348), .B2(n4717), .A(n4696), .ZN(n4697) );
  OAI211_X1 U5852 ( .C1(n4720), .C2(n6351), .A(n4698), .B(n4697), .ZN(U3062)
         );
  NAND2_X1 U5853 ( .A1(n4714), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4701) );
  OAI22_X1 U5854 ( .A1(n5207), .A2(n4715), .B1(n6308), .B2(n6293), .ZN(n4699)
         );
  AOI21_X1 U5855 ( .B1(n6344), .B2(n4717), .A(n4699), .ZN(n4700) );
  OAI211_X1 U5856 ( .C1(n4720), .C2(n6347), .A(n4701), .B(n4700), .ZN(U3061)
         );
  NAND2_X1 U5857 ( .A1(n4714), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4704) );
  OAI22_X1 U5858 ( .A1(n5215), .A2(n4715), .B1(n6415), .B2(n6293), .ZN(n4702)
         );
  AOI21_X1 U5859 ( .B1(n6411), .B2(n4717), .A(n4702), .ZN(n4703) );
  OAI211_X1 U5860 ( .C1(n4720), .C2(n6355), .A(n4704), .B(n4703), .ZN(U3063)
         );
  NAND2_X1 U5861 ( .A1(n4714), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4707) );
  OAI22_X1 U5862 ( .A1(n5219), .A2(n4715), .B1(n6327), .B2(n6293), .ZN(n4705)
         );
  AOI21_X1 U5863 ( .B1(n6371), .B2(n4717), .A(n4705), .ZN(n4706) );
  OAI211_X1 U5864 ( .C1(n4720), .C2(n6375), .A(n4707), .B(n4706), .ZN(U3067)
         );
  NAND2_X1 U5865 ( .A1(n4714), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4710) );
  OAI22_X1 U5866 ( .A1(n5199), .A2(n4715), .B1(n6435), .B2(n6293), .ZN(n4708)
         );
  AOI21_X1 U5867 ( .B1(n6429), .B2(n4717), .A(n4708), .ZN(n4709) );
  OAI211_X1 U5868 ( .C1(n4720), .C2(n6367), .A(n4710), .B(n4709), .ZN(U3066)
         );
  NAND2_X1 U5869 ( .A1(n4714), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4713) );
  OAI22_X1 U5870 ( .A1(n5211), .A2(n4715), .B1(n6427), .B2(n6293), .ZN(n4711)
         );
  AOI21_X1 U5871 ( .B1(n6423), .B2(n4717), .A(n4711), .ZN(n4712) );
  OAI211_X1 U5872 ( .C1(n4720), .C2(n6363), .A(n4713), .B(n4712), .ZN(U3065)
         );
  NAND2_X1 U5873 ( .A1(n4714), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4719) );
  OAI22_X1 U5874 ( .A1(n5203), .A2(n4715), .B1(n6397), .B2(n6293), .ZN(n4716)
         );
  AOI21_X1 U5875 ( .B1(n6380), .B2(n4717), .A(n4716), .ZN(n4718) );
  OAI211_X1 U5876 ( .C1(n4720), .C2(n6343), .A(n4719), .B(n4718), .ZN(U3060)
         );
  OR2_X1 U5877 ( .A1(n4721), .A2(n6383), .ZN(n4723) );
  AOI21_X1 U5878 ( .B1(n6382), .B2(n4723), .A(n4722), .ZN(n4728) );
  NOR2_X1 U5879 ( .A1(n5016), .A2(n4526), .ZN(n5192) );
  NOR2_X1 U5880 ( .A1(n6378), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4726)
         );
  AOI21_X1 U5881 ( .B1(n5844), .B2(n6385), .A(n4726), .ZN(n4729) );
  NAND3_X1 U5882 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6377), .A3(n6460), .ZN(n5843) );
  OAI22_X1 U5883 ( .A1(n4728), .A2(n4729), .B1(n5843), .B2(n6475), .ZN(n4724)
         );
  INV_X1 U5884 ( .A(n6287), .ZN(n5189) );
  INV_X1 U5885 ( .A(n4726), .ZN(n4754) );
  OAI22_X1 U5886 ( .A1(n5229), .A2(n4754), .B1(n6421), .B2(n4753), .ZN(n4727)
         );
  AOI21_X1 U5887 ( .B1(n6417), .B2(n5882), .A(n4727), .ZN(n4734) );
  INV_X1 U5888 ( .A(n5843), .ZN(n4732) );
  INV_X1 U5889 ( .A(n4728), .ZN(n4730) );
  NAND2_X1 U5890 ( .A1(n4730), .A2(n4729), .ZN(n4731) );
  OAI211_X1 U5891 ( .C1(n6338), .C2(n4732), .A(n4731), .B(n6337), .ZN(n4756)
         );
  NAND2_X1 U5892 ( .A1(n4756), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4733) );
  OAI211_X1 U5893 ( .C1(n4759), .C2(n6359), .A(n4734), .B(n4733), .ZN(U3048)
         );
  OAI22_X1 U5894 ( .A1(n5211), .A2(n4754), .B1(n6427), .B2(n4753), .ZN(n4735)
         );
  AOI21_X1 U5895 ( .B1(n6423), .B2(n5882), .A(n4735), .ZN(n4737) );
  NAND2_X1 U5896 ( .A1(n4756), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4736) );
  OAI211_X1 U5897 ( .C1(n4759), .C2(n6363), .A(n4737), .B(n4736), .ZN(U3049)
         );
  OAI22_X1 U5898 ( .A1(n5199), .A2(n4754), .B1(n6435), .B2(n4753), .ZN(n4738)
         );
  AOI21_X1 U5899 ( .B1(n6429), .B2(n5882), .A(n4738), .ZN(n4740) );
  NAND2_X1 U5900 ( .A1(n4756), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4739) );
  OAI211_X1 U5901 ( .C1(n4759), .C2(n6367), .A(n4740), .B(n4739), .ZN(U3050)
         );
  OAI22_X1 U5902 ( .A1(n5219), .A2(n4754), .B1(n6327), .B2(n4753), .ZN(n4741)
         );
  AOI21_X1 U5903 ( .B1(n6371), .B2(n5882), .A(n4741), .ZN(n4743) );
  NAND2_X1 U5904 ( .A1(n4756), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4742) );
  OAI211_X1 U5905 ( .C1(n4759), .C2(n6375), .A(n4743), .B(n4742), .ZN(U3051)
         );
  OAI22_X1 U5906 ( .A1(n5207), .A2(n4754), .B1(n6308), .B2(n4753), .ZN(n4744)
         );
  AOI21_X1 U5907 ( .B1(n6344), .B2(n5882), .A(n4744), .ZN(n4746) );
  NAND2_X1 U5908 ( .A1(n4756), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4745) );
  OAI211_X1 U5909 ( .C1(n4759), .C2(n6347), .A(n4746), .B(n4745), .ZN(U3045)
         );
  OAI22_X1 U5910 ( .A1(n5203), .A2(n4754), .B1(n6397), .B2(n4753), .ZN(n4747)
         );
  AOI21_X1 U5911 ( .B1(n6380), .B2(n5882), .A(n4747), .ZN(n4749) );
  NAND2_X1 U5912 ( .A1(n4756), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4748) );
  OAI211_X1 U5913 ( .C1(n4759), .C2(n6343), .A(n4749), .B(n4748), .ZN(U3044)
         );
  OAI22_X1 U5914 ( .A1(n5215), .A2(n4754), .B1(n6415), .B2(n4753), .ZN(n4750)
         );
  AOI21_X1 U5915 ( .B1(n6411), .B2(n5882), .A(n4750), .ZN(n4752) );
  NAND2_X1 U5916 ( .A1(n4756), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4751) );
  OAI211_X1 U5917 ( .C1(n4759), .C2(n6355), .A(n4752), .B(n4751), .ZN(U3047)
         );
  OAI22_X1 U5918 ( .A1(n5223), .A2(n4754), .B1(n6311), .B2(n4753), .ZN(n4755)
         );
  AOI21_X1 U5919 ( .B1(n6348), .B2(n5882), .A(n4755), .ZN(n4758) );
  NAND2_X1 U5920 ( .A1(n4756), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4757) );
  OAI211_X1 U5921 ( .C1(n4759), .C2(n6351), .A(n4758), .B(n4757), .ZN(U3046)
         );
  INV_X1 U5922 ( .A(n5125), .ZN(n5115) );
  NAND3_X1 U5923 ( .A1(n4760), .A2(n5115), .A3(n6385), .ZN(n4762) );
  INV_X1 U5924 ( .A(n4767), .ZN(n4761) );
  OR2_X1 U5925 ( .A1(n6447), .A2(n4761), .ZN(n4792) );
  NAND2_X1 U5926 ( .A1(n4762), .A2(n4792), .ZN(n4763) );
  AOI22_X1 U5927 ( .A1(n4765), .A2(n4763), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4767), .ZN(n4797) );
  INV_X1 U5928 ( .A(n4763), .ZN(n4764) );
  AOI21_X1 U5929 ( .B1(n4765), .B2(n4764), .A(n6387), .ZN(n4766) );
  OAI21_X1 U5930 ( .B1(n6338), .B2(n4767), .A(n4766), .ZN(n4791) );
  NAND2_X1 U5931 ( .A1(n4791), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4772) );
  OAI22_X1 U5932 ( .A1(n5223), .A2(n4792), .B1(n6311), .B2(n5884), .ZN(n4770)
         );
  AOI21_X1 U5933 ( .B1(n6348), .B2(n4794), .A(n4770), .ZN(n4771) );
  OAI211_X1 U5934 ( .C1(n4797), .C2(n6351), .A(n4772), .B(n4771), .ZN(U3030)
         );
  NAND2_X1 U5935 ( .A1(n4791), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4775) );
  OAI22_X1 U5936 ( .A1(n5229), .A2(n4792), .B1(n6421), .B2(n5884), .ZN(n4773)
         );
  AOI21_X1 U5937 ( .B1(n6417), .B2(n4794), .A(n4773), .ZN(n4774) );
  OAI211_X1 U5938 ( .C1(n4797), .C2(n6359), .A(n4775), .B(n4774), .ZN(U3032)
         );
  NAND2_X1 U5939 ( .A1(n4791), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4778) );
  OAI22_X1 U5940 ( .A1(n5215), .A2(n4792), .B1(n6415), .B2(n5884), .ZN(n4776)
         );
  AOI21_X1 U5941 ( .B1(n6411), .B2(n4794), .A(n4776), .ZN(n4777) );
  OAI211_X1 U5942 ( .C1(n4797), .C2(n6355), .A(n4778), .B(n4777), .ZN(U3031)
         );
  NAND2_X1 U5943 ( .A1(n4791), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4781) );
  OAI22_X1 U5944 ( .A1(n5199), .A2(n4792), .B1(n6435), .B2(n5884), .ZN(n4779)
         );
  AOI21_X1 U5945 ( .B1(n6429), .B2(n4794), .A(n4779), .ZN(n4780) );
  OAI211_X1 U5946 ( .C1(n4797), .C2(n6367), .A(n4781), .B(n4780), .ZN(U3034)
         );
  NAND2_X1 U5947 ( .A1(n4791), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4784) );
  OAI22_X1 U5948 ( .A1(n5203), .A2(n4792), .B1(n6397), .B2(n5884), .ZN(n4782)
         );
  AOI21_X1 U5949 ( .B1(n6380), .B2(n4794), .A(n4782), .ZN(n4783) );
  OAI211_X1 U5950 ( .C1(n4797), .C2(n6343), .A(n4784), .B(n4783), .ZN(U3028)
         );
  NAND2_X1 U5951 ( .A1(n4791), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4787) );
  OAI22_X1 U5952 ( .A1(n5211), .A2(n4792), .B1(n6427), .B2(n5884), .ZN(n4785)
         );
  AOI21_X1 U5953 ( .B1(n6423), .B2(n4794), .A(n4785), .ZN(n4786) );
  OAI211_X1 U5954 ( .C1(n4797), .C2(n6363), .A(n4787), .B(n4786), .ZN(U3033)
         );
  NAND2_X1 U5955 ( .A1(n4791), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4790) );
  OAI22_X1 U5956 ( .A1(n5207), .A2(n4792), .B1(n6308), .B2(n5884), .ZN(n4788)
         );
  AOI21_X1 U5957 ( .B1(n6344), .B2(n4794), .A(n4788), .ZN(n4789) );
  OAI211_X1 U5958 ( .C1(n4797), .C2(n6347), .A(n4790), .B(n4789), .ZN(U3029)
         );
  NAND2_X1 U5959 ( .A1(n4791), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4796) );
  OAI22_X1 U5960 ( .A1(n5219), .A2(n4792), .B1(n6327), .B2(n5884), .ZN(n4793)
         );
  AOI21_X1 U5961 ( .B1(n6371), .B2(n4794), .A(n4793), .ZN(n4795) );
  OAI211_X1 U5962 ( .C1(n4797), .C2(n6375), .A(n4796), .B(n4795), .ZN(U3035)
         );
  NAND3_X1 U5963 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6456), .ZN(n4849) );
  NOR2_X1 U5964 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4849), .ZN(n4834)
         );
  INV_X1 U5965 ( .A(n6289), .ZN(n5840) );
  NAND2_X1 U5966 ( .A1(n5840), .A2(n4798), .ZN(n5124) );
  AOI21_X1 U5967 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5124), .A(n4799), .ZN(
        n5119) );
  OAI211_X1 U5968 ( .C1(n6571), .C2(n4834), .A(n5119), .B(n5841), .ZN(n4804)
         );
  NAND3_X1 U5969 ( .A1(n6434), .A2(n6338), .A3(n4805), .ZN(n4802) );
  AOI22_X1 U5970 ( .A1(n4802), .A2(n5845), .B1(n4801), .B2(n6294), .ZN(n4803)
         );
  INV_X1 U5971 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4809) );
  NAND2_X1 U5972 ( .A1(n5191), .A2(n6382), .ZN(n5126) );
  INV_X1 U5973 ( .A(n6290), .ZN(n5118) );
  OAI22_X1 U5974 ( .A1(n5126), .A2(n4843), .B1(n5118), .B2(n5124), .ZN(n4835)
         );
  AOI22_X1 U5975 ( .A1(n6412), .A2(n4835), .B1(n6410), .B2(n4834), .ZN(n4806)
         );
  OAI21_X1 U5976 ( .B1(n5864), .B2(n6434), .A(n4806), .ZN(n4807) );
  AOI21_X1 U5977 ( .B1(n4899), .B2(n6352), .A(n4807), .ZN(n4808) );
  OAI21_X1 U5978 ( .B1(n4840), .B2(n4809), .A(n4808), .ZN(U3119) );
  INV_X1 U5979 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4813) );
  AOI22_X1 U5980 ( .A1(n6431), .A2(n4835), .B1(n6428), .B2(n4834), .ZN(n4810)
         );
  OAI21_X1 U5981 ( .B1(n5876), .B2(n6434), .A(n4810), .ZN(n4811) );
  AOI21_X1 U5982 ( .B1(n4899), .B2(n6364), .A(n4811), .ZN(n4812) );
  OAI21_X1 U5983 ( .B1(n4840), .B2(n4813), .A(n4812), .ZN(U3122) );
  INV_X1 U5984 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4817) );
  AOI22_X1 U5985 ( .A1(n6424), .A2(n4835), .B1(n6422), .B2(n4834), .ZN(n4814)
         );
  OAI21_X1 U5986 ( .B1(n5872), .B2(n6434), .A(n4814), .ZN(n4815) );
  AOI21_X1 U5987 ( .B1(n4899), .B2(n6360), .A(n4815), .ZN(n4816) );
  OAI21_X1 U5988 ( .B1(n4840), .B2(n4817), .A(n4816), .ZN(U3121) );
  INV_X1 U5989 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4821) );
  AOI22_X1 U5990 ( .A1(n6441), .A2(n4835), .B1(n6437), .B2(n4834), .ZN(n4818)
         );
  OAI21_X1 U5991 ( .B1(n6446), .B2(n6434), .A(n4818), .ZN(n4819) );
  AOI21_X1 U5992 ( .B1(n4899), .B2(n6438), .A(n4819), .ZN(n4820) );
  OAI21_X1 U5993 ( .B1(n4840), .B2(n4821), .A(n4820), .ZN(U3123) );
  INV_X1 U5994 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4825) );
  AOI22_X1 U5995 ( .A1(n6394), .A2(n4835), .B1(n6379), .B2(n4834), .ZN(n4822)
         );
  OAI21_X1 U5996 ( .B1(n5854), .B2(n6434), .A(n4822), .ZN(n4823) );
  AOI21_X1 U5997 ( .B1(n6340), .B2(n4899), .A(n4823), .ZN(n4824) );
  OAI21_X1 U5998 ( .B1(n4840), .B2(n4825), .A(n4824), .ZN(U3116) );
  INV_X1 U5999 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U6000 ( .A1(n6400), .A2(n4835), .B1(n6398), .B2(n4834), .ZN(n4826)
         );
  OAI21_X1 U6001 ( .B1(n6403), .B2(n6434), .A(n4826), .ZN(n4827) );
  AOI21_X1 U6002 ( .B1(n4899), .B2(n6399), .A(n4827), .ZN(n4828) );
  OAI21_X1 U6003 ( .B1(n4840), .B2(n4829), .A(n4828), .ZN(U3117) );
  INV_X1 U6004 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U6005 ( .A1(n6406), .A2(n4835), .B1(n6404), .B2(n4834), .ZN(n4830)
         );
  OAI21_X1 U6006 ( .B1(n6409), .B2(n6434), .A(n4830), .ZN(n4831) );
  AOI21_X1 U6007 ( .B1(n4899), .B2(n6405), .A(n4831), .ZN(n4832) );
  OAI21_X1 U6008 ( .B1(n4840), .B2(n4833), .A(n4832), .ZN(U3118) );
  INV_X1 U6009 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4839) );
  AOI22_X1 U6010 ( .A1(n6418), .A2(n4835), .B1(n6416), .B2(n4834), .ZN(n4836)
         );
  OAI21_X1 U6011 ( .B1(n5868), .B2(n6434), .A(n4836), .ZN(n4837) );
  AOI21_X1 U6012 ( .B1(n4899), .B2(n6356), .A(n4837), .ZN(n4838) );
  OAI21_X1 U6013 ( .B1(n4840), .B2(n4839), .A(n4838), .ZN(U3120) );
  OR2_X1 U6014 ( .A1(n4862), .A2(n4843), .ZN(n4845) );
  NOR2_X1 U6015 ( .A1(n6447), .A2(n4849), .ZN(n4898) );
  INV_X1 U6016 ( .A(n4898), .ZN(n4844) );
  AND2_X1 U6017 ( .A1(n4845), .A2(n4844), .ZN(n4851) );
  INV_X1 U6018 ( .A(n4851), .ZN(n4848) );
  NAND2_X1 U6019 ( .A1(n6382), .A2(n4846), .ZN(n4850) );
  AOI21_X1 U6020 ( .B1(n6388), .B2(n4849), .A(n6387), .ZN(n4847) );
  OAI21_X1 U6021 ( .B1(n4848), .B2(n4850), .A(n4847), .ZN(n4897) );
  OAI22_X1 U6022 ( .A1(n4851), .A2(n4850), .B1(n6475), .B2(n4849), .ZN(n4896)
         );
  AOI22_X1 U6023 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4897), .B1(n6424), 
        .B2(n4896), .ZN(n4853) );
  AOI22_X1 U6024 ( .A1(n4899), .A2(n6423), .B1(n6422), .B2(n4898), .ZN(n4852)
         );
  OAI211_X1 U6025 ( .C1(n5103), .C2(n6427), .A(n4853), .B(n4852), .ZN(U3129)
         );
  AOI22_X1 U6026 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4897), .B1(n6400), 
        .B2(n4896), .ZN(n4855) );
  AOI22_X1 U6027 ( .A1(n4899), .A2(n6344), .B1(n6398), .B2(n4898), .ZN(n4854)
         );
  OAI211_X1 U6028 ( .C1(n5103), .C2(n6308), .A(n4855), .B(n4854), .ZN(U3125)
         );
  AOI22_X1 U6029 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4897), .B1(n6394), 
        .B2(n4896), .ZN(n4857) );
  AOI22_X1 U6030 ( .A1(n6380), .A2(n4899), .B1(n6379), .B2(n4898), .ZN(n4856)
         );
  OAI211_X1 U6031 ( .C1(n5103), .C2(n6397), .A(n4857), .B(n4856), .ZN(U3124)
         );
  AOI22_X1 U6032 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4897), .B1(n6418), 
        .B2(n4896), .ZN(n4859) );
  AOI22_X1 U6033 ( .A1(n4899), .A2(n6417), .B1(n6416), .B2(n4898), .ZN(n4858)
         );
  OAI211_X1 U6034 ( .C1(n5103), .C2(n6421), .A(n4859), .B(n4858), .ZN(U3128)
         );
  NAND2_X1 U6035 ( .A1(n6381), .A2(n4860), .ZN(n4870) );
  INV_X1 U6036 ( .A(n4870), .ZN(n4861) );
  OAI21_X1 U6037 ( .B1(n4870), .B2(n6593), .A(n6382), .ZN(n4867) );
  OR2_X1 U6038 ( .A1(n4862), .A2(n5125), .ZN(n4864) );
  NAND3_X1 U6039 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6460), .A3(n6456), .ZN(n5117) );
  NOR2_X1 U6040 ( .A1(n6447), .A2(n5117), .ZN(n4889) );
  INV_X1 U6041 ( .A(n4889), .ZN(n4863) );
  AND2_X1 U6042 ( .A1(n4864), .A2(n4863), .ZN(n4868) );
  INV_X1 U6043 ( .A(n4868), .ZN(n4866) );
  AOI21_X1 U6044 ( .B1(n6388), .B2(n5117), .A(n6387), .ZN(n4865) );
  OAI21_X1 U6045 ( .B1(n4867), .B2(n4866), .A(n4865), .ZN(n4888) );
  OAI22_X1 U6046 ( .A1(n4868), .A2(n4867), .B1(n6475), .B2(n5117), .ZN(n4887)
         );
  AOI22_X1 U6047 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4888), .B1(n6431), 
        .B2(n4887), .ZN(n4872) );
  NOR2_X2 U6048 ( .A1(n4870), .A2(n4869), .ZN(n5160) );
  AOI22_X1 U6049 ( .A1(n5160), .A2(n6429), .B1(n6428), .B2(n4889), .ZN(n4871)
         );
  OAI211_X1 U6050 ( .C1(n6435), .C2(n5188), .A(n4872), .B(n4871), .ZN(U3098)
         );
  AOI22_X1 U6051 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4897), .B1(n6406), 
        .B2(n4896), .ZN(n4874) );
  AOI22_X1 U6052 ( .A1(n4899), .A2(n6348), .B1(n6404), .B2(n4898), .ZN(n4873)
         );
  OAI211_X1 U6053 ( .C1(n5103), .C2(n6311), .A(n4874), .B(n4873), .ZN(U3126)
         );
  AOI22_X1 U6054 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4888), .B1(n6418), 
        .B2(n4887), .ZN(n4876) );
  AOI22_X1 U6055 ( .A1(n5160), .A2(n6417), .B1(n6416), .B2(n4889), .ZN(n4875)
         );
  OAI211_X1 U6056 ( .C1(n6421), .C2(n5188), .A(n4876), .B(n4875), .ZN(U3096)
         );
  AOI22_X1 U6057 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4888), .B1(n6412), 
        .B2(n4887), .ZN(n4878) );
  AOI22_X1 U6058 ( .A1(n5160), .A2(n6411), .B1(n6410), .B2(n4889), .ZN(n4877)
         );
  OAI211_X1 U6059 ( .C1(n6415), .C2(n5188), .A(n4878), .B(n4877), .ZN(U3095)
         );
  AOI22_X1 U6060 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4888), .B1(n6406), 
        .B2(n4887), .ZN(n4880) );
  AOI22_X1 U6061 ( .A1(n5160), .A2(n6348), .B1(n6404), .B2(n4889), .ZN(n4879)
         );
  OAI211_X1 U6062 ( .C1(n6311), .C2(n5188), .A(n4880), .B(n4879), .ZN(U3094)
         );
  AOI22_X1 U6063 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4888), .B1(n6400), 
        .B2(n4887), .ZN(n4882) );
  AOI22_X1 U6064 ( .A1(n5160), .A2(n6344), .B1(n6398), .B2(n4889), .ZN(n4881)
         );
  OAI211_X1 U6065 ( .C1(n6308), .C2(n5188), .A(n4882), .B(n4881), .ZN(U3093)
         );
  AOI22_X1 U6066 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4888), .B1(n6394), 
        .B2(n4887), .ZN(n4884) );
  AOI22_X1 U6067 ( .A1(n5160), .A2(n6380), .B1(n6379), .B2(n4889), .ZN(n4883)
         );
  OAI211_X1 U6068 ( .C1(n6397), .C2(n5188), .A(n4884), .B(n4883), .ZN(U3092)
         );
  AOI22_X1 U6069 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4888), .B1(n6424), 
        .B2(n4887), .ZN(n4886) );
  AOI22_X1 U6070 ( .A1(n5160), .A2(n6423), .B1(n6422), .B2(n4889), .ZN(n4885)
         );
  OAI211_X1 U6071 ( .C1(n6427), .C2(n5188), .A(n4886), .B(n4885), .ZN(U3097)
         );
  AOI22_X1 U6072 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4888), .B1(n6441), 
        .B2(n4887), .ZN(n4891) );
  AOI22_X1 U6073 ( .A1(n5160), .A2(n6371), .B1(n6437), .B2(n4889), .ZN(n4890)
         );
  OAI211_X1 U6074 ( .C1(n6327), .C2(n5188), .A(n4891), .B(n4890), .ZN(U3099)
         );
  AOI22_X1 U6075 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4897), .B1(n6441), 
        .B2(n4896), .ZN(n4893) );
  AOI22_X1 U6076 ( .A1(n4899), .A2(n6371), .B1(n6437), .B2(n4898), .ZN(n4892)
         );
  OAI211_X1 U6077 ( .C1(n5103), .C2(n6327), .A(n4893), .B(n4892), .ZN(U3131)
         );
  AOI22_X1 U6078 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4897), .B1(n6412), 
        .B2(n4896), .ZN(n4895) );
  AOI22_X1 U6079 ( .A1(n4899), .A2(n6411), .B1(n6410), .B2(n4898), .ZN(n4894)
         );
  OAI211_X1 U6080 ( .C1(n5103), .C2(n6415), .A(n4895), .B(n4894), .ZN(U3127)
         );
  AOI22_X1 U6081 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4897), .B1(n6431), 
        .B2(n4896), .ZN(n4901) );
  AOI22_X1 U6082 ( .A1(n4899), .A2(n6429), .B1(n6428), .B2(n4898), .ZN(n4900)
         );
  OAI211_X1 U6083 ( .C1(n5103), .C2(n6435), .A(n4901), .B(n4900), .ZN(U3130)
         );
  AND2_X1 U6084 ( .A1(n4903), .A2(n4902), .ZN(n4905) );
  AND2_X1 U6085 ( .A1(n4905), .A2(n4904), .ZN(n5106) );
  OAI21_X1 U6086 ( .B1(n5106), .B2(n4906), .A(n4916), .ZN(n6612) );
  OR2_X1 U6087 ( .A1(n5110), .A2(n4907), .ZN(n4908) );
  AND2_X1 U6088 ( .A1(n4919), .A2(n4908), .ZN(n6621) );
  AOI22_X1 U6089 ( .A1(n6621), .A2(n6084), .B1(EBX_REG_14__SCAN_IN), .B2(n5583), .ZN(n4909) );
  OAI21_X1 U6090 ( .B1(n6612), .B2(n6078), .A(n4909), .ZN(U2845) );
  AOI22_X1 U6091 ( .A1(n5173), .A2(DATAI_14_), .B1(n6098), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n4910) );
  OAI21_X1 U6092 ( .B1(n6612), .B2(n5931), .A(n4910), .ZN(U2877) );
  AOI21_X1 U6093 ( .B1(n4955), .B2(n4956), .A(n5105), .ZN(n4999) );
  INV_X1 U6094 ( .A(n4999), .ZN(n4944) );
  AND2_X1 U6095 ( .A1(n6053), .A2(n4911), .ZN(n4912) );
  NOR2_X1 U6096 ( .A1(n4979), .A2(n4912), .ZN(n4993) );
  NOR2_X1 U6097 ( .A1(n6081), .A2(n4940), .ZN(n4913) );
  AOI21_X1 U6098 ( .B1(n4993), .B2(n6084), .A(n4913), .ZN(n4914) );
  OAI21_X1 U6099 ( .B1(n4944), .B2(n6078), .A(n4914), .ZN(U2851) );
  AOI22_X1 U6100 ( .A1(n5173), .A2(DATAI_8_), .B1(n6098), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4915) );
  OAI21_X1 U6101 ( .B1(n4944), .B2(n5931), .A(n4915), .ZN(U2883) );
  OAI21_X1 U6102 ( .B1(n3555), .B2(n3554), .A(n5020), .ZN(n5723) );
  INV_X1 U6103 ( .A(n5024), .ZN(n4918) );
  AOI21_X1 U6104 ( .B1(n4920), .B2(n4919), .A(n4918), .ZN(n5961) );
  AOI22_X1 U6105 ( .A1(n5961), .A2(n6084), .B1(n5583), .B2(EBX_REG_15__SCAN_IN), .ZN(n4921) );
  OAI21_X1 U6106 ( .B1(n5723), .B2(n6078), .A(n4921), .ZN(U2844) );
  AOI22_X1 U6107 ( .A1(n5173), .A2(DATAI_15_), .B1(n6098), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n4922) );
  OAI21_X1 U6108 ( .B1(n5723), .B2(n5931), .A(n4922), .ZN(U2876) );
  NAND2_X1 U6109 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .ZN(
        n4923) );
  NAND2_X1 U6110 ( .A1(n4966), .A2(REIP_REG_2__SCAN_IN), .ZN(n5007) );
  OAI21_X1 U6111 ( .B1(n4923), .B2(n5007), .A(n5899), .ZN(n5530) );
  INV_X1 U6112 ( .A(n5530), .ZN(n4924) );
  AOI21_X1 U6113 ( .B1(n5899), .B2(n4925), .A(n4924), .ZN(n4926) );
  INV_X1 U6114 ( .A(n4926), .ZN(n6043) );
  INV_X1 U6115 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6527) );
  OR2_X1 U6116 ( .A1(n6608), .A2(n4927), .ZN(n5531) );
  NOR2_X1 U6117 ( .A1(n5531), .A2(n6520), .ZN(n6072) );
  INV_X1 U6118 ( .A(n6072), .ZN(n4928) );
  NOR2_X1 U6119 ( .A1(n4928), .A2(n6522), .ZN(n6049) );
  NAND2_X1 U6120 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6049), .ZN(n6064) );
  INV_X1 U6121 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6529) );
  OAI21_X1 U6122 ( .B1(n6527), .B2(n6064), .A(n6529), .ZN(n4942) );
  NOR2_X1 U6123 ( .A1(n4929), .A2(EBX_REG_31__SCAN_IN), .ZN(n4930) );
  NAND2_X1 U6124 ( .A1(n4931), .A2(n4930), .ZN(n4932) );
  NAND2_X1 U6125 ( .A1(n4933), .A2(n4932), .ZN(n4934) );
  NAND2_X1 U6126 ( .A1(n4993), .A2(n6058), .ZN(n4939) );
  NOR2_X1 U6127 ( .A1(n4935), .A2(n6480), .ZN(n4936) );
  INV_X1 U6128 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4995) );
  INV_X1 U6129 ( .A(n4966), .ZN(n5035) );
  NOR2_X1 U6130 ( .A1(n5035), .A2(n5997), .ZN(n6610) );
  INV_X1 U6131 ( .A(n6610), .ZN(n6066) );
  OAI21_X1 U6132 ( .B1(n6619), .B2(n4995), .A(n6066), .ZN(n4937) );
  AOI21_X1 U6133 ( .B1(n6614), .B2(n4998), .A(n4937), .ZN(n4938) );
  OAI211_X1 U6134 ( .C1(n4940), .C2(n6035), .A(n4939), .B(n4938), .ZN(n4941)
         );
  AOI21_X1 U6135 ( .B1(n6043), .B2(n4942), .A(n4941), .ZN(n4943) );
  OAI21_X1 U6136 ( .B1(n6060), .B2(n4944), .A(n4943), .ZN(U2819) );
  INV_X1 U6137 ( .A(n6192), .ZN(n5352) );
  NAND2_X1 U6138 ( .A1(n4134), .A2(n4946), .ZN(n4949) );
  INV_X1 U6139 ( .A(n4947), .ZN(n4948) );
  AOI21_X1 U6140 ( .B1(n4950), .B2(n4949), .A(n4948), .ZN(n6234) );
  NAND2_X1 U6141 ( .A1(n6234), .A2(n6193), .ZN(n4954) );
  AND2_X1 U6142 ( .A1(n6279), .A2(REIP_REG_6__SCAN_IN), .ZN(n6228) );
  INV_X1 U6143 ( .A(n4951), .ZN(n5051) );
  NOR2_X1 U6144 ( .A1(n6197), .A2(n5051), .ZN(n4952) );
  AOI211_X1 U6145 ( .C1(n6187), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6228), 
        .B(n4952), .ZN(n4953) );
  OAI211_X1 U6146 ( .C1(n5352), .C2(n5054), .A(n4954), .B(n4953), .ZN(U2980)
         );
  AND2_X1 U6147 ( .A1(n5105), .A2(n4957), .ZN(n5235) );
  NAND2_X1 U6148 ( .A1(n5105), .A2(n4958), .ZN(n5166) );
  OAI21_X1 U6149 ( .B1(n5235), .B2(n4959), .A(n5166), .ZN(n5351) );
  INV_X1 U6150 ( .A(n5347), .ZN(n4971) );
  INV_X1 U6151 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6634) );
  INV_X1 U6152 ( .A(n4960), .ZN(n4963) );
  INV_X1 U6153 ( .A(n4961), .ZN(n4962) );
  OAI21_X1 U6154 ( .B1(n4963), .B2(n4962), .A(n5170), .ZN(n5114) );
  INV_X1 U6155 ( .A(n5114), .ZN(n6199) );
  AOI22_X1 U6156 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6054), .B1(n6058), 
        .B2(n6199), .ZN(n4964) );
  OAI211_X1 U6157 ( .C1(n6035), .C2(n6634), .A(n4964), .B(n6066), .ZN(n4970)
         );
  INV_X1 U6158 ( .A(n4965), .ZN(n6024) );
  OAI21_X1 U6159 ( .B1(n6608), .B2(n6024), .A(n4966), .ZN(n6028) );
  INV_X1 U6160 ( .A(n6028), .ZN(n5520) );
  AOI21_X1 U6161 ( .B1(n6025), .B2(n4967), .A(REIP_REG_11__SCAN_IN), .ZN(n4968) );
  NOR2_X1 U6162 ( .A1(n5520), .A2(n4968), .ZN(n4969) );
  AOI211_X1 U6163 ( .C1(n6614), .C2(n4971), .A(n4970), .B(n4969), .ZN(n4972)
         );
  OAI21_X1 U6164 ( .B1(n5351), .B2(n6060), .A(n4972), .ZN(U2816) );
  AOI22_X1 U6165 ( .A1(n5173), .A2(DATAI_11_), .B1(n6098), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4973) );
  OAI21_X1 U6166 ( .B1(n5351), .B2(n5931), .A(n4973), .ZN(U2880) );
  NAND2_X1 U6167 ( .A1(n4975), .A2(n4974), .ZN(n4976) );
  NAND2_X1 U6168 ( .A1(n5236), .A2(n4976), .ZN(n5275) );
  INV_X1 U6169 ( .A(DATAI_9_), .ZN(n6787) );
  OAI222_X1 U6170 ( .A1(n5275), .A2(n5931), .B1(n5255), .B2(n6787), .C1(n5586), 
        .C2(n4396), .ZN(U2882) );
  INV_X1 U6171 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4981) );
  NOR2_X1 U6172 ( .A1(n4979), .A2(n4978), .ZN(n4980) );
  OR2_X1 U6173 ( .A1(n4977), .A2(n4980), .ZN(n6205) );
  OAI222_X1 U6174 ( .A1(n5275), .A2(n6078), .B1(n6081), .B2(n4981), .C1(n6077), 
        .C2(n6205), .ZN(U2850) );
  OAI21_X1 U6175 ( .B1(n4984), .B2(n4983), .A(n5269), .ZN(n5002) );
  NOR2_X1 U6176 ( .A1(n6254), .A2(n6529), .ZN(n4997) );
  NAND3_X1 U6177 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n6280), .ZN(n6241) );
  NAND2_X1 U6178 ( .A1(n6250), .A2(n6241), .ZN(n6232) );
  NAND2_X1 U6179 ( .A1(n6270), .A2(n6232), .ZN(n6264) );
  INV_X1 U6180 ( .A(n6264), .ZN(n4985) );
  OAI21_X1 U6181 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6214), .ZN(n4991) );
  AOI22_X1 U6182 ( .A1(n6224), .A2(n4989), .B1(n4988), .B2(n4987), .ZN(n6221)
         );
  OAI22_X1 U6183 ( .A1(n5285), .A2(n4991), .B1(n6221), .B2(n4990), .ZN(n4992)
         );
  AOI211_X1 U6184 ( .C1(n6273), .C2(n4993), .A(n4997), .B(n4992), .ZN(n4994)
         );
  OAI21_X1 U6185 ( .B1(n5002), .B2(n6262), .A(n4994), .ZN(U3010) );
  NOR2_X1 U6186 ( .A1(n5702), .A2(n4995), .ZN(n4996) );
  AOI211_X1 U6187 ( .C1(n5946), .C2(n4998), .A(n4997), .B(n4996), .ZN(n5001)
         );
  NAND2_X1 U6188 ( .A1(n4999), .A2(n6181), .ZN(n5000) );
  OAI211_X1 U6189 ( .C1(n5002), .C2(n6165), .A(n5001), .B(n5000), .ZN(U2978)
         );
  NAND2_X1 U6190 ( .A1(n5006), .A2(n5003), .ZN(n5004) );
  AND2_X1 U6191 ( .A1(n5006), .A2(n5005), .ZN(n5549) );
  AND2_X1 U6192 ( .A1(n6025), .A2(REIP_REG_1__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U6193 ( .A1(n6025), .A2(n6804), .ZN(n5039) );
  INV_X1 U6194 ( .A(n5007), .ZN(n5008) );
  NAND2_X1 U6195 ( .A1(n5039), .A2(n5008), .ZN(n5183) );
  OAI21_X1 U6196 ( .B1(n5009), .B2(REIP_REG_2__SCAN_IN), .A(n5183), .ZN(n5014)
         );
  INV_X1 U6197 ( .A(n6196), .ZN(n5010) );
  AOI22_X1 U6198 ( .A1(n6054), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6614), 
        .B2(n5010), .ZN(n5013) );
  NAND2_X1 U6199 ( .A1(n6058), .A2(n6272), .ZN(n5012) );
  NAND2_X1 U6200 ( .A1(n6611), .A2(EBX_REG_2__SCAN_IN), .ZN(n5011) );
  NAND4_X1 U6201 ( .A1(n5014), .A2(n5013), .A3(n5012), .A4(n5011), .ZN(n5015)
         );
  AOI21_X1 U6202 ( .B1(n5549), .B2(n5016), .A(n5015), .ZN(n5017) );
  OAI21_X1 U6203 ( .B1(n5018), .B2(n6065), .A(n5017), .ZN(U2825) );
  AND2_X1 U6204 ( .A1(n5020), .A2(n5019), .ZN(n5022) );
  OR2_X1 U6205 ( .A1(n5022), .A2(n5244), .ZN(n6094) );
  INV_X1 U6206 ( .A(n5246), .ZN(n5023) );
  AOI21_X1 U6207 ( .B1(n5025), .B2(n5024), .A(n5023), .ZN(n5834) );
  AOI22_X1 U6208 ( .A1(n5834), .A2(n6084), .B1(EBX_REG_16__SCAN_IN), .B2(n5583), .ZN(n5026) );
  OAI21_X1 U6209 ( .B1(n6094), .B2(n6078), .A(n5026), .ZN(U2843) );
  NAND2_X1 U6210 ( .A1(n5711), .A2(n6614), .ZN(n5027) );
  OAI211_X1 U6211 ( .C1(n6619), .C2(n6801), .A(n5027), .B(n6066), .ZN(n5032)
         );
  INV_X1 U6212 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U6213 ( .A1(n5899), .A2(n5028), .ZN(n6622) );
  INV_X1 U6214 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5251) );
  NOR2_X1 U6215 ( .A1(n6540), .A2(n5251), .ZN(n5260) );
  AOI21_X1 U6216 ( .B1(n6540), .B2(n5251), .A(n5260), .ZN(n5029) );
  AOI22_X1 U6217 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6611), .B1(n5259), .B2(n5029), .ZN(n5030) );
  OAI21_X1 U6218 ( .B1(n6540), .B2(n6622), .A(n5030), .ZN(n5031) );
  AOI211_X1 U6219 ( .C1(n5834), .C2(n6058), .A(n5032), .B(n5031), .ZN(n5033)
         );
  OAI21_X1 U6220 ( .B1(n6094), .B2(n6060), .A(n5033), .ZN(U2811) );
  NAND2_X1 U6221 ( .A1(n6058), .A2(n5034), .ZN(n5037) );
  AOI22_X1 U6222 ( .A1(n6054), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5035), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5036) );
  OAI211_X1 U6223 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6075), .A(n5037), 
        .B(n5036), .ZN(n5041) );
  NAND2_X1 U6224 ( .A1(n6611), .A2(EBX_REG_1__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U6225 ( .A1(n5039), .A2(n5038), .ZN(n5040) );
  NOR2_X1 U6226 ( .A1(n5041), .A2(n5040), .ZN(n5043) );
  NAND2_X1 U6227 ( .A1(n5403), .A2(n5549), .ZN(n5042) );
  OAI211_X1 U6228 ( .C1(n5044), .C2(n6065), .A(n5043), .B(n5042), .ZN(U2826)
         );
  OAI21_X1 U6229 ( .B1(n5547), .B2(n5045), .A(n5530), .ZN(n6071) );
  INV_X1 U6230 ( .A(n5046), .ZN(n6229) );
  INV_X1 U6231 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6525) );
  AOI22_X1 U6232 ( .A1(n6058), .A2(n6229), .B1(n6049), .B2(n6525), .ZN(n5047)
         );
  OAI21_X1 U6233 ( .B1(n5048), .B2(n6035), .A(n5047), .ZN(n5049) );
  AOI211_X1 U6234 ( .C1(n6054), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6610), 
        .B(n5049), .ZN(n5050) );
  OAI21_X1 U6235 ( .B1(n6075), .B2(n5051), .A(n5050), .ZN(n5052) );
  AOI21_X1 U6236 ( .B1(n6071), .B2(REIP_REG_6__SCAN_IN), .A(n5052), .ZN(n5053)
         );
  OAI21_X1 U6237 ( .B1(n6060), .B2(n5054), .A(n5053), .ZN(U2821) );
  NOR2_X1 U6238 ( .A1(n6608), .A2(REIP_REG_9__SCAN_IN), .ZN(n6044) );
  AOI22_X1 U6239 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6611), .B1(n5055), .B2(n6044), 
        .ZN(n5056) );
  INV_X1 U6240 ( .A(n5056), .ZN(n5061) );
  INV_X1 U6241 ( .A(n5271), .ZN(n5057) );
  AOI21_X1 U6242 ( .B1(n6614), .B2(n5057), .A(n6610), .ZN(n5059) );
  NAND2_X1 U6243 ( .A1(n6054), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5058)
         );
  OAI211_X1 U6244 ( .C1(n6205), .C2(n6624), .A(n5059), .B(n5058), .ZN(n5060)
         );
  AOI211_X1 U6245 ( .C1(n6043), .C2(REIP_REG_9__SCAN_IN), .A(n5061), .B(n5060), 
        .ZN(n5062) );
  OAI21_X1 U6246 ( .B1(n6060), .B2(n5275), .A(n5062), .ZN(U2818) );
  INV_X1 U6247 ( .A(n5126), .ZN(n5066) );
  INV_X1 U6248 ( .A(n6295), .ZN(n5065) );
  NOR3_X1 U6249 ( .A1(n5118), .A2(n6377), .A3(n5840), .ZN(n5064) );
  AOI21_X1 U6250 ( .B1(n5066), .B2(n5065), .A(n5064), .ZN(n5097) );
  INV_X1 U6251 ( .A(n5067), .ZN(n5068) );
  NOR2_X1 U6252 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5068), .ZN(n5075)
         );
  INV_X1 U6253 ( .A(n5075), .ZN(n5096) );
  OAI22_X1 U6254 ( .A1(n6375), .A2(n5097), .B1(n5219), .B2(n5096), .ZN(n5069)
         );
  AOI21_X1 U6255 ( .B1(n6438), .B2(n5099), .A(n5069), .ZN(n5077) );
  INV_X1 U6256 ( .A(n5103), .ZN(n5070) );
  OAI21_X1 U6257 ( .B1(n5070), .B2(n5099), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5071) );
  NAND3_X1 U6258 ( .A1(n6295), .A2(n6382), .A3(n5071), .ZN(n5074) );
  OAI21_X1 U6259 ( .B1(n6289), .B2(n6475), .A(n5072), .ZN(n6298) );
  NOR3_X1 U6260 ( .A1(n6298), .A2(n6377), .A3(n6299), .ZN(n5073) );
  NAND2_X1 U6261 ( .A1(n5100), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5076)
         );
  OAI211_X1 U6262 ( .C1(n6446), .C2(n5103), .A(n5077), .B(n5076), .ZN(U3139)
         );
  OAI22_X1 U6263 ( .A1(n6367), .A2(n5097), .B1(n5199), .B2(n5096), .ZN(n5078)
         );
  AOI21_X1 U6264 ( .B1(n6364), .B2(n5099), .A(n5078), .ZN(n5080) );
  NAND2_X1 U6265 ( .A1(n5100), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5079)
         );
  OAI211_X1 U6266 ( .C1(n5876), .C2(n5103), .A(n5080), .B(n5079), .ZN(U3138)
         );
  OAI22_X1 U6267 ( .A1(n6355), .A2(n5097), .B1(n5215), .B2(n5096), .ZN(n5081)
         );
  AOI21_X1 U6268 ( .B1(n6352), .B2(n5099), .A(n5081), .ZN(n5083) );
  NAND2_X1 U6269 ( .A1(n5100), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5082)
         );
  OAI211_X1 U6270 ( .C1(n5864), .C2(n5103), .A(n5083), .B(n5082), .ZN(U3135)
         );
  OAI22_X1 U6271 ( .A1(n6351), .A2(n5097), .B1(n5223), .B2(n5096), .ZN(n5084)
         );
  AOI21_X1 U6272 ( .B1(n6405), .B2(n5099), .A(n5084), .ZN(n5086) );
  NAND2_X1 U6273 ( .A1(n5100), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5085)
         );
  OAI211_X1 U6274 ( .C1(n6409), .C2(n5103), .A(n5086), .B(n5085), .ZN(U3134)
         );
  OAI22_X1 U6275 ( .A1(n6347), .A2(n5097), .B1(n5207), .B2(n5096), .ZN(n5087)
         );
  AOI21_X1 U6276 ( .B1(n6399), .B2(n5099), .A(n5087), .ZN(n5089) );
  NAND2_X1 U6277 ( .A1(n5100), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5088)
         );
  OAI211_X1 U6278 ( .C1(n6403), .C2(n5103), .A(n5089), .B(n5088), .ZN(U3133)
         );
  OAI22_X1 U6279 ( .A1(n6343), .A2(n5097), .B1(n5203), .B2(n5096), .ZN(n5090)
         );
  AOI21_X1 U6280 ( .B1(n6340), .B2(n5099), .A(n5090), .ZN(n5092) );
  NAND2_X1 U6281 ( .A1(n5100), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5091)
         );
  OAI211_X1 U6282 ( .C1(n5854), .C2(n5103), .A(n5092), .B(n5091), .ZN(U3132)
         );
  OAI22_X1 U6283 ( .A1(n6363), .A2(n5097), .B1(n5211), .B2(n5096), .ZN(n5093)
         );
  AOI21_X1 U6284 ( .B1(n6360), .B2(n5099), .A(n5093), .ZN(n5095) );
  NAND2_X1 U6285 ( .A1(n5100), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5094)
         );
  OAI211_X1 U6286 ( .C1(n5872), .C2(n5103), .A(n5095), .B(n5094), .ZN(U3137)
         );
  OAI22_X1 U6287 ( .A1(n6359), .A2(n5097), .B1(n5229), .B2(n5096), .ZN(n5098)
         );
  AOI21_X1 U6288 ( .B1(n6356), .B2(n5099), .A(n5098), .ZN(n5102) );
  NAND2_X1 U6289 ( .A1(n5100), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5101)
         );
  OAI211_X1 U6290 ( .C1(n5868), .C2(n5103), .A(n5102), .B(n5101), .ZN(U3136)
         );
  NAND2_X1 U6291 ( .A1(n5105), .A2(n5104), .ZN(n5164) );
  AOI21_X1 U6292 ( .B1(n5107), .B2(n5164), .A(n5106), .ZN(n5527) );
  INV_X1 U6293 ( .A(n5170), .ZN(n5109) );
  AOI21_X1 U6294 ( .B1(n5109), .B2(n5169), .A(n5108), .ZN(n5111) );
  OR2_X1 U6295 ( .A1(n5111), .A2(n5110), .ZN(n5982) );
  OAI22_X1 U6296 ( .A1(n5982), .A2(n6077), .B1(n6645), .B2(n6081), .ZN(n5112)
         );
  AOI21_X1 U6297 ( .B1(n5527), .B2(n6085), .A(n5112), .ZN(n5113) );
  INV_X1 U6298 ( .A(n5113), .ZN(U2846) );
  OAI222_X1 U6299 ( .A1(n5114), .A2(n6077), .B1(n6081), .B2(n6634), .C1(n6078), 
        .C2(n5351), .ZN(U2848) );
  AOI21_X1 U6300 ( .B1(n5115), .B2(n5191), .A(n6388), .ZN(n5123) );
  OAI21_X1 U6301 ( .B1(n5160), .B2(n6368), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5122) );
  NOR2_X1 U6302 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5117), .ZN(n5155)
         );
  OAI21_X1 U6303 ( .B1(n6571), .B2(n5155), .A(n5118), .ZN(n5121) );
  INV_X1 U6304 ( .A(n5119), .ZN(n5120) );
  AOI211_X2 U6305 ( .C1(n5123), .C2(n5122), .A(n5121), .B(n5120), .ZN(n5163)
         );
  INV_X1 U6306 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5130) );
  OAI22_X1 U6307 ( .A1(n5126), .A2(n5125), .B1(n5841), .B2(n5124), .ZN(n5156)
         );
  AOI22_X1 U6308 ( .A1(n6406), .A2(n5156), .B1(n6404), .B2(n5155), .ZN(n5127)
         );
  OAI21_X1 U6309 ( .B1(n6409), .B2(n5158), .A(n5127), .ZN(n5128) );
  AOI21_X1 U6310 ( .B1(n6405), .B2(n5160), .A(n5128), .ZN(n5129) );
  OAI21_X1 U6311 ( .B1(n5163), .B2(n5130), .A(n5129), .ZN(U3086) );
  INV_X1 U6312 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5134) );
  AOI22_X1 U6313 ( .A1(n6431), .A2(n5156), .B1(n6428), .B2(n5155), .ZN(n5131)
         );
  OAI21_X1 U6314 ( .B1(n5876), .B2(n5158), .A(n5131), .ZN(n5132) );
  AOI21_X1 U6315 ( .B1(n6364), .B2(n5160), .A(n5132), .ZN(n5133) );
  OAI21_X1 U6316 ( .B1(n5163), .B2(n5134), .A(n5133), .ZN(U3090) );
  INV_X1 U6317 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5138) );
  AOI22_X1 U6318 ( .A1(n6394), .A2(n5156), .B1(n6379), .B2(n5155), .ZN(n5135)
         );
  OAI21_X1 U6319 ( .B1(n5854), .B2(n5158), .A(n5135), .ZN(n5136) );
  AOI21_X1 U6320 ( .B1(n6340), .B2(n5160), .A(n5136), .ZN(n5137) );
  OAI21_X1 U6321 ( .B1(n5163), .B2(n5138), .A(n5137), .ZN(U3084) );
  INV_X1 U6322 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5142) );
  AOI22_X1 U6323 ( .A1(n6441), .A2(n5156), .B1(n6437), .B2(n5155), .ZN(n5139)
         );
  OAI21_X1 U6324 ( .B1(n6446), .B2(n5158), .A(n5139), .ZN(n5140) );
  AOI21_X1 U6325 ( .B1(n6438), .B2(n5160), .A(n5140), .ZN(n5141) );
  OAI21_X1 U6326 ( .B1(n5163), .B2(n5142), .A(n5141), .ZN(U3091) );
  INV_X1 U6327 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5146) );
  AOI22_X1 U6328 ( .A1(n6418), .A2(n5156), .B1(n6416), .B2(n5155), .ZN(n5143)
         );
  OAI21_X1 U6329 ( .B1(n5868), .B2(n5158), .A(n5143), .ZN(n5144) );
  AOI21_X1 U6330 ( .B1(n6356), .B2(n5160), .A(n5144), .ZN(n5145) );
  OAI21_X1 U6331 ( .B1(n5163), .B2(n5146), .A(n5145), .ZN(U3088) );
  INV_X1 U6332 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5150) );
  AOI22_X1 U6333 ( .A1(n6412), .A2(n5156), .B1(n6410), .B2(n5155), .ZN(n5147)
         );
  OAI21_X1 U6334 ( .B1(n5864), .B2(n5158), .A(n5147), .ZN(n5148) );
  AOI21_X1 U6335 ( .B1(n6352), .B2(n5160), .A(n5148), .ZN(n5149) );
  OAI21_X1 U6336 ( .B1(n5163), .B2(n5150), .A(n5149), .ZN(U3087) );
  INV_X1 U6337 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5154) );
  AOI22_X1 U6338 ( .A1(n6400), .A2(n5156), .B1(n6398), .B2(n5155), .ZN(n5151)
         );
  OAI21_X1 U6339 ( .B1(n6403), .B2(n5158), .A(n5151), .ZN(n5152) );
  AOI21_X1 U6340 ( .B1(n6399), .B2(n5160), .A(n5152), .ZN(n5153) );
  OAI21_X1 U6341 ( .B1(n5163), .B2(n5154), .A(n5153), .ZN(U3085) );
  INV_X1 U6342 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5162) );
  AOI22_X1 U6343 ( .A1(n6424), .A2(n5156), .B1(n6422), .B2(n5155), .ZN(n5157)
         );
  OAI21_X1 U6344 ( .B1(n5872), .B2(n5158), .A(n5157), .ZN(n5159) );
  AOI21_X1 U6345 ( .B1(n6360), .B2(n5160), .A(n5159), .ZN(n5161) );
  OAI21_X1 U6346 ( .B1(n5163), .B2(n5162), .A(n5161), .ZN(U3089) );
  INV_X1 U6347 ( .A(n5164), .ZN(n5165) );
  AOI21_X1 U6348 ( .B1(n5167), .B2(n5166), .A(n5165), .ZN(n6030) );
  INV_X1 U6349 ( .A(n6030), .ZN(n5172) );
  AOI22_X1 U6350 ( .A1(n5173), .A2(DATAI_12_), .B1(n6098), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5168) );
  OAI21_X1 U6351 ( .B1(n5172), .B2(n5931), .A(n5168), .ZN(U2879) );
  XNOR2_X1 U6352 ( .A(n5170), .B(n5169), .ZN(n6027) );
  AOI22_X1 U6353 ( .A1(n6027), .A2(n6084), .B1(EBX_REG_12__SCAN_IN), .B2(n5583), .ZN(n5171) );
  OAI21_X1 U6354 ( .B1(n5172), .B2(n6078), .A(n5171), .ZN(U2847) );
  INV_X1 U6355 ( .A(n5527), .ZN(n5358) );
  AOI22_X1 U6356 ( .A1(n5173), .A2(DATAI_13_), .B1(n6098), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5174) );
  OAI21_X1 U6357 ( .B1(n5358), .B2(n5931), .A(n5174), .ZN(U2878) );
  NAND2_X1 U6358 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  AND2_X1 U6359 ( .A1(n5178), .A2(n5177), .ZN(n6261) );
  NAND2_X1 U6360 ( .A1(n6058), .A2(n6261), .ZN(n5182) );
  INV_X1 U6361 ( .A(n6186), .ZN(n5179) );
  AOI22_X1 U6362 ( .A1(n6054), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6614), 
        .B2(n5179), .ZN(n5181) );
  NAND2_X1 U6363 ( .A1(n6611), .A2(EBX_REG_3__SCAN_IN), .ZN(n5180) );
  NAND3_X1 U6364 ( .A1(n5182), .A2(n5181), .A3(n5180), .ZN(n5186) );
  INV_X1 U6365 ( .A(REIP_REG_3__SCAN_IN), .ZN(n5184) );
  AOI21_X1 U6366 ( .B1(n5184), .B2(n5183), .A(n5530), .ZN(n5185) );
  AOI211_X1 U6367 ( .C1(n5549), .C2(n5191), .A(n5186), .B(n5185), .ZN(n5187)
         );
  OAI21_X1 U6368 ( .B1(n6065), .B2(n6083), .A(n5187), .ZN(U2824) );
  OAI21_X1 U6369 ( .B1(n5231), .B2(n6430), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5190) );
  NAND2_X1 U6370 ( .A1(n5190), .A2(n6338), .ZN(n5197) );
  INV_X1 U6371 ( .A(n5197), .ZN(n5194) );
  AND2_X1 U6372 ( .A1(n5192), .A2(n5191), .ZN(n6386) );
  NOR2_X1 U6373 ( .A1(n5841), .A2(n6377), .ZN(n5193) );
  AOI22_X1 U6374 ( .A1(n5194), .A2(n6386), .B1(n6289), .B2(n5193), .ZN(n5234)
         );
  NAND3_X1 U6375 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6460), .ZN(n6391) );
  NOR2_X1 U6376 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6391), .ZN(n5198)
         );
  OAI22_X1 U6377 ( .A1(n6475), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n6571), .B2(n5198), .ZN(n5195) );
  INV_X1 U6378 ( .A(n5195), .ZN(n5196) );
  NOR2_X1 U6379 ( .A1(n6290), .A2(n6298), .ZN(n5849) );
  OAI211_X1 U6380 ( .C1(n5197), .C2(n6386), .A(n5196), .B(n5849), .ZN(n5227)
         );
  NAND2_X1 U6381 ( .A1(n5227), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5202)
         );
  INV_X1 U6382 ( .A(n5198), .ZN(n5228) );
  OAI22_X1 U6383 ( .A1(n5199), .A2(n5228), .B1(n6435), .B2(n6445), .ZN(n5200)
         );
  AOI21_X1 U6384 ( .B1(n6429), .B2(n5231), .A(n5200), .ZN(n5201) );
  OAI211_X1 U6385 ( .C1(n5234), .C2(n6367), .A(n5202), .B(n5201), .ZN(U3106)
         );
  NAND2_X1 U6386 ( .A1(n5227), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5206)
         );
  OAI22_X1 U6387 ( .A1(n5203), .A2(n5228), .B1(n6397), .B2(n6445), .ZN(n5204)
         );
  AOI21_X1 U6388 ( .B1(n6380), .B2(n5231), .A(n5204), .ZN(n5205) );
  OAI211_X1 U6389 ( .C1(n5234), .C2(n6343), .A(n5206), .B(n5205), .ZN(U3100)
         );
  NAND2_X1 U6390 ( .A1(n5227), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5210)
         );
  OAI22_X1 U6391 ( .A1(n5207), .A2(n5228), .B1(n6308), .B2(n6445), .ZN(n5208)
         );
  AOI21_X1 U6392 ( .B1(n6344), .B2(n5231), .A(n5208), .ZN(n5209) );
  OAI211_X1 U6393 ( .C1(n5234), .C2(n6347), .A(n5210), .B(n5209), .ZN(U3101)
         );
  NAND2_X1 U6394 ( .A1(n5227), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5214)
         );
  OAI22_X1 U6395 ( .A1(n5211), .A2(n5228), .B1(n6427), .B2(n6445), .ZN(n5212)
         );
  AOI21_X1 U6396 ( .B1(n6423), .B2(n5231), .A(n5212), .ZN(n5213) );
  OAI211_X1 U6397 ( .C1(n5234), .C2(n6363), .A(n5214), .B(n5213), .ZN(U3105)
         );
  NAND2_X1 U6398 ( .A1(n5227), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5218)
         );
  OAI22_X1 U6399 ( .A1(n5215), .A2(n5228), .B1(n6415), .B2(n6445), .ZN(n5216)
         );
  AOI21_X1 U6400 ( .B1(n6411), .B2(n5231), .A(n5216), .ZN(n5217) );
  OAI211_X1 U6401 ( .C1(n5234), .C2(n6355), .A(n5218), .B(n5217), .ZN(U3103)
         );
  NAND2_X1 U6402 ( .A1(n5227), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5222)
         );
  OAI22_X1 U6403 ( .A1(n5219), .A2(n5228), .B1(n6327), .B2(n6445), .ZN(n5220)
         );
  AOI21_X1 U6404 ( .B1(n6371), .B2(n5231), .A(n5220), .ZN(n5221) );
  OAI211_X1 U6405 ( .C1(n5234), .C2(n6375), .A(n5222), .B(n5221), .ZN(U3107)
         );
  NAND2_X1 U6406 ( .A1(n5227), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5226)
         );
  OAI22_X1 U6407 ( .A1(n5223), .A2(n5228), .B1(n6311), .B2(n6445), .ZN(n5224)
         );
  AOI21_X1 U6408 ( .B1(n6348), .B2(n5231), .A(n5224), .ZN(n5225) );
  OAI211_X1 U6409 ( .C1(n5234), .C2(n6351), .A(n5226), .B(n5225), .ZN(U3102)
         );
  NAND2_X1 U6410 ( .A1(n5227), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5233)
         );
  OAI22_X1 U6411 ( .A1(n5229), .A2(n5228), .B1(n6421), .B2(n6445), .ZN(n5230)
         );
  AOI21_X1 U6412 ( .B1(n6417), .B2(n5231), .A(n5230), .ZN(n5232) );
  OAI211_X1 U6413 ( .C1(n5234), .C2(n6359), .A(n5233), .B(n5232), .ZN(U3104)
         );
  AOI21_X1 U6414 ( .B1(n5237), .B2(n5236), .A(n5235), .ZN(n6042) );
  OR2_X1 U6415 ( .A1(n4977), .A2(n5238), .ZN(n5239) );
  NAND2_X1 U6416 ( .A1(n4960), .A2(n5239), .ZN(n6037) );
  OAI22_X1 U6417 ( .A1(n6037), .A2(n6077), .B1(n6036), .B2(n6081), .ZN(n5240)
         );
  AOI21_X1 U6418 ( .B1(n6042), .B2(n6085), .A(n5240), .ZN(n5241) );
  INV_X1 U6419 ( .A(n5241), .ZN(U2849) );
  NOR2_X1 U6420 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  OR2_X1 U6421 ( .A1(n5242), .A2(n5245), .ZN(n5945) );
  AOI21_X1 U6422 ( .B1(n5247), .B2(n5246), .A(n5331), .ZN(n5822) );
  AOI22_X1 U6423 ( .A1(n5822), .A2(n6084), .B1(n5583), .B2(EBX_REG_17__SCAN_IN), .ZN(n5248) );
  OAI21_X1 U6424 ( .B1(n5945), .B2(n6078), .A(n5248), .ZN(U2842) );
  AOI21_X1 U6425 ( .B1(n6054), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6610), 
        .ZN(n5249) );
  OAI21_X1 U6426 ( .B1(n6075), .B2(n5719), .A(n5249), .ZN(n5253) );
  AOI22_X1 U6427 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6611), .B1(n5259), .B2(n5251), .ZN(n5250) );
  OAI21_X1 U6428 ( .B1(n5251), .B2(n6622), .A(n5250), .ZN(n5252) );
  AOI211_X1 U6429 ( .C1(n5961), .C2(n6058), .A(n5253), .B(n5252), .ZN(n5254)
         );
  OAI21_X1 U6430 ( .B1(n5723), .B2(n6060), .A(n5254), .ZN(U2812) );
  INV_X1 U6431 ( .A(n6042), .ZN(n5256) );
  INV_X1 U6432 ( .A(DATAI_10_), .ZN(n6777) );
  OAI222_X1 U6433 ( .A1(n5256), .A2(n5931), .B1(n5255), .B2(n6777), .C1(n5586), 
        .C2(n4313), .ZN(U2881) );
  INV_X1 U6434 ( .A(n5947), .ZN(n5258) );
  AOI21_X1 U6435 ( .B1(n6611), .B2(EBX_REG_17__SCAN_IN), .A(n6610), .ZN(n5257)
         );
  OAI21_X1 U6436 ( .B1(n5258), .B2(n6075), .A(n5257), .ZN(n5266) );
  AOI21_X1 U6437 ( .B1(n5260), .B2(n5259), .A(REIP_REG_17__SCAN_IN), .ZN(n5264) );
  NOR2_X1 U6438 ( .A1(n5547), .A2(n5261), .ZN(n6016) );
  INV_X1 U6439 ( .A(n6016), .ZN(n5263) );
  OAI22_X1 U6440 ( .A1(n5264), .A2(n5263), .B1(n5262), .B2(n6619), .ZN(n5265)
         );
  AOI211_X1 U6441 ( .C1(n6058), .C2(n5822), .A(n5266), .B(n5265), .ZN(n5267)
         );
  OAI21_X1 U6442 ( .B1(n5945), .B2(n6060), .A(n5267), .ZN(U2810) );
  NAND2_X1 U6443 ( .A1(n5269), .A2(n5268), .ZN(n5277) );
  NAND2_X1 U6444 ( .A1(n5278), .A2(n5276), .ZN(n5270) );
  XNOR2_X1 U6445 ( .A(n5277), .B(n5270), .ZN(n6209) );
  NAND2_X1 U6446 ( .A1(n6209), .A2(n6193), .ZN(n5274) );
  AND2_X1 U6447 ( .A1(n6279), .A2(REIP_REG_9__SCAN_IN), .ZN(n6206) );
  NOR2_X1 U6448 ( .A1(n6197), .A2(n5271), .ZN(n5272) );
  AOI211_X1 U6449 ( .C1(n6187), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6206), 
        .B(n5272), .ZN(n5273) );
  OAI211_X1 U6450 ( .C1(n5352), .C2(n5275), .A(n5274), .B(n5273), .ZN(U2977)
         );
  NAND2_X1 U6451 ( .A1(n5342), .A2(n5340), .ZN(n5280) );
  NAND2_X1 U6452 ( .A1(n5277), .A2(n5276), .ZN(n5279) );
  NAND2_X1 U6453 ( .A1(n5279), .A2(n5278), .ZN(n5341) );
  XOR2_X1 U6454 ( .A(n5280), .B(n5341), .Z(n5290) );
  AOI22_X1 U6455 ( .A1(n6187), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6279), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5281) );
  OAI21_X1 U6456 ( .B1(n6197), .B2(n5282), .A(n5281), .ZN(n5283) );
  AOI21_X1 U6457 ( .B1(n6042), .B2(n6181), .A(n5283), .ZN(n5284) );
  OAI21_X1 U6458 ( .B1(n5290), .B2(n6165), .A(n5284), .ZN(U2976) );
  OAI21_X1 U6459 ( .B1(n5369), .B2(n5285), .A(n6221), .ZN(n6208) );
  OAI22_X1 U6460 ( .A1(n6037), .A2(n6255), .B1(n6532), .B2(n6254), .ZN(n5288)
         );
  NAND2_X1 U6461 ( .A1(n5285), .A2(n6214), .ZN(n6212) );
  AOI221_X1 U6462 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n4159), .C2(n5286), .A(n6212), 
        .ZN(n5287) );
  AOI211_X1 U6463 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6208), .A(n5288), .B(n5287), .ZN(n5289) );
  OAI21_X1 U6464 ( .B1(n5290), .B2(n6262), .A(n5289), .ZN(U3008) );
  CLKBUF_X1 U6465 ( .A(n5291), .Z(n5296) );
  INV_X1 U6466 ( .A(n5292), .ZN(n5293) );
  NOR2_X1 U6467 ( .A1(n5294), .A2(n5293), .ZN(n5295) );
  XNOR2_X1 U6468 ( .A(n5296), .B(n5295), .ZN(n5305) );
  OAI221_X1 U6469 ( .B1(n5297), .B2(n6250), .C1(n5297), .C2(n5793), .A(n6204), 
        .ZN(n5298) );
  OAI221_X1 U6470 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .C1(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .C2(n6200), .A(n5298), .ZN(n5300) );
  NOR2_X1 U6471 ( .A1(n6254), .A2(n6534), .ZN(n5302) );
  AOI21_X1 U6472 ( .B1(n6027), .B2(n6273), .A(n5302), .ZN(n5299) );
  OAI211_X1 U6473 ( .C1(n5305), .C2(n6262), .A(n5300), .B(n5299), .ZN(U3006)
         );
  AND2_X1 U6474 ( .A1(n6187), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5301)
         );
  AOI211_X1 U6475 ( .C1(n5946), .C2(n6029), .A(n5302), .B(n5301), .ZN(n5304)
         );
  NAND2_X1 U6476 ( .A1(n6030), .A2(n6181), .ZN(n5303) );
  OAI211_X1 U6477 ( .C1(n5305), .C2(n6165), .A(n5304), .B(n5303), .ZN(U2974)
         );
  INV_X1 U6478 ( .A(n5336), .ZN(n5309) );
  INV_X1 U6479 ( .A(n5307), .ZN(n5308) );
  OAI21_X1 U6480 ( .B1(n5309), .B2(n5308), .A(n5689), .ZN(n5707) );
  INV_X1 U6481 ( .A(n5310), .ZN(n5313) );
  INV_X1 U6482 ( .A(n5311), .ZN(n5799) );
  MUX2_X1 U6483 ( .A(n5313), .B(n5799), .S(n5312), .Z(n5330) );
  NAND2_X1 U6484 ( .A1(n5331), .A2(n5330), .ZN(n5333) );
  INV_X1 U6485 ( .A(n5314), .ZN(n5315) );
  XNOR2_X1 U6486 ( .A(n5333), .B(n5315), .ZN(n5812) );
  INV_X1 U6487 ( .A(n5812), .ZN(n5322) );
  AOI21_X1 U6488 ( .B1(n6614), .B2(n5704), .A(n6610), .ZN(n5316) );
  OAI21_X1 U6489 ( .B1(n6619), .B2(n5701), .A(n5316), .ZN(n5321) );
  OAI21_X1 U6490 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5317), .ZN(n5319) );
  AOI22_X1 U6491 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6611), .B1(
        REIP_REG_19__SCAN_IN), .B2(n6016), .ZN(n5318) );
  OAI21_X1 U6492 ( .B1(n6018), .B2(n5319), .A(n5318), .ZN(n5320) );
  AOI211_X1 U6493 ( .C1(n6058), .C2(n5322), .A(n5321), .B(n5320), .ZN(n5323)
         );
  OAI21_X1 U6494 ( .B1(n5707), .B2(n6060), .A(n5323), .ZN(U2808) );
  NOR2_X2 U6495 ( .A1(n6098), .A2(n5324), .ZN(n6095) );
  AOI22_X1 U6496 ( .A1(n6095), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6098), .ZN(n5328) );
  AND2_X1 U6497 ( .A1(n3012), .A2(n5325), .ZN(n5326) );
  NAND2_X1 U6498 ( .A1(n6099), .A2(DATAI_3_), .ZN(n5327) );
  OAI211_X1 U6499 ( .C1(n5707), .C2(n5931), .A(n5328), .B(n5327), .ZN(U2872)
         );
  INV_X1 U6500 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5329) );
  OAI222_X1 U6501 ( .A1(n6078), .A2(n5707), .B1(n6077), .B2(n5812), .C1(n5329), 
        .C2(n6081), .ZN(U2840) );
  OR2_X1 U6502 ( .A1(n5331), .A2(n5330), .ZN(n5332) );
  INV_X1 U6503 ( .A(n6020), .ZN(n5339) );
  OR2_X1 U6504 ( .A1(n5242), .A2(n5334), .ZN(n5335) );
  AND2_X1 U6505 ( .A1(n5336), .A2(n5335), .ZN(n6088) );
  INV_X1 U6506 ( .A(n6088), .ZN(n5337) );
  OAI222_X1 U6507 ( .A1(n6077), .A2(n5339), .B1(n6081), .B2(n5338), .C1(n6078), 
        .C2(n5337), .ZN(U2841) );
  NAND2_X1 U6508 ( .A1(n5341), .A2(n5340), .ZN(n5343) );
  NAND2_X1 U6509 ( .A1(n5343), .A2(n5342), .ZN(n5345) );
  XNOR2_X1 U6510 ( .A(n5818), .B(n6792), .ZN(n5344) );
  XNOR2_X1 U6511 ( .A(n5345), .B(n5344), .ZN(n6201) );
  NAND2_X1 U6512 ( .A1(n6201), .A2(n6193), .ZN(n5350) );
  INV_X1 U6513 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5346) );
  NOR2_X1 U6514 ( .A1(n6254), .A2(n5346), .ZN(n6198) );
  NOR2_X1 U6515 ( .A1(n6197), .A2(n5347), .ZN(n5348) );
  AOI211_X1 U6516 ( .C1(n6187), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6198), 
        .B(n5348), .ZN(n5349) );
  OAI211_X1 U6517 ( .C1(n5352), .C2(n5351), .A(n5350), .B(n5349), .ZN(U2975)
         );
  XNOR2_X1 U6518 ( .A(n3021), .B(n5354), .ZN(n5988) );
  NAND2_X1 U6519 ( .A1(n5988), .A2(n6193), .ZN(n5357) );
  AND2_X1 U6520 ( .A1(n6279), .A2(REIP_REG_13__SCAN_IN), .ZN(n5983) );
  NOR2_X1 U6521 ( .A1(n6197), .A2(n5521), .ZN(n5355) );
  AOI211_X1 U6522 ( .C1(n6187), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5983), 
        .B(n5355), .ZN(n5356) );
  OAI211_X1 U6523 ( .C1(n5352), .C2(n5358), .A(n5357), .B(n5356), .ZN(U2973)
         );
  INV_X1 U6524 ( .A(n5360), .ZN(n5362) );
  NOR2_X1 U6525 ( .A1(n5362), .A2(n5361), .ZN(n5363) );
  XNOR2_X1 U6526 ( .A(n5359), .B(n5363), .ZN(n5977) );
  NAND2_X1 U6527 ( .A1(n5977), .A2(n6193), .ZN(n5366) );
  OAI22_X1 U6528 ( .A1(n5702), .A2(n6620), .B1(n6254), .B2(n6623), .ZN(n5364)
         );
  AOI21_X1 U6529 ( .B1(n5946), .B2(n6613), .A(n5364), .ZN(n5365) );
  OAI211_X1 U6530 ( .C1(n5352), .C2(n6612), .A(n5366), .B(n5365), .ZN(U2972)
         );
  OAI21_X1 U6531 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5369), .A(n5368), 
        .ZN(n5374) );
  INV_X1 U6532 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6533 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5370) );
  OAI21_X1 U6534 ( .B1(n5378), .B2(n6262), .A(n5377), .ZN(U2987) );
  INV_X1 U6535 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5379) );
  OAI22_X1 U6536 ( .A1(n5380), .A2(n6077), .B1(n5379), .B2(n6081), .ZN(U2828)
         );
  INV_X1 U6537 ( .A(n5398), .ZN(n5381) );
  AOI21_X1 U6538 ( .B1(n5408), .B2(n5381), .A(n6578), .ZN(n5389) );
  AOI22_X1 U6539 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5383), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5382), .ZN(n5405) );
  INV_X1 U6540 ( .A(n5405), .ZN(n5387) );
  NOR2_X1 U6541 ( .A1(n6480), .A2(n5384), .ZN(n5404) );
  INV_X1 U6542 ( .A(n5408), .ZN(n6574) );
  NOR2_X1 U6543 ( .A1(n6574), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5386)
         );
  AOI222_X1 U6544 ( .A1(n5387), .A2(n5404), .B1(n5398), .B2(n5386), .C1(n5385), 
        .C2(n6489), .ZN(n5388) );
  OAI22_X1 U6545 ( .A1(n5389), .A2(n3204), .B1(n6578), .B2(n5388), .ZN(U3459)
         );
  AOI21_X1 U6546 ( .B1(n6448), .B2(n6489), .A(n6578), .ZN(n5396) );
  AND2_X1 U6547 ( .A1(n5390), .A2(n5395), .ZN(n5391) );
  AOI21_X1 U6548 ( .B1(n6385), .B2(n5402), .A(n5391), .ZN(n6450) );
  OAI21_X1 U6549 ( .B1(n6450), .B2(STATE2_REG_3__SCAN_IN), .A(n6480), .ZN(
        n5393) );
  INV_X1 U6550 ( .A(n5404), .ZN(n5392) );
  AOI22_X1 U6551 ( .A1(n5393), .A2(n5392), .B1(n5408), .B2(n5395), .ZN(n5394)
         );
  OAI22_X1 U6552 ( .A1(n5396), .A2(n5395), .B1(n6578), .B2(n5394), .ZN(U3461)
         );
  INV_X1 U6553 ( .A(n6448), .ZN(n5397) );
  NOR2_X1 U6554 ( .A1(n5397), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5401)
         );
  NOR3_X1 U6555 ( .A1(n5399), .A2(n4509), .A3(n5398), .ZN(n5400) );
  AOI211_X1 U6556 ( .C1(n5403), .C2(n5402), .A(n5401), .B(n5400), .ZN(n6451)
         );
  INV_X1 U6557 ( .A(n6489), .ZN(n6576) );
  AOI22_X1 U6558 ( .A1(n5406), .A2(n5408), .B1(n5405), .B2(n5404), .ZN(n5407)
         );
  OAI21_X1 U6559 ( .B1(n6451), .B2(n6576), .A(n5407), .ZN(n5410) );
  AOI22_X1 U6560 ( .A1(n5412), .A2(n5410), .B1(n5409), .B2(n5408), .ZN(n5411)
         );
  OAI21_X1 U6561 ( .B1(n5413), .B2(n5412), .A(n5411), .ZN(U3460) );
  INV_X1 U6562 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5697) );
  OAI21_X1 U6563 ( .B1(n5414), .B2(n5697), .A(n5818), .ZN(n5415) );
  AND2_X2 U6564 ( .A1(n5696), .A2(n5415), .ZN(n5685) );
  XNOR2_X1 U6565 ( .A(n5818), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5684)
         );
  NAND2_X2 U6566 ( .A1(n5685), .A2(n5684), .ZN(n5659) );
  OR2_X1 U6567 ( .A1(n5625), .A2(n5416), .ZN(n5417) );
  INV_X1 U6568 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5789) );
  XNOR2_X1 U6569 ( .A(n5818), .B(n5789), .ZN(n5678) );
  NOR2_X1 U6570 ( .A1(n5818), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5669)
         );
  NAND2_X1 U6571 ( .A1(n5676), .A2(n5669), .ZN(n5661) );
  INV_X1 U6572 ( .A(n5676), .ZN(n5418) );
  NAND3_X1 U6573 ( .A1(n5625), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5419) );
  XNOR2_X1 U6574 ( .A(n5420), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5436)
         );
  NOR2_X1 U6575 ( .A1(n5508), .A2(n5422), .ZN(n5423) );
  OR2_X1 U6576 ( .A1(n5421), .A2(n5423), .ZN(n5574) );
  INV_X1 U6577 ( .A(n5574), .ZN(n5502) );
  INV_X1 U6578 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5498) );
  NOR2_X1 U6579 ( .A1(n6254), .A2(n5498), .ZN(n5432) );
  AOI21_X1 U6580 ( .B1(n5770), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5425) );
  INV_X1 U6581 ( .A(n5761), .ZN(n5424) );
  NOR2_X1 U6582 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  AOI211_X1 U6583 ( .C1(n6273), .C2(n5502), .A(n5432), .B(n5426), .ZN(n5427)
         );
  OAI21_X1 U6584 ( .B1(n5436), .B2(n6262), .A(n5427), .ZN(U2994) );
  INV_X1 U6585 ( .A(n5428), .ZN(n5431) );
  INV_X1 U6586 ( .A(n5429), .ZN(n5430) );
  AOI21_X1 U6587 ( .B1(n5431), .B2(n5430), .A(n5484), .ZN(n5494) );
  AOI21_X1 U6588 ( .B1(n6187), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5432), 
        .ZN(n5433) );
  OAI21_X1 U6589 ( .B1(n6197), .B2(n5495), .A(n5433), .ZN(n5434) );
  AOI21_X1 U6590 ( .B1(n5494), .B2(n6181), .A(n5434), .ZN(n5435) );
  OAI21_X1 U6591 ( .B1(n5436), .B2(n6165), .A(n5435), .ZN(U2962) );
  NOR3_X1 U6592 ( .A1(n5437), .A2(REIP_REG_30__SCAN_IN), .A3(n6557), .ZN(n5442) );
  NAND2_X1 U6593 ( .A1(n5552), .A2(n6058), .ZN(n5440) );
  AOI22_X1 U6594 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6054), .B1(n6614), 
        .B2(n5438), .ZN(n5439) );
  OAI211_X1 U6595 ( .C1(n5554), .C2(n6035), .A(n5440), .B(n5439), .ZN(n5441)
         );
  OAI21_X1 U6596 ( .B1(n5593), .B2(n6060), .A(n5444), .ZN(U2797) );
  NAND2_X1 U6597 ( .A1(n5458), .A2(n5446), .ZN(n5447) );
  XNOR2_X1 U6598 ( .A(n5459), .B(n5449), .ZN(n5725) );
  INV_X1 U6599 ( .A(n5725), .ZN(n5555) );
  OAI22_X1 U6600 ( .A1(n6654), .A2(n6619), .B1(n6075), .B2(n5621), .ZN(n5450)
         );
  AOI21_X1 U6601 ( .B1(EBX_REG_29__SCAN_IN), .B2(n6611), .A(n5450), .ZN(n5451)
         );
  OAI21_X1 U6602 ( .B1(n5464), .B2(n6557), .A(n5451), .ZN(n5452) );
  AOI21_X1 U6603 ( .B1(n5555), .B2(n6058), .A(n5452), .ZN(n5454) );
  OAI211_X1 U6604 ( .C1(n5596), .C2(n6060), .A(n5454), .B(n5453), .ZN(U2798)
         );
  OR2_X1 U6605 ( .A1(n5558), .A2(n5456), .ZN(n5457) );
  AND2_X1 U6606 ( .A1(n5458), .A2(n5457), .ZN(n5635) );
  INV_X1 U6607 ( .A(n5635), .ZN(n5599) );
  OAI21_X1 U6608 ( .B1(n5564), .B2(n5460), .A(n5459), .ZN(n5733) );
  INV_X1 U6609 ( .A(n5733), .ZN(n5467) );
  INV_X1 U6610 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6763) );
  OAI22_X1 U6611 ( .A1(n5461), .A2(n6619), .B1(n6075), .B2(n5633), .ZN(n5462)
         );
  AOI21_X1 U6612 ( .B1(n6611), .B2(EBX_REG_28__SCAN_IN), .A(n5462), .ZN(n5463)
         );
  OAI21_X1 U6613 ( .B1(n5464), .B2(n6763), .A(n5463), .ZN(n5466) );
  INV_X1 U6614 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6555) );
  NOR3_X1 U6615 ( .A1(n5896), .A2(REIP_REG_28__SCAN_IN), .A3(n6555), .ZN(n5465) );
  AOI211_X1 U6616 ( .C1(n6058), .C2(n5467), .A(n5466), .B(n5465), .ZN(n5468)
         );
  OAI21_X1 U6617 ( .B1(n5599), .B2(n6060), .A(n5468), .ZN(U2799) );
  INV_X1 U6618 ( .A(n5482), .ZN(n5471) );
  INV_X1 U6619 ( .A(n5469), .ZN(n5470) );
  OAI21_X1 U6620 ( .B1(n5471), .B2(n5470), .A(n5559), .ZN(n5651) );
  INV_X1 U6621 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U6622 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5486), .ZN(n5489) );
  INV_X1 U6623 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6641) );
  OAI21_X1 U6624 ( .B1(n6803), .B2(n5489), .A(n6641), .ZN(n5477) );
  NAND2_X1 U6625 ( .A1(n5481), .A2(n5472), .ZN(n5473) );
  NAND2_X1 U6626 ( .A1(n5562), .A2(n5473), .ZN(n5750) );
  OAI22_X1 U6627 ( .A1(n5568), .A2(n6035), .B1(n5647), .B2(n6075), .ZN(n5474)
         );
  AOI21_X1 U6628 ( .B1(n6054), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5474), 
        .ZN(n5475) );
  OAI21_X1 U6629 ( .B1(n5750), .B2(n6624), .A(n5475), .ZN(n5476) );
  AOI21_X1 U6630 ( .B1(n5477), .B2(n5889), .A(n5476), .ZN(n5478) );
  OAI21_X1 U6631 ( .B1(n5651), .B2(n6060), .A(n5478), .ZN(U2801) );
  OR2_X1 U6632 ( .A1(n5421), .A2(n5479), .ZN(n5480) );
  NAND2_X1 U6633 ( .A1(n5481), .A2(n5480), .ZN(n5757) );
  OAI21_X1 U6634 ( .B1(n5484), .B2(n5483), .A(n5482), .ZN(n5654) );
  INV_X1 U6635 ( .A(n5654), .ZN(n5485) );
  NAND2_X1 U6636 ( .A1(n5485), .A2(n6615), .ZN(n5493) );
  NAND2_X1 U6637 ( .A1(n6054), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5488)
         );
  INV_X1 U6638 ( .A(n5499), .ZN(n5513) );
  AND2_X1 U6639 ( .A1(n5498), .A2(n5486), .ZN(n5500) );
  OAI21_X1 U6640 ( .B1(n5513), .B2(n5500), .A(REIP_REG_25__SCAN_IN), .ZN(n5487) );
  OAI211_X1 U6641 ( .C1(REIP_REG_25__SCAN_IN), .C2(n5489), .A(n5488), .B(n5487), .ZN(n5491) );
  NOR2_X1 U6642 ( .A1(n6035), .A2(n5571), .ZN(n5490) );
  AOI211_X1 U6643 ( .C1(n6614), .C2(n5657), .A(n5491), .B(n5490), .ZN(n5492)
         );
  OAI211_X1 U6644 ( .C1(n6624), .C2(n5757), .A(n5493), .B(n5492), .ZN(U2802)
         );
  INV_X1 U6645 ( .A(n5494), .ZN(n5609) );
  OAI22_X1 U6646 ( .A1(n6806), .A2(n6619), .B1(n6075), .B2(n5495), .ZN(n5496)
         );
  AOI21_X1 U6647 ( .B1(EBX_REG_24__SCAN_IN), .B2(n6611), .A(n5496), .ZN(n5497)
         );
  OAI21_X1 U6648 ( .B1(n5499), .B2(n5498), .A(n5497), .ZN(n5501) );
  AOI211_X1 U6649 ( .C1(n6058), .C2(n5502), .A(n5501), .B(n5500), .ZN(n5503)
         );
  OAI21_X1 U6650 ( .B1(n5609), .B2(n6060), .A(n5503), .ZN(U2803) );
  INV_X1 U6651 ( .A(n5504), .ZN(n5506) );
  INV_X1 U6652 ( .A(n5505), .ZN(n5580) );
  AOI21_X1 U6653 ( .B1(n5506), .B2(n5580), .A(n5429), .ZN(n5667) );
  INV_X1 U6654 ( .A(n5667), .ZN(n5612) );
  INV_X1 U6655 ( .A(n5582), .ZN(n5782) );
  AOI21_X1 U6656 ( .B1(n5782), .B2(n5581), .A(n5507), .ZN(n5509) );
  NOR2_X1 U6657 ( .A1(n5509), .A2(n5508), .ZN(n5765) );
  INV_X1 U6658 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5577) );
  OAI22_X1 U6659 ( .A1(n5577), .A2(n6035), .B1(n5510), .B2(n6619), .ZN(n5512)
         );
  NOR2_X1 U6660 ( .A1(n6075), .A2(n5665), .ZN(n5511) );
  AOI211_X1 U6661 ( .C1(n5765), .C2(n6058), .A(n5512), .B(n5511), .ZN(n5516)
         );
  NAND2_X1 U6662 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5903) );
  INV_X1 U6663 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6548) );
  OAI21_X1 U6664 ( .B1(n5903), .B2(n5915), .A(n6548), .ZN(n5514) );
  NAND2_X1 U6665 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  OAI211_X1 U6666 ( .C1(n5612), .C2(n6060), .A(n5516), .B(n5515), .ZN(U2804)
         );
  INV_X1 U6667 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5519) );
  INV_X1 U6668 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6779) );
  NAND3_X1 U6669 ( .A1(n6025), .A2(n6779), .A3(n5517), .ZN(n5518) );
  OAI211_X1 U6670 ( .C1(n6619), .C2(n5519), .A(n6066), .B(n5518), .ZN(n5526)
         );
  OAI21_X1 U6671 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6608), .A(n5520), .ZN(n5523) );
  OAI22_X1 U6672 ( .A1(n6035), .A2(n6645), .B1(n6075), .B2(n5521), .ZN(n5522)
         );
  AOI21_X1 U6673 ( .B1(n5523), .B2(REIP_REG_13__SCAN_IN), .A(n5522), .ZN(n5524) );
  OAI21_X1 U6674 ( .B1(n5982), .B2(n6624), .A(n5524), .ZN(n5525) );
  AOI211_X1 U6675 ( .C1(n5527), .C2(n6615), .A(n5526), .B(n5525), .ZN(n5528)
         );
  INV_X1 U6676 ( .A(n5528), .ZN(U2814) );
  INV_X1 U6677 ( .A(n5529), .ZN(n5534) );
  OAI221_X1 U6678 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5531), .C1(n6520), .C2(
        n5530), .A(n6066), .ZN(n5532) );
  AOI21_X1 U6679 ( .B1(n6054), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5532), 
        .ZN(n5533) );
  OAI21_X1 U6680 ( .B1(n6075), .B2(n5534), .A(n5533), .ZN(n5535) );
  AOI21_X1 U6681 ( .B1(n6611), .B2(EBX_REG_4__SCAN_IN), .A(n5535), .ZN(n5536)
         );
  OAI21_X1 U6682 ( .B1(n6624), .B2(n6256), .A(n5536), .ZN(n5537) );
  AOI21_X1 U6683 ( .B1(n5549), .B2(n5538), .A(n5537), .ZN(n5539) );
  OAI21_X1 U6684 ( .B1(n5540), .B2(n6065), .A(n5539), .ZN(U2823) );
  AOI21_X1 U6685 ( .B1(n6619), .B2(n6075), .A(n5541), .ZN(n5542) );
  AOI21_X1 U6686 ( .B1(n6611), .B2(EBX_REG_0__SCAN_IN), .A(n5542), .ZN(n5545)
         );
  NAND2_X1 U6687 ( .A1(n6058), .A2(n5543), .ZN(n5544) );
  OAI211_X1 U6688 ( .C1(n5547), .C2(n5546), .A(n5545), .B(n5544), .ZN(n5548)
         );
  AOI21_X1 U6689 ( .B1(n6385), .B2(n5549), .A(n5548), .ZN(n5550) );
  OAI21_X1 U6690 ( .B1(n5551), .B2(n6065), .A(n5550), .ZN(U2827) );
  INV_X1 U6691 ( .A(n5552), .ZN(n5553) );
  OAI222_X1 U6692 ( .A1(n6078), .A2(n5593), .B1(n6081), .B2(n5554), .C1(n5553), 
        .C2(n6077), .ZN(U2829) );
  AOI22_X1 U6693 ( .A1(n5555), .A2(n6084), .B1(n5583), .B2(EBX_REG_29__SCAN_IN), .ZN(n5556) );
  OAI21_X1 U6694 ( .B1(n5596), .B2(n6078), .A(n5556), .ZN(U2830) );
  OAI222_X1 U6695 ( .A1(n5557), .A2(n6081), .B1(n6077), .B2(n5733), .C1(n5599), 
        .C2(n6078), .ZN(U2831) );
  AOI21_X1 U6696 ( .B1(n5560), .B2(n5559), .A(n5558), .ZN(n5894) );
  INV_X1 U6697 ( .A(n5894), .ZN(n5602) );
  AND2_X1 U6698 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  OR2_X1 U6699 ( .A1(n5564), .A2(n5563), .ZN(n5892) );
  INV_X1 U6700 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5565) );
  OAI22_X1 U6701 ( .A1(n5892), .A2(n6077), .B1(n5565), .B2(n6081), .ZN(n5566)
         );
  INV_X1 U6702 ( .A(n5566), .ZN(n5567) );
  OAI21_X1 U6703 ( .B1(n5602), .B2(n6078), .A(n5567), .ZN(U2832) );
  OAI22_X1 U6704 ( .A1(n5750), .A2(n6077), .B1(n5568), .B2(n6081), .ZN(n5569)
         );
  INV_X1 U6705 ( .A(n5569), .ZN(n5570) );
  OAI21_X1 U6706 ( .B1(n5651), .B2(n6078), .A(n5570), .ZN(U2833) );
  OAI22_X1 U6707 ( .A1(n5757), .A2(n6077), .B1(n5571), .B2(n6081), .ZN(n5572)
         );
  INV_X1 U6708 ( .A(n5572), .ZN(n5573) );
  OAI21_X1 U6709 ( .B1(n5654), .B2(n6078), .A(n5573), .ZN(U2834) );
  INV_X1 U6710 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5575) );
  OAI222_X1 U6711 ( .A1(n6078), .A2(n5609), .B1(n6081), .B2(n5575), .C1(n5574), 
        .C2(n6077), .ZN(U2835) );
  INV_X1 U6712 ( .A(n5765), .ZN(n5576) );
  OAI222_X1 U6713 ( .A1(n6078), .A2(n5612), .B1(n6081), .B2(n5577), .C1(n5576), 
        .C2(n6077), .ZN(U2836) );
  OAI21_X1 U6714 ( .B1(n5691), .B2(n5681), .A(n5578), .ZN(n5579) );
  INV_X1 U6715 ( .A(n5902), .ZN(n5615) );
  XNOR2_X1 U6716 ( .A(n5582), .B(n5581), .ZN(n5901) );
  AOI22_X1 U6717 ( .A1(n5901), .A2(n6084), .B1(EBX_REG_22__SCAN_IN), .B2(n5583), .ZN(n5584) );
  OAI21_X1 U6718 ( .B1(n5615), .B2(n6078), .A(n5584), .ZN(U2837) );
  NAND2_X1 U6719 ( .A1(n5588), .A2(n5587), .ZN(n5590) );
  AOI22_X1 U6720 ( .A1(n6095), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6098), .ZN(n5589) );
  NAND2_X1 U6721 ( .A1(n5590), .A2(n5589), .ZN(U2860) );
  AOI22_X1 U6722 ( .A1(n6095), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6098), .ZN(n5592) );
  NAND2_X1 U6723 ( .A1(n6099), .A2(DATAI_14_), .ZN(n5591) );
  OAI211_X1 U6724 ( .C1(n5593), .C2(n5931), .A(n5592), .B(n5591), .ZN(U2861)
         );
  AOI22_X1 U6725 ( .A1(n6095), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6098), .ZN(n5595) );
  NAND2_X1 U6726 ( .A1(n6099), .A2(DATAI_13_), .ZN(n5594) );
  OAI211_X1 U6727 ( .C1(n5596), .C2(n5931), .A(n5595), .B(n5594), .ZN(U2862)
         );
  AOI22_X1 U6728 ( .A1(n6095), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6098), .ZN(n5598) );
  NAND2_X1 U6729 ( .A1(n6099), .A2(DATAI_12_), .ZN(n5597) );
  OAI211_X1 U6730 ( .C1(n5599), .C2(n5931), .A(n5598), .B(n5597), .ZN(U2863)
         );
  AOI22_X1 U6731 ( .A1(n6099), .A2(DATAI_11_), .B1(n6098), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U6732 ( .A1(n6095), .A2(DATAI_27_), .ZN(n5600) );
  OAI211_X1 U6733 ( .C1(n5602), .C2(n5931), .A(n5601), .B(n5600), .ZN(U2864)
         );
  AOI22_X1 U6734 ( .A1(n6095), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6098), .ZN(n5604) );
  NAND2_X1 U6735 ( .A1(n6099), .A2(DATAI_10_), .ZN(n5603) );
  OAI211_X1 U6736 ( .C1(n5651), .C2(n5931), .A(n5604), .B(n5603), .ZN(U2865)
         );
  AOI22_X1 U6737 ( .A1(n6095), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6098), .ZN(n5606) );
  NAND2_X1 U6738 ( .A1(n6099), .A2(DATAI_9_), .ZN(n5605) );
  OAI211_X1 U6739 ( .C1(n5654), .C2(n5931), .A(n5606), .B(n5605), .ZN(U2866)
         );
  AOI22_X1 U6740 ( .A1(n6095), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6098), .ZN(n5608) );
  NAND2_X1 U6741 ( .A1(n6099), .A2(DATAI_8_), .ZN(n5607) );
  OAI211_X1 U6742 ( .C1(n5609), .C2(n5931), .A(n5608), .B(n5607), .ZN(U2867)
         );
  AOI22_X1 U6743 ( .A1(n6095), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6098), .ZN(n5611) );
  NAND2_X1 U6744 ( .A1(n6099), .A2(DATAI_7_), .ZN(n5610) );
  OAI211_X1 U6745 ( .C1(n5612), .C2(n5931), .A(n5611), .B(n5610), .ZN(U2868)
         );
  AOI22_X1 U6746 ( .A1(n6099), .A2(DATAI_6_), .B1(n6098), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U6747 ( .A1(n6095), .A2(DATAI_22_), .ZN(n5613) );
  OAI211_X1 U6748 ( .C1(n5615), .C2(n5931), .A(n5614), .B(n5613), .ZN(U2869)
         );
  INV_X1 U6749 ( .A(n5616), .ZN(n5618) );
  NAND2_X1 U6750 ( .A1(n5618), .A2(n3033), .ZN(n5619) );
  XNOR2_X1 U6751 ( .A(n5619), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5731)
         );
  NAND2_X1 U6752 ( .A1(n6279), .A2(REIP_REG_29__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U6753 ( .A1(n6187), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5620)
         );
  OAI211_X1 U6754 ( .C1(n6197), .C2(n5621), .A(n5724), .B(n5620), .ZN(n5622)
         );
  AOI21_X1 U6755 ( .B1(n5623), .B2(n6181), .A(n5622), .ZN(n5624) );
  OAI21_X1 U6756 ( .B1(n5731), .B2(n6165), .A(n5624), .ZN(U2957) );
  NAND3_X1 U6757 ( .A1(n3014), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5625), .ZN(n5630) );
  NAND2_X1 U6758 ( .A1(n5643), .A2(n5627), .ZN(n5628) );
  OR2_X1 U6759 ( .A1(n5626), .A2(n5628), .ZN(n5637) );
  AOI22_X1 U6760 ( .A1(n5630), .A2(n5637), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5629), .ZN(n5631) );
  XNOR2_X1 U6761 ( .A(n5631), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5740)
         );
  NAND2_X1 U6762 ( .A1(n6279), .A2(REIP_REG_28__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U6763 ( .A1(n6187), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5632)
         );
  OAI211_X1 U6764 ( .C1(n6197), .C2(n5633), .A(n5732), .B(n5632), .ZN(n5634)
         );
  AOI21_X1 U6765 ( .B1(n5635), .B2(n6181), .A(n5634), .ZN(n5636) );
  OAI21_X1 U6766 ( .B1(n5740), .B2(n6165), .A(n5636), .ZN(U2958) );
  NAND2_X1 U6767 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  XNOR2_X1 U6768 ( .A(n5639), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5748)
         );
  NAND2_X1 U6769 ( .A1(n5946), .A2(n5885), .ZN(n5640) );
  NAND2_X1 U6770 ( .A1(n6279), .A2(REIP_REG_27__SCAN_IN), .ZN(n5741) );
  OAI211_X1 U6771 ( .C1(n5702), .C2(n5887), .A(n5640), .B(n5741), .ZN(n5641)
         );
  AOI21_X1 U6772 ( .B1(n5894), .B2(n6181), .A(n5641), .ZN(n5642) );
  OAI21_X1 U6773 ( .B1(n5748), .B2(n6165), .A(n5642), .ZN(U2959) );
  NOR2_X1 U6774 ( .A1(n5644), .A2(n5643), .ZN(n5645) );
  XNOR2_X1 U6775 ( .A(n3014), .B(n5645), .ZN(n5749) );
  NAND2_X1 U6776 ( .A1(n5749), .A2(n6193), .ZN(n5650) );
  NOR2_X1 U6777 ( .A1(n6254), .A2(n6641), .ZN(n5752) );
  NOR2_X1 U6778 ( .A1(n6197), .A2(n5647), .ZN(n5648) );
  AOI211_X1 U6779 ( .C1(n6187), .C2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5752), 
        .B(n5648), .ZN(n5649) );
  OAI211_X1 U6780 ( .C1(n5352), .C2(n5651), .A(n5650), .B(n5649), .ZN(U2960)
         );
  AOI21_X1 U6781 ( .B1(n5652), .B2(n5626), .A(n4180), .ZN(n5763) );
  OR2_X1 U6782 ( .A1(n6254), .A2(n6803), .ZN(n5756) );
  OAI21_X1 U6783 ( .B1(n5702), .B2(n5653), .A(n5756), .ZN(n5656) );
  NOR2_X1 U6784 ( .A1(n5654), .A2(n5352), .ZN(n5655) );
  AOI211_X1 U6785 ( .C1(n5946), .C2(n5657), .A(n5656), .B(n5655), .ZN(n5658)
         );
  OAI21_X1 U6786 ( .B1(n5763), .B2(n6165), .A(n5658), .ZN(U2961) );
  NAND2_X1 U6787 ( .A1(n5805), .A2(n5660), .ZN(n5662) );
  OAI21_X1 U6788 ( .B1(n5659), .B2(n5662), .A(n5661), .ZN(n5663) );
  XNOR2_X1 U6789 ( .A(n5663), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5772)
         );
  NOR2_X1 U6790 ( .A1(n6254), .A2(n6548), .ZN(n5764) );
  AOI21_X1 U6791 ( .B1(n6187), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5764), 
        .ZN(n5664) );
  OAI21_X1 U6792 ( .B1(n6197), .B2(n5665), .A(n5664), .ZN(n5666) );
  AOI21_X1 U6793 ( .B1(n5667), .B2(n6181), .A(n5666), .ZN(n5668) );
  OAI21_X1 U6794 ( .B1(n5772), .B2(n6165), .A(n5668), .ZN(U2963) );
  AOI21_X1 U6795 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5818), .A(n5669), 
        .ZN(n5670) );
  XNOR2_X1 U6796 ( .A(n5671), .B(n5670), .ZN(n5781) );
  INV_X1 U6797 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5672) );
  NOR2_X1 U6798 ( .A1(n6254), .A2(n5672), .ZN(n5775) );
  AOI21_X1 U6799 ( .B1(n6187), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5775), 
        .ZN(n5673) );
  OAI21_X1 U6800 ( .B1(n6197), .B2(n5897), .A(n5673), .ZN(n5674) );
  AOI21_X1 U6801 ( .B1(n5902), .B2(n6181), .A(n5674), .ZN(n5675) );
  OAI21_X1 U6802 ( .B1(n5781), .B2(n6165), .A(n5675), .ZN(U2964) );
  AOI21_X1 U6803 ( .B1(n5678), .B2(n5677), .A(n5676), .ZN(n5792) );
  INV_X1 U6804 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5679) );
  NOR2_X1 U6805 ( .A1(n6254), .A2(n5679), .ZN(n5785) );
  NOR2_X1 U6806 ( .A1(n5702), .A2(n5910), .ZN(n5680) );
  AOI211_X1 U6807 ( .C1(n5946), .C2(n5912), .A(n5785), .B(n5680), .ZN(n5683)
         );
  XOR2_X1 U6808 ( .A(n5681), .B(n5691), .Z(n5932) );
  NAND2_X1 U6809 ( .A1(n5932), .A2(n6181), .ZN(n5682) );
  OAI211_X1 U6810 ( .C1(n5792), .C2(n6165), .A(n5683), .B(n5682), .ZN(U2965)
         );
  OAI21_X1 U6811 ( .B1(n5685), .B2(n5684), .A(n5659), .ZN(n5809) );
  INV_X1 U6812 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5686) );
  OR2_X1 U6813 ( .A1(n6254), .A2(n5686), .ZN(n5803) );
  OAI21_X1 U6814 ( .B1(n5702), .B2(n5687), .A(n5803), .ZN(n5693) );
  NAND2_X1 U6815 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  NAND2_X1 U6816 ( .A1(n5691), .A2(n5690), .ZN(n5935) );
  NOR2_X1 U6817 ( .A1(n5935), .A2(n5352), .ZN(n5692) );
  AOI211_X1 U6818 ( .C1(n5946), .C2(n5919), .A(n5693), .B(n5692), .ZN(n5694)
         );
  OAI21_X1 U6819 ( .B1(n5809), .B2(n6165), .A(n5694), .ZN(U2966) );
  INV_X1 U6820 ( .A(n5695), .ZN(n5698) );
  OAI21_X1 U6821 ( .B1(n5698), .B2(n5697), .A(n5696), .ZN(n5699) );
  XNOR2_X1 U6822 ( .A(n5699), .B(n3024), .ZN(n5810) );
  NAND2_X1 U6823 ( .A1(n5810), .A2(n6193), .ZN(n5706) );
  INV_X1 U6824 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5700) );
  OR2_X1 U6825 ( .A1(n6254), .A2(n5700), .ZN(n5811) );
  OAI21_X1 U6826 ( .B1(n5702), .B2(n5701), .A(n5811), .ZN(n5703) );
  AOI21_X1 U6827 ( .B1(n5704), .B2(n5946), .A(n5703), .ZN(n5705) );
  OAI211_X1 U6828 ( .C1(n5352), .C2(n5707), .A(n5706), .B(n5705), .ZN(U2967)
         );
  XNOR2_X1 U6829 ( .A(n5818), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5710)
         );
  XNOR2_X1 U6830 ( .A(n5709), .B(n5710), .ZN(n5836) );
  AOI22_X1 U6831 ( .A1(n6187), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6279), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U6832 ( .A1(n5711), .A2(n5946), .ZN(n5712) );
  OAI211_X1 U6833 ( .C1(n6094), .C2(n5352), .A(n5713), .B(n5712), .ZN(n5714)
         );
  INV_X1 U6834 ( .A(n5714), .ZN(n5715) );
  OAI21_X1 U6835 ( .B1(n5836), .B2(n6165), .A(n5715), .ZN(U2970) );
  XNOR2_X1 U6836 ( .A(n5818), .B(n5717), .ZN(n5718) );
  XNOR2_X1 U6837 ( .A(n5716), .B(n5718), .ZN(n5964) );
  NAND2_X1 U6838 ( .A1(n5964), .A2(n6193), .ZN(n5722) );
  NOR2_X1 U6839 ( .A1(n6254), .A2(n5251), .ZN(n5960) );
  NOR2_X1 U6840 ( .A1(n5719), .A2(n6197), .ZN(n5720) );
  AOI211_X1 U6841 ( .C1(n6187), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5960), 
        .B(n5720), .ZN(n5721) );
  OAI211_X1 U6842 ( .C1(n5352), .C2(n5723), .A(n5722), .B(n5721), .ZN(U2971)
         );
  OAI21_X1 U6843 ( .B1(n5725), .B2(n6255), .A(n5724), .ZN(n5726) );
  AOI21_X1 U6844 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5727), .A(n5726), 
        .ZN(n5730) );
  NAND3_X1 U6845 ( .A1(n5746), .A2(n4253), .A3(n5728), .ZN(n5729) );
  OAI211_X1 U6846 ( .C1(n5731), .C2(n6262), .A(n5730), .B(n5729), .ZN(U2989)
         );
  INV_X1 U6847 ( .A(n5742), .ZN(n5738) );
  OAI21_X1 U6848 ( .B1(n5733), .B2(n6255), .A(n5732), .ZN(n5737) );
  INV_X1 U6849 ( .A(n5746), .ZN(n5735) );
  NOR3_X1 U6850 ( .A1(n5735), .A2(n5734), .A3(n4253), .ZN(n5736) );
  AOI211_X1 U6851 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5738), .A(n5737), .B(n5736), .ZN(n5739) );
  OAI21_X1 U6852 ( .B1(n5740), .B2(n6262), .A(n5739), .ZN(U2990) );
  INV_X1 U6853 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5745) );
  OAI21_X1 U6854 ( .B1(n5892), .B2(n6255), .A(n5741), .ZN(n5744) );
  NOR2_X1 U6855 ( .A1(n5742), .A2(n5745), .ZN(n5743) );
  AOI211_X1 U6856 ( .C1(n5746), .C2(n5745), .A(n5744), .B(n5743), .ZN(n5747)
         );
  OAI21_X1 U6857 ( .B1(n5748), .B2(n6262), .A(n5747), .ZN(U2991) );
  XNOR2_X1 U6858 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U6859 ( .A1(n5749), .A2(n6277), .ZN(n5754) );
  NOR2_X1 U6860 ( .A1(n5750), .A2(n6255), .ZN(n5751) );
  AOI211_X1 U6861 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5761), .A(n5752), .B(n5751), .ZN(n5753) );
  OAI211_X1 U6862 ( .C1(n5758), .C2(n5755), .A(n5754), .B(n5753), .ZN(U2992)
         );
  OAI21_X1 U6863 ( .B1(n5757), .B2(n6255), .A(n5756), .ZN(n5760) );
  NOR2_X1 U6864 ( .A1(n5758), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5759)
         );
  AOI211_X1 U6865 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5761), .A(n5760), .B(n5759), .ZN(n5762) );
  OAI21_X1 U6866 ( .B1(n5763), .B2(n6262), .A(n5762), .ZN(U2993) );
  AOI21_X1 U6867 ( .B1(n5765), .B2(n6273), .A(n5764), .ZN(n5766) );
  OAI21_X1 U6868 ( .B1(n5767), .B2(n5769), .A(n5766), .ZN(n5768) );
  AOI21_X1 U6869 ( .B1(n5770), .B2(n5769), .A(n5768), .ZN(n5771) );
  OAI21_X1 U6870 ( .B1(n5772), .B2(n6262), .A(n5771), .ZN(U2995) );
  INV_X1 U6871 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5773) );
  NOR2_X1 U6872 ( .A1(n5787), .A2(n5773), .ZN(n5774) );
  AOI211_X1 U6873 ( .C1(n6273), .C2(n5901), .A(n5775), .B(n5774), .ZN(n5780)
         );
  INV_X1 U6874 ( .A(n5776), .ZN(n5777) );
  NAND3_X1 U6875 ( .A1(n5790), .A2(n5778), .A3(n5777), .ZN(n5779) );
  OAI211_X1 U6876 ( .C1(n5781), .C2(n6262), .A(n5780), .B(n5779), .ZN(U2996)
         );
  AOI21_X1 U6877 ( .B1(n5784), .B2(n5783), .A(n5782), .ZN(n5924) );
  AOI21_X1 U6878 ( .B1(n5924), .B2(n6273), .A(n5785), .ZN(n5786) );
  OAI21_X1 U6879 ( .B1(n5787), .B2(n5789), .A(n5786), .ZN(n5788) );
  AOI21_X1 U6880 ( .B1(n5790), .B2(n5789), .A(n5788), .ZN(n5791) );
  OAI21_X1 U6881 ( .B1(n5792), .B2(n6262), .A(n5791), .ZN(U2997) );
  AOI21_X1 U6882 ( .B1(n5794), .B2(n5793), .A(INSTADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n5795) );
  INV_X1 U6883 ( .A(n5795), .ZN(n5796) );
  AND2_X1 U6884 ( .A1(n5824), .A2(n5796), .ZN(n5958) );
  NAND2_X1 U6885 ( .A1(n6227), .A2(n5957), .ZN(n5797) );
  NAND2_X1 U6886 ( .A1(n5958), .A2(n5797), .ZN(n5814) );
  MUX2_X1 U6887 ( .A(n5800), .B(n5799), .S(n5798), .Z(n5802) );
  XNOR2_X1 U6888 ( .A(n5802), .B(n5801), .ZN(n5927) );
  OAI21_X1 U6889 ( .B1(n5927), .B2(n6255), .A(n5803), .ZN(n5807) );
  NOR3_X1 U6890 ( .A1(n5817), .A2(n5805), .A3(n5804), .ZN(n5806) );
  AOI211_X1 U6891 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5814), .A(n5807), .B(n5806), .ZN(n5808) );
  OAI21_X1 U6892 ( .B1(n5809), .B2(n6262), .A(n5808), .ZN(U2998) );
  NAND2_X1 U6893 ( .A1(n5810), .A2(n6277), .ZN(n5816) );
  OAI21_X1 U6894 ( .B1(n5812), .B2(n6255), .A(n5811), .ZN(n5813) );
  AOI21_X1 U6895 ( .B1(n5814), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5813), 
        .ZN(n5815) );
  OAI211_X1 U6896 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5817), .A(n5816), .B(n5815), .ZN(U2999) );
  NOR3_X1 U6897 ( .A1(n5709), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5818), 
        .ZN(n5941) );
  AND2_X1 U6898 ( .A1(n5818), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5819)
         );
  NAND2_X1 U6899 ( .A1(n5709), .A2(n5819), .ZN(n5939) );
  INV_X1 U6900 ( .A(n5939), .ZN(n5820) );
  NOR2_X1 U6901 ( .A1(n5941), .A2(n5820), .ZN(n5821) );
  XNOR2_X1 U6902 ( .A(n5821), .B(n5952), .ZN(n5950) );
  INV_X1 U6903 ( .A(n5951), .ZN(n5826) );
  AOI22_X1 U6904 ( .A1(n5822), .A2(n6273), .B1(n6279), .B2(
        REIP_REG_17__SCAN_IN), .ZN(n5823) );
  OAI21_X1 U6905 ( .B1(n5824), .B2(n5952), .A(n5823), .ZN(n5825) );
  AOI21_X1 U6906 ( .B1(n5826), .B2(n5952), .A(n5825), .ZN(n5827) );
  OAI21_X1 U6907 ( .B1(n5950), .B2(n6262), .A(n5827), .ZN(U3001) );
  OAI211_X1 U6908 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5959), .B(n5828), .ZN(n5829) );
  OAI21_X1 U6909 ( .B1(n6254), .B2(n6540), .A(n5829), .ZN(n5833) );
  AOI21_X1 U6910 ( .B1(n5830), .B2(n6227), .A(n5970), .ZN(n5962) );
  NOR2_X1 U6911 ( .A1(n5962), .A2(n5831), .ZN(n5832) );
  AOI211_X1 U6912 ( .C1(n6273), .C2(n5834), .A(n5833), .B(n5832), .ZN(n5835)
         );
  OAI21_X1 U6913 ( .B1(n5836), .B2(n6262), .A(n5835), .ZN(U3002) );
  OAI211_X1 U6914 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3022), .A(n6383), .B(
        n6382), .ZN(n5837) );
  OAI21_X1 U6915 ( .B1(n5838), .B2(n4526), .A(n5837), .ZN(n5839) );
  MUX2_X1 U6916 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5839), .S(n6285), 
        .Z(U3464) );
  NOR3_X1 U6917 ( .A1(n5841), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5840), 
        .ZN(n5842) );
  AOI21_X1 U6918 ( .B1(n5844), .B2(n6338), .A(n5842), .ZN(n5880) );
  NOR2_X1 U6919 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5843), .ZN(n5878)
         );
  INV_X1 U6920 ( .A(n5844), .ZN(n5848) );
  INV_X1 U6921 ( .A(n5884), .ZN(n5846) );
  OAI21_X1 U6922 ( .B1(n5882), .B2(n5846), .A(n5845), .ZN(n5847) );
  NAND2_X1 U6923 ( .A1(n5848), .A2(n5847), .ZN(n5850) );
  OAI221_X1 U6924 ( .B1(n5878), .B2(n6571), .C1(n5878), .C2(n5850), .A(n5849), 
        .ZN(n5877) );
  AOI22_X1 U6925 ( .A1(n6379), .A2(n5878), .B1(INSTQUEUE_REG_2__0__SCAN_IN), 
        .B2(n5877), .ZN(n5851) );
  OAI21_X1 U6926 ( .B1(n6343), .B2(n5880), .A(n5851), .ZN(n5852) );
  AOI21_X1 U6927 ( .B1(n6340), .B2(n5882), .A(n5852), .ZN(n5853) );
  OAI21_X1 U6928 ( .B1(n5854), .B2(n5884), .A(n5853), .ZN(U3036) );
  AOI22_X1 U6929 ( .A1(n6398), .A2(n5878), .B1(INSTQUEUE_REG_2__1__SCAN_IN), 
        .B2(n5877), .ZN(n5855) );
  OAI21_X1 U6930 ( .B1(n6347), .B2(n5880), .A(n5855), .ZN(n5856) );
  AOI21_X1 U6931 ( .B1(n6399), .B2(n5882), .A(n5856), .ZN(n5857) );
  OAI21_X1 U6932 ( .B1(n6403), .B2(n5884), .A(n5857), .ZN(U3037) );
  AOI22_X1 U6933 ( .A1(n6404), .A2(n5878), .B1(INSTQUEUE_REG_2__2__SCAN_IN), 
        .B2(n5877), .ZN(n5858) );
  OAI21_X1 U6934 ( .B1(n6351), .B2(n5880), .A(n5858), .ZN(n5859) );
  AOI21_X1 U6935 ( .B1(n6405), .B2(n5882), .A(n5859), .ZN(n5860) );
  OAI21_X1 U6936 ( .B1(n6409), .B2(n5884), .A(n5860), .ZN(U3038) );
  AOI22_X1 U6937 ( .A1(n6410), .A2(n5878), .B1(INSTQUEUE_REG_2__3__SCAN_IN), 
        .B2(n5877), .ZN(n5861) );
  OAI21_X1 U6938 ( .B1(n6355), .B2(n5880), .A(n5861), .ZN(n5862) );
  AOI21_X1 U6939 ( .B1(n6352), .B2(n5882), .A(n5862), .ZN(n5863) );
  OAI21_X1 U6940 ( .B1(n5864), .B2(n5884), .A(n5863), .ZN(U3039) );
  AOI22_X1 U6941 ( .A1(n6416), .A2(n5878), .B1(INSTQUEUE_REG_2__4__SCAN_IN), 
        .B2(n5877), .ZN(n5865) );
  OAI21_X1 U6942 ( .B1(n6359), .B2(n5880), .A(n5865), .ZN(n5866) );
  AOI21_X1 U6943 ( .B1(n6356), .B2(n5882), .A(n5866), .ZN(n5867) );
  OAI21_X1 U6944 ( .B1(n5868), .B2(n5884), .A(n5867), .ZN(U3040) );
  AOI22_X1 U6945 ( .A1(n6422), .A2(n5878), .B1(INSTQUEUE_REG_2__5__SCAN_IN), 
        .B2(n5877), .ZN(n5869) );
  OAI21_X1 U6946 ( .B1(n6363), .B2(n5880), .A(n5869), .ZN(n5870) );
  AOI21_X1 U6947 ( .B1(n6360), .B2(n5882), .A(n5870), .ZN(n5871) );
  OAI21_X1 U6948 ( .B1(n5872), .B2(n5884), .A(n5871), .ZN(U3041) );
  AOI22_X1 U6949 ( .A1(n6428), .A2(n5878), .B1(INSTQUEUE_REG_2__6__SCAN_IN), 
        .B2(n5877), .ZN(n5873) );
  OAI21_X1 U6950 ( .B1(n6367), .B2(n5880), .A(n5873), .ZN(n5874) );
  AOI21_X1 U6951 ( .B1(n6364), .B2(n5882), .A(n5874), .ZN(n5875) );
  OAI21_X1 U6952 ( .B1(n5876), .B2(n5884), .A(n5875), .ZN(U3042) );
  AOI22_X1 U6953 ( .A1(n6437), .A2(n5878), .B1(INSTQUEUE_REG_2__7__SCAN_IN), 
        .B2(n5877), .ZN(n5879) );
  OAI21_X1 U6954 ( .B1(n6375), .B2(n5880), .A(n5879), .ZN(n5881) );
  AOI21_X1 U6955 ( .B1(n6438), .B2(n5882), .A(n5881), .ZN(n5883) );
  OAI21_X1 U6956 ( .B1(n6446), .B2(n5884), .A(n5883), .ZN(U3043) );
  AND2_X1 U6957 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n6132), .ZN(U2892) );
  INV_X1 U6958 ( .A(n5885), .ZN(n5886) );
  OAI22_X1 U6959 ( .A1(n5887), .A2(n6619), .B1(n6075), .B2(n5886), .ZN(n5888)
         );
  AOI21_X1 U6960 ( .B1(n6611), .B2(EBX_REG_27__SCAN_IN), .A(n5888), .ZN(n5891)
         );
  NAND2_X1 U6961 ( .A1(n5889), .A2(REIP_REG_27__SCAN_IN), .ZN(n5890) );
  OAI211_X1 U6962 ( .C1(n5892), .C2(n6624), .A(n5891), .B(n5890), .ZN(n5893)
         );
  AOI21_X1 U6963 ( .B1(n5894), .B2(n6615), .A(n5893), .ZN(n5895) );
  OAI21_X1 U6964 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5896), .A(n5895), .ZN(U2800) );
  AOI22_X1 U6965 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6611), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6054), .ZN(n5908) );
  INV_X1 U6966 ( .A(n5897), .ZN(n5900) );
  AND2_X1 U6967 ( .A1(n5899), .A2(n5898), .ZN(n5917) );
  AOI22_X1 U6968 ( .A1(n5900), .A2(n6614), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5917), .ZN(n5907) );
  AOI22_X1 U6969 ( .A1(n5902), .A2(n6615), .B1(n6058), .B2(n5901), .ZN(n5906)
         );
  INV_X1 U6970 ( .A(n5915), .ZN(n5904) );
  OAI211_X1 U6971 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5904), .B(n5903), .ZN(n5905) );
  NAND4_X1 U6972 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(U2805)
         );
  AOI22_X1 U6973 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6611), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5917), .ZN(n5909) );
  OAI21_X1 U6974 ( .B1(n5910), .B2(n6619), .A(n5909), .ZN(n5911) );
  AOI21_X1 U6975 ( .B1(n5912), .B2(n6614), .A(n5911), .ZN(n5914) );
  AOI22_X1 U6976 ( .A1(n5932), .A2(n6615), .B1(n5924), .B2(n6058), .ZN(n5913)
         );
  OAI211_X1 U6977 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5915), .A(n5914), .B(n5913), .ZN(U2806) );
  AOI22_X1 U6978 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6611), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6054), .ZN(n5923) );
  OAI22_X1 U6979 ( .A1(n5935), .A2(n6060), .B1(n5927), .B2(n6624), .ZN(n5916)
         );
  INV_X1 U6980 ( .A(n5916), .ZN(n5922) );
  OAI21_X1 U6981 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5918), .A(n5917), .ZN(n5921) );
  NAND2_X1 U6982 ( .A1(n5919), .A2(n6614), .ZN(n5920) );
  NAND4_X1 U6983 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(U2807)
         );
  INV_X1 U6984 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5926) );
  AOI22_X1 U6985 ( .A1(n5932), .A2(n6085), .B1(n5924), .B2(n6084), .ZN(n5925)
         );
  OAI21_X1 U6986 ( .B1(n5926), .B2(n6081), .A(n5925), .ZN(U2838) );
  INV_X1 U6987 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5930) );
  OAI22_X1 U6988 ( .A1(n5935), .A2(n6078), .B1(n5927), .B2(n6077), .ZN(n5928)
         );
  INV_X1 U6989 ( .A(n5928), .ZN(n5929) );
  OAI21_X1 U6990 ( .B1(n5930), .B2(n6081), .A(n5929), .ZN(U2839) );
  INV_X1 U6991 ( .A(n5931), .ZN(n6096) );
  AOI22_X1 U6992 ( .A1(n5932), .A2(n6096), .B1(n6095), .B2(DATAI_21_), .ZN(
        n5934) );
  AOI22_X1 U6993 ( .A1(n6099), .A2(DATAI_5_), .B1(n6098), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U6994 ( .A1(n5934), .A2(n5933), .ZN(U2870) );
  INV_X1 U6995 ( .A(n5935), .ZN(n5936) );
  AOI22_X1 U6996 ( .A1(n5936), .A2(n6096), .B1(n6095), .B2(DATAI_20_), .ZN(
        n5938) );
  AOI22_X1 U6997 ( .A1(n6099), .A2(DATAI_4_), .B1(n6098), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U6998 ( .A1(n5938), .A2(n5937), .ZN(U2871) );
  AOI22_X1 U6999 ( .A1(n6279), .A2(REIP_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6187), .ZN(n5944) );
  NOR2_X1 U7000 ( .A1(n5939), .A2(n5952), .ZN(n5940) );
  AOI21_X1 U7001 ( .B1(n5941), .B2(n5952), .A(n5940), .ZN(n5942) );
  XNOR2_X1 U7002 ( .A(n5942), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5954)
         );
  AOI22_X1 U7003 ( .A1(n5954), .A2(n6193), .B1(n6192), .B2(n6088), .ZN(n5943)
         );
  OAI211_X1 U7004 ( .C1(n6197), .C2(n6023), .A(n5944), .B(n5943), .ZN(U2968)
         );
  AOI22_X1 U7005 ( .A1(n6279), .A2(REIP_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6187), .ZN(n5949) );
  INV_X1 U7006 ( .A(n5945), .ZN(n6091) );
  AOI22_X1 U7007 ( .A1(n6091), .A2(n6181), .B1(n5947), .B2(n5946), .ZN(n5948)
         );
  OAI211_X1 U7008 ( .C1(n5950), .C2(n6165), .A(n5949), .B(n5948), .ZN(U2969)
         );
  NOR3_X1 U7009 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5952), .A3(n5951), 
        .ZN(n5953) );
  AOI21_X1 U7010 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6279), .A(n5953), .ZN(n5956) );
  AOI22_X1 U7011 ( .A1(n5954), .A2(n6277), .B1(n6273), .B2(n6020), .ZN(n5955)
         );
  OAI211_X1 U7012 ( .C1(n5958), .C2(n5957), .A(n5956), .B(n5955), .ZN(U3000)
         );
  INV_X1 U7013 ( .A(n5959), .ZN(n5967) );
  AOI21_X1 U7014 ( .B1(n5961), .B2(n6273), .A(n5960), .ZN(n5966) );
  INV_X1 U7015 ( .A(n5962), .ZN(n5963) );
  AOI22_X1 U7016 ( .A1(n5964), .A2(n6277), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5963), .ZN(n5965) );
  OAI211_X1 U7017 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n5967), .A(n5966), .B(n5965), .ZN(U3003) );
  NOR3_X1 U7018 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5968), .A3(n5971), 
        .ZN(n5986) );
  NOR3_X1 U7019 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5969), .A3(n5971), 
        .ZN(n5985) );
  AOI21_X1 U7020 ( .B1(n5972), .B2(n5971), .A(n5970), .ZN(n5973) );
  OAI21_X1 U7021 ( .B1(n5975), .B2(n5974), .A(n5973), .ZN(n5987) );
  AOI211_X1 U7022 ( .C1(n5976), .C2(n5986), .A(n5985), .B(n5987), .ZN(n5979)
         );
  AOI222_X1 U7023 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6279), .B1(n6273), .B2(
        n6621), .C1(n6277), .C2(n5977), .ZN(n5978) );
  OAI221_X1 U7024 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5981), .C1(
        n5980), .C2(n5979), .A(n5978), .ZN(U3004) );
  INV_X1 U7025 ( .A(n5982), .ZN(n5984) );
  AOI21_X1 U7026 ( .B1(n5984), .B2(n6273), .A(n5983), .ZN(n5991) );
  AOI21_X1 U7027 ( .B1(n5986), .B2(n6280), .A(n5985), .ZN(n5990) );
  AOI22_X1 U7028 ( .A1(n5988), .A2(n6277), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5987), .ZN(n5989) );
  NAND3_X1 U7029 ( .A1(n5991), .A2(n5990), .A3(n5989), .ZN(U3005) );
  INV_X1 U7030 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6515) );
  AOI21_X1 U7031 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6515), .A(n6509), .ZN(n5999) );
  INV_X1 U7032 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7033 ( .A1(n6509), .A2(STATE_REG_1__SCAN_IN), .ZN(n6550) );
  INV_X1 U7034 ( .A(n6550), .ZN(n6553) );
  AOI21_X1 U7035 ( .B1(n5999), .B2(n5992), .A(n6553), .ZN(U2789) );
  INV_X1 U7036 ( .A(n5993), .ZN(n5995) );
  OAI21_X1 U7037 ( .B1(n5995), .B2(n5994), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5996) );
  OAI21_X1 U7038 ( .B1(n5997), .B2(n6596), .A(n5996), .ZN(U2790) );
  INV_X1 U7039 ( .A(n6553), .ZN(n6606) );
  NOR2_X1 U7040 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6000) );
  OAI21_X1 U7041 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6000), .A(n6606), .ZN(n5998)
         );
  OAI21_X1 U7042 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6606), .A(n5998), .ZN(
        U2791) );
  NOR2_X1 U7043 ( .A1(n6553), .A2(n5999), .ZN(n6498) );
  OAI21_X1 U7044 ( .B1(BS16_N), .B2(n6000), .A(n6498), .ZN(n6565) );
  OAI21_X1 U7045 ( .B1(n6498), .B2(n6593), .A(n6565), .ZN(U2792) );
  OAI21_X1 U7046 ( .B1(n6002), .B2(n6001), .A(n6165), .ZN(U2793) );
  NOR4_X1 U7047 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n6006) );
  NOR4_X1 U7048 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6005) );
  NOR4_X1 U7049 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6004) );
  NOR4_X1 U7050 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6003) );
  NAND4_X1 U7051 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n6012)
         );
  NOR4_X1 U7052 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6010) );
  AOI211_X1 U7053 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_27__SCAN_IN), .B(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6009) );
  NOR4_X1 U7054 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6008)
         );
  NOR4_X1 U7055 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6007) );
  NAND4_X1 U7056 ( .A1(n6010), .A2(n6009), .A3(n6008), .A4(n6007), .ZN(n6011)
         );
  NOR2_X1 U7057 ( .A1(n6012), .A2(n6011), .ZN(n6588) );
  INV_X1 U7058 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6658) );
  NOR3_X1 U7059 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6014) );
  OAI21_X1 U7060 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6014), .A(n6588), .ZN(n6013)
         );
  OAI21_X1 U7061 ( .B1(n6588), .B2(n6658), .A(n6013), .ZN(U2794) );
  INV_X1 U7062 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6786) );
  NOR2_X1 U7063 ( .A1(REIP_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n6582) );
  OAI21_X1 U7064 ( .B1(n6014), .B2(n6582), .A(n6588), .ZN(n6015) );
  OAI21_X1 U7065 ( .B1(n6588), .B2(n6786), .A(n6015), .ZN(U2795) );
  AOI22_X1 U7066 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6611), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6016), .ZN(n6017) );
  OAI21_X1 U7067 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6018), .A(n6017), .ZN(n6019) );
  AOI211_X1 U7068 ( .C1(n6054), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6610), 
        .B(n6019), .ZN(n6022) );
  AOI22_X1 U7069 ( .A1(n6088), .A2(n6615), .B1(n6020), .B2(n6058), .ZN(n6021)
         );
  OAI211_X1 U7070 ( .C1(n6023), .C2(n6075), .A(n6022), .B(n6021), .ZN(U2809)
         );
  AND3_X1 U7071 ( .A1(n6025), .A2(n6024), .A3(n6534), .ZN(n6026) );
  AOI21_X1 U7072 ( .B1(n6027), .B2(n6058), .A(n6026), .ZN(n6034) );
  AOI22_X1 U7073 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6054), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6028), .ZN(n6033) );
  AOI21_X1 U7074 ( .B1(n6611), .B2(EBX_REG_12__SCAN_IN), .A(n6610), .ZN(n6032)
         );
  AOI22_X1 U7075 ( .A1(n6030), .A2(n6615), .B1(n6614), .B2(n6029), .ZN(n6031)
         );
  NAND4_X1 U7076 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(U2815)
         );
  OAI22_X1 U7077 ( .A1(n6037), .A2(n6624), .B1(n6036), .B2(n6035), .ZN(n6038)
         );
  INV_X1 U7078 ( .A(n6038), .ZN(n6048) );
  NOR3_X1 U7079 ( .A1(n6608), .A2(REIP_REG_10__SCAN_IN), .A3(n6039), .ZN(n6040) );
  AOI211_X1 U7080 ( .C1(n6054), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6610), 
        .B(n6040), .ZN(n6047) );
  AOI22_X1 U7081 ( .A1(n6042), .A2(n6615), .B1(n6614), .B2(n6041), .ZN(n6046)
         );
  OAI21_X1 U7082 ( .B1(n6044), .B2(n6043), .A(REIP_REG_10__SCAN_IN), .ZN(n6045) );
  NAND4_X1 U7083 ( .A1(n6048), .A2(n6047), .A3(n6046), .A4(n6045), .ZN(U2817)
         );
  AOI21_X1 U7084 ( .B1(n6049), .B2(n6525), .A(n6071), .ZN(n6063) );
  NAND2_X1 U7085 ( .A1(n6051), .A2(n6050), .ZN(n6052) );
  NAND2_X1 U7086 ( .A1(n6053), .A2(n6052), .ZN(n6076) );
  INV_X1 U7087 ( .A(n6076), .ZN(n6213) );
  NAND2_X1 U7088 ( .A1(n6611), .A2(EBX_REG_7__SCAN_IN), .ZN(n6056) );
  AOI21_X1 U7089 ( .B1(n6054), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6610), 
        .ZN(n6055) );
  OAI211_X1 U7090 ( .C1(n6075), .C2(n6169), .A(n6056), .B(n6055), .ZN(n6057)
         );
  AOI21_X1 U7091 ( .B1(n6213), .B2(n6058), .A(n6057), .ZN(n6059) );
  OAI21_X1 U7092 ( .B1(n6164), .B2(n6060), .A(n6059), .ZN(n6061) );
  INV_X1 U7093 ( .A(n6061), .ZN(n6062) );
  OAI221_X1 U7094 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6064), .C1(n6527), .C2(
        n6063), .A(n6062), .ZN(U2820) );
  INV_X1 U7095 ( .A(n6065), .ZN(n6070) );
  INV_X1 U7096 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6780) );
  OAI21_X1 U7097 ( .B1(n6619), .B2(n6780), .A(n6066), .ZN(n6067) );
  AOI21_X1 U7098 ( .B1(n6611), .B2(EBX_REG_5__SCAN_IN), .A(n6067), .ZN(n6068)
         );
  OAI21_X1 U7099 ( .B1(n6624), .B2(n6239), .A(n6068), .ZN(n6069) );
  AOI21_X1 U7100 ( .B1(n6173), .B2(n6070), .A(n6069), .ZN(n6074) );
  OAI21_X1 U7101 ( .B1(REIP_REG_5__SCAN_IN), .B2(n6072), .A(n6071), .ZN(n6073)
         );
  OAI211_X1 U7102 ( .C1(n6075), .C2(n6176), .A(n6074), .B(n6073), .ZN(U2822)
         );
  INV_X1 U7103 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6082) );
  OAI22_X1 U7104 ( .A1(n6164), .A2(n6078), .B1(n6077), .B2(n6076), .ZN(n6079)
         );
  INV_X1 U7105 ( .A(n6079), .ZN(n6080) );
  OAI21_X1 U7106 ( .B1(n6082), .B2(n6081), .A(n6080), .ZN(U2852) );
  INV_X1 U7107 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6087) );
  INV_X1 U7108 ( .A(n6083), .ZN(n6182) );
  AOI22_X1 U7109 ( .A1(n6182), .A2(n6085), .B1(n6084), .B2(n6261), .ZN(n6086)
         );
  OAI21_X1 U7110 ( .B1(n6087), .B2(n6081), .A(n6086), .ZN(U2856) );
  AOI22_X1 U7111 ( .A1(n6088), .A2(n6096), .B1(n6095), .B2(DATAI_18_), .ZN(
        n6090) );
  AOI22_X1 U7112 ( .A1(n6099), .A2(DATAI_2_), .B1(n6098), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7113 ( .A1(n6090), .A2(n6089), .ZN(U2873) );
  AOI22_X1 U7114 ( .A1(n6091), .A2(n6096), .B1(n6095), .B2(DATAI_17_), .ZN(
        n6093) );
  AOI22_X1 U7115 ( .A1(n6099), .A2(DATAI_1_), .B1(n6098), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7116 ( .A1(n6093), .A2(n6092), .ZN(U2874) );
  INV_X1 U7117 ( .A(n6094), .ZN(n6097) );
  AOI22_X1 U7118 ( .A1(n6097), .A2(n6096), .B1(n6095), .B2(DATAI_16_), .ZN(
        n6101) );
  AOI22_X1 U7119 ( .A1(n6099), .A2(DATAI_0_), .B1(n6098), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7120 ( .A1(n6101), .A2(n6100), .ZN(U2875) );
  INV_X1 U7121 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6764) );
  INV_X1 U7122 ( .A(n6102), .ZN(n6107) );
  AOI22_X1 U7123 ( .A1(n6132), .A2(DATAO_REG_29__SCAN_IN), .B1(n6107), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6103) );
  OAI21_X1 U7124 ( .B1(n6764), .B2(n6106), .A(n6103), .ZN(U2894) );
  INV_X1 U7125 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U7126 ( .A1(n6132), .A2(DATAO_REG_27__SCAN_IN), .B1(n6107), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6104) );
  OAI21_X1 U7127 ( .B1(n6655), .B2(n6106), .A(n6104), .ZN(U2896) );
  AOI22_X1 U7128 ( .A1(n6132), .A2(DATAO_REG_21__SCAN_IN), .B1(n6107), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6105) );
  OAI21_X1 U7129 ( .B1(n4328), .B2(n6106), .A(n6105), .ZN(U2902) );
  INV_X1 U7130 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n6807) );
  AOI22_X1 U7131 ( .A1(n6107), .A2(EAX_REG_16__SCAN_IN), .B1(
        UWORD_REG_0__SCAN_IN), .B2(n4374), .ZN(n6108) );
  OAI21_X1 U7132 ( .B1(n6807), .B2(n6118), .A(n6108), .ZN(U2907) );
  INV_X1 U7133 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6160) );
  AOI22_X1 U7134 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U7135 ( .B1(n6160), .B2(n6135), .A(n6109), .ZN(U2908) );
  INV_X1 U7136 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6111) );
  AOI22_X1 U7137 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6110) );
  OAI21_X1 U7138 ( .B1(n6111), .B2(n6135), .A(n6110), .ZN(U2909) );
  INV_X1 U7139 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6113) );
  AOI22_X1 U7140 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7141 ( .B1(n6113), .B2(n6135), .A(n6112), .ZN(U2910) );
  INV_X1 U7142 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6115) );
  AOI22_X1 U7143 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6114) );
  OAI21_X1 U7144 ( .B1(n6115), .B2(n6135), .A(n6114), .ZN(U2911) );
  INV_X1 U7145 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6757) );
  AOI22_X1 U7146 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6116), .B1(
        LWORD_REG_11__SCAN_IN), .B2(n4374), .ZN(n6117) );
  OAI21_X1 U7147 ( .B1(n6757), .B2(n6118), .A(n6117), .ZN(U2912) );
  AOI22_X1 U7148 ( .A1(DATAO_REG_10__SCAN_IN), .A2(n6132), .B1(
        LWORD_REG_10__SCAN_IN), .B2(n4374), .ZN(n6119) );
  OAI21_X1 U7149 ( .B1(n4313), .B2(n6135), .A(n6119), .ZN(U2913) );
  AOI22_X1 U7150 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6120) );
  OAI21_X1 U7151 ( .B1(n4396), .B2(n6135), .A(n6120), .ZN(U2914) );
  INV_X1 U7152 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6122) );
  AOI22_X1 U7153 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6121) );
  OAI21_X1 U7154 ( .B1(n6122), .B2(n6135), .A(n6121), .ZN(U2915) );
  AOI22_X1 U7155 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7156 ( .B1(n6124), .B2(n6135), .A(n6123), .ZN(U2916) );
  AOI22_X1 U7157 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6125) );
  OAI21_X1 U7158 ( .B1(n4412), .B2(n6135), .A(n6125), .ZN(U2917) );
  AOI22_X1 U7159 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6126) );
  OAI21_X1 U7160 ( .B1(n3533), .B2(n6135), .A(n6126), .ZN(U2918) );
  AOI22_X1 U7161 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6127) );
  OAI21_X1 U7162 ( .B1(n4393), .B2(n6135), .A(n6127), .ZN(U2919) );
  AOI22_X1 U7163 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6128) );
  OAI21_X1 U7164 ( .B1(n6129), .B2(n6135), .A(n6128), .ZN(U2920) );
  AOI22_X1 U7165 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6130) );
  OAI21_X1 U7166 ( .B1(n4315), .B2(n6135), .A(n6130), .ZN(U2921) );
  AOI22_X1 U7167 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6131) );
  OAI21_X1 U7168 ( .B1(n4404), .B2(n6135), .A(n6131), .ZN(U2922) );
  AOI22_X1 U7169 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n4374), .B1(n6132), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6134) );
  OAI21_X1 U7170 ( .B1(n6136), .B2(n6135), .A(n6134), .ZN(U2923) );
  AOI22_X1 U7171 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6153), .B1(n6156), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7172 ( .A1(n6157), .A2(DATAI_8_), .ZN(n6145) );
  NAND2_X1 U7173 ( .A1(n6137), .A2(n6145), .ZN(U2932) );
  NAND2_X1 U7174 ( .A1(n6157), .A2(DATAI_11_), .ZN(n6147) );
  INV_X1 U7175 ( .A(n6147), .ZN(n6138) );
  AOI21_X1 U7176 ( .B1(n6153), .B2(EAX_REG_27__SCAN_IN), .A(n6138), .ZN(n6139)
         );
  OAI21_X1 U7177 ( .B1(n6655), .B2(n6143), .A(n6139), .ZN(U2935) );
  AOI22_X1 U7178 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6153), .B1(n6156), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7179 ( .A1(n6157), .A2(DATAI_12_), .ZN(n6149) );
  NAND2_X1 U7180 ( .A1(n6140), .A2(n6149), .ZN(U2936) );
  NAND2_X1 U7181 ( .A1(n6157), .A2(DATAI_13_), .ZN(n6151) );
  INV_X1 U7182 ( .A(n6151), .ZN(n6141) );
  AOI21_X1 U7183 ( .B1(n6153), .B2(EAX_REG_29__SCAN_IN), .A(n6141), .ZN(n6142)
         );
  OAI21_X1 U7184 ( .B1(n6764), .B2(n6143), .A(n6142), .ZN(U2937) );
  AOI22_X1 U7185 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6153), .B1(n6156), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7186 ( .A1(n6157), .A2(DATAI_14_), .ZN(n6154) );
  NAND2_X1 U7187 ( .A1(n6144), .A2(n6154), .ZN(U2938) );
  AOI22_X1 U7188 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6153), .B1(n6156), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7189 ( .A1(n6146), .A2(n6145), .ZN(U2947) );
  AOI22_X1 U7190 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6153), .B1(n6156), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7191 ( .A1(n6148), .A2(n6147), .ZN(U2950) );
  AOI22_X1 U7192 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6153), .B1(n6156), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7193 ( .A1(n6150), .A2(n6149), .ZN(U2951) );
  AOI22_X1 U7194 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6153), .B1(n6156), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7195 ( .A1(n6152), .A2(n6151), .ZN(U2952) );
  AOI22_X1 U7196 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6153), .B1(
        LWORD_REG_14__SCAN_IN), .B2(n6156), .ZN(n6155) );
  NAND2_X1 U7197 ( .A1(n6155), .A2(n6154), .ZN(U2953) );
  AOI22_X1 U7198 ( .A1(n6157), .A2(DATAI_15_), .B1(n6156), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6158) );
  OAI21_X1 U7199 ( .B1(n6160), .B2(n6159), .A(n6158), .ZN(U2954) );
  AOI22_X1 U7200 ( .A1(n6279), .A2(REIP_REG_7__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n6187), .ZN(n6168) );
  OAI21_X1 U7201 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(n6216) );
  OAI22_X1 U7202 ( .A1(n6216), .A2(n6165), .B1(n5352), .B2(n6164), .ZN(n6166)
         );
  INV_X1 U7203 ( .A(n6166), .ZN(n6167) );
  OAI211_X1 U7204 ( .C1(n6197), .C2(n6169), .A(n6168), .B(n6167), .ZN(U2979)
         );
  AOI22_X1 U7205 ( .A1(n6279), .A2(REIP_REG_5__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n6187), .ZN(n6175) );
  NAND2_X1 U7206 ( .A1(n6170), .A2(n6171), .ZN(n6172) );
  NAND2_X1 U7207 ( .A1(n4134), .A2(n6172), .ZN(n6244) );
  AOI22_X1 U7208 ( .A1(n6244), .A2(n6193), .B1(n6173), .B2(n6181), .ZN(n6174)
         );
  OAI211_X1 U7209 ( .C1(n6197), .C2(n6176), .A(n6175), .B(n6174), .ZN(U2981)
         );
  AOI22_X1 U7210 ( .A1(n6279), .A2(REIP_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6187), .ZN(n6185) );
  OR2_X1 U7211 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  NAND2_X1 U7212 ( .A1(n6180), .A2(n6179), .ZN(n6263) );
  INV_X1 U7213 ( .A(n6263), .ZN(n6183) );
  AOI22_X1 U7214 ( .A1(n6183), .A2(n6193), .B1(n6182), .B2(n6181), .ZN(n6184)
         );
  OAI211_X1 U7215 ( .C1(n6197), .C2(n6186), .A(n6185), .B(n6184), .ZN(U2983)
         );
  AOI22_X1 U7216 ( .A1(n6279), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6187), .ZN(n6195) );
  XOR2_X1 U7217 ( .A(n6188), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6190) );
  XNOR2_X1 U7218 ( .A(n6190), .B(n6189), .ZN(n6278) );
  AOI22_X1 U7219 ( .A1(n6278), .A2(n6193), .B1(n6192), .B2(n6191), .ZN(n6194)
         );
  OAI211_X1 U7220 ( .C1(n6197), .C2(n6196), .A(n6195), .B(n6194), .ZN(U2984)
         );
  AOI21_X1 U7221 ( .B1(n6199), .B2(n6273), .A(n6198), .ZN(n6203) );
  AOI22_X1 U7222 ( .A1(n6201), .A2(n6277), .B1(n6200), .B2(n6792), .ZN(n6202)
         );
  OAI211_X1 U7223 ( .C1(n6204), .C2(n6792), .A(n6203), .B(n6202), .ZN(U3007)
         );
  INV_X1 U7224 ( .A(n6205), .ZN(n6207) );
  AOI21_X1 U7225 ( .B1(n6207), .B2(n6273), .A(n6206), .ZN(n6211) );
  AOI22_X1 U7226 ( .A1(n6209), .A2(n6277), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6208), .ZN(n6210) );
  OAI211_X1 U7227 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6212), .A(n6211), 
        .B(n6210), .ZN(U3009) );
  AOI22_X1 U7228 ( .A1(n6213), .A2(n6273), .B1(n6279), .B2(REIP_REG_7__SCAN_IN), .ZN(n6219) );
  INV_X1 U7229 ( .A(n6214), .ZN(n6215) );
  OAI22_X1 U7230 ( .A1(n6216), .A2(n6262), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6215), .ZN(n6217) );
  INV_X1 U7231 ( .A(n6217), .ZN(n6218) );
  OAI211_X1 U7232 ( .C1(n6221), .C2(n6220), .A(n6219), .B(n6218), .ZN(U3011)
         );
  NAND2_X1 U7233 ( .A1(n6250), .A2(n6222), .ZN(n6226) );
  NAND2_X1 U7234 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7235 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  NAND2_X1 U7236 ( .A1(n6226), .A2(n6225), .ZN(n6276) );
  AOI221_X1 U7237 ( .B1(n6231), .B2(n6227), .C1(n6230), .C2(n6227), .A(n6276), 
        .ZN(n6248) );
  AOI21_X1 U7238 ( .B1(n6229), .B2(n6273), .A(n6228), .ZN(n6236) );
  NOR3_X1 U7239 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6231), .A3(n6230), 
        .ZN(n6233) );
  AOI22_X1 U7240 ( .A1(n6234), .A2(n6277), .B1(n6233), .B2(n6232), .ZN(n6235)
         );
  OAI211_X1 U7241 ( .C1(n6248), .C2(n6237), .A(n6236), .B(n6235), .ZN(U3012)
         );
  NOR2_X1 U7242 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6238), .ZN(n6247)
         );
  INV_X1 U7243 ( .A(n6239), .ZN(n6240) );
  AOI22_X1 U7244 ( .A1(n6240), .A2(n6273), .B1(n6279), .B2(REIP_REG_5__SCAN_IN), .ZN(n6246) );
  NOR3_X1 U7245 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6242), .A3(n6241), 
        .ZN(n6243) );
  AOI21_X1 U7246 ( .B1(n6244), .B2(n6277), .A(n6243), .ZN(n6245) );
  OAI211_X1 U7247 ( .C1(n6248), .C2(n6247), .A(n6246), .B(n6245), .ZN(U3013)
         );
  INV_X1 U7248 ( .A(n6276), .ZN(n6249) );
  OAI21_X1 U7249 ( .B1(n6250), .B2(n6270), .A(n6249), .ZN(n6251) );
  INV_X1 U7250 ( .A(n6251), .ZN(n6269) );
  AOI211_X1 U7251 ( .C1(n6800), .C2(n6268), .A(n6252), .B(n6264), .ZN(n6259)
         );
  NOR2_X1 U7252 ( .A1(n6253), .A2(n6262), .ZN(n6258) );
  OAI22_X1 U7253 ( .A1(n6256), .A2(n6255), .B1(n6520), .B2(n6254), .ZN(n6257)
         );
  NOR3_X1 U7254 ( .A1(n6259), .A2(n6258), .A3(n6257), .ZN(n6260) );
  OAI21_X1 U7255 ( .B1(n6269), .B2(n6800), .A(n6260), .ZN(U3014) );
  AOI22_X1 U7256 ( .A1(n6273), .A2(n6261), .B1(n6279), .B2(REIP_REG_3__SCAN_IN), .ZN(n6267) );
  OAI22_X1 U7257 ( .A1(n6264), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6263), 
        .B2(n6262), .ZN(n6265) );
  INV_X1 U7258 ( .A(n6265), .ZN(n6266) );
  OAI211_X1 U7259 ( .C1(n6269), .C2(n6268), .A(n6267), .B(n6266), .ZN(U3015)
         );
  OAI21_X1 U7260 ( .B1(n6271), .B2(n4102), .A(n6270), .ZN(n6274) );
  AOI22_X1 U7261 ( .A1(n6275), .A2(n6274), .B1(n6273), .B2(n6272), .ZN(n6284)
         );
  AOI22_X1 U7262 ( .A1(n6278), .A2(n6277), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6276), .ZN(n6283) );
  NAND2_X1 U7263 ( .A1(n6279), .A2(REIP_REG_2__SCAN_IN), .ZN(n6282) );
  NAND3_X1 U7264 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4102), .A3(n6280), 
        .ZN(n6281) );
  NAND4_X1 U7265 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(U3016)
         );
  INV_X1 U7266 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6286) );
  NOR2_X1 U7267 ( .A1(n6286), .A2(n6285), .ZN(U3019) );
  NAND3_X1 U7268 ( .A1(n6290), .A2(n6289), .A3(n6377), .ZN(n6291) );
  OAI21_X1 U7269 ( .B1(n6292), .B2(n6295), .A(n6291), .ZN(n6321) );
  AND2_X1 U7270 ( .A1(n6447), .A2(n6339), .ZN(n6320) );
  AOI22_X1 U7271 ( .A1(n6394), .A2(n6321), .B1(n6379), .B2(n6320), .ZN(n6305)
         );
  NOR3_X1 U7272 ( .A1(n6322), .A2(n6370), .A3(n6388), .ZN(n6297) );
  OR2_X1 U7273 ( .A1(n6295), .A2(n6294), .ZN(n6330) );
  OAI21_X1 U7274 ( .B1(n6297), .B2(n6296), .A(n6330), .ZN(n6303) );
  INV_X1 U7275 ( .A(n6298), .ZN(n6302) );
  INV_X1 U7276 ( .A(n6320), .ZN(n6300) );
  AOI211_X1 U7277 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6300), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6299), .ZN(n6301) );
  NAND3_X1 U7278 ( .A1(n6303), .A2(n6302), .A3(n6301), .ZN(n6323) );
  AOI22_X1 U7279 ( .A1(n6323), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6380), 
        .B2(n6322), .ZN(n6304) );
  OAI211_X1 U7280 ( .C1(n6397), .C2(n6326), .A(n6305), .B(n6304), .ZN(U3068)
         );
  AOI22_X1 U7281 ( .A1(n6400), .A2(n6321), .B1(n6398), .B2(n6320), .ZN(n6307)
         );
  AOI22_X1 U7282 ( .A1(n6323), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6344), 
        .B2(n6322), .ZN(n6306) );
  OAI211_X1 U7283 ( .C1(n6308), .C2(n6326), .A(n6307), .B(n6306), .ZN(U3069)
         );
  AOI22_X1 U7284 ( .A1(n6406), .A2(n6321), .B1(n6404), .B2(n6320), .ZN(n6310)
         );
  AOI22_X1 U7285 ( .A1(n6323), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6348), 
        .B2(n6322), .ZN(n6309) );
  OAI211_X1 U7286 ( .C1(n6311), .C2(n6326), .A(n6310), .B(n6309), .ZN(U3070)
         );
  AOI22_X1 U7287 ( .A1(n6412), .A2(n6321), .B1(n6410), .B2(n6320), .ZN(n6313)
         );
  AOI22_X1 U7288 ( .A1(n6323), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6411), 
        .B2(n6322), .ZN(n6312) );
  OAI211_X1 U7289 ( .C1(n6415), .C2(n6326), .A(n6313), .B(n6312), .ZN(U3071)
         );
  AOI22_X1 U7290 ( .A1(n6418), .A2(n6321), .B1(n6416), .B2(n6320), .ZN(n6315)
         );
  AOI22_X1 U7291 ( .A1(n6323), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6417), 
        .B2(n6322), .ZN(n6314) );
  OAI211_X1 U7292 ( .C1(n6421), .C2(n6326), .A(n6315), .B(n6314), .ZN(U3072)
         );
  AOI22_X1 U7293 ( .A1(n6424), .A2(n6321), .B1(n6422), .B2(n6320), .ZN(n6317)
         );
  AOI22_X1 U7294 ( .A1(n6323), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6423), 
        .B2(n6322), .ZN(n6316) );
  OAI211_X1 U7295 ( .C1(n6427), .C2(n6326), .A(n6317), .B(n6316), .ZN(U3073)
         );
  AOI22_X1 U7296 ( .A1(n6431), .A2(n6321), .B1(n6428), .B2(n6320), .ZN(n6319)
         );
  AOI22_X1 U7297 ( .A1(n6323), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6429), 
        .B2(n6322), .ZN(n6318) );
  OAI211_X1 U7298 ( .C1(n6435), .C2(n6326), .A(n6319), .B(n6318), .ZN(U3074)
         );
  AOI22_X1 U7299 ( .A1(n6441), .A2(n6321), .B1(n6437), .B2(n6320), .ZN(n6325)
         );
  AOI22_X1 U7300 ( .A1(n6323), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6371), 
        .B2(n6322), .ZN(n6324) );
  OAI211_X1 U7301 ( .C1(n6327), .C2(n6326), .A(n6325), .B(n6324), .ZN(U3075)
         );
  NOR2_X1 U7302 ( .A1(n6328), .A2(n6388), .ZN(n6335) );
  OR2_X1 U7303 ( .A1(n6330), .A2(n6329), .ZN(n6331) );
  AND2_X1 U7304 ( .A1(n6331), .A2(n6333), .ZN(n6334) );
  INV_X1 U7305 ( .A(n6334), .ZN(n6332) );
  AOI22_X1 U7306 ( .A1(n6335), .A2(n6332), .B1(n6339), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n6376) );
  INV_X1 U7307 ( .A(n6333), .ZN(n6369) );
  AOI22_X1 U7308 ( .A1(n6379), .A2(n6369), .B1(n6370), .B2(n6380), .ZN(n6342)
         );
  NAND2_X1 U7309 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  OAI211_X1 U7310 ( .C1(n6339), .C2(n6338), .A(n6337), .B(n6336), .ZN(n6372)
         );
  AOI22_X1 U7311 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6372), .B1(n6340), 
        .B2(n6368), .ZN(n6341) );
  OAI211_X1 U7312 ( .C1(n6376), .C2(n6343), .A(n6342), .B(n6341), .ZN(U3076)
         );
  AOI22_X1 U7313 ( .A1(n6398), .A2(n6369), .B1(n6370), .B2(n6344), .ZN(n6346)
         );
  AOI22_X1 U7314 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6372), .B1(n6399), 
        .B2(n6368), .ZN(n6345) );
  OAI211_X1 U7315 ( .C1(n6376), .C2(n6347), .A(n6346), .B(n6345), .ZN(U3077)
         );
  AOI22_X1 U7316 ( .A1(n6404), .A2(n6369), .B1(n6370), .B2(n6348), .ZN(n6350)
         );
  AOI22_X1 U7317 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6372), .B1(n6405), 
        .B2(n6368), .ZN(n6349) );
  OAI211_X1 U7318 ( .C1(n6376), .C2(n6351), .A(n6350), .B(n6349), .ZN(U3078)
         );
  AOI22_X1 U7319 ( .A1(n6410), .A2(n6369), .B1(n6368), .B2(n6352), .ZN(n6354)
         );
  AOI22_X1 U7320 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6372), .B1(n6411), 
        .B2(n6370), .ZN(n6353) );
  OAI211_X1 U7321 ( .C1(n6376), .C2(n6355), .A(n6354), .B(n6353), .ZN(U3079)
         );
  AOI22_X1 U7322 ( .A1(n6416), .A2(n6369), .B1(n6368), .B2(n6356), .ZN(n6358)
         );
  AOI22_X1 U7323 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6372), .B1(n6417), 
        .B2(n6370), .ZN(n6357) );
  OAI211_X1 U7324 ( .C1(n6376), .C2(n6359), .A(n6358), .B(n6357), .ZN(U3080)
         );
  AOI22_X1 U7325 ( .A1(n6422), .A2(n6369), .B1(n6368), .B2(n6360), .ZN(n6362)
         );
  AOI22_X1 U7326 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6372), .B1(n6423), 
        .B2(n6370), .ZN(n6361) );
  OAI211_X1 U7327 ( .C1(n6376), .C2(n6363), .A(n6362), .B(n6361), .ZN(U3081)
         );
  AOI22_X1 U7328 ( .A1(n6428), .A2(n6369), .B1(n6370), .B2(n6429), .ZN(n6366)
         );
  AOI22_X1 U7329 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6372), .B1(n6364), 
        .B2(n6368), .ZN(n6365) );
  OAI211_X1 U7330 ( .C1(n6376), .C2(n6367), .A(n6366), .B(n6365), .ZN(U3082)
         );
  AOI22_X1 U7331 ( .A1(n6437), .A2(n6369), .B1(n6368), .B2(n6438), .ZN(n6374)
         );
  AOI22_X1 U7332 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6372), .B1(n6371), 
        .B2(n6370), .ZN(n6373) );
  OAI211_X1 U7333 ( .C1(n6376), .C2(n6375), .A(n6374), .B(n6373), .ZN(U3083)
         );
  NOR2_X1 U7334 ( .A1(n6378), .A2(n6377), .ZN(n6436) );
  AOI22_X1 U7335 ( .A1(n6430), .A2(n6380), .B1(n6379), .B2(n6436), .ZN(n6396)
         );
  INV_X1 U7336 ( .A(n6381), .ZN(n6384) );
  OAI21_X1 U7337 ( .B1(n6384), .B2(n6383), .A(n6382), .ZN(n6393) );
  AOI21_X1 U7338 ( .B1(n6386), .B2(n6385), .A(n6436), .ZN(n6392) );
  INV_X1 U7339 ( .A(n6392), .ZN(n6390) );
  AOI21_X1 U7340 ( .B1(n6388), .B2(n6391), .A(n6387), .ZN(n6389) );
  OAI21_X1 U7341 ( .B1(n6393), .B2(n6390), .A(n6389), .ZN(n6442) );
  OAI22_X1 U7342 ( .A1(n6393), .A2(n6392), .B1(n6391), .B2(n6475), .ZN(n6440)
         );
  AOI22_X1 U7343 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6442), .B1(n6394), 
        .B2(n6440), .ZN(n6395) );
  OAI211_X1 U7344 ( .C1(n6397), .C2(n6434), .A(n6396), .B(n6395), .ZN(U3108)
         );
  INV_X1 U7345 ( .A(n6434), .ZN(n6439) );
  AOI22_X1 U7346 ( .A1(n6439), .A2(n6399), .B1(n6398), .B2(n6436), .ZN(n6402)
         );
  AOI22_X1 U7347 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6442), .B1(n6400), 
        .B2(n6440), .ZN(n6401) );
  OAI211_X1 U7348 ( .C1(n6403), .C2(n6445), .A(n6402), .B(n6401), .ZN(U3109)
         );
  AOI22_X1 U7349 ( .A1(n6439), .A2(n6405), .B1(n6404), .B2(n6436), .ZN(n6408)
         );
  AOI22_X1 U7350 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6442), .B1(n6406), 
        .B2(n6440), .ZN(n6407) );
  OAI211_X1 U7351 ( .C1(n6409), .C2(n6445), .A(n6408), .B(n6407), .ZN(U3110)
         );
  AOI22_X1 U7352 ( .A1(n6430), .A2(n6411), .B1(n6410), .B2(n6436), .ZN(n6414)
         );
  AOI22_X1 U7353 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6442), .B1(n6412), 
        .B2(n6440), .ZN(n6413) );
  OAI211_X1 U7354 ( .C1(n6415), .C2(n6434), .A(n6414), .B(n6413), .ZN(U3111)
         );
  AOI22_X1 U7355 ( .A1(n6430), .A2(n6417), .B1(n6416), .B2(n6436), .ZN(n6420)
         );
  AOI22_X1 U7356 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6442), .B1(n6418), 
        .B2(n6440), .ZN(n6419) );
  OAI211_X1 U7357 ( .C1(n6421), .C2(n6434), .A(n6420), .B(n6419), .ZN(U3112)
         );
  AOI22_X1 U7358 ( .A1(n6430), .A2(n6423), .B1(n6422), .B2(n6436), .ZN(n6426)
         );
  AOI22_X1 U7359 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6442), .B1(n6424), 
        .B2(n6440), .ZN(n6425) );
  OAI211_X1 U7360 ( .C1(n6427), .C2(n6434), .A(n6426), .B(n6425), .ZN(U3113)
         );
  AOI22_X1 U7361 ( .A1(n6430), .A2(n6429), .B1(n6428), .B2(n6436), .ZN(n6433)
         );
  AOI22_X1 U7362 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6442), .B1(n6431), 
        .B2(n6440), .ZN(n6432) );
  OAI211_X1 U7363 ( .C1(n6435), .C2(n6434), .A(n6433), .B(n6432), .ZN(U3114)
         );
  AOI22_X1 U7364 ( .A1(n6439), .A2(n6438), .B1(n6437), .B2(n6436), .ZN(n6444)
         );
  AOI22_X1 U7365 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6442), .B1(n6441), 
        .B2(n6440), .ZN(n6443) );
  OAI211_X1 U7366 ( .C1(n6446), .C2(n6445), .A(n6444), .B(n6443), .ZN(U3115)
         );
  INV_X1 U7367 ( .A(n6461), .ZN(n6458) );
  AOI21_X1 U7368 ( .B1(n6448), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n6447), 
        .ZN(n6449) );
  AND2_X1 U7369 ( .A1(n6450), .A2(n6449), .ZN(n6453) );
  INV_X1 U7370 ( .A(n6453), .ZN(n6455) );
  AOI211_X1 U7371 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6453), .A(n6452), .B(n6451), .ZN(n6454) );
  AOI21_X1 U7372 ( .B1(n6456), .B2(n6455), .A(n6454), .ZN(n6457) );
  OAI21_X1 U7373 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6458), .A(n6457), 
        .ZN(n6459) );
  OAI21_X1 U7374 ( .B1(n6461), .B2(n6460), .A(n6459), .ZN(n6463) );
  INV_X1 U7375 ( .A(n6463), .ZN(n6466) );
  INV_X1 U7376 ( .A(n6465), .ZN(n6462) );
  AOI21_X1 U7377 ( .B1(n6463), .B2(n6462), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n6464) );
  AOI21_X1 U7378 ( .B1(n6466), .B2(n6465), .A(n6464), .ZN(n6474) );
  NOR2_X1 U7379 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6468) );
  OAI21_X1 U7380 ( .B1(n6469), .B2(n6468), .A(n6467), .ZN(n6470) );
  NOR3_X1 U7381 ( .A1(n6472), .A2(n6471), .A3(n6470), .ZN(n6473) );
  OAI21_X1 U7382 ( .B1(n6474), .B2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n6473), 
        .ZN(n6483) );
  NOR3_X1 U7383 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6475), .A3(n6590), .ZN(
        n6476) );
  OAI22_X1 U7384 ( .A1(n6479), .A2(n6478), .B1(n6477), .B2(n6476), .ZN(n6494)
         );
  AOI221_X1 U7385 ( .B1(n6480), .B2(n6596), .C1(n6480), .C2(n6483), .A(n6494), 
        .ZN(n6481) );
  INV_X1 U7386 ( .A(n6481), .ZN(n6572) );
  OAI21_X1 U7387 ( .B1(n6595), .B2(n6574), .A(n6572), .ZN(n6486) );
  AOI221_X1 U7388 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6572), .C1(n6590), .C2(
        n6572), .A(n6596), .ZN(n6488) );
  AOI211_X1 U7389 ( .C1(n6490), .C2(n6483), .A(n6482), .B(n6488), .ZN(n6484)
         );
  OAI221_X1 U7390 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6486), .C1(n6596), .C2(
        n6485), .A(n6484), .ZN(U3148) );
  AOI21_X1 U7391 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6488), .A(n6487), .ZN(
        n6492) );
  NOR2_X1 U7392 ( .A1(READY_N), .A2(n6596), .ZN(n6495) );
  OAI221_X1 U7393 ( .B1(n6490), .B2(n6489), .C1(n6490), .C2(n6495), .A(n6572), 
        .ZN(n6491) );
  OAI211_X1 U7394 ( .C1(n6494), .C2(n6493), .A(n6492), .B(n6491), .ZN(U3149)
         );
  OAI211_X1 U7395 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6495), .A(n6569), .B(
        n6595), .ZN(n6496) );
  NAND2_X1 U7396 ( .A1(n6497), .A2(n6496), .ZN(U3150) );
  INV_X1 U7397 ( .A(n6498), .ZN(n6567) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6567), .ZN(U3151) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6567), .ZN(U3152) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6567), .ZN(U3153) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6567), .ZN(U3154) );
  AND2_X1 U7402 ( .A1(n6567), .A2(DATAWIDTH_REG_27__SCAN_IN), .ZN(U3155) );
  AND2_X1 U7403 ( .A1(n6567), .A2(DATAWIDTH_REG_26__SCAN_IN), .ZN(U3156) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6567), .ZN(U3157) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6567), .ZN(U3158) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6567), .ZN(U3159) );
  INV_X1 U7407 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6630) );
  NOR2_X1 U7408 ( .A1(n6498), .A2(n6630), .ZN(U3160) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6567), .ZN(U3161) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6567), .ZN(U3162) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6567), .ZN(U3163) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6567), .ZN(U3164) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6567), .ZN(U3165) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6567), .ZN(U3166) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6567), .ZN(U3167) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6567), .ZN(U3168) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6567), .ZN(U3169) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6567), .ZN(U3170) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6567), .ZN(U3171) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6567), .ZN(U3172) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6567), .ZN(U3173) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6567), .ZN(U3174) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6567), .ZN(U3175) );
  AND2_X1 U7424 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6567), .ZN(U3176) );
  AND2_X1 U7425 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6567), .ZN(U3177) );
  AND2_X1 U7426 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6567), .ZN(U3178) );
  AND2_X1 U7427 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6567), .ZN(U3179) );
  AND2_X1 U7428 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6567), .ZN(U3180) );
  NOR2_X1 U7429 ( .A1(n6515), .A2(n6505), .ZN(n6506) );
  AOI22_X1 U7430 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6514) );
  AND2_X1 U7431 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6502) );
  INV_X1 U7432 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6500) );
  INV_X1 U7433 ( .A(NA_N), .ZN(n6507) );
  AOI221_X1 U7434 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6507), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6511) );
  AOI221_X1 U7435 ( .B1(n6502), .B2(n6606), .C1(n6500), .C2(n6606), .A(n6511), 
        .ZN(n6499) );
  OAI21_X1 U7436 ( .B1(n6506), .B2(n6514), .A(n6499), .ZN(U3181) );
  NOR2_X1 U7437 ( .A1(n6509), .A2(n6500), .ZN(n6508) );
  NAND2_X1 U7438 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6501) );
  OAI21_X1 U7439 ( .B1(n6508), .B2(n6502), .A(n6501), .ZN(n6503) );
  OAI211_X1 U7440 ( .C1(n6505), .C2(n6590), .A(n6504), .B(n6503), .ZN(U3182)
         );
  AOI21_X1 U7441 ( .B1(n6508), .B2(n6507), .A(n6506), .ZN(n6513) );
  AOI221_X1 U7442 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6590), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6510) );
  AOI221_X1 U7443 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6510), .C2(HOLD), .A(n6509), .ZN(n6512) );
  OAI22_X1 U7444 ( .A1(n6514), .A2(n6513), .B1(n6512), .B2(n6511), .ZN(U3183)
         );
  NOR2_X2 U7445 ( .A1(n6515), .A2(n6606), .ZN(n6558) );
  INV_X1 U7446 ( .A(n6558), .ZN(n6563) );
  NAND2_X1 U7447 ( .A1(n6515), .A2(n6553), .ZN(n6560) );
  INV_X1 U7448 ( .A(n6560), .ZN(n6561) );
  AOI22_X1 U7449 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6550), .ZN(n6516) );
  OAI21_X1 U7450 ( .B1(n6804), .B2(n6563), .A(n6516), .ZN(U3184) );
  INV_X1 U7451 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6518) );
  AOI22_X1 U7452 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6550), .ZN(n6517) );
  OAI21_X1 U7453 ( .B1(n6518), .B2(n6563), .A(n6517), .ZN(U3185) );
  AOI22_X1 U7454 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6550), .ZN(n6519) );
  OAI21_X1 U7455 ( .B1(n6520), .B2(n6560), .A(n6519), .ZN(U3186) );
  AOI22_X1 U7456 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6550), .ZN(n6521) );
  OAI21_X1 U7457 ( .B1(n6522), .B2(n6560), .A(n6521), .ZN(U3187) );
  AOI22_X1 U7458 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6550), .ZN(n6523) );
  OAI21_X1 U7459 ( .B1(n6525), .B2(n6560), .A(n6523), .ZN(U3188) );
  AOI22_X1 U7460 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6550), .ZN(n6524) );
  OAI21_X1 U7461 ( .B1(n6525), .B2(n6563), .A(n6524), .ZN(U3189) );
  AOI22_X1 U7462 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6550), .ZN(n6526) );
  OAI21_X1 U7463 ( .B1(n6527), .B2(n6563), .A(n6526), .ZN(U3190) );
  AOI22_X1 U7464 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6550), .ZN(n6528) );
  OAI21_X1 U7465 ( .B1(n6529), .B2(n6563), .A(n6528), .ZN(U3191) );
  AOI22_X1 U7466 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6550), .ZN(n6530) );
  OAI21_X1 U7467 ( .B1(n6532), .B2(n6560), .A(n6530), .ZN(U3192) );
  AOI22_X1 U7468 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6550), .ZN(n6531) );
  OAI21_X1 U7469 ( .B1(n6532), .B2(n6563), .A(n6531), .ZN(U3193) );
  AOI22_X1 U7470 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6550), .ZN(n6533) );
  OAI21_X1 U7471 ( .B1(n6534), .B2(n6560), .A(n6533), .ZN(U3194) );
  AOI22_X1 U7472 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6606), .ZN(n6535) );
  OAI21_X1 U7473 ( .B1(n6779), .B2(n6560), .A(n6535), .ZN(U3195) );
  AOI22_X1 U7474 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6550), .ZN(n6536) );
  OAI21_X1 U7475 ( .B1(n6623), .B2(n6560), .A(n6536), .ZN(U3196) );
  AOI22_X1 U7476 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6550), .ZN(n6537) );
  OAI21_X1 U7477 ( .B1(n6623), .B2(n6563), .A(n6537), .ZN(U3197) );
  AOI22_X1 U7478 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6550), .ZN(n6538) );
  OAI21_X1 U7479 ( .B1(n6540), .B2(n6560), .A(n6538), .ZN(U3198) );
  AOI22_X1 U7480 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6550), .ZN(n6539) );
  OAI21_X1 U7481 ( .B1(n6540), .B2(n6563), .A(n6539), .ZN(U3199) );
  INV_X1 U7482 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6543) );
  AOI22_X1 U7483 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6550), .ZN(n6541) );
  OAI21_X1 U7484 ( .B1(n6543), .B2(n6560), .A(n6541), .ZN(U3200) );
  AOI22_X1 U7485 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6550), .ZN(n6542) );
  OAI21_X1 U7486 ( .B1(n6543), .B2(n6563), .A(n6542), .ZN(U3201) );
  AOI22_X1 U7487 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6550), .ZN(n6544) );
  OAI21_X1 U7488 ( .B1(n5700), .B2(n6563), .A(n6544), .ZN(U3202) );
  AOI22_X1 U7489 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6550), .ZN(n6545) );
  OAI21_X1 U7490 ( .B1(n5679), .B2(n6560), .A(n6545), .ZN(U3203) );
  AOI22_X1 U7491 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6550), .ZN(n6546) );
  OAI21_X1 U7492 ( .B1(n5679), .B2(n6563), .A(n6546), .ZN(U3204) );
  AOI22_X1 U7493 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6550), .ZN(n6547) );
  OAI21_X1 U7494 ( .B1(n6548), .B2(n6560), .A(n6547), .ZN(U3205) );
  AOI22_X1 U7495 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6550), .ZN(n6549) );
  OAI21_X1 U7496 ( .B1(n5498), .B2(n6560), .A(n6549), .ZN(U3206) );
  AOI22_X1 U7497 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6550), .ZN(n6551) );
  OAI21_X1 U7498 ( .B1(n5498), .B2(n6563), .A(n6551), .ZN(U3207) );
  AOI22_X1 U7499 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6606), .ZN(n6552) );
  OAI21_X1 U7500 ( .B1(n6803), .B2(n6563), .A(n6552), .ZN(U3208) );
  INV_X1 U7501 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6770) );
  OAI222_X1 U7502 ( .A1(n6563), .A2(n6641), .B1(n6770), .B2(n6553), .C1(n6555), 
        .C2(n6560), .ZN(U3209) );
  AOI22_X1 U7503 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6606), .ZN(n6554) );
  OAI21_X1 U7504 ( .B1(n6555), .B2(n6563), .A(n6554), .ZN(U3210) );
  AOI22_X1 U7505 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6606), .ZN(n6556) );
  OAI21_X1 U7506 ( .B1(n6557), .B2(n6560), .A(n6556), .ZN(U3211) );
  AOI22_X1 U7507 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6558), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6606), .ZN(n6559) );
  OAI21_X1 U7508 ( .B1(n6564), .B2(n6560), .A(n6559), .ZN(U3212) );
  AOI22_X1 U7509 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6561), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6606), .ZN(n6562) );
  OAI21_X1 U7510 ( .B1(n6564), .B2(n6563), .A(n6562), .ZN(U3213) );
  MUX2_X1 U7511 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6606), .Z(U3445) );
  MUX2_X1 U7512 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6606), .Z(U3446) );
  MUX2_X1 U7513 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6606), .Z(U3447) );
  MUX2_X1 U7514 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6606), .Z(U3448) );
  INV_X1 U7515 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6581) );
  INV_X1 U7516 ( .A(n6565), .ZN(n6566) );
  AOI21_X1 U7517 ( .B1(n6581), .B2(n6567), .A(n6566), .ZN(U3451) );
  AOI21_X1 U7518 ( .B1(n6567), .B2(DATAWIDTH_REG_1__SCAN_IN), .A(n6566), .ZN(
        n6568) );
  INV_X1 U7519 ( .A(n6568), .ZN(U3452) );
  OAI211_X1 U7520 ( .C1(n6572), .C2(n6571), .A(n6570), .B(n6569), .ZN(U3453)
         );
  INV_X1 U7521 ( .A(n6573), .ZN(n6577) );
  OAI22_X1 U7522 ( .A1(n6577), .A2(n6576), .B1(n6575), .B2(n6574), .ZN(n6579)
         );
  MUX2_X1 U7523 ( .A(n6579), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6578), 
        .Z(U3456) );
  NOR3_X1 U7524 ( .A1(n6581), .A2(REIP_REG_0__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6580) );
  AOI221_X1 U7525 ( .B1(n6582), .B2(n6581), .C1(REIP_REG_1__SCAN_IN), .C2(
        REIP_REG_0__SCAN_IN), .A(n6580), .ZN(n6584) );
  INV_X1 U7526 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6583) );
  INV_X1 U7527 ( .A(n6588), .ZN(n6585) );
  AOI22_X1 U7528 ( .A1(n6588), .A2(n6584), .B1(n6583), .B2(n6585), .ZN(U3468)
         );
  NOR2_X1 U7529 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6587) );
  INV_X1 U7530 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6586) );
  AOI22_X1 U7531 ( .A1(n6588), .A2(n6587), .B1(n6586), .B2(n6585), .ZN(U3469)
         );
  NAND2_X1 U7532 ( .A1(n6606), .A2(W_R_N_REG_SCAN_IN), .ZN(n6589) );
  OAI21_X1 U7533 ( .B1(n6606), .B2(READREQUEST_REG_SCAN_IN), .A(n6589), .ZN(
        U3470) );
  NAND2_X1 U7534 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6590), .ZN(n6602) );
  INV_X1 U7535 ( .A(n6591), .ZN(n6592) );
  AOI211_X1 U7536 ( .C1(n6594), .C2(n6593), .A(n6602), .B(n6592), .ZN(n6597)
         );
  OAI21_X1 U7537 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(n6605) );
  INV_X1 U7538 ( .A(n6598), .ZN(n6601) );
  INV_X1 U7539 ( .A(n6599), .ZN(n6600) );
  OAI211_X1 U7540 ( .C1(n6603), .C2(n6602), .A(n6601), .B(n6600), .ZN(n6604)
         );
  MUX2_X1 U7541 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(n6605), .S(n6604), .Z(
        U3472) );
  MUX2_X1 U7542 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6606), .Z(U3473) );
  NOR3_X1 U7543 ( .A1(n6608), .A2(REIP_REG_14__SCAN_IN), .A3(n6607), .ZN(n6609) );
  AOI211_X1 U7544 ( .C1(n6611), .C2(EBX_REG_14__SCAN_IN), .A(n6610), .B(n6609), 
        .ZN(n6618) );
  INV_X1 U7545 ( .A(n6612), .ZN(n6616) );
  AOI22_X1 U7546 ( .A1(n6616), .A2(n6615), .B1(n6614), .B2(n6613), .ZN(n6617)
         );
  OAI211_X1 U7547 ( .C1(n6620), .C2(n6619), .A(n6618), .B(n6617), .ZN(n6627)
         );
  INV_X1 U7548 ( .A(n6621), .ZN(n6625) );
  OAI22_X1 U7549 ( .A1(n6625), .A2(n6624), .B1(n6623), .B2(n6622), .ZN(n6626)
         );
  NOR2_X1 U7550 ( .A1(n6627), .A2(n6626), .ZN(n6824) );
  AOI22_X1 U7551 ( .A1(n6757), .A2(keyinput94), .B1(n6780), .B2(keyinput118), 
        .ZN(n6628) );
  OAI221_X1 U7552 ( .B1(n6757), .B2(keyinput94), .C1(n6780), .C2(keyinput118), 
        .A(n6628), .ZN(n6638) );
  AOI22_X1 U7553 ( .A1(n6630), .A2(keyinput115), .B1(keyinput127), .B2(n6807), 
        .ZN(n6629) );
  OAI221_X1 U7554 ( .B1(n6630), .B2(keyinput115), .C1(n6807), .C2(keyinput127), 
        .A(n6629), .ZN(n6637) );
  AOI22_X1 U7555 ( .A1(n4817), .A2(keyinput67), .B1(keyinput95), .B2(n6632), 
        .ZN(n6631) );
  OAI221_X1 U7556 ( .B1(n4817), .B2(keyinput67), .C1(n6632), .C2(keyinput95), 
        .A(n6631), .ZN(n6636) );
  AOI22_X1 U7557 ( .A1(n6634), .A2(keyinput76), .B1(keyinput96), .B2(n6792), 
        .ZN(n6633) );
  OAI221_X1 U7558 ( .B1(n6634), .B2(keyinput76), .C1(n6792), .C2(keyinput96), 
        .A(n6633), .ZN(n6635) );
  NOR4_X1 U7559 ( .A1(n6638), .A2(n6637), .A3(n6636), .A4(n6635), .ZN(n6682)
         );
  AOI22_X1 U7560 ( .A1(n6763), .A2(keyinput89), .B1(keyinput126), .B2(n6777), 
        .ZN(n6639) );
  OAI221_X1 U7561 ( .B1(n6763), .B2(keyinput89), .C1(n6777), .C2(keyinput126), 
        .A(n6639), .ZN(n6649) );
  INV_X1 U7562 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6808) );
  AOI22_X1 U7563 ( .A1(n6808), .A2(keyinput125), .B1(keyinput120), .B2(n4328), 
        .ZN(n6640) );
  OAI221_X1 U7564 ( .B1(n6808), .B2(keyinput125), .C1(n4328), .C2(keyinput120), 
        .A(n6640), .ZN(n6648) );
  XOR2_X1 U7565 ( .A(n6641), .B(keyinput122), .Z(n6644) );
  XNOR2_X1 U7566 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .B(keyinput90), .ZN(n6643) );
  XNOR2_X1 U7567 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput121), .ZN(
        n6642) );
  NAND3_X1 U7568 ( .A1(n6644), .A2(n6643), .A3(n6642), .ZN(n6647) );
  XNOR2_X1 U7569 ( .A(n6645), .B(keyinput87), .ZN(n6646) );
  NOR4_X1 U7570 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n6681)
         );
  AOI22_X1 U7571 ( .A1(n6651), .A2(keyinput85), .B1(n4102), .B2(keyinput104), 
        .ZN(n6650) );
  OAI221_X1 U7572 ( .B1(n6651), .B2(keyinput85), .C1(n4102), .C2(keyinput104), 
        .A(n6650), .ZN(n6652) );
  INV_X1 U7573 ( .A(n6652), .ZN(n6665) );
  AOI22_X1 U7574 ( .A1(n6655), .A2(keyinput69), .B1(n6654), .B2(keyinput103), 
        .ZN(n6653) );
  OAI221_X1 U7575 ( .B1(n6655), .B2(keyinput69), .C1(n6654), .C2(keyinput103), 
        .A(n6653), .ZN(n6656) );
  INV_X1 U7576 ( .A(n6656), .ZN(n6664) );
  INV_X1 U7577 ( .A(keyinput83), .ZN(n6657) );
  XNOR2_X1 U7578 ( .A(n6658), .B(n6657), .ZN(n6663) );
  XNOR2_X1 U7579 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .B(keyinput88), .ZN(n6661)
         );
  XNOR2_X1 U7580 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .B(keyinput99), .ZN(n6660)
         );
  XNOR2_X1 U7581 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .B(keyinput105), .ZN(
        n6659) );
  AND3_X1 U7582 ( .A1(n6661), .A2(n6660), .A3(n6659), .ZN(n6662) );
  AND4_X1 U7583 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6680)
         );
  INV_X1 U7584 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6667) );
  AOI22_X1 U7585 ( .A1(n6667), .A2(keyinput107), .B1(keyinput75), .B2(n6764), 
        .ZN(n6666) );
  OAI221_X1 U7586 ( .B1(n6667), .B2(keyinput107), .C1(n6764), .C2(keyinput75), 
        .A(n6666), .ZN(n6678) );
  INV_X1 U7587 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6756) );
  INV_X1 U7588 ( .A(BS16_N), .ZN(n6789) );
  AOI22_X1 U7589 ( .A1(n6756), .A2(keyinput106), .B1(keyinput70), .B2(n6789), 
        .ZN(n6668) );
  OAI221_X1 U7590 ( .B1(n6756), .B2(keyinput106), .C1(n6789), .C2(keyinput70), 
        .A(n6668), .ZN(n6677) );
  INV_X1 U7591 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U7592 ( .A1(n6671), .A2(keyinput64), .B1(n6670), .B2(keyinput78), 
        .ZN(n6669) );
  OAI221_X1 U7593 ( .B1(n6671), .B2(keyinput64), .C1(n6670), .C2(keyinput78), 
        .A(n6669), .ZN(n6676) );
  INV_X1 U7594 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6672) );
  XOR2_X1 U7595 ( .A(n6672), .B(keyinput77), .Z(n6674) );
  XNOR2_X1 U7596 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput80), .ZN(
        n6673) );
  NAND2_X1 U7597 ( .A1(n6674), .A2(n6673), .ZN(n6675) );
  NOR4_X1 U7598 ( .A1(n6678), .A2(n6677), .A3(n6676), .A4(n6675), .ZN(n6679)
         );
  AND4_X1 U7599 ( .A1(n6682), .A2(n6681), .A3(n6680), .A4(n6679), .ZN(n6822)
         );
  OAI22_X1 U7600 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(keyinput117), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput82), .ZN(n6683) );
  AOI221_X1 U7601 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput117), 
        .C1(keyinput82), .C2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6683), .ZN(
        n6690) );
  OAI22_X1 U7602 ( .A1(REIP_REG_1__SCAN_IN), .A2(keyinput100), .B1(
        DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput74), .ZN(n6684) );
  AOI221_X1 U7603 ( .B1(REIP_REG_1__SCAN_IN), .B2(keyinput100), .C1(keyinput74), .C2(DATAWIDTH_REG_26__SCAN_IN), .A(n6684), .ZN(n6689) );
  OAI22_X1 U7604 ( .A1(EBX_REG_20__SCAN_IN), .A2(keyinput119), .B1(keyinput93), 
        .B2(ADDRESS_REG_25__SCAN_IN), .ZN(n6685) );
  AOI221_X1 U7605 ( .B1(EBX_REG_20__SCAN_IN), .B2(keyinput119), .C1(
        ADDRESS_REG_25__SCAN_IN), .C2(keyinput93), .A(n6685), .ZN(n6688) );
  OAI22_X1 U7606 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(keyinput68), .B1(
        DATAI_9_), .B2(keyinput114), .ZN(n6686) );
  AOI221_X1 U7607 ( .B1(INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput68), .C1(
        keyinput114), .C2(DATAI_9_), .A(n6686), .ZN(n6687) );
  NAND4_X1 U7608 ( .A1(n6690), .A2(n6689), .A3(n6688), .A4(n6687), .ZN(n6718)
         );
  OAI22_X1 U7609 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(keyinput116), .B1(
        EAX_REG_25__SCAN_IN), .B2(keyinput84), .ZN(n6691) );
  AOI221_X1 U7610 ( .B1(INSTQUEUE_REG_2__2__SCAN_IN), .B2(keyinput116), .C1(
        keyinput84), .C2(EAX_REG_25__SCAN_IN), .A(n6691), .ZN(n6698) );
  OAI22_X1 U7611 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(keyinput91), .B1(
        DATAI_16_), .B2(keyinput73), .ZN(n6692) );
  AOI221_X1 U7612 ( .B1(INSTQUEUE_REG_2__0__SCAN_IN), .B2(keyinput91), .C1(
        keyinput73), .C2(DATAI_16_), .A(n6692), .ZN(n6697) );
  OAI22_X1 U7613 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(keyinput113), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput72), .ZN(n6693) );
  AOI221_X1 U7614 ( .B1(INSTQUEUE_REG_6__5__SCAN_IN), .B2(keyinput113), .C1(
        keyinput72), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6693), .ZN(n6696) );
  OAI22_X1 U7615 ( .A1(DATAI_6_), .A2(keyinput66), .B1(keyinput124), .B2(
        BYTEENABLE_REG_3__SCAN_IN), .ZN(n6694) );
  AOI221_X1 U7616 ( .B1(DATAI_6_), .B2(keyinput66), .C1(
        BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput124), .A(n6694), .ZN(n6695) );
  NAND4_X1 U7617 ( .A1(n6698), .A2(n6697), .A3(n6696), .A4(n6695), .ZN(n6717)
         );
  OAI22_X1 U7618 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(keyinput123), .B1(
        REIP_REG_13__SCAN_IN), .B2(keyinput86), .ZN(n6699) );
  AOI221_X1 U7619 ( .B1(INSTQUEUE_REG_13__3__SCAN_IN), .B2(keyinput123), .C1(
        keyinput86), .C2(REIP_REG_13__SCAN_IN), .A(n6699), .ZN(n6706) );
  OAI22_X1 U7620 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput92), .B1(
        LWORD_REG_7__SCAN_IN), .B2(keyinput108), .ZN(n6700) );
  AOI221_X1 U7621 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput92), .C1(
        keyinput108), .C2(LWORD_REG_7__SCAN_IN), .A(n6700), .ZN(n6705) );
  INV_X1 U7622 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6791) );
  OAI22_X1 U7623 ( .A1(n6791), .A2(keyinput97), .B1(keyinput98), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6701) );
  AOI221_X1 U7624 ( .B1(n6791), .B2(keyinput97), .C1(LWORD_REG_14__SCAN_IN), 
        .C2(keyinput98), .A(n6701), .ZN(n6704) );
  OAI22_X1 U7625 ( .A1(n6801), .A2(keyinput101), .B1(keyinput112), .B2(
        REIP_REG_21__SCAN_IN), .ZN(n6702) );
  AOI221_X1 U7626 ( .B1(n6801), .B2(keyinput101), .C1(REIP_REG_21__SCAN_IN), 
        .C2(keyinput112), .A(n6702), .ZN(n6703) );
  NAND4_X1 U7627 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(n6716)
         );
  OAI22_X1 U7628 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(keyinput102), .B1(
        REIP_REG_2__SCAN_IN), .B2(keyinput109), .ZN(n6707) );
  AOI221_X1 U7629 ( .B1(INSTQUEUE_REG_11__1__SCAN_IN), .B2(keyinput102), .C1(
        keyinput109), .C2(REIP_REG_2__SCAN_IN), .A(n6707), .ZN(n6714) );
  OAI22_X1 U7630 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(keyinput65), .B1(
        REIP_REG_25__SCAN_IN), .B2(keyinput111), .ZN(n6708) );
  AOI221_X1 U7631 ( .B1(INSTQUEUE_REG_14__0__SCAN_IN), .B2(keyinput65), .C1(
        keyinput111), .C2(REIP_REG_25__SCAN_IN), .A(n6708), .ZN(n6713) );
  OAI22_X1 U7632 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput81), .B1(
        keyinput71), .B2(DATAO_REG_10__SCAN_IN), .ZN(n6709) );
  AOI221_X1 U7633 ( .B1(PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput81), .C1(
        DATAO_REG_10__SCAN_IN), .C2(keyinput71), .A(n6709), .ZN(n6712) );
  OAI22_X1 U7634 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(keyinput79), .B1(
        DATAO_REG_31__SCAN_IN), .B2(keyinput110), .ZN(n6710) );
  AOI221_X1 U7635 ( .B1(DATAWIDTH_REG_27__SCAN_IN), .B2(keyinput79), .C1(
        keyinput110), .C2(DATAO_REG_31__SCAN_IN), .A(n6710), .ZN(n6711) );
  NAND4_X1 U7636 ( .A1(n6714), .A2(n6713), .A3(n6712), .A4(n6711), .ZN(n6715)
         );
  NOR4_X1 U7637 ( .A1(n6718), .A2(n6717), .A3(n6716), .A4(n6715), .ZN(n6821)
         );
  AOI22_X1 U7638 ( .A1(EBX_REG_13__SCAN_IN), .A2(keyinput23), .B1(
        INSTADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput0), .ZN(n6719) );
  OAI221_X1 U7639 ( .B1(EBX_REG_13__SCAN_IN), .B2(keyinput23), .C1(
        INSTADDRPOINTER_REG_24__SCAN_IN), .C2(keyinput0), .A(n6719), .ZN(n6726) );
  AOI22_X1 U7640 ( .A1(DATAI_1_), .A2(keyinput21), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput39), .ZN(n6720) );
  OAI221_X1 U7641 ( .B1(DATAI_1_), .B2(keyinput21), .C1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .C2(keyinput39), .A(n6720), .ZN(n6725) );
  AOI22_X1 U7642 ( .A1(UWORD_REG_5__SCAN_IN), .A2(keyinput56), .B1(
        INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput4), .ZN(n6721) );
  OAI221_X1 U7643 ( .B1(UWORD_REG_5__SCAN_IN), .B2(keyinput56), .C1(
        INSTQUEUE_REG_9__3__SCAN_IN), .C2(keyinput4), .A(n6721), .ZN(n6724) );
  AOI22_X1 U7644 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(keyinput26), .B1(
        INSTQUEUE_REG_14__0__SCAN_IN), .B2(keyinput1), .ZN(n6722) );
  OAI221_X1 U7645 ( .B1(INSTQUEUE_REG_15__6__SCAN_IN), .B2(keyinput26), .C1(
        INSTQUEUE_REG_14__0__SCAN_IN), .C2(keyinput1), .A(n6722), .ZN(n6723)
         );
  NOR4_X1 U7646 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6754)
         );
  AOI22_X1 U7647 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(keyinput51), .B1(
        DATAO_REG_10__SCAN_IN), .B2(keyinput7), .ZN(n6727) );
  OAI221_X1 U7648 ( .B1(DATAWIDTH_REG_22__SCAN_IN), .B2(keyinput51), .C1(
        DATAO_REG_10__SCAN_IN), .C2(keyinput7), .A(n6727), .ZN(n6734) );
  AOI22_X1 U7649 ( .A1(REIP_REG_26__SCAN_IN), .A2(keyinput58), .B1(
        INSTQUEUE_REG_12__5__SCAN_IN), .B2(keyinput3), .ZN(n6728) );
  OAI221_X1 U7650 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput58), .C1(
        INSTQUEUE_REG_12__5__SCAN_IN), .C2(keyinput3), .A(n6728), .ZN(n6733)
         );
  AOI22_X1 U7651 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput19), .B1(
        EBX_REG_11__SCAN_IN), .B2(keyinput12), .ZN(n6729) );
  OAI221_X1 U7652 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput19), .C1(
        EBX_REG_11__SCAN_IN), .C2(keyinput12), .A(n6729), .ZN(n6732) );
  AOI22_X1 U7653 ( .A1(EBX_REG_1__SCAN_IN), .A2(keyinput31), .B1(
        INSTQUEUE_REG_5__4__SCAN_IN), .B2(keyinput14), .ZN(n6730) );
  OAI221_X1 U7654 ( .B1(EBX_REG_1__SCAN_IN), .B2(keyinput31), .C1(
        INSTQUEUE_REG_5__4__SCAN_IN), .C2(keyinput14), .A(n6730), .ZN(n6731)
         );
  NOR4_X1 U7655 ( .A1(n6734), .A2(n6733), .A3(n6732), .A4(n6731), .ZN(n6753)
         );
  AOI22_X1 U7656 ( .A1(REIP_REG_2__SCAN_IN), .A2(keyinput45), .B1(
        INSTQUEUE_REG_15__5__SCAN_IN), .B2(keyinput13), .ZN(n6735) );
  OAI221_X1 U7657 ( .B1(REIP_REG_2__SCAN_IN), .B2(keyinput45), .C1(
        INSTQUEUE_REG_15__5__SCAN_IN), .C2(keyinput13), .A(n6735), .ZN(n6742)
         );
  AOI22_X1 U7658 ( .A1(UWORD_REG_11__SCAN_IN), .A2(keyinput5), .B1(
        DATAWIDTH_REG_27__SCAN_IN), .B2(keyinput15), .ZN(n6736) );
  OAI221_X1 U7659 ( .B1(UWORD_REG_11__SCAN_IN), .B2(keyinput5), .C1(
        DATAWIDTH_REG_27__SCAN_IN), .C2(keyinput15), .A(n6736), .ZN(n6741) );
  AOI22_X1 U7660 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(keyinput38), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(keyinput16), .ZN(n6737) );
  OAI221_X1 U7661 ( .B1(INSTQUEUE_REG_11__1__SCAN_IN), .B2(keyinput38), .C1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(keyinput16), .A(n6737), .ZN(
        n6740) );
  AOI22_X1 U7662 ( .A1(LWORD_REG_14__SCAN_IN), .A2(keyinput34), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput8), .ZN(n6738) );
  OAI221_X1 U7663 ( .B1(LWORD_REG_14__SCAN_IN), .B2(keyinput34), .C1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .C2(keyinput8), .A(n6738), .ZN(n6739)
         );
  NOR4_X1 U7664 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n6752)
         );
  AOI22_X1 U7665 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput48), .B1(
        EBX_REG_20__SCAN_IN), .B2(keyinput55), .ZN(n6743) );
  OAI221_X1 U7666 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput48), .C1(
        EBX_REG_20__SCAN_IN), .C2(keyinput55), .A(n6743), .ZN(n6750) );
  AOI22_X1 U7667 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(keyinput10), .B1(
        STATEBS16_REG_SCAN_IN), .B2(keyinput28), .ZN(n6744) );
  OAI221_X1 U7668 ( .B1(DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput10), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput28), .A(n6744), .ZN(n6749) );
  AOI22_X1 U7669 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(keyinput24), .B1(
        INSTQUEUE_REG_1__1__SCAN_IN), .B2(keyinput43), .ZN(n6745) );
  OAI221_X1 U7670 ( .B1(INSTQUEUE_REG_8__7__SCAN_IN), .B2(keyinput24), .C1(
        INSTQUEUE_REG_1__1__SCAN_IN), .C2(keyinput43), .A(n6745), .ZN(n6748)
         );
  AOI22_X1 U7671 ( .A1(DATAO_REG_31__SCAN_IN), .A2(keyinput46), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput53), .ZN(n6746) );
  OAI221_X1 U7672 ( .B1(DATAO_REG_31__SCAN_IN), .B2(keyinput46), .C1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .C2(keyinput53), .A(n6746), .ZN(n6747) );
  NOR4_X1 U7673 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n6751)
         );
  NAND4_X1 U7674 ( .A1(n6754), .A2(n6753), .A3(n6752), .A4(n6751), .ZN(n6820)
         );
  AOI22_X1 U7675 ( .A1(n6757), .A2(keyinput30), .B1(n6756), .B2(keyinput42), 
        .ZN(n6755) );
  OAI221_X1 U7676 ( .B1(n6757), .B2(keyinput30), .C1(n6756), .C2(keyinput42), 
        .A(n6755), .ZN(n6768) );
  AOI22_X1 U7677 ( .A1(n4102), .A2(keyinput40), .B1(keyinput20), .B2(n4311), 
        .ZN(n6758) );
  OAI221_X1 U7678 ( .B1(n4102), .B2(keyinput40), .C1(n4311), .C2(keyinput20), 
        .A(n6758), .ZN(n6767) );
  INV_X1 U7679 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6761) );
  INV_X1 U7680 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6760) );
  AOI22_X1 U7681 ( .A1(n6761), .A2(keyinput52), .B1(n6760), .B2(keyinput27), 
        .ZN(n6759) );
  OAI221_X1 U7682 ( .B1(n6761), .B2(keyinput52), .C1(n6760), .C2(keyinput27), 
        .A(n6759), .ZN(n6766) );
  AOI22_X1 U7683 ( .A1(n6764), .A2(keyinput11), .B1(n6763), .B2(keyinput25), 
        .ZN(n6762) );
  OAI221_X1 U7684 ( .B1(n6764), .B2(keyinput11), .C1(n6763), .C2(keyinput25), 
        .A(n6762), .ZN(n6765) );
  NOR4_X1 U7685 ( .A1(n6768), .A2(n6767), .A3(n6766), .A4(n6765), .ZN(n6818)
         );
  INV_X1 U7686 ( .A(DATAI_16_), .ZN(n6771) );
  AOI22_X1 U7687 ( .A1(n6771), .A2(keyinput9), .B1(keyinput29), .B2(n6770), 
        .ZN(n6769) );
  OAI221_X1 U7688 ( .B1(n6771), .B2(keyinput9), .C1(n6770), .C2(keyinput29), 
        .A(n6769), .ZN(n6784) );
  INV_X1 U7689 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6774) );
  AOI22_X1 U7690 ( .A1(n6774), .A2(keyinput59), .B1(keyinput17), .B2(n6773), 
        .ZN(n6772) );
  OAI221_X1 U7691 ( .B1(n6774), .B2(keyinput59), .C1(n6773), .C2(keyinput17), 
        .A(n6772), .ZN(n6783) );
  AOI22_X1 U7692 ( .A1(n6777), .A2(keyinput62), .B1(keyinput2), .B2(n6776), 
        .ZN(n6775) );
  OAI221_X1 U7693 ( .B1(n6777), .B2(keyinput62), .C1(n6776), .C2(keyinput2), 
        .A(n6775), .ZN(n6782) );
  AOI22_X1 U7694 ( .A1(n6780), .A2(keyinput54), .B1(keyinput22), .B2(n6779), 
        .ZN(n6778) );
  OAI221_X1 U7695 ( .B1(n6780), .B2(keyinput54), .C1(n6779), .C2(keyinput22), 
        .A(n6778), .ZN(n6781) );
  NOR4_X1 U7696 ( .A1(n6784), .A2(n6783), .A3(n6782), .A4(n6781), .ZN(n6817)
         );
  AOI22_X1 U7697 ( .A1(n6787), .A2(keyinput50), .B1(keyinput60), .B2(n6786), 
        .ZN(n6785) );
  OAI221_X1 U7698 ( .B1(n6787), .B2(keyinput50), .C1(n6786), .C2(keyinput60), 
        .A(n6785), .ZN(n6798) );
  AOI22_X1 U7699 ( .A1(n6789), .A2(keyinput6), .B1(n4325), .B2(keyinput44), 
        .ZN(n6788) );
  OAI221_X1 U7700 ( .B1(n6789), .B2(keyinput6), .C1(n4325), .C2(keyinput44), 
        .A(n6788), .ZN(n6797) );
  AOI22_X1 U7701 ( .A1(n6792), .A2(keyinput32), .B1(n6791), .B2(keyinput33), 
        .ZN(n6790) );
  OAI221_X1 U7702 ( .B1(n6792), .B2(keyinput32), .C1(n6791), .C2(keyinput33), 
        .A(n6790), .ZN(n6796) );
  XNOR2_X1 U7703 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput57), .ZN(
        n6794) );
  XNOR2_X1 U7704 ( .A(keyinput49), .B(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6793)
         );
  NAND2_X1 U7705 ( .A1(n6794), .A2(n6793), .ZN(n6795) );
  NOR4_X1 U7706 ( .A1(n6798), .A2(n6797), .A3(n6796), .A4(n6795), .ZN(n6816)
         );
  AOI22_X1 U7707 ( .A1(n6801), .A2(keyinput37), .B1(n6800), .B2(keyinput41), 
        .ZN(n6799) );
  OAI221_X1 U7708 ( .B1(n6801), .B2(keyinput37), .C1(n6800), .C2(keyinput41), 
        .A(n6799), .ZN(n6814) );
  AOI22_X1 U7709 ( .A1(n6804), .A2(keyinput36), .B1(n6803), .B2(keyinput47), 
        .ZN(n6802) );
  OAI221_X1 U7710 ( .B1(n6804), .B2(keyinput36), .C1(n6803), .C2(keyinput47), 
        .A(n6802), .ZN(n6813) );
  AOI22_X1 U7711 ( .A1(n6807), .A2(keyinput63), .B1(n6806), .B2(keyinput18), 
        .ZN(n6805) );
  OAI221_X1 U7712 ( .B1(n6807), .B2(keyinput63), .C1(n6806), .C2(keyinput18), 
        .A(n6805), .ZN(n6812) );
  XOR2_X1 U7713 ( .A(n6808), .B(keyinput61), .Z(n6810) );
  XNOR2_X1 U7714 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .B(keyinput35), .ZN(n6809)
         );
  NAND2_X1 U7715 ( .A1(n6810), .A2(n6809), .ZN(n6811) );
  NOR4_X1 U7716 ( .A1(n6814), .A2(n6813), .A3(n6812), .A4(n6811), .ZN(n6815)
         );
  NAND4_X1 U7717 ( .A1(n6818), .A2(n6817), .A3(n6816), .A4(n6815), .ZN(n6819)
         );
  AOI211_X1 U7718 ( .C1(n6822), .C2(n6821), .A(n6820), .B(n6819), .ZN(n6823)
         );
  XNOR2_X1 U7719 ( .A(n6824), .B(n6823), .ZN(U2813) );
  AND4_X1 U3973 ( .A1(n3118), .A2(n3117), .A3(n3116), .A4(n3115), .ZN(n3124)
         );
  CLKBUF_X2 U34720 ( .A(n3128), .Z(n3789) );
  CLKBUF_X1 U34730 ( .A(n3145), .Z(n3865) );
  AND2_X4 U3894 ( .A1(n4479), .A2(n5398), .ZN(n3145) );
  BUF_X2 U3491 ( .A(n3076), .Z(n3864) );
  CLKBUF_X1 U3492 ( .A(n3214), .Z(n3863) );
  AND4_X1 U3503 ( .A1(n3102), .A2(n3101), .A3(n3100), .A4(n3099), .ZN(n3103)
         );
  AND4_X1 U3508 ( .A1(n3080), .A2(n3079), .A3(n3078), .A4(n3077), .ZN(n3086)
         );
  BUF_X1 U3531 ( .A(n3178), .Z(n4185) );
  OR2_X1 U3550 ( .A1(n3151), .A2(n3150), .ZN(n4235) );
  CLKBUF_X1 U3558 ( .A(n5455), .Z(n5558) );
  CLKBUF_X1 U3606 ( .A(n5306), .Z(n5336) );
  CLKBUF_X1 U3649 ( .A(n3866), .Z(n4483) );
  CLKBUF_X1 U3658 ( .A(n3193), .Z(n4538) );
  CLKBUF_X1 U3723 ( .A(n3164), .Z(n3012) );
  CLKBUF_X1 U3770 ( .A(n4519), .Z(n3022) );
  CLKBUF_X1 U3796 ( .A(n4466), .Z(n5191) );
  CLKBUF_X1 U3815 ( .A(n4041), .Z(n5459) );
endmodule

