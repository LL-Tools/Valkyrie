

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, 
        keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, 
        keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, 
        keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, 
        keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, 
        keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, 
        keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, 
        keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, 
        keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, 
        keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, 
        keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525;

  INV_X1 U2241 ( .A(n3191), .ZN(n3261) );
  CLKBUF_X2 U2242 ( .A(n2459), .Z(n3434) );
  AND2_X2 U2243 ( .A1(n2303), .A2(n2302), .ZN(n3196) );
  CLKBUF_X3 U2244 ( .A(n2498), .Z(n3218) );
  NAND2_X1 U2245 ( .A1(n3768), .A2(n3705), .ZN(n2198) );
  NAND2_X1 U2246 ( .A1(n3552), .A2(n3491), .ZN(n2587) );
  NAND3_X1 U2247 ( .A1(n2040), .A2(n2039), .A3(n2151), .ZN(n3031) );
  AOI21_X1 U2248 ( .B1(n2561), .B2(n2049), .A(n2048), .ZN(n2717) );
  OAI21_X1 U2249 ( .B1(n3159), .B2(n2022), .A(n2044), .ZN(n3307) );
  NAND2_X1 U2250 ( .A1(n2062), .A2(n2061), .ZN(n2572) );
  XNOR2_X2 U2251 ( .A(n2868), .B(n2881), .ZN(n2870) );
  AND2_X2 U2252 ( .A1(n2108), .A2(n2107), .ZN(n2868) );
  XNOR2_X2 U2253 ( .A(n2110), .B(n2400), .ZN(n2395) );
  XNOR2_X2 U2254 ( .A(n2385), .B(n2676), .ZN(n2387) );
  AND2_X1 U2255 ( .A1(n2303), .A2(n2302), .ZN(n1999) );
  NAND2_X4 U2256 ( .A1(n2530), .A2(n2587), .ZN(n2423) );
  NAND2_X2 U2257 ( .A1(n2281), .A2(n2243), .ZN(n2530) );
  AOI21_X2 U2258 ( .B1(n3787), .B2(n3703), .A(n3702), .ZN(n3768) );
  OAI21_X1 U2259 ( .B1(n3066), .B2(n3065), .A(n3231), .ZN(n3067) );
  AND2_X1 U2260 ( .A1(n2922), .A2(n2921), .ZN(n2923) );
  AOI21_X1 U2261 ( .B1(n2514), .B2(n2513), .A(n2512), .ZN(n2522) );
  INV_X2 U2262 ( .A(n4284), .ZN(n2000) );
  OR2_X1 U2263 ( .A1(n2423), .A2(n4356), .ZN(n2498) );
  AND2_X1 U2264 ( .A1(n2197), .A2(n2011), .ZN(n3737) );
  OAI21_X1 U2265 ( .B1(n3239), .B2(n3184), .A(n3185), .ZN(n3333) );
  OR2_X1 U2266 ( .A1(n3239), .A2(n3182), .ZN(n2224) );
  NAND2_X1 U2267 ( .A1(n3159), .A2(n3158), .ZN(n3240) );
  OAI211_X1 U2268 ( .C1(n3315), .C2(n3403), .A(n3316), .B(n3401), .ZN(n3089)
         );
  NAND2_X1 U2269 ( .A1(n2046), .A2(n3083), .ZN(n3401) );
  NAND2_X1 U2270 ( .A1(n3067), .A2(n2047), .ZN(n2046) );
  OAI21_X1 U2271 ( .B1(n2895), .B2(n3517), .A(n3510), .ZN(n2983) );
  OAI21_X1 U2272 ( .B1(n2778), .B2(n2777), .A(n2776), .ZN(n2922) );
  NAND2_X1 U2273 ( .A1(n2540), .A2(n2541), .ZN(n2561) );
  NAND2_X1 U2274 ( .A1(n2539), .A2(n2538), .ZN(n2540) );
  NAND2_X1 U2275 ( .A1(n2522), .A2(n2521), .ZN(n2539) );
  AND2_X1 U2276 ( .A1(n2538), .A2(n2520), .ZN(n2521) );
  AOI21_X1 U2277 ( .B1(n2179), .B2(n2634), .A(n2002), .ZN(n2178) );
  INV_X1 U2278 ( .A(n2572), .ZN(n2463) );
  NAND2_X2 U2279 ( .A1(n2586), .A2(n4304), .ZN(n4284) );
  INV_X1 U2280 ( .A(n2498), .ZN(n3263) );
  INV_X2 U2281 ( .A(n3435), .ZN(n3282) );
  INV_X2 U2282 ( .A(n2009), .ZN(n3285) );
  NAND2_X4 U2283 ( .A1(n2087), .A2(n2086), .ZN(n3436) );
  NAND2_X2 U2284 ( .A1(n2493), .A2(n2587), .ZN(n3191) );
  INV_X1 U2285 ( .A(n2302), .ZN(n2301) );
  NAND2_X1 U2286 ( .A1(n2289), .A2(IR_REG_31__SCAN_IN), .ZN(n2290) );
  NAND2_X1 U2287 ( .A1(n2286), .A2(n4388), .ZN(n2289) );
  INV_X1 U2288 ( .A(n2455), .ZN(n3491) );
  XNOR2_X1 U2289 ( .A(n2269), .B(n2268), .ZN(n3552) );
  AND2_X1 U2290 ( .A1(n2042), .A2(n2041), .ZN(n2286) );
  AND2_X1 U2291 ( .A1(n2043), .A2(n2210), .ZN(n2042) );
  AND2_X1 U2292 ( .A1(n2093), .A2(n2019), .ZN(n2041) );
  AND2_X1 U2293 ( .A1(n2230), .A2(n4386), .ZN(n2094) );
  AND2_X1 U2294 ( .A1(n2212), .A2(n2211), .ZN(n2210) );
  AND4_X1 U2295 ( .A1(n2229), .A2(n2228), .A3(n2227), .A4(n2226), .ZN(n2230)
         );
  NOR2_X1 U2296 ( .A1(IR_REG_14__SCAN_IN), .A2(n2017), .ZN(n2212) );
  INV_X1 U2297 ( .A(IR_REG_3__SCAN_IN), .ZN(n2336) );
  INV_X1 U2298 ( .A(IR_REG_22__SCAN_IN), .ZN(n2277) );
  NOR2_X1 U2299 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2226)
         );
  NOR2_X1 U2300 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2227)
         );
  INV_X1 U2301 ( .A(IR_REG_1__SCAN_IN), .ZN(n2131) );
  NOR2_X1 U2302 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2228)
         );
  NOR2_X1 U2303 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2229)
         );
  INV_X1 U2304 ( .A(IR_REG_0__SCAN_IN), .ZN(n2038) );
  OAI21_X2 U2305 ( .B1(n3392), .B2(n3285), .A(n3200), .ZN(n3775) );
  AOI211_X2 U2306 ( .C1(n3355), .C2(n3064), .A(n3361), .B(n3063), .ZN(n3066)
         );
  INV_X1 U2307 ( .A(n3469), .ZN(n2203) );
  AOI21_X1 U2308 ( .B1(n3999), .B2(n3680), .A(n3679), .ZN(n3976) );
  AND2_X1 U2309 ( .A1(n3678), .A2(n3981), .ZN(n3679) );
  NAND2_X1 U2310 ( .A1(n2919), .A2(n2918), .ZN(n2925) );
  INV_X1 U2311 ( .A(n2927), .ZN(n2154) );
  INV_X1 U2312 ( .A(n2469), .ZN(n3435) );
  AND2_X1 U2313 ( .A1(n3568), .A2(n3452), .ZN(n3695) );
  NOR2_X1 U2314 ( .A1(n3005), .A2(n2209), .ZN(n2208) );
  INV_X1 U2315 ( .A(n2907), .ZN(n2209) );
  NAND2_X1 U2316 ( .A1(n2575), .A2(n2574), .ZN(n2603) );
  NAND2_X1 U2317 ( .A1(n2499), .A2(n2572), .ZN(n3489) );
  AND2_X1 U2318 ( .A1(n2236), .A2(n2070), .ZN(n2043) );
  INV_X1 U2319 ( .A(n2213), .ZN(n2070) );
  NOR2_X1 U2320 ( .A1(IR_REG_25__SCAN_IN), .A2(n2235), .ZN(n2236) );
  OAI22_X1 U2321 ( .A1(n3218), .A2(n2463), .B1(n2499), .B2(n3204), .ZN(n2510)
         );
  XNOR2_X1 U2322 ( .A(n2497), .B(n3191), .ZN(n2511) );
  OAI22_X1 U2323 ( .A1(n2463), .A2(n3081), .B1(n2499), .B2(n2423), .ZN(n2497)
         );
  AOI21_X1 U2324 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2424), .A(n2494), .ZN(n2496)
         );
  NAND2_X1 U2325 ( .A1(n2420), .A2(n2419), .ZN(n2421) );
  NAND2_X1 U2326 ( .A1(n2424), .A2(IR_REG_0__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U2327 ( .A1(n3258), .A2(n2478), .ZN(n2419) );
  OR2_X1 U2328 ( .A1(n2454), .A2(n4171), .ZN(n2493) );
  NOR2_X1 U2329 ( .A1(n2303), .A2(n2301), .ZN(n2459) );
  NOR2_X1 U2330 ( .A1(n2242), .A2(n2435), .ZN(n2243) );
  OR2_X1 U2331 ( .A1(n2079), .A2(n2546), .ZN(n2078) );
  INV_X1 U2332 ( .A(n2342), .ZN(n2079) );
  XNOR2_X1 U2333 ( .A(n2340), .B(n4201), .ZN(n4195) );
  NOR2_X1 U2334 ( .A1(n2013), .A2(n2194), .ZN(n2193) );
  OR2_X1 U2335 ( .A1(n2195), .A2(n2013), .ZN(n2192) );
  AND2_X1 U2336 ( .A1(n2011), .A2(n3709), .ZN(n2195) );
  AND2_X1 U2337 ( .A1(n3816), .A2(n3797), .ZN(n3702) );
  AND2_X1 U2338 ( .A1(n3688), .A2(n3687), .ZN(n3689) );
  AOI21_X1 U2339 ( .B1(n3676), .B2(n3675), .A(n3674), .ZN(n3999) );
  AND2_X1 U2340 ( .A1(n3578), .A2(n2478), .ZN(n2465) );
  INV_X1 U2341 ( .A(n2573), .ZN(n2499) );
  NAND2_X1 U2342 ( .A1(n2530), .A2(n4312), .ZN(n2582) );
  OAI211_X1 U2343 ( .C1(IR_REG_31__SCAN_IN), .C2(IR_REG_29__SCAN_IN), .A(n2289), .B(n2066), .ZN(n2302) );
  OR2_X1 U2344 ( .A1(n2286), .A2(n2067), .ZN(n2066) );
  NAND2_X1 U2345 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2067) );
  INV_X1 U2346 ( .A(n2326), .ZN(n2327) );
  INV_X1 U2347 ( .A(n3571), .ZN(n2948) );
  INV_X1 U2348 ( .A(n2702), .ZN(n2631) );
  NAND2_X1 U2349 ( .A1(n2091), .A2(IR_REG_28__SCAN_IN), .ZN(n2090) );
  NAND2_X1 U2350 ( .A1(n3258), .A2(n2012), .ZN(n2174) );
  NAND2_X1 U2351 ( .A1(n3258), .A2(n2173), .ZN(n2172) );
  AOI21_X1 U2352 ( .B1(n2168), .B2(n2165), .A(n2164), .ZN(n2163) );
  INV_X1 U2353 ( .A(n2170), .ZN(n2165) );
  INV_X1 U2354 ( .A(n3250), .ZN(n2164) );
  INV_X1 U2355 ( .A(n2168), .ZN(n2166) );
  AND2_X1 U2356 ( .A1(n2943), .A2(n2924), .ZN(n2152) );
  INV_X1 U2357 ( .A(n2963), .ZN(n2964) );
  INV_X1 U2358 ( .A(n2655), .ZN(n2158) );
  AND2_X1 U2359 ( .A1(n3430), .A2(n3429), .ZN(n3655) );
  AND2_X1 U2360 ( .A1(n3449), .A2(n3752), .ZN(n3659) );
  AND2_X1 U2361 ( .A1(n3600), .A2(n3599), .ZN(n3601) );
  OR2_X1 U2362 ( .A1(n3186), .A2(n3309), .ZN(n3194) );
  NAND2_X1 U2363 ( .A1(n3753), .A2(n3659), .ZN(n2060) );
  NAND2_X1 U2364 ( .A1(n3770), .A2(n3657), .ZN(n3753) );
  OAI21_X1 U2365 ( .B1(n3977), .B2(n2135), .A(n3685), .ZN(n2134) );
  AND2_X1 U2366 ( .A1(n3420), .A2(n3459), .ZN(n3524) );
  AND2_X1 U2367 ( .A1(n2007), .A2(n3706), .ZN(n2098) );
  AND2_X1 U2368 ( .A1(n2101), .A2(n3004), .ZN(n2100) );
  AND2_X1 U2369 ( .A1(n2917), .A2(n2841), .ZN(n2101) );
  NAND2_X1 U2370 ( .A1(n2232), .A2(IR_REG_31__SCAN_IN), .ZN(n2246) );
  NAND2_X1 U2371 ( .A1(n2268), .A2(n2266), .ZN(n2216) );
  INV_X1 U2372 ( .A(IR_REG_20__SCAN_IN), .ZN(n2268) );
  INV_X1 U2373 ( .A(IR_REG_19__SCAN_IN), .ZN(n2266) );
  INV_X1 U2374 ( .A(IR_REG_17__SCAN_IN), .ZN(n2211) );
  AOI21_X1 U2375 ( .B1(n2170), .B2(n3105), .A(n2169), .ZN(n2168) );
  INV_X1 U2376 ( .A(n3379), .ZN(n2169) );
  NAND2_X1 U2377 ( .A1(n2219), .A2(n3180), .ZN(n2218) );
  INV_X1 U2378 ( .A(n3335), .ZN(n2219) );
  NAND2_X1 U2379 ( .A1(n2654), .A2(n2653), .ZN(n2655) );
  INV_X1 U2380 ( .A(n2652), .ZN(n2654) );
  AND2_X1 U2381 ( .A1(n2562), .A2(n2560), .ZN(n2159) );
  NOR2_X1 U2382 ( .A1(n2923), .A2(n2154), .ZN(n2153) );
  NAND2_X1 U2383 ( .A1(n2085), .A2(n2084), .ZN(n2478) );
  OAI21_X1 U2384 ( .B1(n2088), .B2(n2089), .A(DATAI_0_), .ZN(n2084) );
  AND2_X1 U2385 ( .A1(n2511), .A2(n2510), .ZN(n2512) );
  AND2_X1 U2386 ( .A1(n3070), .A2(n3069), .ZN(n3403) );
  NOR2_X1 U2387 ( .A1(n2388), .A2(n2106), .ZN(n2105) );
  NOR2_X1 U2388 ( .A1(n2388), .A2(n2373), .ZN(n2104) );
  OR2_X1 U2389 ( .A1(n2369), .A2(n2368), .ZN(n2380) );
  NAND2_X1 U2390 ( .A1(n4209), .A2(n2025), .ZN(n2871) );
  OR2_X1 U2391 ( .A1(n4233), .A2(n2887), .ZN(n2076) );
  NAND2_X1 U2392 ( .A1(n2076), .A2(n2075), .ZN(n3600) );
  INV_X1 U2393 ( .A(n2890), .ZN(n2075) );
  XNOR2_X1 U2394 ( .A(n3601), .B(n4317), .ZN(n4243) );
  OR2_X1 U2395 ( .A1(n2008), .A2(n4258), .ZN(n2127) );
  OR2_X1 U2396 ( .A1(n4243), .A2(n2128), .ZN(n2126) );
  OR2_X1 U2397 ( .A1(n4258), .A2(n4244), .ZN(n2128) );
  OR2_X1 U2398 ( .A1(n4243), .A2(n4244), .ZN(n2129) );
  NOR2_X1 U2399 ( .A1(n4261), .A2(n3612), .ZN(n3620) );
  NAND2_X1 U2400 ( .A1(n4269), .A2(n2102), .ZN(n3623) );
  NAND2_X1 U2401 ( .A1(n4282), .A2(n2103), .ZN(n2102) );
  NOR2_X1 U2402 ( .A1(n3623), .A2(n3624), .ZN(n3638) );
  OR2_X1 U2403 ( .A1(n3220), .A2(n3277), .ZN(n3648) );
  NOR2_X1 U2404 ( .A1(n3194), .A2(n3393), .ZN(n3208) );
  NAND2_X1 U2405 ( .A1(n3707), .A2(n2024), .ZN(n2194) );
  AND2_X1 U2406 ( .A1(n3215), .A2(n3214), .ZN(n3759) );
  AND3_X1 U2407 ( .A1(n3179), .A2(n3178), .A3(n3177), .ZN(n3816) );
  AOI21_X1 U2408 ( .B1(n2139), .B2(n2004), .A(n2140), .ZN(n3827) );
  INV_X1 U2409 ( .A(n3902), .ZN(n2139) );
  AOI21_X1 U2410 ( .B1(n2144), .B2(n2146), .A(n2143), .ZN(n2142) );
  INV_X1 U2411 ( .A(n3694), .ZN(n2143) );
  INV_X1 U2412 ( .A(n2149), .ZN(n2144) );
  NOR2_X1 U2413 ( .A1(n2150), .A2(n3693), .ZN(n2149) );
  INV_X1 U2414 ( .A(n3691), .ZN(n2150) );
  OR2_X1 U2415 ( .A1(n3949), .A2(n3957), .ZN(n3686) );
  NOR2_X1 U2416 ( .A1(n3048), .A2(n3406), .ZN(n3071) );
  NAND2_X1 U2417 ( .A1(n2054), .A2(n3650), .ZN(n3960) );
  NAND2_X1 U2418 ( .A1(n3978), .A2(n3649), .ZN(n2054) );
  INV_X1 U2419 ( .A(n3683), .ZN(n3979) );
  NAND2_X1 U2420 ( .A1(n2974), .A2(REG3_REG_12__SCAN_IN), .ZN(n2989) );
  AOI21_X1 U2421 ( .B1(n2201), .B2(n2200), .A(n2026), .ZN(n2199) );
  INV_X1 U2422 ( .A(n2208), .ZN(n2200) );
  INV_X1 U2423 ( .A(n2206), .ZN(n2205) );
  OAI22_X1 U2424 ( .A1(n3005), .A2(n2207), .B1(n3004), .B2(n3017), .ZN(n2206)
         );
  NAND2_X1 U2425 ( .A1(n2907), .A2(n2908), .ZN(n2207) );
  NAND2_X1 U2426 ( .A1(n2909), .A2(n2208), .ZN(n2204) );
  AND2_X1 U2427 ( .A1(n3417), .A2(n3007), .ZN(n3469) );
  NOR2_X1 U2428 ( .A1(n2828), .A2(n2947), .ZN(n2897) );
  NAND2_X1 U2429 ( .A1(n2824), .A2(n3507), .ZN(n2895) );
  NOR2_X1 U2430 ( .A1(n3730), .A2(n3716), .ZN(n4029) );
  NAND2_X1 U2431 ( .A1(n3744), .A2(n3731), .ZN(n3730) );
  AND2_X1 U2432 ( .A1(n3021), .A2(n3040), .ZN(n4012) );
  NAND2_X1 U2433 ( .A1(n2812), .A2(n4329), .ZN(n4354) );
  XNOR2_X1 U2434 ( .A(n2278), .B(n2277), .ZN(n2454) );
  NAND2_X1 U2435 ( .A1(n2276), .A2(IR_REG_31__SCAN_IN), .ZN(n2278) );
  INV_X1 U2436 ( .A(IR_REG_4__SCAN_IN), .ZN(n2138) );
  INV_X1 U2437 ( .A(n3577), .ZN(n2593) );
  OAI21_X1 U2438 ( .B1(n3436), .B2(n2367), .A(n2462), .ZN(n2573) );
  INV_X1 U2439 ( .A(n2478), .ZN(n2507) );
  INV_X1 U2440 ( .A(n3570), .ZN(n3017) );
  AND2_X1 U2441 ( .A1(n2456), .A2(n4304), .ZN(n3394) );
  OR2_X1 U2442 ( .A1(n2501), .A2(n4168), .ZN(n3407) );
  OR2_X1 U2443 ( .A1(n2501), .A2(n3579), .ZN(n3408) );
  INV_X1 U2444 ( .A(n3925), .ZN(n3890) );
  OR2_X1 U2445 ( .A1(n2789), .A2(n2788), .ZN(n3571) );
  NAND2_X1 U2446 ( .A1(n2176), .A2(n2177), .ZN(n2702) );
  NAND2_X1 U2447 ( .A1(n2459), .A2(REG0_REG_1__SCAN_IN), .ZN(n2062) );
  OR2_X1 U2448 ( .A1(n2416), .A2(n2415), .ZN(n3578) );
  NAND2_X1 U2449 ( .A1(n2111), .A2(n2348), .ZN(n3593) );
  OR2_X1 U2450 ( .A1(n3595), .A2(n3590), .ZN(n2111) );
  INV_X1 U2451 ( .A(n2077), .ZN(n2345) );
  OAI21_X1 U2452 ( .B1(n4195), .B2(n2546), .A(n2341), .ZN(n2077) );
  XNOR2_X1 U2453 ( .A(n2871), .B(n4222), .ZN(n4219) );
  NAND2_X1 U2454 ( .A1(n4219), .A2(REG2_REG_10__SCAN_IN), .ZN(n4218) );
  OAI21_X1 U2455 ( .B1(n4247), .B2(n2113), .A(n2112), .ZN(n4261) );
  NAND2_X1 U2456 ( .A1(n2114), .A2(REG2_REG_14__SCAN_IN), .ZN(n2113) );
  NAND2_X1 U2457 ( .A1(n3611), .A2(n2114), .ZN(n2112) );
  INV_X1 U2458 ( .A(n4262), .ZN(n2114) );
  NAND2_X1 U2459 ( .A1(n4270), .A2(n4271), .ZN(n4269) );
  OAI21_X1 U2460 ( .B1(n3635), .B2(n2120), .A(n2119), .ZN(n2118) );
  NAND2_X1 U2461 ( .A1(n2121), .A2(n4276), .ZN(n2120) );
  INV_X1 U2462 ( .A(n2074), .ZN(n3635) );
  INV_X1 U2463 ( .A(n2187), .ZN(n2186) );
  OR2_X1 U2464 ( .A1(n2582), .A2(n2487), .ZN(n4304) );
  NAND2_X1 U2465 ( .A1(n2175), .A2(n3258), .ZN(n2171) );
  INV_X1 U2466 ( .A(n3738), .ZN(n2057) );
  NAND2_X1 U2467 ( .A1(n2214), .A2(n2215), .ZN(n2213) );
  INV_X1 U2468 ( .A(n2216), .ZN(n2214) );
  NOR2_X1 U2469 ( .A1(n2322), .A2(IR_REG_27__SCAN_IN), .ZN(n2089) );
  OAI21_X1 U2470 ( .B1(n2284), .B2(n2082), .A(n2003), .ZN(n2088) );
  NAND2_X1 U2471 ( .A1(IR_REG_28__SCAN_IN), .A2(n2083), .ZN(n2082) );
  INV_X1 U2472 ( .A(n2089), .ZN(n2086) );
  INV_X1 U2473 ( .A(n2088), .ZN(n2087) );
  INV_X1 U2474 ( .A(n2464), .ZN(n3473) );
  OR2_X1 U2475 ( .A1(n3175), .A2(n3337), .ZN(n3186) );
  INV_X1 U2476 ( .A(IR_REG_18__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U2477 ( .A1(n3593), .A2(n2016), .ZN(n2110) );
  NAND2_X1 U2478 ( .A1(n2335), .A2(n2334), .ZN(n2340) );
  OAI21_X1 U2479 ( .B1(n2405), .B2(n2404), .A(n2023), .ZN(n2072) );
  AND2_X1 U2480 ( .A1(n2117), .A2(n2116), .ZN(n2886) );
  NAND2_X1 U2481 ( .A1(n2966), .A2(REG1_REG_11__SCAN_IN), .ZN(n2116) );
  AND3_X1 U2482 ( .A1(n2127), .A2(n2126), .A3(n2036), .ZN(n3627) );
  NAND2_X1 U2483 ( .A1(n4272), .A2(n2123), .ZN(n2122) );
  NAND2_X1 U2484 ( .A1(n4282), .A2(n4083), .ZN(n2123) );
  NAND2_X1 U2485 ( .A1(n2055), .A2(n2058), .ZN(n3663) );
  INV_X1 U2486 ( .A(n3660), .ZN(n2058) );
  NAND2_X1 U2487 ( .A1(n2060), .A2(n2056), .ZN(n2055) );
  NOR2_X1 U2488 ( .A1(n3658), .A2(n2057), .ZN(n2056) );
  NAND2_X1 U2489 ( .A1(n2064), .A2(n3655), .ZN(n3789) );
  INV_X1 U2490 ( .A(n3697), .ZN(n2141) );
  NAND2_X1 U2491 ( .A1(n3946), .A2(n2063), .ZN(n3810) );
  AND2_X1 U2492 ( .A1(n2065), .A2(n3652), .ZN(n2063) );
  AND2_X1 U2493 ( .A1(n3571), .A2(n2917), .ZN(n3517) );
  NAND2_X1 U2494 ( .A1(n2593), .A2(n2617), .ZN(n3493) );
  NAND2_X1 U2495 ( .A1(n3496), .A2(n3493), .ZN(n2591) );
  INV_X1 U2496 ( .A(n3815), .ZN(n3715) );
  AND2_X1 U2497 ( .A1(n2577), .A2(n2630), .ZN(n2096) );
  INV_X1 U2498 ( .A(n2616), .ZN(n2097) );
  XNOR2_X1 U2499 ( .A(n2464), .B(n3488), .ZN(n2482) );
  INV_X1 U2500 ( .A(IR_REG_27__SCAN_IN), .ZN(n2343) );
  AND2_X1 U2501 ( .A1(n2234), .A2(n2277), .ZN(n2238) );
  AND2_X1 U2502 ( .A1(n2251), .A2(n2225), .ZN(n2037) );
  OR3_X1 U2503 ( .A1(n2825), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2850) );
  AND2_X1 U2504 ( .A1(n2032), .A2(n3104), .ZN(n2170) );
  OAI22_X1 U2505 ( .A1(n2479), .A2(n3081), .B1(n2507), .B2(n2423), .ZN(n2494)
         );
  NAND2_X1 U2506 ( .A1(n2161), .A2(n2160), .ZN(n3343) );
  AOI21_X1 U2507 ( .B1(n2163), .B2(n2166), .A(n2027), .ZN(n2160) );
  AND2_X1 U2508 ( .A1(n3062), .A2(n3061), .ZN(n3360) );
  AND2_X1 U2509 ( .A1(n2969), .A2(n2968), .ZN(n3029) );
  AOI21_X1 U2510 ( .B1(n2943), .B2(n2154), .A(n2029), .ZN(n2151) );
  NAND2_X1 U2511 ( .A1(n2925), .A2(n2152), .ZN(n2040) );
  AND2_X1 U2512 ( .A1(n2159), .A2(n2674), .ZN(n2049) );
  INV_X1 U2513 ( .A(n2157), .ZN(n2048) );
  AOI21_X1 U2514 ( .B1(n2158), .B2(n2674), .A(n2223), .ZN(n2157) );
  AND3_X1 U2515 ( .A1(n2585), .A2(n2579), .A3(n2583), .ZN(n2457) );
  AND2_X1 U2516 ( .A1(n3156), .A2(n3155), .ZN(n3699) );
  AND4_X1 U2517 ( .A1(n2994), .A2(n2993), .A3(n2992), .A4(n2991), .ZN(n3677)
         );
  NOR2_X1 U2518 ( .A1(n3285), .A2(REG3_REG_3__SCAN_IN), .ZN(n2175) );
  OAI21_X1 U2519 ( .B1(n3282), .B2(n2305), .A(n2304), .ZN(n2173) );
  OAI21_X1 U2520 ( .B1(n2458), .B2(n2469), .A(n2051), .ZN(n2050) );
  NAND2_X1 U2521 ( .A1(n1999), .A2(REG2_REG_1__SCAN_IN), .ZN(n2051) );
  NAND2_X1 U2522 ( .A1(n2009), .A2(REG3_REG_0__SCAN_IN), .ZN(n2411) );
  AOI21_X1 U2523 ( .B1(n2395), .B2(REG2_REG_3__SCAN_IN), .A(n2109), .ZN(n2350)
         );
  AND2_X1 U2524 ( .A1(n2110), .A2(n2535), .ZN(n2109) );
  XNOR2_X1 U2525 ( .A(n2072), .B(n2881), .ZN(n2406) );
  NAND2_X1 U2526 ( .A1(n4175), .A2(REG2_REG_7__SCAN_IN), .ZN(n2107) );
  NAND2_X1 U2527 ( .A1(n2880), .A2(n2071), .ZN(n2882) );
  OR2_X1 U2528 ( .A1(n2072), .A2(n2881), .ZN(n2071) );
  NOR2_X1 U2529 ( .A1(n4204), .A2(n2124), .ZN(n2884) );
  AND2_X1 U2530 ( .A1(n2883), .A2(REG1_REG_9__SCAN_IN), .ZN(n2124) );
  OR2_X1 U2531 ( .A1(n4225), .A2(n4224), .ZN(n2117) );
  XNOR2_X1 U2532 ( .A(n2886), .B(n4318), .ZN(n4234) );
  NAND2_X1 U2533 ( .A1(n4273), .A2(n4274), .ZN(n4272) );
  NAND2_X1 U2534 ( .A1(n2122), .A2(n3630), .ZN(n2121) );
  OR2_X1 U2535 ( .A1(n2122), .A2(n3630), .ZN(n2074) );
  NOR2_X1 U2536 ( .A1(n2190), .A2(n2184), .ZN(n2183) );
  INV_X1 U2537 ( .A(n3705), .ZN(n2184) );
  NAND2_X1 U2538 ( .A1(n3720), .A2(n2192), .ZN(n2190) );
  OAI21_X1 U2539 ( .B1(n2188), .B2(n3722), .A(n2196), .ZN(n2187) );
  OR2_X1 U2540 ( .A1(n3743), .A2(n3731), .ZN(n2196) );
  NAND2_X1 U2541 ( .A1(n2189), .A2(n2192), .ZN(n2188) );
  INV_X1 U2542 ( .A(n2193), .ZN(n2189) );
  AND2_X1 U2543 ( .A1(n3648), .A2(n3221), .ZN(n3732) );
  INV_X1 U2544 ( .A(n3663), .ZN(n3723) );
  AND2_X1 U2545 ( .A1(n2060), .A2(n2059), .ZN(n3739) );
  NOR2_X1 U2546 ( .A1(n3148), .A2(n3374), .ZN(n3162) );
  NAND2_X1 U2547 ( .A1(n3162), .A2(REG3_REG_23__SCAN_IN), .ZN(n3175) );
  AND2_X1 U2548 ( .A1(n3812), .A2(n3478), .ZN(n3830) );
  AND4_X1 U2549 ( .A1(n3143), .A2(n3142), .A3(n3141), .A4(n3140), .ZN(n3859)
         );
  NAND2_X1 U2550 ( .A1(n3127), .A2(REG3_REG_20__SCAN_IN), .ZN(n3138) );
  AND4_X1 U2551 ( .A1(n3132), .A2(n3131), .A3(n3130), .A4(n3129), .ZN(n3888)
         );
  NOR2_X1 U2552 ( .A1(n3106), .A2(n4511), .ZN(n3107) );
  OR2_X1 U2553 ( .A1(n3091), .A2(n3090), .ZN(n3106) );
  NAND2_X1 U2554 ( .A1(n3946), .A2(n3652), .ZN(n3924) );
  NAND2_X1 U2555 ( .A1(n3958), .A2(n3651), .ZN(n3948) );
  OR2_X1 U2556 ( .A1(n3986), .A2(n3713), .ZN(n3964) );
  NAND2_X1 U2557 ( .A1(n3682), .A2(n2136), .ZN(n2132) );
  INV_X1 U2558 ( .A(n2134), .ZN(n2133) );
  NAND2_X1 U2559 ( .A1(n3940), .A2(n3939), .ZN(n3938) );
  OR2_X1 U2560 ( .A1(n3046), .A2(n3045), .ZN(n3048) );
  INV_X1 U2561 ( .A(n3713), .ZN(n3965) );
  NAND2_X1 U2562 ( .A1(n2053), .A2(n2052), .ZN(n3958) );
  INV_X1 U2563 ( .A(n3970), .ZN(n2052) );
  INV_X1 U2564 ( .A(n3960), .ZN(n2053) );
  NAND2_X1 U2565 ( .A1(n3421), .A2(n3524), .ZN(n3978) );
  NAND2_X1 U2566 ( .A1(n2984), .A2(n3520), .ZN(n3415) );
  NAND2_X1 U2567 ( .A1(n2983), .A2(n3512), .ZN(n2984) );
  INV_X1 U2568 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2947) );
  NAND2_X1 U2569 ( .A1(n2721), .A2(REG3_REG_8__SCAN_IN), .ZN(n2783) );
  OAI21_X1 U2570 ( .B1(n2797), .B2(n2796), .A(n3508), .ZN(n2823) );
  OR2_X1 U2571 ( .A1(n2506), .A2(n3552), .ZN(n4001) );
  NAND2_X1 U2572 ( .A1(n2069), .A2(n3504), .ZN(n2797) );
  NAND2_X1 U2573 ( .A1(n2755), .A2(n3515), .ZN(n2069) );
  AND2_X1 U2574 ( .A1(n3505), .A2(n3508), .ZN(n3468) );
  AND2_X1 U2575 ( .A1(n2481), .A2(n3556), .ZN(n4010) );
  AND2_X1 U2576 ( .A1(n4168), .A2(n2474), .ZN(n4006) );
  OAI21_X1 U2577 ( .B1(n2700), .B2(n2637), .A(n3502), .ZN(n2739) );
  NAND2_X1 U2578 ( .A1(n2181), .A2(n2697), .ZN(n2699) );
  INV_X1 U2579 ( .A(n2696), .ZN(n2181) );
  INV_X1 U2580 ( .A(n2701), .ZN(n2709) );
  NAND2_X1 U2581 ( .A1(n2068), .A2(n3498), .ZN(n2700) );
  NAND2_X1 U2582 ( .A1(n2636), .A2(n3471), .ZN(n2068) );
  AND2_X1 U2583 ( .A1(n3498), .A2(n3495), .ZN(n3471) );
  INV_X1 U2584 ( .A(n4006), .ZN(n3954) );
  OR2_X1 U2585 ( .A1(n3488), .A2(n2464), .ZN(n2590) );
  INV_X1 U2586 ( .A(n2591), .ZN(n3472) );
  AND2_X1 U2587 ( .A1(n3805), .A2(n2035), .ZN(n3744) );
  NAND2_X1 U2588 ( .A1(n3805), .A2(n2098), .ZN(n3762) );
  NAND2_X1 U2589 ( .A1(n3805), .A2(n2007), .ZN(n3781) );
  AND2_X1 U2590 ( .A1(n3805), .A2(n3797), .ZN(n3799) );
  NOR2_X1 U2591 ( .A1(n4061), .A2(n3715), .ZN(n3805) );
  OR2_X1 U2592 ( .A1(n2001), .A2(n3836), .ZN(n4061) );
  NOR2_X1 U2593 ( .A1(n3932), .A2(n2005), .ZN(n3872) );
  NOR3_X1 U2594 ( .A1(n3932), .A2(n3714), .A3(n3911), .ZN(n3893) );
  NOR2_X1 U2595 ( .A1(n3964), .A2(n3942), .ZN(n3941) );
  NAND2_X1 U2596 ( .A1(n3941), .A2(n3930), .ZN(n3932) );
  OR2_X1 U2597 ( .A1(n4014), .A2(n3984), .ZN(n3986) );
  NAND2_X1 U2598 ( .A1(n4012), .A2(n4011), .ZN(n4014) );
  AND2_X1 U2599 ( .A1(n2805), .A2(n2031), .ZN(n3021) );
  NAND2_X1 U2600 ( .A1(n2805), .A2(n2100), .ZN(n3020) );
  NAND2_X1 U2601 ( .A1(n2805), .A2(n2101), .ZN(n2910) );
  NOR2_X1 U2602 ( .A1(n2760), .A2(n2802), .ZN(n2805) );
  AND2_X1 U2603 ( .A1(n2805), .A2(n2841), .ZN(n2838) );
  OR2_X1 U2604 ( .A1(n2745), .A2(n2766), .ZN(n2760) );
  NAND2_X1 U2605 ( .A1(n2097), .A2(n2577), .ZN(n2614) );
  AND3_X1 U2606 ( .A1(n2491), .A2(n2490), .A3(n2489), .ZN(n2613) );
  XNOR2_X1 U2607 ( .A(n2272), .B(n2215), .ZN(n2455) );
  NOR2_X1 U2608 ( .A1(n2850), .A2(IR_REG_9__SCAN_IN), .ZN(n2866) );
  NAND2_X1 U2609 ( .A1(n3436), .A2(DATAI_23_), .ZN(n3815) );
  AND4_X1 U2610 ( .A1(n2902), .A2(n2901), .A3(n2900), .A4(n2899), .ZN(n3008)
         );
  NAND2_X1 U2611 ( .A1(n2162), .A2(n2168), .ZN(n3249) );
  NAND2_X1 U2612 ( .A1(n3325), .A2(n2170), .ZN(n2162) );
  XNOR2_X1 U2613 ( .A(n2511), .B(n2500), .ZN(n2513) );
  NAND2_X1 U2614 ( .A1(n3342), .A2(n3346), .ZN(n3296) );
  INV_X1 U2615 ( .A(n2045), .ZN(n2044) );
  OAI21_X1 U2616 ( .B1(n2022), .B2(n3158), .A(n2217), .ZN(n2045) );
  AOI22_X1 U2617 ( .A1(n3182), .A2(n3335), .B1(n3184), .B2(n3185), .ZN(n2217)
         );
  AND4_X1 U2618 ( .A1(n2550), .A2(n2549), .A3(n2548), .A4(n2547), .ZN(n2658)
         );
  NAND2_X1 U2619 ( .A1(n2656), .A2(n2655), .ZN(n2675) );
  AND4_X1 U2620 ( .A1(n3113), .A2(n3112), .A3(n3111), .A4(n3110), .ZN(n3925)
         );
  INV_X1 U2621 ( .A(n3792), .ZN(n3797) );
  NAND2_X1 U2622 ( .A1(n2159), .A2(n2561), .ZN(n2656) );
  AND4_X1 U2623 ( .A1(n2726), .A2(n2725), .A3(n2724), .A4(n2723), .ZN(n2929)
         );
  AND2_X1 U2624 ( .A1(n2156), .A2(n2155), .ZN(n2926) );
  INV_X1 U2625 ( .A(n2923), .ZN(n2156) );
  INV_X1 U2626 ( .A(n3836), .ZN(n3698) );
  AND4_X1 U2627 ( .A1(n3096), .A2(n3095), .A3(n3094), .A4(n3093), .ZN(n3950)
         );
  NAND2_X1 U2628 ( .A1(n2167), .A2(n3104), .ZN(n3381) );
  OR2_X1 U2629 ( .A1(n3325), .A2(n3105), .ZN(n2167) );
  AND4_X1 U2630 ( .A1(n2568), .A2(n2567), .A3(n2566), .A4(n2565), .ZN(n2732)
         );
  AND4_X1 U2631 ( .A1(n2691), .A2(n2690), .A3(n2689), .A4(n2688), .ZN(n2799)
         );
  NAND2_X1 U2632 ( .A1(n2534), .A2(n2533), .ZN(n3397) );
  AND2_X1 U2633 ( .A1(n3258), .A2(n2445), .ZN(n3560) );
  INV_X1 U2634 ( .A(n3759), .ZN(n3726) );
  INV_X1 U2635 ( .A(n3816), .ZN(n3774) );
  INV_X1 U2636 ( .A(n3699), .ZN(n3846) );
  INV_X1 U2637 ( .A(n3888), .ZN(n3568) );
  INV_X1 U2638 ( .A(n3950), .ZN(n3688) );
  OR2_X1 U2639 ( .A1(n2318), .A2(n2317), .ZN(n3683) );
  INV_X1 U2640 ( .A(n3677), .ZN(n3981) );
  OR2_X1 U2641 ( .A1(n2979), .A2(n2978), .ZN(n4005) );
  OR2_X1 U2642 ( .A1(n2833), .A2(n2832), .ZN(n3570) );
  INV_X1 U2643 ( .A(n2929), .ZN(n3572) );
  OR2_X1 U2644 ( .A1(n2643), .A2(n2642), .ZN(n3574) );
  INV_X1 U2645 ( .A(n2732), .ZN(n3575) );
  INV_X1 U2646 ( .A(n2658), .ZN(n3576) );
  NAND2_X1 U2647 ( .A1(n2473), .A2(n2010), .ZN(n3577) );
  NAND2_X1 U2648 ( .A1(n2091), .A2(n2131), .ZN(n2130) );
  XNOR2_X1 U2649 ( .A(n2367), .B(REG1_REG_1__SCAN_IN), .ZN(n2360) );
  NOR3_X2 U2650 ( .A1(n2361), .A2(n2347), .A3(n2038), .ZN(n3595) );
  AOI21_X1 U2651 ( .B1(n2387), .B2(REG2_REG_6__SCAN_IN), .A(n2034), .ZN(n2389)
         );
  OR2_X1 U2652 ( .A1(n2406), .A2(n2818), .ZN(n2880) );
  AND2_X1 U2653 ( .A1(n2882), .A2(n2125), .ZN(n4204) );
  INV_X1 U2654 ( .A(n4205), .ZN(n2125) );
  INV_X1 U2655 ( .A(n2882), .ZN(n4206) );
  XNOR2_X1 U2656 ( .A(n2884), .B(n4222), .ZN(n4215) );
  NAND2_X1 U2657 ( .A1(n4218), .A2(n2872), .ZN(n4229) );
  INV_X1 U2658 ( .A(n2117), .ZN(n4223) );
  INV_X1 U2659 ( .A(n2076), .ZN(n2891) );
  XNOR2_X1 U2660 ( .A(n2115), .B(n4251), .ZN(n4247) );
  NOR2_X1 U2661 ( .A1(n4247), .A2(n4248), .ZN(n4246) );
  NAND2_X1 U2662 ( .A1(n2127), .A2(n2126), .ZN(n4257) );
  NAND2_X1 U2663 ( .A1(n3621), .A2(n3622), .ZN(n4270) );
  AOI21_X1 U2664 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4172), .A(n3638), .ZN(n3640) );
  AND2_X1 U2665 ( .A1(n2074), .A2(n2073), .ZN(n3637) );
  NAND2_X1 U2666 ( .A1(n4172), .A2(REG1_REG_18__SCAN_IN), .ZN(n2073) );
  NAND2_X1 U2667 ( .A1(n2185), .A2(n2192), .ZN(n3721) );
  NAND2_X1 U2668 ( .A1(n2198), .A2(n2193), .ZN(n2185) );
  AND2_X1 U2669 ( .A1(n3209), .A2(n3220), .ZN(n3746) );
  INV_X1 U2670 ( .A(n2194), .ZN(n2191) );
  OAI21_X1 U2671 ( .B1(n3902), .B2(n2145), .A(n2142), .ZN(n3851) );
  NAND2_X1 U2672 ( .A1(n2148), .A2(n3692), .ZN(n3870) );
  NAND2_X1 U2673 ( .A1(n3902), .A2(n2149), .ZN(n2148) );
  NAND2_X1 U2674 ( .A1(n3902), .A2(n3691), .ZN(n3882) );
  NAND2_X1 U2675 ( .A1(n3975), .A2(n3682), .ZN(n3971) );
  NAND2_X1 U2676 ( .A1(n2204), .A2(n2201), .ZN(n3013) );
  NAND2_X1 U2677 ( .A1(n2204), .A2(n2205), .ZN(n3011) );
  OAI21_X1 U2678 ( .B1(n2909), .B2(n2908), .A(n2907), .ZN(n3006) );
  AND2_X1 U2679 ( .A1(n4284), .A2(n2626), .ZN(n3972) );
  OR2_X1 U2680 ( .A1(n2464), .A2(n2465), .ZN(n2466) );
  NAND2_X1 U2681 ( .A1(n2508), .A2(n2033), .ZN(n4300) );
  INV_X1 U2682 ( .A(n4369), .ZN(n4367) );
  INV_X1 U2683 ( .A(n4036), .ZN(n2081) );
  INV_X1 U2684 ( .A(n4035), .ZN(n2080) );
  AND2_X2 U2685 ( .A1(n2613), .A2(n2612), .ZN(n4362) );
  INV_X1 U2686 ( .A(n3579), .ZN(n4168) );
  NAND2_X1 U2687 ( .A1(n2244), .A2(IR_REG_31__SCAN_IN), .ZN(n2233) );
  INV_X1 U2688 ( .A(n2454), .ZN(n3562) );
  XNOR2_X1 U2689 ( .A(n2441), .B(IR_REG_19__SCAN_IN), .ZN(n4171) );
  INV_X1 U2690 ( .A(n2247), .ZN(n2137) );
  XNOR2_X1 U2691 ( .A(n2339), .B(IR_REG_4__SCAN_IN), .ZN(n4201) );
  NAND2_X1 U2692 ( .A1(n2327), .A2(IR_REG_31__SCAN_IN), .ZN(n2330) );
  OAI22_X1 U2693 ( .A1(n3407), .A2(n2463), .B1(n3394), .B2(n2507), .ZN(n2460)
         );
  OAI22_X1 U2694 ( .A1(n3408), .A2(n2463), .B1(n3394), .B2(n2577), .ZN(n2526)
         );
  INV_X1 U2695 ( .A(n2118), .ZN(n3632) );
  OR3_X1 U2696 ( .A1(n3932), .A2(n2005), .A3(n3845), .ZN(n2001) );
  AND2_X1 U2697 ( .A1(n2945), .A2(n2942), .ZN(n2943) );
  NAND2_X1 U2698 ( .A1(n2137), .A2(n2020), .ZN(n2250) );
  AND2_X1 U2699 ( .A1(n2732), .A2(n2731), .ZN(n2002) );
  INV_X1 U2700 ( .A(IR_REG_14__SCAN_IN), .ZN(n2231) );
  AND2_X1 U2701 ( .A1(n2018), .A2(n2090), .ZN(n2003) );
  AND2_X1 U2702 ( .A1(n2146), .A2(n3697), .ZN(n2004) );
  OR3_X1 U2703 ( .A1(n3714), .A2(n3911), .A3(n3452), .ZN(n2005) );
  AND2_X1 U2704 ( .A1(n2097), .A2(n2096), .ZN(n2006) );
  AND2_X1 U2705 ( .A1(n3797), .A2(n3779), .ZN(n2007) );
  INV_X1 U2706 ( .A(n2423), .ZN(n3120) );
  NAND2_X1 U2707 ( .A1(n2530), .A2(n2418), .ZN(n2422) );
  OR2_X1 U2708 ( .A1(n3601), .A2(n4317), .ZN(n2008) );
  NAND2_X1 U2709 ( .A1(n2042), .A2(n2093), .ZN(n2284) );
  AND2_X1 U2710 ( .A1(n2303), .A2(n2301), .ZN(n2009) );
  AND3_X1 U2711 ( .A1(n2472), .A2(n2471), .A3(n2470), .ZN(n2010) );
  OR2_X1 U2712 ( .A1(n3775), .A2(n3760), .ZN(n2011) );
  AND2_X1 U2713 ( .A1(n3434), .A2(REG0_REG_3__SCAN_IN), .ZN(n2012) );
  AND2_X1 U2714 ( .A1(n3726), .A2(n3745), .ZN(n2013) );
  AND2_X1 U2715 ( .A1(n2009), .A2(REG3_REG_1__SCAN_IN), .ZN(n2014) );
  NOR2_X1 U2716 ( .A1(n4246), .A2(n3611), .ZN(n2015) );
  NAND2_X1 U2717 ( .A1(n2093), .A2(n2210), .ZN(n2265) );
  INV_X1 U2718 ( .A(n3658), .ZN(n2059) );
  OR2_X1 U2719 ( .A1(n3587), .A2(n2349), .ZN(n2016) );
  OR2_X1 U2720 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2017)
         );
  INV_X1 U2721 ( .A(n2202), .ZN(n2201) );
  NAND2_X1 U2722 ( .A1(n2205), .A2(n2203), .ZN(n2202) );
  INV_X1 U2723 ( .A(n3720), .ZN(n3722) );
  NAND2_X1 U2724 ( .A1(n2326), .A2(n2225), .ZN(n2247) );
  NAND2_X1 U2725 ( .A1(n2092), .A2(IR_REG_27__SCAN_IN), .ZN(n2018) );
  INV_X1 U2726 ( .A(IR_REG_26__SCAN_IN), .ZN(n2083) );
  AND3_X1 U2727 ( .A1(n2092), .A2(n2083), .A3(n2343), .ZN(n2019) );
  AND2_X1 U2728 ( .A1(n2336), .A2(n2138), .ZN(n2020) );
  AND2_X1 U2729 ( .A1(n2129), .A2(n2008), .ZN(n2021) );
  INV_X1 U2730 ( .A(IR_REG_28__SCAN_IN), .ZN(n2092) );
  XNOR2_X1 U2731 ( .A(n2233), .B(IR_REG_24__SCAN_IN), .ZN(n2281) );
  AND2_X1 U2732 ( .A1(n2255), .A2(n2230), .ZN(n2855) );
  NAND2_X1 U2733 ( .A1(n2925), .A2(n2924), .ZN(n2155) );
  NAND2_X1 U2734 ( .A1(n2855), .A2(n2231), .ZN(n3054) );
  NAND2_X1 U2735 ( .A1(n3172), .A2(n2218), .ZN(n2022) );
  AND2_X1 U2736 ( .A1(n2210), .A2(n2855), .ZN(n3099) );
  OR2_X1 U2737 ( .A1(n4175), .A2(REG1_REG_7__SCAN_IN), .ZN(n2023) );
  OAI21_X1 U2738 ( .B1(n2909), .B2(n2202), .A(n2199), .ZN(n3676) );
  OR2_X1 U2739 ( .A1(n3704), .A2(n3779), .ZN(n2024) );
  INV_X1 U2740 ( .A(n3692), .ZN(n2147) );
  INV_X1 U2741 ( .A(n3014), .ZN(n3023) );
  INV_X1 U2742 ( .A(IR_REG_21__SCAN_IN), .ZN(n2215) );
  NAND2_X1 U2743 ( .A1(n3976), .A2(n3977), .ZN(n3975) );
  OR2_X1 U2744 ( .A1(n4323), .A2(n4484), .ZN(n2025) );
  INV_X1 U2745 ( .A(n2099), .ZN(n3904) );
  NOR2_X1 U2746 ( .A1(n3932), .A2(n3911), .ZN(n2099) );
  AND2_X1 U2747 ( .A1(n3008), .A2(n3023), .ZN(n2026) );
  NOR2_X1 U2748 ( .A1(n3126), .A2(n3125), .ZN(n2027) );
  NAND2_X1 U2749 ( .A1(n3859), .A2(n3852), .ZN(n2028) );
  INV_X1 U2750 ( .A(n2146), .ZN(n2145) );
  NOR2_X1 U2751 ( .A1(n3695), .A2(n2147), .ZN(n2146) );
  INV_X1 U2752 ( .A(n3682), .ZN(n2135) );
  OAI21_X1 U2753 ( .B1(n2142), .B2(n2141), .A(n2028), .ZN(n2140) );
  AND2_X1 U2754 ( .A1(n2962), .A2(n2964), .ZN(n2029) );
  OR2_X1 U2755 ( .A1(n3863), .A2(n3423), .ZN(n3653) );
  INV_X1 U2756 ( .A(n3653), .ZN(n2065) );
  AND2_X1 U2757 ( .A1(n2096), .A2(n2731), .ZN(n2030) );
  AND2_X1 U2758 ( .A1(n2100), .A2(n3023), .ZN(n2031) );
  INV_X1 U2759 ( .A(n3684), .ZN(n2136) );
  NAND2_X1 U2760 ( .A1(n3502), .A2(n3499), .ZN(n2697) );
  INV_X1 U2761 ( .A(n2697), .ZN(n2179) );
  XNOR2_X1 U2762 ( .A(n2237), .B(IR_REG_26__SCAN_IN), .ZN(n4169) );
  NAND2_X1 U2763 ( .A1(n2699), .A2(n2634), .ZN(n2733) );
  NAND2_X1 U2764 ( .A1(n2855), .A2(n2212), .ZN(n3097) );
  INV_X1 U2765 ( .A(n3845), .ZN(n3852) );
  AND2_X1 U2766 ( .A1(n3436), .A2(DATAI_21_), .ZN(n3845) );
  INV_X1 U2767 ( .A(IR_REG_31__SCAN_IN), .ZN(n2091) );
  NAND2_X1 U2768 ( .A1(n3116), .A2(n3117), .ZN(n2032) );
  OR2_X1 U2769 ( .A1(n4002), .A2(n2463), .ZN(n2033) );
  AND2_X1 U2770 ( .A1(n2386), .A2(n2676), .ZN(n2034) );
  OAI21_X1 U2771 ( .B1(n2284), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2322) );
  AND2_X1 U2772 ( .A1(n2098), .A2(n3708), .ZN(n2035) );
  INV_X1 U2773 ( .A(n2095), .ZN(n2708) );
  INV_X1 U2774 ( .A(n3706), .ZN(n3760) );
  NAND2_X1 U2775 ( .A1(n4315), .A2(REG1_REG_15__SCAN_IN), .ZN(n2036) );
  INV_X1 U2776 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2103) );
  INV_X1 U2777 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2106) );
  AOI21_X1 U2778 ( .B1(n4268), .B2(ADDR_REG_18__SCAN_IN), .A(n3631), .ZN(n2119) );
  AND3_X2 U2779 ( .A1(n2020), .A2(n2326), .A3(n2037), .ZN(n2255) );
  AND2_X2 U2780 ( .A1(n2038), .A2(n2131), .ZN(n2326) );
  AOI21_X2 U2781 ( .B1(n3031), .B2(n3030), .A(n3029), .ZN(n3355) );
  NAND2_X1 U2782 ( .A1(n2923), .A2(n2943), .ZN(n2039) );
  AOI21_X1 U2783 ( .B1(n3307), .B2(n3303), .A(n3305), .ZN(n3387) );
  NOR2_X1 U2784 ( .A1(n2046), .A2(n3083), .ZN(n3315) );
  NAND2_X1 U2785 ( .A1(n3066), .A2(n3065), .ZN(n2047) );
  NOR2_X1 U2786 ( .A1(n2014), .A2(n2050), .ZN(n2061) );
  OR2_X1 U2787 ( .A1(n2303), .A2(n2302), .ZN(n2469) );
  NAND2_X1 U2788 ( .A1(n3810), .A2(n3654), .ZN(n2064) );
  OAI22_X1 U2789 ( .A1(n4195), .A2(n2078), .B1(n2079), .B2(n2341), .ZN(n2369)
         );
  NOR2_X1 U2790 ( .A1(n4214), .A2(n2885), .ZN(n4225) );
  OAI211_X2 U2791 ( .C1(n2325), .C2(n2131), .A(n2327), .B(n2130), .ZN(n2367)
         );
  OAI211_X1 U2792 ( .C1(n4093), .C2(n2081), .A(n2080), .B(n4037), .ZN(n4116)
         );
  AOI21_X1 U2793 ( .B1(n3716), .B2(n3730), .A(n4029), .ZN(n4036) );
  NAND3_X1 U2794 ( .A1(n2087), .A2(n2086), .A3(IR_REG_0__SCAN_IN), .ZN(n2085)
         );
  AND2_X2 U2795 ( .A1(n2094), .A2(n2255), .ZN(n2093) );
  NAND3_X1 U2796 ( .A1(n2097), .A2(n2709), .A3(n2096), .ZN(n2095) );
  NAND3_X1 U2797 ( .A1(n2097), .A2(n2709), .A3(n2030), .ZN(n2745) );
  AOI22_X1 U2798 ( .A1(n2387), .A2(n2105), .B1(n2386), .B2(n2104), .ZN(n2108)
         );
  INV_X1 U2799 ( .A(n2108), .ZN(n2401) );
  INV_X1 U2800 ( .A(n3610), .ZN(n2115) );
  AOI21_X2 U2801 ( .B1(REG2_REG_5__SCAN_IN), .B2(n2371), .A(n2370), .ZN(n2385)
         );
  INV_X1 U2802 ( .A(n2129), .ZN(n4242) );
  OAI22_X1 U2803 ( .A1(n3976), .A2(n2132), .B1(n3684), .B2(n2133), .ZN(n3940)
         );
  NAND2_X1 U2804 ( .A1(n2944), .A2(n2943), .ZN(n2965) );
  NAND2_X1 U2805 ( .A1(n2153), .A2(n2155), .ZN(n2944) );
  NAND2_X1 U2806 ( .A1(n3325), .A2(n2163), .ZN(n2161) );
  NOR2_X1 U2807 ( .A1(n2173), .A2(n2012), .ZN(n2176) );
  NAND4_X1 U2808 ( .A1(n2174), .A2(n2536), .A3(n2172), .A4(n2171), .ZN(n2537)
         );
  INV_X1 U2809 ( .A(n2175), .ZN(n2177) );
  NAND2_X1 U2810 ( .A1(n2696), .A2(n2634), .ZN(n2180) );
  NAND2_X1 U2811 ( .A1(n2180), .A2(n2178), .ZN(n2736) );
  NAND2_X1 U2812 ( .A1(n3768), .A2(n2183), .ZN(n2182) );
  NAND2_X1 U2813 ( .A1(n2182), .A2(n2186), .ZN(n3711) );
  AND2_X1 U2814 ( .A1(n2198), .A2(n2024), .ZN(n3751) );
  NAND2_X1 U2815 ( .A1(n2198), .A2(n2191), .ZN(n2197) );
  NAND2_X1 U2816 ( .A1(n3489), .A2(n2589), .ZN(n2464) );
  OR2_X1 U2817 ( .A1(n2265), .A2(n2216), .ZN(n2271) );
  NOR2_X1 U2818 ( .A1(n2265), .A2(n2213), .ZN(n2275) );
  AND2_X2 U2819 ( .A1(n3240), .A2(n3172), .ZN(n3239) );
  NAND2_X1 U2820 ( .A1(n3436), .A2(DATAI_1_), .ZN(n2462) );
  OR2_X1 U2821 ( .A1(n3282), .A2(n4051), .ZN(n3188) );
  NAND2_X1 U2822 ( .A1(n2009), .A2(REG3_REG_2__SCAN_IN), .ZN(n2471) );
  AND2_X1 U2823 ( .A1(n3919), .A2(n4356), .ZN(n4294) );
  AOI21_X2 U2824 ( .B1(n2717), .B2(n2716), .A(n2715), .ZN(n2720) );
  NAND2_X1 U2825 ( .A1(n2275), .A2(n2277), .ZN(n2232) );
  NAND2_X1 U2826 ( .A1(n2519), .A2(n2518), .ZN(n2520) );
  AOI21_X2 U2827 ( .B1(n3808), .B2(n3701), .A(n2221), .ZN(n3787) );
  INV_X1 U2828 ( .A(n3258), .ZN(n3216) );
  AND4_X1 U2829 ( .A1(n3052), .A2(n3051), .A3(n3050), .A4(n3049), .ZN(n4003)
         );
  OAI211_X1 U2830 ( .C1(n3308), .C2(n3285), .A(n3189), .B(n3188), .ZN(n3793)
         );
  INV_X1 U2831 ( .A(n3793), .ZN(n3704) );
  OR2_X1 U2832 ( .A1(n3699), .A2(n3698), .ZN(n2220) );
  AND2_X1 U2833 ( .A1(n3831), .A2(n3715), .ZN(n2221) );
  AND2_X1 U2834 ( .A1(n3268), .A2(n3267), .ZN(n2222) );
  AND2_X1 U2835 ( .A1(n2673), .A2(n2672), .ZN(n2223) );
  NAND2_X1 U2836 ( .A1(n2517), .A2(n2516), .ZN(n2538) );
  INV_X1 U2837 ( .A(n3468), .ZN(n2769) );
  INV_X1 U2838 ( .A(IR_REG_2__SCAN_IN), .ZN(n2225) );
  AND2_X1 U2839 ( .A1(n3809), .A2(n3541), .ZN(n3654) );
  INV_X1 U2840 ( .A(n3185), .ZN(n3180) );
  OAI22_X1 U2841 ( .A1(n2593), .A2(n3204), .B1(n2577), .B2(n2423), .ZN(n2515)
         );
  AND2_X1 U2842 ( .A1(n3454), .A2(n3788), .ZN(n3656) );
  NAND2_X1 U2843 ( .A1(n3087), .A2(n3086), .ZN(n3088) );
  INV_X1 U2844 ( .A(n3984), .ZN(n3681) );
  AND2_X1 U2845 ( .A1(n3107), .A2(REG3_REG_19__SCAN_IN), .ZN(n3127) );
  INV_X1 U2846 ( .A(n3372), .ZN(n3158) );
  OR2_X1 U2847 ( .A1(n3138), .A2(n3297), .ZN(n3148) );
  OR2_X1 U2848 ( .A1(n3890), .A2(n3911), .ZN(n3691) );
  NAND2_X1 U2849 ( .A1(n4003), .A2(n3681), .ZN(n3682) );
  AND2_X1 U2850 ( .A1(n3448), .A2(n3447), .ZN(n3710) );
  INV_X1 U2851 ( .A(n2931), .ZN(n2917) );
  AND2_X1 U2852 ( .A1(n3579), .A2(n2474), .ZN(n3912) );
  INV_X1 U2853 ( .A(n2510), .ZN(n2500) );
  INV_X1 U2854 ( .A(n3942), .ZN(n3949) );
  INV_X1 U2855 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2782) );
  INV_X1 U2856 ( .A(n3831), .ZN(n3700) );
  INV_X1 U2857 ( .A(n2799), .ZN(n4370) );
  INV_X1 U2858 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2988) );
  OR2_X1 U2859 ( .A1(n3661), .A2(n3481), .ZN(n3720) );
  INV_X1 U2860 ( .A(n3745), .ZN(n3708) );
  AND2_X1 U2861 ( .A1(n3979), .A2(n3965), .ZN(n3684) );
  NAND2_X1 U2862 ( .A1(n2576), .A2(n2591), .ZN(n2601) );
  AND2_X1 U2863 ( .A1(n2242), .A2(n2436), .ZN(n2437) );
  AND2_X1 U2864 ( .A1(n3436), .A2(DATAI_27_), .ZN(n3745) );
  INV_X1 U2865 ( .A(n3673), .ZN(n3040) );
  INV_X1 U2866 ( .A(n3912), .ZN(n4002) );
  AND2_X1 U2867 ( .A1(n2293), .A2(n4169), .ZN(n2440) );
  NOR2_X1 U2868 ( .A1(n2685), .A2(n2307), .ZN(n2721) );
  AND2_X1 U2869 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2564) );
  OR2_X1 U2870 ( .A1(n2783), .A2(n2782), .ZN(n2828) );
  OR2_X1 U2871 ( .A1(n2989), .A2(n2988), .ZN(n3046) );
  AND2_X1 U2872 ( .A1(n2897), .A2(REG3_REG_11__SCAN_IN), .ZN(n2974) );
  NAND2_X1 U2873 ( .A1(n2564), .A2(REG3_REG_5__SCAN_IN), .ZN(n2685) );
  OR2_X1 U2874 ( .A1(n3195), .A2(n3208), .ZN(n3392) );
  AND4_X1 U2875 ( .A1(n3076), .A2(n3075), .A3(n3074), .A4(n3073), .ZN(n3957)
         );
  INV_X1 U2876 ( .A(n4245), .ZN(n4278) );
  INV_X1 U2877 ( .A(n4001), .ZN(n4031) );
  INV_X1 U2878 ( .A(n3830), .ZN(n3826) );
  OR2_X1 U2879 ( .A1(n2312), .A2(n2311), .ZN(n3913) );
  AND2_X1 U2880 ( .A1(n4284), .A2(n3643), .ZN(n3919) );
  INV_X1 U2881 ( .A(n4010), .ZN(n3945) );
  AOI21_X1 U2882 ( .B1(n2440), .B2(n2438), .A(n2437), .ZN(n2579) );
  AND2_X1 U2883 ( .A1(n2417), .A2(n3552), .ZN(n4356) );
  AND2_X1 U2884 ( .A1(n4299), .A2(n2454), .ZN(n4339) );
  AND2_X1 U2885 ( .A1(n2864), .A2(n2863), .ZN(n2966) );
  NAND2_X1 U2886 ( .A1(n2457), .A2(n2443), .ZN(n3399) );
  NAND2_X1 U2887 ( .A1(n3226), .A2(n3225), .ZN(n3669) );
  OR2_X1 U2888 ( .A1(n3167), .A2(n3166), .ZN(n3831) );
  INV_X1 U2889 ( .A(n4003), .ZN(n3963) );
  OR2_X1 U2890 ( .A1(n4188), .A2(n3559), .ZN(n4245) );
  OR2_X1 U2891 ( .A1(n4188), .A2(n4168), .ZN(n4281) );
  OR2_X1 U2892 ( .A1(n4188), .A2(n4186), .ZN(n4256) );
  INV_X1 U2893 ( .A(n4294), .ZN(n4015) );
  NAND2_X1 U2894 ( .A1(n4369), .A2(n4356), .ZN(n4110) );
  AND2_X2 U2895 ( .A1(n2613), .A2(n2579), .ZN(n4369) );
  NAND2_X1 U2896 ( .A1(n4362), .A2(n4356), .ZN(n4166) );
  INV_X1 U2897 ( .A(n4362), .ZN(n4361) );
  INV_X1 U2898 ( .A(n4311), .ZN(n4310) );
  NAND2_X1 U2899 ( .A1(n2295), .A2(n2294), .ZN(n4311) );
  AND2_X1 U2900 ( .A1(n2529), .A2(STATE_REG_SCAN_IN), .ZN(n4312) );
  OR2_X1 U2901 ( .A1(n3056), .A2(n3055), .ZN(n4317) );
  INV_X1 U2902 ( .A(n3573), .ZN(U4043) );
  INV_X1 U2903 ( .A(IR_REG_23__SCAN_IN), .ZN(n2245) );
  NAND2_X1 U2904 ( .A1(n2246), .A2(n2245), .ZN(n2244) );
  NOR2_X1 U2905 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2234)
         );
  INV_X1 U2906 ( .A(n2238), .ZN(n2235) );
  NAND2_X1 U2907 ( .A1(n2284), .A2(IR_REG_31__SCAN_IN), .ZN(n2237) );
  INV_X1 U2908 ( .A(n4169), .ZN(n2242) );
  NAND2_X1 U2909 ( .A1(n2275), .A2(n2238), .ZN(n2239) );
  NAND2_X1 U2910 ( .A1(n2239), .A2(IR_REG_31__SCAN_IN), .ZN(n2240) );
  MUX2_X1 U2911 ( .A(IR_REG_31__SCAN_IN), .B(n2240), .S(IR_REG_25__SCAN_IN), 
        .Z(n2241) );
  NAND2_X1 U2912 ( .A1(n2241), .A2(n2284), .ZN(n2435) );
  OAI21_X1 U2913 ( .B1(n2246), .B2(n2245), .A(n2244), .ZN(n2529) );
  INV_X1 U2914 ( .A(n4312), .ZN(n2297) );
  OR2_X2 U2915 ( .A1(n2530), .A2(n2297), .ZN(n3573) );
  INV_X2 U2916 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2917 ( .A(DATAI_3_), .ZN(n2248) );
  NAND2_X1 U2918 ( .A1(n2247), .A2(IR_REG_31__SCAN_IN), .ZN(n2337) );
  XNOR2_X1 U2919 ( .A(n2337), .B(IR_REG_3__SCAN_IN), .ZN(n2535) );
  INV_X1 U2920 ( .A(n2535), .ZN(n2400) );
  MUX2_X1 U2921 ( .A(n2248), .B(n2400), .S(STATE_REG_SCAN_IN), .Z(n2249) );
  INV_X1 U2922 ( .A(n2249), .ZN(U3349) );
  NAND2_X1 U2923 ( .A1(n2250), .A2(IR_REG_31__SCAN_IN), .ZN(n2252) );
  INV_X1 U2924 ( .A(IR_REG_5__SCAN_IN), .ZN(n2251) );
  XNOR2_X1 U2925 ( .A(n2252), .B(n2251), .ZN(n2635) );
  INV_X1 U2926 ( .A(DATAI_5_), .ZN(n2253) );
  MUX2_X1 U2927 ( .A(n2635), .B(n2253), .S(U3149), .Z(n2254) );
  INV_X1 U2928 ( .A(n2254), .ZN(U3347) );
  OR2_X1 U2929 ( .A1(n2255), .A2(n2091), .ZN(n2256) );
  XNOR2_X1 U2930 ( .A(n2256), .B(IR_REG_6__SCAN_IN), .ZN(n2676) );
  INV_X1 U2931 ( .A(n2676), .ZN(n2373) );
  INV_X1 U2932 ( .A(DATAI_6_), .ZN(n2257) );
  MUX2_X1 U2933 ( .A(n2373), .B(n2257), .S(U3149), .Z(n2258) );
  INV_X1 U2934 ( .A(n2258), .ZN(U3346) );
  INV_X1 U2935 ( .A(DATAI_8_), .ZN(n4409) );
  INV_X1 U2936 ( .A(IR_REG_6__SCAN_IN), .ZN(n2259) );
  NAND2_X1 U2937 ( .A1(n2255), .A2(n2259), .ZN(n2825) );
  NAND2_X1 U2938 ( .A1(n2825), .A2(IR_REG_31__SCAN_IN), .ZN(n2378) );
  INV_X1 U2939 ( .A(IR_REG_7__SCAN_IN), .ZN(n2260) );
  NAND2_X1 U2940 ( .A1(n2378), .A2(n2260), .ZN(n2261) );
  NAND2_X1 U2941 ( .A1(n2261), .A2(IR_REG_31__SCAN_IN), .ZN(n2263) );
  INV_X1 U2942 ( .A(IR_REG_8__SCAN_IN), .ZN(n2262) );
  XNOR2_X1 U2943 ( .A(n2263), .B(n2262), .ZN(n2881) );
  MUX2_X1 U2944 ( .A(n4409), .B(n2881), .S(STATE_REG_SCAN_IN), .Z(n2264) );
  INV_X1 U2945 ( .A(n2264), .ZN(U3344) );
  INV_X1 U2946 ( .A(DATAI_20_), .ZN(n4402) );
  NAND2_X1 U2947 ( .A1(n2265), .A2(IR_REG_31__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U2948 ( .A1(n2441), .A2(n2266), .ZN(n2267) );
  NAND2_X1 U2949 ( .A1(n2267), .A2(IR_REG_31__SCAN_IN), .ZN(n2269) );
  INV_X1 U2950 ( .A(n3552), .ZN(n2480) );
  NAND2_X1 U2951 ( .A1(n2480), .A2(STATE_REG_SCAN_IN), .ZN(n2270) );
  OAI21_X1 U2952 ( .B1(STATE_REG_SCAN_IN), .B2(n4402), .A(n2270), .ZN(U3332)
         );
  INV_X1 U2953 ( .A(DATAI_21_), .ZN(n2274) );
  NAND2_X1 U2954 ( .A1(n2271), .A2(IR_REG_31__SCAN_IN), .ZN(n2272) );
  NAND2_X1 U2955 ( .A1(n3491), .A2(STATE_REG_SCAN_IN), .ZN(n2273) );
  OAI21_X1 U2956 ( .B1(STATE_REG_SCAN_IN), .B2(n2274), .A(n2273), .ZN(U3331)
         );
  INV_X1 U2957 ( .A(DATAI_22_), .ZN(n2280) );
  INV_X1 U2958 ( .A(n2275), .ZN(n2276) );
  NAND2_X1 U2959 ( .A1(n3562), .A2(STATE_REG_SCAN_IN), .ZN(n2279) );
  OAI21_X1 U2960 ( .B1(STATE_REG_SCAN_IN), .B2(n2280), .A(n2279), .ZN(U3330)
         );
  INV_X1 U2961 ( .A(DATAI_24_), .ZN(n2283) );
  NAND2_X1 U2962 ( .A1(n2281), .A2(STATE_REG_SCAN_IN), .ZN(n2282) );
  OAI21_X1 U2963 ( .B1(STATE_REG_SCAN_IN), .B2(n2283), .A(n2282), .ZN(U3328)
         );
  INV_X1 U2964 ( .A(DATAI_31_), .ZN(n4400) );
  INV_X1 U2965 ( .A(IR_REG_29__SCAN_IN), .ZN(n4388) );
  OR4_X1 U2966 ( .A1(n2289), .A2(IR_REG_30__SCAN_IN), .A3(n2091), .A4(U3149), 
        .ZN(n2285) );
  OAI21_X1 U2967 ( .B1(STATE_REG_SCAN_IN), .B2(n4400), .A(n2285), .ZN(U3321)
         );
  INV_X1 U2968 ( .A(DATAI_29_), .ZN(n2288) );
  NAND2_X1 U2969 ( .A1(n2301), .A2(STATE_REG_SCAN_IN), .ZN(n2287) );
  OAI21_X1 U2970 ( .B1(STATE_REG_SCAN_IN), .B2(n2288), .A(n2287), .ZN(U3323)
         );
  INV_X1 U2971 ( .A(DATAI_30_), .ZN(n4399) );
  XNOR2_X2 U2972 ( .A(n2290), .B(IR_REG_30__SCAN_IN), .ZN(n2303) );
  NAND2_X1 U2973 ( .A1(n2303), .A2(STATE_REG_SCAN_IN), .ZN(n2291) );
  OAI21_X1 U2974 ( .B1(STATE_REG_SCAN_IN), .B2(n4399), .A(n2291), .ZN(U3322)
         );
  NAND2_X1 U2975 ( .A1(n2435), .A2(B_REG_SCAN_IN), .ZN(n2292) );
  MUX2_X1 U2976 ( .A(n2292), .B(B_REG_SCAN_IN), .S(n2281), .Z(n2293) );
  INV_X1 U2977 ( .A(n2440), .ZN(n2295) );
  INV_X1 U2978 ( .A(n2582), .ZN(n2294) );
  INV_X1 U2979 ( .A(D_REG_1__SCAN_IN), .ZN(n2439) );
  INV_X1 U2980 ( .A(n2435), .ZN(n4170) );
  NOR3_X1 U2981 ( .A1(n2297), .A2(n4169), .A3(n4170), .ZN(n2296) );
  AOI21_X1 U2982 ( .B1(n4311), .B2(n2439), .A(n2296), .ZN(U3459) );
  INV_X1 U2983 ( .A(D_REG_0__SCAN_IN), .ZN(n2438) );
  NOR2_X1 U2984 ( .A1(n2297), .A2(n2281), .ZN(n2298) );
  AOI22_X1 U2985 ( .A1(n4311), .A2(n2438), .B1(n2298), .B2(n2242), .ZN(U3458)
         );
  OR2_X1 U2986 ( .A1(n2529), .A2(U3149), .ZN(n3564) );
  NAND2_X1 U2987 ( .A1(n2582), .A2(n3564), .ZN(n2320) );
  INV_X1 U2988 ( .A(n2320), .ZN(n2300) );
  NAND2_X1 U2989 ( .A1(n3562), .A2(n3491), .ZN(n2450) );
  INV_X1 U2990 ( .A(n2450), .ZN(n2474) );
  NAND2_X1 U2991 ( .A1(n2529), .A2(n2474), .ZN(n2299) );
  AND2_X1 U2992 ( .A1(n3436), .A2(n2299), .ZN(n2321) );
  NOR2_X2 U2993 ( .A1(n2300), .A2(n2321), .ZN(n4268) );
  NOR2_X1 U2994 ( .A1(n4268), .A2(U4043), .ZN(U3148) );
  INV_X1 U2995 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4509) );
  INV_X1 U2996 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2305) );
  NAND2_X1 U2997 ( .A1(n3196), .A2(REG2_REG_3__SCAN_IN), .ZN(n2304) );
  NAND2_X1 U2998 ( .A1(n2702), .A2(U4043), .ZN(n2306) );
  OAI21_X1 U2999 ( .B1(U4043), .B2(n4509), .A(n2306), .ZN(U3553) );
  INV_X1 U3000 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U3001 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2307) );
  INV_X1 U3002 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3045) );
  INV_X1 U3003 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3406) );
  NAND2_X1 U3004 ( .A1(n3071), .A2(REG3_REG_16__SCAN_IN), .ZN(n3091) );
  INV_X1 U3005 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3090) );
  INV_X1 U3006 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4511) );
  NOR2_X1 U3007 ( .A1(n3107), .A2(REG3_REG_19__SCAN_IN), .ZN(n2308) );
  OR2_X1 U3008 ( .A1(n3127), .A2(n2308), .ZN(n3251) );
  INV_X1 U3009 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4076) );
  OAI22_X1 U3010 ( .A1(n3285), .A2(n3251), .B1(n3282), .B2(n4076), .ZN(n2312)
         );
  NAND2_X1 U3011 ( .A1(n3196), .A2(REG2_REG_19__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U3012 ( .A1(n3434), .A2(REG0_REG_19__SCAN_IN), .ZN(n2309) );
  NAND2_X1 U3013 ( .A1(n2310), .A2(n2309), .ZN(n2311) );
  NAND2_X1 U3014 ( .A1(n3913), .A2(U4043), .ZN(n2313) );
  OAI21_X1 U3015 ( .B1(U4043), .B2(n4506), .A(n2313), .ZN(U3569) );
  INV_X1 U3016 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4508) );
  AND2_X1 U3017 ( .A1(n3048), .A2(n3406), .ZN(n2314) );
  OR2_X1 U3018 ( .A1(n2314), .A2(n3071), .ZN(n3967) );
  INV_X1 U3019 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3602) );
  OAI22_X1 U3020 ( .A1(n3285), .A2(n3967), .B1(n3282), .B2(n3602), .ZN(n2318)
         );
  NAND2_X1 U3021 ( .A1(n3196), .A2(REG2_REG_15__SCAN_IN), .ZN(n2316) );
  NAND2_X1 U3022 ( .A1(n3434), .A2(REG0_REG_15__SCAN_IN), .ZN(n2315) );
  NAND2_X1 U3023 ( .A1(n2316), .A2(n2315), .ZN(n2317) );
  NAND2_X1 U3024 ( .A1(n3683), .A2(U4043), .ZN(n2319) );
  OAI21_X1 U3025 ( .B1(U4043), .B2(n4508), .A(n2319), .ZN(U3565) );
  NAND2_X1 U3026 ( .A1(n2321), .A2(n2320), .ZN(n4188) );
  NAND2_X1 U3027 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2323) );
  NAND2_X1 U3028 ( .A1(n2322), .A2(n2323), .ZN(n2324) );
  XNOR2_X1 U3029 ( .A(n2324), .B(IR_REG_28__SCAN_IN), .ZN(n3579) );
  NAND2_X1 U3030 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2325)
         );
  AND2_X1 U3031 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2359)
         );
  NAND2_X1 U3032 ( .A1(n2360), .A2(n2359), .ZN(n2329) );
  INV_X1 U3033 ( .A(n2367), .ZN(n4177) );
  NAND2_X1 U3034 ( .A1(n4177), .A2(REG1_REG_1__SCAN_IN), .ZN(n2328) );
  NAND2_X1 U3035 ( .A1(n2329), .A2(n2328), .ZN(n3586) );
  XNOR2_X2 U3036 ( .A(n2330), .B(IR_REG_2__SCAN_IN), .ZN(n4176) );
  INV_X1 U3037 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2468) );
  XNOR2_X1 U3038 ( .A(n4176), .B(n2468), .ZN(n3585) );
  NAND2_X1 U3039 ( .A1(n3586), .A2(n3585), .ZN(n2332) );
  NAND2_X1 U3040 ( .A1(n4176), .A2(REG1_REG_2__SCAN_IN), .ZN(n2331) );
  NAND2_X1 U3041 ( .A1(n2332), .A2(n2331), .ZN(n2333) );
  XNOR2_X1 U3042 ( .A(n2333), .B(n2400), .ZN(n2394) );
  NAND2_X1 U3043 ( .A1(n2394), .A2(REG1_REG_3__SCAN_IN), .ZN(n2335) );
  NAND2_X1 U3044 ( .A1(n2333), .A2(n2535), .ZN(n2334) );
  NAND2_X1 U3045 ( .A1(n2337), .A2(n2336), .ZN(n2338) );
  NAND2_X1 U3046 ( .A1(n2338), .A2(IR_REG_31__SCAN_IN), .ZN(n2339) );
  INV_X1 U3047 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U3048 ( .A1(n2340), .A2(n4201), .ZN(n2341) );
  INV_X1 U3049 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4461) );
  MUX2_X1 U3050 ( .A(REG1_REG_5__SCAN_IN), .B(n4461), .S(n2635), .Z(n2344) );
  MUX2_X1 U3051 ( .A(n4461), .B(REG1_REG_5__SCAN_IN), .S(n2635), .Z(n2342) );
  XNOR2_X1 U3052 ( .A(n2322), .B(n2343), .ZN(n3665) );
  INV_X1 U3053 ( .A(n3665), .ZN(n4186) );
  AOI211_X1 U3054 ( .C1(n2345), .C2(n2344), .A(n2369), .B(n4256), .ZN(n2356)
         );
  INV_X1 U3055 ( .A(n4176), .ZN(n3587) );
  INV_X1 U3056 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2349) );
  INV_X1 U3057 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2346) );
  MUX2_X1 U3058 ( .A(REG2_REG_1__SCAN_IN), .B(n2346), .S(n2367), .Z(n2361) );
  INV_X1 U3059 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2347) );
  NOR2_X1 U3060 ( .A1(n2367), .A2(n2346), .ZN(n3590) );
  MUX2_X1 U3061 ( .A(REG2_REG_2__SCAN_IN), .B(n2349), .S(n4176), .Z(n2348) );
  XNOR2_X1 U3062 ( .A(n2350), .B(n4201), .ZN(n4196) );
  INV_X1 U3063 ( .A(n2350), .ZN(n2351) );
  AOI22_X1 U3064 ( .A1(n4196), .A2(REG2_REG_4__SCAN_IN), .B1(n4201), .B2(n2351), .ZN(n2354) );
  INV_X1 U3065 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2352) );
  MUX2_X1 U3066 ( .A(REG2_REG_5__SCAN_IN), .B(n2352), .S(n2635), .Z(n2353) );
  NOR2_X1 U3067 ( .A1(n2354), .A2(n2353), .ZN(n2370) );
  OR2_X1 U3068 ( .A1(n3579), .A2(n3665), .ZN(n3559) );
  AOI211_X1 U3069 ( .C1(n2354), .C2(n2353), .A(n2370), .B(n4245), .ZN(n2355)
         );
  NOR2_X1 U3070 ( .A1(n2356), .A2(n2355), .ZN(n2358) );
  AND2_X1 U3071 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2660) );
  AOI21_X1 U3072 ( .B1(n4268), .B2(ADDR_REG_5__SCAN_IN), .A(n2660), .ZN(n2357)
         );
  OAI211_X1 U3073 ( .C1(n2635), .C2(n4281), .A(n2358), .B(n2357), .ZN(U3245)
         );
  INV_X1 U3074 ( .A(n4256), .ZN(n4276) );
  XOR2_X1 U3075 ( .A(n2360), .B(n2359), .Z(n2364) );
  NOR2_X1 U3076 ( .A1(n2038), .A2(n2347), .ZN(n3581) );
  INV_X1 U3077 ( .A(n3581), .ZN(n2362) );
  AOI211_X1 U3078 ( .C1(n2362), .C2(n2361), .A(n3595), .B(n4245), .ZN(n2363)
         );
  AOI21_X1 U3079 ( .B1(n4276), .B2(n2364), .A(n2363), .ZN(n2366) );
  AOI22_X1 U3080 ( .A1(n4268), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n2365) );
  OAI211_X1 U3081 ( .C1(n2367), .C2(n4281), .A(n2366), .B(n2365), .ZN(U3241)
         );
  NOR2_X1 U3082 ( .A1(n2635), .A2(n4461), .ZN(n2368) );
  XNOR2_X1 U3083 ( .A(n2380), .B(n2373), .ZN(n2379) );
  XNOR2_X1 U3084 ( .A(n2379), .B(REG1_REG_6__SCAN_IN), .ZN(n2377) );
  INV_X1 U3085 ( .A(n2635), .ZN(n2371) );
  XOR2_X1 U3086 ( .A(REG2_REG_6__SCAN_IN), .B(n2387), .Z(n2375) );
  AND2_X1 U3087 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n2693) );
  AOI21_X1 U3088 ( .B1(n4268), .B2(ADDR_REG_6__SCAN_IN), .A(n2693), .ZN(n2372)
         );
  OAI21_X1 U3089 ( .B1(n2373), .B2(n4281), .A(n2372), .ZN(n2374) );
  AOI21_X1 U3090 ( .B1(n2375), .B2(n4278), .A(n2374), .ZN(n2376) );
  OAI21_X1 U3091 ( .B1(n2377), .B2(n4256), .A(n2376), .ZN(U3246) );
  INV_X1 U3092 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4462) );
  XNOR2_X1 U3093 ( .A(n2378), .B(IR_REG_7__SCAN_IN), .ZN(n4175) );
  MUX2_X1 U3094 ( .A(n4462), .B(REG1_REG_7__SCAN_IN), .S(n4175), .Z(n2383) );
  NAND2_X1 U3095 ( .A1(n2379), .A2(REG1_REG_6__SCAN_IN), .ZN(n2382) );
  NAND2_X1 U3096 ( .A1(n2380), .A2(n2676), .ZN(n2381) );
  NAND2_X1 U3097 ( .A1(n2382), .A2(n2381), .ZN(n2405) );
  XOR2_X1 U3098 ( .A(n2383), .B(n2405), .Z(n2393) );
  INV_X1 U3099 ( .A(n4281), .ZN(n4252) );
  AND2_X1 U3100 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n2728) );
  AOI21_X1 U3101 ( .B1(n4268), .B2(ADDR_REG_7__SCAN_IN), .A(n2728), .ZN(n2384)
         );
  INV_X1 U3102 ( .A(n2384), .ZN(n2391) );
  INV_X1 U3103 ( .A(n2385), .ZN(n2386) );
  INV_X1 U3104 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2763) );
  MUX2_X1 U3105 ( .A(n2763), .B(REG2_REG_7__SCAN_IN), .S(n4175), .Z(n2388) );
  AOI211_X1 U3106 ( .C1(n2389), .C2(n2388), .A(n4245), .B(n2401), .ZN(n2390)
         );
  AOI211_X1 U3107 ( .C1(n4252), .C2(n4175), .A(n2391), .B(n2390), .ZN(n2392)
         );
  OAI21_X1 U3108 ( .B1(n4256), .B2(n2393), .A(n2392), .ZN(U3247) );
  XOR2_X1 U3109 ( .A(REG1_REG_3__SCAN_IN), .B(n2394), .Z(n2397) );
  INV_X1 U3110 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2597) );
  XNOR2_X1 U3111 ( .A(n2395), .B(n2597), .ZN(n2396) );
  AOI22_X1 U3112 ( .A1(n4276), .A2(n2397), .B1(n4278), .B2(n2396), .ZN(n2399)
         );
  INV_X1 U3113 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4416) );
  NOR2_X1 U3114 ( .A1(STATE_REG_SCAN_IN), .A2(n4416), .ZN(n2552) );
  AOI21_X1 U3115 ( .B1(n4268), .B2(ADDR_REG_3__SCAN_IN), .A(n2552), .ZN(n2398)
         );
  OAI211_X1 U3116 ( .C1(n2400), .C2(n4281), .A(n2399), .B(n2398), .ZN(U3243)
         );
  XOR2_X1 U3117 ( .A(REG2_REG_8__SCAN_IN), .B(n2870), .Z(n2410) );
  INV_X1 U3118 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2402) );
  NOR2_X1 U3119 ( .A1(n2402), .A2(STATE_REG_SCAN_IN), .ZN(n2790) );
  NOR2_X1 U3120 ( .A1(n4281), .A2(n2881), .ZN(n2403) );
  AOI211_X1 U3121 ( .C1(n4268), .C2(ADDR_REG_8__SCAN_IN), .A(n2790), .B(n2403), 
        .ZN(n2409) );
  AND2_X1 U3122 ( .A1(n4175), .A2(REG1_REG_7__SCAN_IN), .ZN(n2404) );
  INV_X1 U3123 ( .A(n2406), .ZN(n2407) );
  INV_X1 U3124 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2818) );
  OAI211_X1 U3125 ( .C1(n2407), .C2(REG1_REG_8__SCAN_IN), .A(n4276), .B(n2880), 
        .ZN(n2408) );
  OAI211_X1 U3126 ( .C1(n2410), .C2(n4245), .A(n2409), .B(n2408), .ZN(U3248)
         );
  NAND2_X1 U3127 ( .A1(n2459), .A2(REG0_REG_0__SCAN_IN), .ZN(n2412) );
  INV_X1 U3128 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4303) );
  NAND2_X1 U3129 ( .A1(n2412), .A2(n2411), .ZN(n2416) );
  INV_X1 U3130 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U3131 ( .A1(n3196), .A2(REG2_REG_0__SCAN_IN), .ZN(n2413) );
  OAI21_X1 U3132 ( .B1(n2414), .B2(n2469), .A(n2413), .ZN(n2415) );
  NAND2_X1 U3133 ( .A1(n2454), .A2(n2455), .ZN(n2506) );
  INV_X1 U3134 ( .A(n2506), .ZN(n2417) );
  INV_X1 U3135 ( .A(n2530), .ZN(n2424) );
  INV_X1 U3136 ( .A(n2587), .ZN(n2418) );
  INV_X2 U3137 ( .A(n2422), .ZN(n3258) );
  AOI21_X1 U3138 ( .B1(n3578), .B2(n3263), .A(n2421), .ZN(n2495) );
  INV_X1 U3139 ( .A(n3578), .ZN(n2479) );
  INV_X2 U3140 ( .A(n3258), .ZN(n3081) );
  XNOR2_X1 U3141 ( .A(n2495), .B(n2496), .ZN(n3580) );
  NOR4_X1 U3142 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2428) );
  NOR4_X1 U3143 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2427) );
  NOR4_X1 U3144 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2426) );
  NOR4_X1 U3145 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2425) );
  NAND4_X1 U3146 ( .A1(n2428), .A2(n2427), .A3(n2426), .A4(n2425), .ZN(n2434)
         );
  NOR2_X1 U3147 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_17__SCAN_IN), .ZN(n2432) );
  NOR4_X1 U31480 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2431) );
  NOR4_X1 U31490 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2430) );
  NOR4_X1 U3150 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2429) );
  NAND4_X1 U3151 ( .A1(n2432), .A2(n2431), .A3(n2430), .A4(n2429), .ZN(n2433)
         );
  OAI21_X1 U3152 ( .B1(n2434), .B2(n2433), .A(n2440), .ZN(n2489) );
  NAND2_X1 U3153 ( .A1(n2242), .A2(n2435), .ZN(n2486) );
  AND2_X1 U3154 ( .A1(n2489), .A2(n2486), .ZN(n2585) );
  INV_X1 U3155 ( .A(n2281), .ZN(n2436) );
  NAND2_X1 U3156 ( .A1(n2440), .A2(n2439), .ZN(n2583) );
  INV_X1 U3157 ( .A(n4171), .ZN(n3643) );
  AND2_X1 U3158 ( .A1(n3552), .A2(n3643), .ZN(n2449) );
  OR2_X1 U3159 ( .A1(n2506), .A2(n2449), .ZN(n2442) );
  NAND2_X1 U3160 ( .A1(n2442), .A2(n2450), .ZN(n2446) );
  NOR2_X1 U3161 ( .A1(n2582), .A2(n2446), .ZN(n2443) );
  INV_X1 U3162 ( .A(n2457), .ZN(n2448) );
  INV_X1 U3163 ( .A(n2493), .ZN(n2444) );
  AND2_X1 U3164 ( .A1(n4312), .A2(n2444), .ZN(n2445) );
  NAND2_X1 U3165 ( .A1(n2448), .A2(n3560), .ZN(n2533) );
  INV_X1 U3166 ( .A(n2533), .ZN(n2452) );
  NAND2_X1 U3167 ( .A1(n2446), .A2(n4001), .ZN(n2447) );
  NAND2_X1 U3168 ( .A1(n2448), .A2(n2447), .ZN(n2451) );
  OR2_X1 U3169 ( .A1(n2450), .A2(n2449), .ZN(n2580) );
  NAND2_X1 U3170 ( .A1(n2451), .A2(n2580), .ZN(n2532) );
  NOR3_X1 U3171 ( .A1(n2452), .A2(n2532), .A3(n2582), .ZN(n2524) );
  INV_X1 U3172 ( .A(n2524), .ZN(n2502) );
  NOR2_X1 U3173 ( .A1(n2582), .A2(n4001), .ZN(n2453) );
  NAND2_X1 U3174 ( .A1(n2457), .A2(n2453), .ZN(n2456) );
  AND2_X1 U3175 ( .A1(n3552), .A2(n4171), .ZN(n4299) );
  NAND2_X1 U3176 ( .A1(n4339), .A2(n2455), .ZN(n2487) );
  NAND2_X1 U3177 ( .A1(n2457), .A2(n3560), .ZN(n2501) );
  INV_X1 U3178 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2458) );
  AOI21_X1 U3179 ( .B1(n2502), .B2(REG3_REG_0__SCAN_IN), .A(n2460), .ZN(n2461)
         );
  OAI21_X1 U3180 ( .B1(n3580), .B2(n3399), .A(n2461), .ZN(U3229) );
  NAND2_X1 U3181 ( .A1(n2463), .A2(n2573), .ZN(n2589) );
  NAND2_X1 U3182 ( .A1(n2464), .A2(n2465), .ZN(n2575) );
  NAND2_X1 U3183 ( .A1(n2575), .A2(n2466), .ZN(n2666) );
  XNOR2_X1 U3184 ( .A(n3562), .B(n2587), .ZN(n2467) );
  NAND2_X1 U3185 ( .A1(n2467), .A2(n3643), .ZN(n2812) );
  NAND2_X1 U3186 ( .A1(n2459), .A2(REG0_REG_2__SCAN_IN), .ZN(n2473) );
  OR2_X1 U3187 ( .A1(n2469), .A2(n2468), .ZN(n2472) );
  NAND2_X1 U3188 ( .A1(n3196), .A2(REG2_REG_2__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3189 ( .A1(n2573), .A2(n4031), .ZN(n2476) );
  NAND2_X1 U3190 ( .A1(n3578), .A2(n4006), .ZN(n2475) );
  OAI211_X1 U3191 ( .C1(n2593), .C2(n4002), .A(n2476), .B(n2475), .ZN(n2477)
         );
  INV_X1 U3192 ( .A(n2477), .ZN(n2484) );
  NAND2_X1 U3193 ( .A1(n2479), .A2(n2478), .ZN(n3488) );
  NAND2_X1 U3194 ( .A1(n3562), .A2(n4171), .ZN(n2481) );
  NAND2_X1 U3195 ( .A1(n2480), .A2(n3491), .ZN(n3556) );
  NAND2_X1 U3196 ( .A1(n2482), .A2(n3945), .ZN(n2483) );
  OAI211_X1 U3197 ( .C1(n2666), .C2(n2812), .A(n2484), .B(n2483), .ZN(n2664)
         );
  INV_X1 U3198 ( .A(n4339), .ZN(n4329) );
  INV_X1 U3199 ( .A(n4356), .ZN(n4093) );
  NAND2_X1 U3200 ( .A1(n2499), .A2(n2507), .ZN(n2616) );
  OAI21_X1 U3201 ( .B1(n2507), .B2(n2499), .A(n2616), .ZN(n2670) );
  OAI22_X1 U3202 ( .A1(n2666), .A2(n4329), .B1(n4093), .B2(n2670), .ZN(n2485)
         );
  NOR2_X1 U3203 ( .A1(n2664), .A2(n2485), .ZN(n4328) );
  NAND2_X1 U3204 ( .A1(n2583), .A2(n2486), .ZN(n2491) );
  NAND2_X1 U3205 ( .A1(n2487), .A2(n2580), .ZN(n2488) );
  NOR2_X1 U3206 ( .A1(n2582), .A2(n2488), .ZN(n2490) );
  NAND2_X1 U3207 ( .A1(n4367), .A2(REG1_REG_1__SCAN_IN), .ZN(n2492) );
  OAI21_X1 U3208 ( .B1(n4328), .B2(n4367), .A(n2492), .ZN(U3519) );
  OAI22_X1 U3209 ( .A1(n2496), .A2(n2495), .B1(n3191), .B2(n2494), .ZN(n2514)
         );
  INV_X2 U32100 ( .A(n3258), .ZN(n3204) );
  XNOR2_X1 U32110 ( .A(n2514), .B(n2513), .ZN(n2505) );
  INV_X1 U32120 ( .A(n3394), .ZN(n3410) );
  INV_X1 U32130 ( .A(n3408), .ZN(n3318) );
  AOI22_X1 U32140 ( .A1(n2573), .A2(n3410), .B1(n3318), .B2(n3578), .ZN(n2504)
         );
  INV_X1 U32150 ( .A(n3407), .ZN(n3319) );
  AOI22_X1 U32160 ( .A1(n2502), .A2(REG3_REG_1__SCAN_IN), .B1(n3319), .B2(
        n3577), .ZN(n2503) );
  OAI211_X1 U32170 ( .C1(n2505), .C2(n3399), .A(n2504), .B(n2503), .ZN(U3219)
         );
  NAND2_X1 U32180 ( .A1(n3578), .A2(n2507), .ZN(n3490) );
  NAND2_X1 U32190 ( .A1(n3488), .A2(n3490), .ZN(n4306) );
  NOR2_X1 U32200 ( .A1(n2507), .A2(n2506), .ZN(n4302) );
  INV_X1 U32210 ( .A(n2812), .ZN(n4000) );
  OAI21_X1 U32220 ( .B1(n4000), .B2(n3945), .A(n4306), .ZN(n2508) );
  AOI211_X1 U32230 ( .C1(n4339), .C2(n4306), .A(n4302), .B(n4300), .ZN(n4326)
         );
  NAND2_X1 U32240 ( .A1(n4367), .A2(REG1_REG_0__SCAN_IN), .ZN(n2509) );
  OAI21_X1 U32250 ( .B1(n4326), .B2(n4367), .A(n2509), .ZN(U3518) );
  MUX2_X1 U32260 ( .A(n4176), .B(DATAI_2_), .S(n3436), .Z(n2617) );
  INV_X1 U32270 ( .A(n2617), .ZN(n2577) );
  XNOR2_X1 U32280 ( .A(n2515), .B(n3191), .ZN(n2519) );
  INV_X1 U32290 ( .A(n2519), .ZN(n2517) );
  OAI22_X1 U32300 ( .A1(n2593), .A2(n3218), .B1(n3204), .B2(n2577), .ZN(n2518)
         );
  INV_X1 U32310 ( .A(n2518), .ZN(n2516) );
  OAI21_X1 U32320 ( .B1(n2522), .B2(n2521), .A(n2539), .ZN(n2527) );
  INV_X1 U32330 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2523) );
  OAI22_X1 U32340 ( .A1(n2524), .A2(n2523), .B1(n2631), .B2(n3407), .ZN(n2525)
         );
  AOI211_X1 U32350 ( .C1(n2527), .C2(n3267), .A(n2526), .B(n2525), .ZN(n2528)
         );
  INV_X1 U32360 ( .A(n2528), .ZN(U3234) );
  NAND2_X1 U32370 ( .A1(n2530), .A2(n2529), .ZN(n2531) );
  OAI21_X1 U32380 ( .B1(n2532), .B2(n2531), .A(STATE_REG_SCAN_IN), .ZN(n2534)
         );
  INV_X1 U32390 ( .A(n3397), .ZN(n3413) );
  MUX2_X1 U32400 ( .A(n2535), .B(DATAI_3_), .S(n3436), .Z(n2627) );
  NAND2_X1 U32410 ( .A1(n2627), .A2(n3120), .ZN(n2536) );
  XNOR2_X1 U32420 ( .A(n2537), .B(n3191), .ZN(n2555) );
  INV_X1 U32430 ( .A(n2627), .ZN(n2630) );
  OAI22_X1 U32440 ( .A1(n2631), .A2(n3218), .B1(n3216), .B2(n2630), .ZN(n2556)
         );
  XOR2_X1 U32450 ( .A(n2555), .B(n2556), .Z(n2541) );
  OAI21_X1 U32460 ( .B1(n2541), .B2(n2540), .A(n2561), .ZN(n2542) );
  NAND2_X1 U32470 ( .A1(n2542), .A2(n3267), .ZN(n2554) );
  NAND2_X1 U32480 ( .A1(n3196), .A2(REG2_REG_4__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32490 ( .A1(n2459), .A2(REG0_REG_4__SCAN_IN), .ZN(n2549) );
  INV_X1 U32500 ( .A(n2564), .ZN(n2545) );
  INV_X1 U32510 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U32520 ( .A1(n4416), .A2(n2543), .ZN(n2544) );
  NAND2_X1 U32530 ( .A1(n2545), .A2(n2544), .ZN(n2710) );
  OR2_X1 U32540 ( .A1(n3285), .A2(n2710), .ZN(n2548) );
  OR2_X1 U32550 ( .A1(n3282), .A2(n2546), .ZN(n2547) );
  OAI22_X1 U32560 ( .A1(n2593), .A2(n3408), .B1(n3407), .B2(n2658), .ZN(n2551)
         );
  AOI211_X1 U32570 ( .C1(n2627), .C2(n3410), .A(n2552), .B(n2551), .ZN(n2553)
         );
  OAI211_X1 U32580 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3413), .A(n2554), .B(n2553), .ZN(U3215) );
  INV_X1 U32590 ( .A(n2555), .ZN(n2558) );
  INV_X1 U32600 ( .A(n2556), .ZN(n2557) );
  NAND2_X1 U32610 ( .A1(n2558), .A2(n2557), .ZN(n2560) );
  AND2_X1 U32620 ( .A1(n2561), .A2(n2560), .ZN(n2563) );
  MUX2_X1 U32630 ( .A(n4201), .B(DATAI_4_), .S(n3436), .Z(n2701) );
  OAI22_X1 U32640 ( .A1(n2658), .A2(n3081), .B1(n2709), .B2(n2423), .ZN(n2559)
         );
  XNOR2_X1 U32650 ( .A(n2559), .B(n3261), .ZN(n2652) );
  OAI22_X1 U32660 ( .A1(n2658), .A2(n3218), .B1(n2709), .B2(n3204), .ZN(n2653)
         );
  XNOR2_X1 U32670 ( .A(n2652), .B(n2653), .ZN(n2562) );
  OAI211_X1 U32680 ( .C1(n2563), .C2(n2562), .A(n3267), .B(n2656), .ZN(n2571)
         );
  AND2_X1 U32690 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4193) );
  NAND2_X1 U32700 ( .A1(n3196), .A2(REG2_REG_5__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U32710 ( .A1(n3434), .A2(REG0_REG_5__SCAN_IN), .ZN(n2567) );
  OAI21_X1 U32720 ( .B1(n2564), .B2(REG3_REG_5__SCAN_IN), .A(n2685), .ZN(n2663) );
  OR2_X1 U32730 ( .A1(n3285), .A2(n2663), .ZN(n2566) );
  OR2_X1 U32740 ( .A1(n3282), .A2(n4461), .ZN(n2565) );
  OAI22_X1 U32750 ( .A1(n2732), .A2(n3407), .B1(n3408), .B2(n2631), .ZN(n2569)
         );
  AOI211_X1 U32760 ( .C1(n2701), .C2(n3410), .A(n4193), .B(n2569), .ZN(n2570)
         );
  OAI211_X1 U32770 ( .C1(n3413), .C2(n2710), .A(n2571), .B(n2570), .ZN(U3227)
         );
  NAND2_X1 U32780 ( .A1(n2572), .A2(n2573), .ZN(n2574) );
  INV_X1 U32790 ( .A(n2603), .ZN(n2576) );
  NAND2_X1 U32800 ( .A1(n3577), .A2(n2577), .ZN(n3496) );
  NAND2_X1 U32810 ( .A1(n2593), .A2(n2577), .ZN(n2578) );
  NAND2_X1 U32820 ( .A1(n2601), .A2(n2578), .ZN(n2629) );
  NAND2_X1 U32830 ( .A1(n2631), .A2(n2627), .ZN(n3498) );
  NAND2_X1 U32840 ( .A1(n2702), .A2(n2630), .ZN(n3495) );
  XNOR2_X1 U32850 ( .A(n2629), .B(n3471), .ZN(n4330) );
  INV_X1 U32860 ( .A(n2579), .ZN(n2612) );
  INV_X1 U32870 ( .A(n2580), .ZN(n2581) );
  NOR2_X1 U32880 ( .A1(n2582), .A2(n2581), .ZN(n2584) );
  NAND4_X1 U32890 ( .A1(n2612), .A2(n2585), .A3(n2584), .A4(n2583), .ZN(n2586)
         );
  OR2_X1 U32900 ( .A1(n2587), .A2(n3643), .ZN(n2625) );
  INV_X1 U32910 ( .A(n2625), .ZN(n2588) );
  NAND2_X1 U32920 ( .A1(n4284), .A2(n2588), .ZN(n2714) );
  NAND2_X1 U32930 ( .A1(n2590), .A2(n2589), .ZN(n2605) );
  NAND2_X1 U32940 ( .A1(n2605), .A2(n3472), .ZN(n2604) );
  NAND2_X1 U32950 ( .A1(n2604), .A2(n3493), .ZN(n2636) );
  XNOR2_X1 U32960 ( .A(n2636), .B(n3471), .ZN(n2595) );
  AOI22_X1 U32970 ( .A1(n3576), .A2(n3912), .B1(n4031), .B2(n2627), .ZN(n2592)
         );
  OAI21_X1 U32980 ( .B1(n2593), .B2(n3954), .A(n2592), .ZN(n2594) );
  AOI21_X1 U32990 ( .B1(n2595), .B2(n3945), .A(n2594), .ZN(n2596) );
  OAI21_X1 U33000 ( .B1(n4330), .B2(n2812), .A(n2596), .ZN(n4331) );
  NAND2_X1 U33010 ( .A1(n4331), .A2(n4284), .ZN(n2600) );
  AOI21_X1 U33020 ( .B1(n2627), .B2(n2614), .A(n2006), .ZN(n4333) );
  OAI22_X1 U33030 ( .A1(n4284), .A2(n2597), .B1(n4304), .B2(
        REG3_REG_3__SCAN_IN), .ZN(n2598) );
  AOI21_X1 U33040 ( .B1(n4333), .B2(n4294), .A(n2598), .ZN(n2599) );
  OAI211_X1 U33050 ( .C1(n4330), .C2(n2714), .A(n2600), .B(n2599), .ZN(U3287)
         );
  INV_X1 U33060 ( .A(n2601), .ZN(n2602) );
  AOI21_X1 U33070 ( .B1(n3472), .B2(n2603), .A(n2602), .ZN(n2607) );
  INV_X1 U33080 ( .A(n2607), .ZN(n4295) );
  OAI21_X1 U33090 ( .B1(n3472), .B2(n2605), .A(n2604), .ZN(n2610) );
  AOI22_X1 U33100 ( .A1(n2572), .A2(n4006), .B1(n2617), .B2(n4031), .ZN(n2606)
         );
  OAI21_X1 U33110 ( .B1(n2631), .B2(n4002), .A(n2606), .ZN(n2609) );
  NOR2_X1 U33120 ( .A1(n2607), .A2(n2812), .ZN(n2608) );
  AOI211_X1 U33130 ( .C1(n3945), .C2(n2610), .A(n2609), .B(n2608), .ZN(n4298)
         );
  INV_X1 U33140 ( .A(n4298), .ZN(n2611) );
  AOI21_X1 U33150 ( .B1(n4339), .B2(n4295), .A(n2611), .ZN(n2624) );
  INV_X1 U33160 ( .A(n2614), .ZN(n2615) );
  AOI21_X1 U33170 ( .B1(n2617), .B2(n2616), .A(n2615), .ZN(n4293) );
  INV_X1 U33180 ( .A(n4166), .ZN(n2620) );
  INV_X1 U33190 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2618) );
  NOR2_X1 U33200 ( .A1(n4362), .A2(n2618), .ZN(n2619) );
  AOI21_X1 U33210 ( .B1(n4293), .B2(n2620), .A(n2619), .ZN(n2621) );
  OAI21_X1 U33220 ( .B1(n2624), .B2(n4361), .A(n2621), .ZN(U3471) );
  INV_X1 U33230 ( .A(n4110), .ZN(n2622) );
  AOI22_X1 U33240 ( .A1(n4293), .A2(n2622), .B1(REG1_REG_2__SCAN_IN), .B2(
        n4367), .ZN(n2623) );
  OAI21_X1 U33250 ( .B1(n2624), .B2(n4367), .A(n2623), .ZN(U3520) );
  NAND2_X1 U33260 ( .A1(n2812), .A2(n2625), .ZN(n2626) );
  INV_X1 U33270 ( .A(n3972), .ZN(n3991) );
  NAND2_X1 U33280 ( .A1(n2702), .A2(n2627), .ZN(n2628) );
  NAND2_X1 U33290 ( .A1(n2629), .A2(n2628), .ZN(n2633) );
  NAND2_X1 U33300 ( .A1(n2631), .A2(n2630), .ZN(n2632) );
  NAND2_X1 U33310 ( .A1(n2633), .A2(n2632), .ZN(n2696) );
  NAND2_X1 U33320 ( .A1(n3576), .A2(n2709), .ZN(n3502) );
  NAND2_X1 U33330 ( .A1(n2658), .A2(n2701), .ZN(n3499) );
  NAND2_X1 U33340 ( .A1(n3576), .A2(n2701), .ZN(n2634) );
  MUX2_X1 U33350 ( .A(n2635), .B(n2253), .S(n3436), .Z(n2731) );
  AND2_X1 U33360 ( .A1(n3575), .A2(n2731), .ZN(n2738) );
  INV_X1 U33370 ( .A(n2738), .ZN(n3501) );
  INV_X1 U33380 ( .A(n2731), .ZN(n2734) );
  NAND2_X1 U33390 ( .A1(n2732), .A2(n2734), .ZN(n3516) );
  NAND2_X1 U33400 ( .A1(n3501), .A2(n3516), .ZN(n3462) );
  XNOR2_X1 U33410 ( .A(n2733), .B(n3462), .ZN(n4343) );
  INV_X1 U33420 ( .A(n3499), .ZN(n2637) );
  XNOR2_X1 U33430 ( .A(n2739), .B(n3462), .ZN(n2646) );
  INV_X1 U33440 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2638) );
  XNOR2_X1 U33450 ( .A(n2685), .B(n2638), .ZN(n4283) );
  INV_X1 U33460 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2639) );
  OAI22_X1 U33470 ( .A1(n3285), .A2(n4283), .B1(n3282), .B2(n2639), .ZN(n2643)
         );
  NAND2_X1 U33480 ( .A1(n3196), .A2(REG2_REG_6__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U33490 ( .A1(n3434), .A2(REG0_REG_6__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U33500 ( .A1(n2641), .A2(n2640), .ZN(n2642) );
  AOI22_X1 U33510 ( .A1(n3574), .A2(n3912), .B1(n2734), .B2(n4031), .ZN(n2644)
         );
  OAI21_X1 U33520 ( .B1(n2658), .B2(n3954), .A(n2644), .ZN(n2645) );
  AOI21_X1 U3353 ( .B1(n2646), .B2(n3945), .A(n2645), .ZN(n4344) );
  MUX2_X1 U33540 ( .A(n4344), .B(n2352), .S(n2000), .Z(n2650) );
  OR2_X1 U3355 ( .A1(n2708), .A2(n2731), .ZN(n2647) );
  AND2_X1 U3356 ( .A1(n2745), .A2(n2647), .ZN(n4347) );
  INV_X1 U3357 ( .A(n2663), .ZN(n2648) );
  INV_X1 U3358 ( .A(n4304), .ZN(n4292) );
  AOI22_X1 U3359 ( .A1(n4347), .A2(n4294), .B1(n2648), .B2(n4292), .ZN(n2649)
         );
  OAI211_X1 U3360 ( .C1(n3991), .C2(n4343), .A(n2650), .B(n2649), .ZN(U3285)
         );
  OAI22_X1 U3361 ( .A1(n2732), .A2(n3204), .B1(n2731), .B2(n2423), .ZN(n2651)
         );
  XNOR2_X1 U3362 ( .A(n2651), .B(n3261), .ZN(n2671) );
  OAI22_X1 U3363 ( .A1(n2732), .A2(n3218), .B1(n2731), .B2(n3216), .ZN(n2672)
         );
  XNOR2_X1 U3364 ( .A(n2671), .B(n2672), .ZN(n2674) );
  XOR2_X1 U3365 ( .A(n2674), .B(n2675), .Z(n2657) );
  NAND2_X1 U3366 ( .A1(n2657), .A2(n3267), .ZN(n2662) );
  INV_X1 U3367 ( .A(n3574), .ZN(n2737) );
  OAI22_X1 U3368 ( .A1(n2658), .A2(n3408), .B1(n3407), .B2(n2737), .ZN(n2659)
         );
  AOI211_X1 U3369 ( .C1(n2734), .C2(n3410), .A(n2660), .B(n2659), .ZN(n2661)
         );
  OAI211_X1 U3370 ( .C1(n3413), .C2(n2663), .A(n2662), .B(n2661), .ZN(U3224)
         );
  MUX2_X1 U3371 ( .A(n2664), .B(REG2_REG_1__SCAN_IN), .S(n2000), .Z(n2665) );
  INV_X1 U3372 ( .A(n2665), .ZN(n2669) );
  INV_X1 U3373 ( .A(n2666), .ZN(n2667) );
  INV_X1 U3374 ( .A(n2714), .ZN(n4307) );
  AOI22_X1 U3375 ( .A1(n2667), .A2(n4307), .B1(REG3_REG_1__SCAN_IN), .B2(n4292), .ZN(n2668) );
  OAI211_X1 U3376 ( .C1(n4015), .C2(n2670), .A(n2669), .B(n2668), .ZN(U3289)
         );
  INV_X1 U3377 ( .A(n2671), .ZN(n2673) );
  NAND2_X1 U3378 ( .A1(n3574), .A2(n3258), .ZN(n2678) );
  MUX2_X1 U3379 ( .A(n2676), .B(DATAI_6_), .S(n3436), .Z(n2766) );
  NAND2_X1 U3380 ( .A1(n2766), .A2(n3120), .ZN(n2677) );
  NAND2_X1 U3381 ( .A1(n2678), .A2(n2677), .ZN(n2679) );
  XNOR2_X1 U3382 ( .A(n2679), .B(n3261), .ZN(n2681) );
  AOI22_X1 U3383 ( .A1(n3574), .A2(n3263), .B1(n2766), .B2(n3258), .ZN(n2680)
         );
  OR2_X1 U3384 ( .A1(n2681), .A2(n2680), .ZN(n2716) );
  INV_X1 U3385 ( .A(n2716), .ZN(n2682) );
  AND2_X1 U3386 ( .A1(n2681), .A2(n2680), .ZN(n2715) );
  NOR2_X1 U3387 ( .A1(n2682), .A2(n2715), .ZN(n2683) );
  XNOR2_X1 U3388 ( .A(n2717), .B(n2683), .ZN(n2684) );
  NAND2_X1 U3389 ( .A1(n2684), .A2(n3267), .ZN(n2695) );
  NAND2_X1 U3390 ( .A1(n3196), .A2(REG2_REG_7__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U3391 ( .A1(n3434), .A2(REG0_REG_7__SCAN_IN), .ZN(n2690) );
  INV_X1 U3392 ( .A(n2685), .ZN(n2686) );
  AOI21_X1 U3393 ( .B1(n2686), .B2(REG3_REG_6__SCAN_IN), .A(
        REG3_REG_7__SCAN_IN), .ZN(n2687) );
  OR2_X1 U3394 ( .A1(n2687), .A2(n2721), .ZN(n2762) );
  OR2_X1 U3395 ( .A1(n3285), .A2(n2762), .ZN(n2689) );
  OR2_X1 U3396 ( .A1(n3282), .A2(n4462), .ZN(n2688) );
  OAI22_X1 U3397 ( .A1(n2732), .A2(n3408), .B1(n3407), .B2(n2799), .ZN(n2692)
         );
  AOI211_X1 U3398 ( .C1(n2766), .C2(n3410), .A(n2693), .B(n2692), .ZN(n2694)
         );
  OAI211_X1 U3399 ( .C1(n3413), .C2(n4283), .A(n2695), .B(n2694), .ZN(U3236)
         );
  NAND2_X1 U3400 ( .A1(n2696), .A2(n2179), .ZN(n2698) );
  NAND2_X1 U3401 ( .A1(n2699), .A2(n2698), .ZN(n4335) );
  XNOR2_X1 U3402 ( .A(n2700), .B(n2179), .ZN(n2706) );
  AOI22_X1 U3403 ( .A1(n2702), .A2(n4006), .B1(n2701), .B2(n4031), .ZN(n2704)
         );
  NAND2_X1 U3404 ( .A1(n3575), .A2(n3912), .ZN(n2703) );
  OAI211_X1 U3405 ( .C1(n4335), .C2(n2812), .A(n2704), .B(n2703), .ZN(n2705)
         );
  AOI21_X1 U3406 ( .B1(n2706), .B2(n3945), .A(n2705), .ZN(n2707) );
  INV_X1 U3407 ( .A(n2707), .ZN(n4337) );
  OAI211_X1 U3408 ( .C1(n2006), .C2(n2709), .A(n2095), .B(n4356), .ZN(n4336)
         );
  OAI22_X1 U3409 ( .A1(n4336), .A2(n4171), .B1(n4304), .B2(n2710), .ZN(n2711)
         );
  OAI21_X1 U3410 ( .B1(n4337), .B2(n2711), .A(n4284), .ZN(n2713) );
  NAND2_X1 U3411 ( .A1(n2000), .A2(REG2_REG_4__SCAN_IN), .ZN(n2712) );
  OAI211_X1 U3412 ( .C1(n4335), .C2(n2714), .A(n2713), .B(n2712), .ZN(U3286)
         );
  MUX2_X1 U3413 ( .A(n4175), .B(DATAI_7_), .S(n3436), .Z(n2802) );
  INV_X1 U3414 ( .A(n2802), .ZN(n2754) );
  OAI22_X1 U3415 ( .A1(n2799), .A2(n3081), .B1(n2754), .B2(n2423), .ZN(n2718)
         );
  XNOR2_X1 U3416 ( .A(n2718), .B(n3191), .ZN(n2775) );
  OAI22_X1 U3417 ( .A1(n2799), .A2(n3218), .B1(n2754), .B2(n3204), .ZN(n2774)
         );
  XOR2_X1 U3418 ( .A(n2775), .B(n2774), .Z(n2719) );
  NAND2_X1 U3419 ( .A1(n2720), .A2(n2719), .ZN(n2776) );
  OAI211_X1 U3420 ( .C1(n2720), .C2(n2719), .A(n2776), .B(n3267), .ZN(n2730)
         );
  NAND2_X1 U3421 ( .A1(n3196), .A2(REG2_REG_8__SCAN_IN), .ZN(n2726) );
  NAND2_X1 U3422 ( .A1(n3434), .A2(REG0_REG_8__SCAN_IN), .ZN(n2725) );
  OR2_X1 U3423 ( .A1(n2721), .A2(REG3_REG_8__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U3424 ( .A1(n2783), .A2(n2722), .ZN(n2781) );
  OR2_X1 U3425 ( .A1(n3285), .A2(n2781), .ZN(n2724) );
  OR2_X1 U3426 ( .A1(n3282), .A2(n2818), .ZN(n2723) );
  OAI22_X1 U3427 ( .A1(n2929), .A2(n3407), .B1(n3408), .B2(n2737), .ZN(n2727)
         );
  AOI211_X1 U3428 ( .C1(n2802), .C2(n3410), .A(n2728), .B(n2727), .ZN(n2729)
         );
  OAI211_X1 U3429 ( .C1(n3413), .C2(n2762), .A(n2730), .B(n2729), .ZN(U3210)
         );
  NAND2_X1 U3430 ( .A1(n3575), .A2(n2734), .ZN(n2735) );
  NAND2_X1 U3431 ( .A1(n2736), .A2(n2735), .ZN(n2768) );
  NAND2_X1 U3432 ( .A1(n2737), .A2(n2766), .ZN(n3504) );
  INV_X1 U3433 ( .A(n2766), .ZN(n2746) );
  NAND2_X1 U3434 ( .A1(n3574), .A2(n2746), .ZN(n3515) );
  NAND2_X1 U3435 ( .A1(n3504), .A2(n3515), .ZN(n3483) );
  XOR2_X1 U3436 ( .A(n2768), .B(n3483), .Z(n4288) );
  INV_X1 U3437 ( .A(n4288), .ZN(n2744) );
  OAI21_X1 U3438 ( .B1(n2739), .B2(n2738), .A(n3516), .ZN(n2755) );
  XNOR2_X1 U3439 ( .A(n2755), .B(n3483), .ZN(n2742) );
  OAI22_X1 U3440 ( .A1(n2799), .A2(n4002), .B1(n2746), .B2(n4001), .ZN(n2740)
         );
  AOI21_X1 U3441 ( .B1(n4006), .B2(n3575), .A(n2740), .ZN(n2741) );
  OAI21_X1 U3442 ( .B1(n2742), .B2(n4010), .A(n2741), .ZN(n2743) );
  AOI21_X1 U3443 ( .B1(n4288), .B2(n4000), .A(n2743), .ZN(n4291) );
  OAI21_X1 U3444 ( .B1(n4329), .B2(n2744), .A(n4291), .ZN(n2752) );
  INV_X1 U3445 ( .A(n2745), .ZN(n2747) );
  OAI21_X1 U3446 ( .B1(n2747), .B2(n2746), .A(n2760), .ZN(n4286) );
  INV_X1 U3447 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2748) );
  OAI22_X1 U3448 ( .A1(n4286), .A2(n4166), .B1(n4362), .B2(n2748), .ZN(n2749)
         );
  AOI21_X1 U3449 ( .B1(n2752), .B2(n4362), .A(n2749), .ZN(n2750) );
  INV_X1 U3450 ( .A(n2750), .ZN(U3479) );
  OAI22_X1 U3451 ( .A1(n4286), .A2(n4110), .B1(n4369), .B2(n2639), .ZN(n2751)
         );
  AOI21_X1 U3452 ( .B1(n2752), .B2(n4369), .A(n2751), .ZN(n2753) );
  INV_X1 U3453 ( .A(n2753), .ZN(U3524) );
  OAI22_X1 U3454 ( .A1(n2929), .A2(n4002), .B1(n2754), .B2(n4001), .ZN(n2758)
         );
  NAND2_X1 U3455 ( .A1(n2799), .A2(n2802), .ZN(n3505) );
  NAND2_X1 U3456 ( .A1(n4370), .A2(n2754), .ZN(n3508) );
  XOR2_X1 U3457 ( .A(n3468), .B(n2797), .Z(n2756) );
  NOR2_X1 U34580 ( .A1(n2756), .A2(n4010), .ZN(n2757) );
  AOI211_X1 U34590 ( .C1(n4006), .C2(n3574), .A(n2758), .B(n2757), .ZN(n4352)
         );
  NAND2_X1 U3460 ( .A1(n2760), .A2(n2802), .ZN(n2759) );
  NAND2_X1 U3461 ( .A1(n2759), .A2(n4356), .ZN(n2761) );
  OR2_X1 U3462 ( .A1(n2761), .A2(n2805), .ZN(n4351) );
  INV_X1 U3463 ( .A(n4351), .ZN(n2765) );
  OAI22_X1 U3464 ( .A1(n4284), .A2(n2763), .B1(n2762), .B2(n4304), .ZN(n2764)
         );
  AOI21_X1 U3465 ( .B1(n2765), .B2(n3919), .A(n2764), .ZN(n2773) );
  AND2_X1 U3466 ( .A1(n3574), .A2(n2766), .ZN(n2767) );
  OAI22_X1 U34670 ( .A1(n2768), .A2(n2767), .B1(n2766), .B2(n3574), .ZN(n2771)
         );
  INV_X1 U3468 ( .A(n2771), .ZN(n2770) );
  NAND2_X1 U34690 ( .A1(n2770), .A2(n2769), .ZN(n2804) );
  NAND2_X1 U3470 ( .A1(n2771), .A2(n3468), .ZN(n4349) );
  NAND3_X1 U34710 ( .A1(n2804), .A2(n4349), .A3(n3972), .ZN(n2772) );
  OAI211_X1 U3472 ( .C1(n4352), .C2(n2000), .A(n2773), .B(n2772), .ZN(U3283)
         );
  INV_X1 U34730 ( .A(n2774), .ZN(n2778) );
  INV_X1 U3474 ( .A(n2775), .ZN(n2777) );
  MUX2_X1 U34750 ( .A(n2881), .B(n4409), .S(n3436), .Z(n2841) );
  OAI22_X1 U3476 ( .A1(n2929), .A2(n3081), .B1(n2841), .B2(n2423), .ZN(n2779)
         );
  XOR2_X1 U34770 ( .A(n2779), .B(n3191), .Z(n2920) );
  INV_X1 U3478 ( .A(n2841), .ZN(n2844) );
  AOI22_X1 U34790 ( .A1(n3572), .A2(n3263), .B1(n2844), .B2(n3258), .ZN(n2918)
         );
  INV_X1 U3480 ( .A(n2918), .ZN(n2921) );
  XNOR2_X1 U34810 ( .A(n2920), .B(n2921), .ZN(n2780) );
  XNOR2_X1 U3482 ( .A(n2922), .B(n2780), .ZN(n2795) );
  INV_X1 U34830 ( .A(n2781), .ZN(n2807) );
  NAND2_X1 U3484 ( .A1(n2783), .A2(n2782), .ZN(n2784) );
  NAND2_X1 U34850 ( .A1(n2828), .A2(n2784), .ZN(n2934) );
  INV_X1 U3486 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2785) );
  OAI22_X1 U34870 ( .A1(n3285), .A2(n2934), .B1(n3282), .B2(n2785), .ZN(n2789)
         );
  NAND2_X1 U3488 ( .A1(n3196), .A2(REG2_REG_9__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U34890 ( .A1(n3434), .A2(REG0_REG_9__SCAN_IN), .ZN(n2786) );
  NAND2_X1 U3490 ( .A1(n2787), .A2(n2786), .ZN(n2788) );
  AOI22_X1 U34910 ( .A1(n3318), .A2(n4370), .B1(n3319), .B2(n3571), .ZN(n2792)
         );
  INV_X1 U3492 ( .A(n2790), .ZN(n2791) );
  OAI211_X1 U34930 ( .C1(n3394), .C2(n2841), .A(n2792), .B(n2791), .ZN(n2793)
         );
  AOI21_X1 U3494 ( .B1(n2807), .B2(n3397), .A(n2793), .ZN(n2794) );
  OAI21_X1 U34950 ( .B1(n2795), .B2(n3399), .A(n2794), .ZN(U3218) );
  INV_X1 U3496 ( .A(n3505), .ZN(n2796) );
  NAND2_X1 U34970 ( .A1(n2929), .A2(n2844), .ZN(n3509) );
  NAND2_X1 U3498 ( .A1(n3572), .A2(n2841), .ZN(n3507) );
  NAND2_X1 U34990 ( .A1(n3509), .A2(n3507), .ZN(n3463) );
  XNOR2_X1 U3500 ( .A(n2823), .B(n3463), .ZN(n2801) );
  AOI22_X1 U35010 ( .A1(n3571), .A2(n3912), .B1(n2844), .B2(n4031), .ZN(n2798)
         );
  OAI21_X1 U3502 ( .B1(n2799), .B2(n3954), .A(n2798), .ZN(n2800) );
  AOI21_X1 U35030 ( .B1(n2801), .B2(n3945), .A(n2800), .ZN(n2813) );
  NAND2_X1 U3504 ( .A1(n4370), .A2(n2802), .ZN(n2803) );
  NAND2_X1 U35050 ( .A1(n2804), .A2(n2803), .ZN(n2843) );
  XNOR2_X1 U35060 ( .A(n2843), .B(n3463), .ZN(n2814) );
  INV_X1 U35070 ( .A(n2814), .ZN(n2810) );
  NOR2_X1 U35080 ( .A1(n2805), .A2(n2841), .ZN(n2806) );
  OR2_X1 U35090 ( .A1(n2838), .A2(n2806), .ZN(n2819) );
  AOI22_X1 U35100 ( .A1(n2000), .A2(REG2_REG_8__SCAN_IN), .B1(n2807), .B2(
        n4292), .ZN(n2808) );
  OAI21_X1 U35110 ( .B1(n2819), .B2(n4015), .A(n2808), .ZN(n2809) );
  AOI21_X1 U35120 ( .B1(n2810), .B2(n3972), .A(n2809), .ZN(n2811) );
  OAI21_X1 U35130 ( .B1(n2000), .B2(n2813), .A(n2811), .ZN(U3282) );
  INV_X1 U35140 ( .A(n4354), .ZN(n4342) );
  OAI21_X1 U35150 ( .B1(n2814), .B2(n4342), .A(n2813), .ZN(n2821) );
  INV_X1 U35160 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2815) );
  OAI22_X1 U35170 ( .A1(n2819), .A2(n4166), .B1(n4362), .B2(n2815), .ZN(n2816)
         );
  AOI21_X1 U35180 ( .B1(n2821), .B2(n4362), .A(n2816), .ZN(n2817) );
  INV_X1 U35190 ( .A(n2817), .ZN(U3483) );
  OAI22_X1 U35200 ( .A1(n2819), .A2(n4110), .B1(n4369), .B2(n2818), .ZN(n2820)
         );
  AOI21_X1 U35210 ( .B1(n2821), .B2(n4369), .A(n2820), .ZN(n2822) );
  INV_X1 U35220 ( .A(n2822), .ZN(U3526) );
  NAND2_X1 U35230 ( .A1(n2823), .A2(n3509), .ZN(n2824) );
  NAND2_X1 U35240 ( .A1(n2850), .A2(IR_REG_31__SCAN_IN), .ZN(n2826) );
  XNOR2_X1 U35250 ( .A(n2826), .B(IR_REG_9__SCAN_IN), .ZN(n2883) );
  MUX2_X1 U35260 ( .A(n2883), .B(DATAI_9_), .S(n3436), .Z(n2931) );
  INV_X1 U35270 ( .A(n3517), .ZN(n2827) );
  NAND2_X1 U35280 ( .A1(n2948), .A2(n2931), .ZN(n3510) );
  NAND2_X1 U35290 ( .A1(n2827), .A2(n3510), .ZN(n3484) );
  XNOR2_X1 U35300 ( .A(n2895), .B(n3484), .ZN(n2837) );
  AND2_X1 U35310 ( .A1(n2828), .A2(n2947), .ZN(n2829) );
  OR2_X1 U35320 ( .A1(n2829), .A2(n2897), .ZN(n2952) );
  INV_X1 U35330 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4464) );
  OAI22_X1 U35340 ( .A1(n3285), .A2(n2952), .B1(n3282), .B2(n4464), .ZN(n2833)
         );
  NAND2_X1 U35350 ( .A1(n3196), .A2(REG2_REG_10__SCAN_IN), .ZN(n2831) );
  NAND2_X1 U35360 ( .A1(n3434), .A2(REG0_REG_10__SCAN_IN), .ZN(n2830) );
  NAND2_X1 U35370 ( .A1(n2831), .A2(n2830), .ZN(n2832) );
  NAND2_X1 U35380 ( .A1(n3570), .A2(n3912), .ZN(n2835) );
  NAND2_X1 U35390 ( .A1(n2931), .A2(n4031), .ZN(n2834) );
  OAI211_X1 U35400 ( .C1(n2929), .C2(n3954), .A(n2835), .B(n2834), .ZN(n2836)
         );
  AOI21_X1 U35410 ( .B1(n2837), .B2(n3945), .A(n2836), .ZN(n4360) );
  OR2_X1 U35420 ( .A1(n2838), .A2(n2917), .ZN(n2839) );
  AND2_X1 U35430 ( .A1(n2910), .A2(n2839), .ZN(n4357) );
  INV_X1 U35440 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4484) );
  OAI22_X1 U35450 ( .A1(n4284), .A2(n4484), .B1(n2934), .B2(n4304), .ZN(n2840)
         );
  AOI21_X1 U35460 ( .B1(n4357), .B2(n4294), .A(n2840), .ZN(n2849) );
  NAND2_X1 U35470 ( .A1(n2929), .A2(n2841), .ZN(n2842) );
  NAND2_X1 U35480 ( .A1(n2843), .A2(n2842), .ZN(n2846) );
  NAND2_X1 U35490 ( .A1(n3572), .A2(n2844), .ZN(n2845) );
  NAND2_X1 U35500 ( .A1(n2846), .A2(n2845), .ZN(n2909) );
  INV_X1 U35510 ( .A(n3484), .ZN(n2847) );
  XNOR2_X1 U35520 ( .A(n2909), .B(n2847), .ZN(n4355) );
  NAND2_X1 U35530 ( .A1(n4355), .A2(n3972), .ZN(n2848) );
  OAI211_X1 U35540 ( .C1(n4360), .C2(n2000), .A(n2849), .B(n2848), .ZN(U3281)
         );
  INV_X1 U35550 ( .A(n2866), .ZN(n2853) );
  INV_X1 U35560 ( .A(IR_REG_10__SCAN_IN), .ZN(n2858) );
  INV_X1 U35570 ( .A(IR_REG_11__SCAN_IN), .ZN(n2861) );
  INV_X1 U35580 ( .A(IR_REG_12__SCAN_IN), .ZN(n2851) );
  NAND3_X1 U35590 ( .A1(n2858), .A2(n2861), .A3(n2851), .ZN(n2852) );
  OAI21_X1 U35600 ( .B1(n2853), .B2(n2852), .A(IR_REG_31__SCAN_IN), .ZN(n2854)
         );
  MUX2_X1 U35610 ( .A(IR_REG_31__SCAN_IN), .B(n2854), .S(IR_REG_13__SCAN_IN), 
        .Z(n2857) );
  INV_X1 U35620 ( .A(n2855), .ZN(n2856) );
  NAND2_X1 U35630 ( .A1(n2857), .A2(n2856), .ZN(n3059) );
  NAND2_X1 U35640 ( .A1(n2866), .A2(n2858), .ZN(n2859) );
  NAND2_X1 U35650 ( .A1(n2859), .A2(IR_REG_31__SCAN_IN), .ZN(n2862) );
  NAND2_X1 U35660 ( .A1(n2862), .A2(n2861), .ZN(n2864) );
  NAND2_X1 U35670 ( .A1(n2864), .A2(IR_REG_31__SCAN_IN), .ZN(n2860) );
  XNOR2_X1 U35680 ( .A(n2860), .B(IR_REG_12__SCAN_IN), .ZN(n2986) );
  OR2_X1 U35690 ( .A1(n2862), .A2(n2861), .ZN(n2863) );
  NAND2_X1 U35700 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2966), .ZN(n2873) );
  INV_X1 U35710 ( .A(n2966), .ZN(n4319) );
  INV_X1 U35720 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2865) );
  AOI22_X1 U35730 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2966), .B1(n4319), .B2(
        n2865), .ZN(n4230) );
  OR2_X1 U35740 ( .A1(n2866), .A2(n2091), .ZN(n2867) );
  XNOR2_X1 U35750 ( .A(n2867), .B(IR_REG_10__SCAN_IN), .ZN(n4320) );
  INV_X1 U35760 ( .A(n2883), .ZN(n4323) );
  AOI22_X1 U35770 ( .A1(n2883), .A2(REG2_REG_9__SCAN_IN), .B1(n4484), .B2(
        n4323), .ZN(n4211) );
  INV_X1 U35780 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2869) );
  OAI22_X1 U35790 ( .A1(n2870), .A2(n2869), .B1(n2868), .B2(n2881), .ZN(n4210)
         );
  NAND2_X1 U35800 ( .A1(n4211), .A2(n4210), .ZN(n4209) );
  NAND2_X1 U35810 ( .A1(n4320), .A2(n2871), .ZN(n2872) );
  INV_X1 U3582 ( .A(n4320), .ZN(n4222) );
  NAND2_X1 U3583 ( .A1(n4230), .A2(n4229), .ZN(n4228) );
  NAND2_X1 U3584 ( .A1(n2873), .A2(n4228), .ZN(n2874) );
  NAND2_X1 U3585 ( .A1(n2986), .A2(n2874), .ZN(n2875) );
  INV_X1 U3586 ( .A(n2986), .ZN(n4318) );
  XNOR2_X1 U3587 ( .A(n2874), .B(n4318), .ZN(n4239) );
  NAND2_X1 U3588 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4239), .ZN(n4238) );
  NAND2_X1 U3589 ( .A1(n2875), .A2(n4238), .ZN(n3608) );
  INV_X1 U3590 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2876) );
  MUX2_X1 U3591 ( .A(REG2_REG_13__SCAN_IN), .B(n2876), .S(n3059), .Z(n2877) );
  INV_X1 U3592 ( .A(n2877), .ZN(n2879) );
  AOI21_X1 U3593 ( .B1(n2879), .B2(n3608), .A(n4245), .ZN(n2878) );
  OAI21_X1 U3594 ( .B1(n3608), .B2(n2879), .A(n2878), .ZN(n2894) );
  NOR2_X1 U3595 ( .A1(STATE_REG_SCAN_IN), .A2(n2988), .ZN(n3367) );
  AOI22_X1 U3596 ( .A1(n2883), .A2(n2785), .B1(REG1_REG_9__SCAN_IN), .B2(n4323), .ZN(n4205) );
  NOR2_X1 U3597 ( .A1(n2884), .A2(n4222), .ZN(n2885) );
  NOR2_X1 U3598 ( .A1(n4464), .A2(n4215), .ZN(n4214) );
  INV_X1 U3599 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U3600 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4319), .B1(n2966), .B2(
        n4108), .ZN(n4224) );
  NOR2_X1 U3601 ( .A1(n2886), .A2(n4318), .ZN(n2887) );
  INV_X1 U3602 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4465) );
  NOR2_X1 U3603 ( .A1(n4465), .A2(n4234), .ZN(n4233) );
  INV_X1 U3604 ( .A(n3059), .ZN(n4174) );
  NAND2_X1 U3605 ( .A1(n4174), .A2(REG1_REG_13__SCAN_IN), .ZN(n3599) );
  INV_X1 U3606 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U3607 ( .A1(n3059), .A2(n4099), .ZN(n2888) );
  NAND2_X1 U3608 ( .A1(n3599), .A2(n2888), .ZN(n2890) );
  INV_X1 U3609 ( .A(n3600), .ZN(n2889) );
  AOI211_X1 U3610 ( .C1(n2891), .C2(n2890), .A(n2889), .B(n4256), .ZN(n2892)
         );
  AOI211_X1 U3611 ( .C1(n4268), .C2(ADDR_REG_13__SCAN_IN), .A(n3367), .B(n2892), .ZN(n2893) );
  OAI211_X1 U3612 ( .C1(n4281), .C2(n3059), .A(n2894), .B(n2893), .ZN(U3253)
         );
  MUX2_X1 U3613 ( .A(n4320), .B(DATAI_10_), .S(n3436), .Z(n3003) );
  NAND2_X1 U3614 ( .A1(n3017), .A2(n3003), .ZN(n3520) );
  INV_X1 U3615 ( .A(n3003), .ZN(n3004) );
  NAND2_X1 U3616 ( .A1(n3570), .A2(n3004), .ZN(n3512) );
  NAND2_X1 U3617 ( .A1(n3520), .A2(n3512), .ZN(n3460) );
  INV_X1 U3618 ( .A(n3460), .ZN(n2896) );
  XNOR2_X1 U3619 ( .A(n2983), .B(n2896), .ZN(n2906) );
  NAND2_X1 U3620 ( .A1(n3196), .A2(REG2_REG_11__SCAN_IN), .ZN(n2902) );
  NAND2_X1 U3621 ( .A1(n3434), .A2(REG0_REG_11__SCAN_IN), .ZN(n2901) );
  NOR2_X1 U3622 ( .A1(n2897), .A2(REG3_REG_11__SCAN_IN), .ZN(n2898) );
  OR2_X1 U3623 ( .A1(n2974), .A2(n2898), .ZN(n3025) );
  OR2_X1 U3624 ( .A1(n3285), .A2(n3025), .ZN(n2900) );
  OR2_X1 U3625 ( .A1(n3282), .A2(n4108), .ZN(n2899) );
  NAND2_X1 U3626 ( .A1(n3003), .A2(n4031), .ZN(n2904) );
  NAND2_X1 U3627 ( .A1(n3571), .A2(n4006), .ZN(n2903) );
  OAI211_X1 U3628 ( .C1(n3008), .C2(n4002), .A(n2904), .B(n2903), .ZN(n2905)
         );
  AOI21_X1 U3629 ( .B1(n2906), .B2(n3945), .A(n2905), .ZN(n2955) );
  AND2_X1 U3630 ( .A1(n3571), .A2(n2931), .ZN(n2908) );
  NAND2_X1 U3631 ( .A1(n2948), .A2(n2917), .ZN(n2907) );
  XNOR2_X1 U3632 ( .A(n3006), .B(n3460), .ZN(n2953) );
  NAND2_X1 U3633 ( .A1(n2910), .A2(n3003), .ZN(n2911) );
  NAND2_X1 U3634 ( .A1(n3020), .A2(n2911), .ZN(n2961) );
  NOR2_X1 U3635 ( .A1(n2961), .A2(n4015), .ZN(n2914) );
  INV_X1 U3636 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2912) );
  OAI22_X1 U3637 ( .A1(n4284), .A2(n2912), .B1(n2952), .B2(n4304), .ZN(n2913)
         );
  AOI211_X1 U3638 ( .C1(n2953), .C2(n3972), .A(n2914), .B(n2913), .ZN(n2915)
         );
  OAI21_X1 U3639 ( .B1(n2000), .B2(n2955), .A(n2915), .ZN(U3280) );
  OAI22_X1 U3640 ( .A1(n2948), .A2(n3081), .B1(n2423), .B2(n2917), .ZN(n2916)
         );
  XNOR2_X1 U3641 ( .A(n2916), .B(n3191), .ZN(n2935) );
  OAI22_X1 U3642 ( .A1(n2948), .A2(n3218), .B1(n3204), .B2(n2917), .ZN(n2936)
         );
  XOR2_X1 U3643 ( .A(n2935), .B(n2936), .Z(n2927) );
  INV_X1 U3644 ( .A(n2922), .ZN(n2919) );
  INV_X1 U3645 ( .A(n2920), .ZN(n2924) );
  OAI21_X1 U3646 ( .B1(n2927), .B2(n2926), .A(n2944), .ZN(n2928) );
  NAND2_X1 U3647 ( .A1(n2928), .A2(n3267), .ZN(n2933) );
  NOR2_X1 U3648 ( .A1(STATE_REG_SCAN_IN), .A2(n2782), .ZN(n4207) );
  OAI22_X1 U3649 ( .A1(n2929), .A2(n3408), .B1(n3407), .B2(n3017), .ZN(n2930)
         );
  AOI211_X1 U3650 ( .C1(n2931), .C2(n3410), .A(n4207), .B(n2930), .ZN(n2932)
         );
  OAI211_X1 U3651 ( .C1(n3413), .C2(n2934), .A(n2933), .B(n2932), .ZN(U3228)
         );
  INV_X1 U3652 ( .A(n2935), .ZN(n2938) );
  INV_X1 U3653 ( .A(n2936), .ZN(n2937) );
  NAND2_X1 U3654 ( .A1(n2938), .A2(n2937), .ZN(n2942) );
  AND2_X1 U3655 ( .A1(n2944), .A2(n2942), .ZN(n2946) );
  NAND2_X1 U3656 ( .A1(n3570), .A2(n3258), .ZN(n2940) );
  NAND2_X1 U3657 ( .A1(n3003), .A2(n3120), .ZN(n2939) );
  NAND2_X1 U3658 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  XNOR2_X1 U3659 ( .A(n2941), .B(n3191), .ZN(n2962) );
  AOI22_X1 U3660 ( .A1(n3570), .A2(n3263), .B1(n3003), .B2(n3258), .ZN(n2963)
         );
  XNOR2_X1 U3661 ( .A(n2962), .B(n2963), .ZN(n2945) );
  OAI211_X1 U3662 ( .C1(n2946), .C2(n2945), .A(n3267), .B(n2965), .ZN(n2951)
         );
  NOR2_X1 U3663 ( .A1(STATE_REG_SCAN_IN), .A2(n2947), .ZN(n4216) );
  OAI22_X1 U3664 ( .A1(n2948), .A2(n3408), .B1(n3407), .B2(n3008), .ZN(n2949)
         );
  AOI211_X1 U3665 ( .C1(n3003), .C2(n3410), .A(n4216), .B(n2949), .ZN(n2950)
         );
  OAI211_X1 U3666 ( .C1(n3413), .C2(n2952), .A(n2951), .B(n2950), .ZN(U3214)
         );
  NAND2_X1 U3667 ( .A1(n2953), .A2(n4354), .ZN(n2954) );
  NAND2_X1 U3668 ( .A1(n2955), .A2(n2954), .ZN(n2958) );
  MUX2_X1 U3669 ( .A(n2958), .B(REG1_REG_10__SCAN_IN), .S(n4367), .Z(n2956) );
  INV_X1 U3670 ( .A(n2956), .ZN(n2957) );
  OAI21_X1 U3671 ( .B1(n4110), .B2(n2961), .A(n2957), .ZN(U3528) );
  MUX2_X1 U3672 ( .A(REG0_REG_10__SCAN_IN), .B(n2958), .S(n4362), .Z(n2959) );
  INV_X1 U3673 ( .A(n2959), .ZN(n2960) );
  OAI21_X1 U3674 ( .B1(n2961), .B2(n4166), .A(n2960), .ZN(U3487) );
  MUX2_X1 U3675 ( .A(n2966), .B(DATAI_11_), .S(n3436), .Z(n3014) );
  OAI22_X1 U3676 ( .A1(n3008), .A2(n3081), .B1(n3023), .B2(n2423), .ZN(n2967)
         );
  XNOR2_X1 U3677 ( .A(n2967), .B(n3191), .ZN(n2969) );
  OAI22_X1 U3678 ( .A1(n3008), .A2(n3218), .B1(n3023), .B2(n3204), .ZN(n2968)
         );
  INV_X1 U3679 ( .A(n3029), .ZN(n2970) );
  OR2_X1 U3680 ( .A1(n2969), .A2(n2968), .ZN(n3030) );
  NAND2_X1 U3681 ( .A1(n2970), .A2(n3030), .ZN(n2971) );
  XNOR2_X1 U3682 ( .A(n3031), .B(n2971), .ZN(n2972) );
  NAND2_X1 U3683 ( .A1(n2972), .A2(n3267), .ZN(n2982) );
  INV_X1 U3684 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2973) );
  NOR2_X1 U3685 ( .A1(STATE_REG_SCAN_IN), .A2(n2973), .ZN(n4226) );
  OR2_X1 U3686 ( .A1(n2974), .A2(REG3_REG_12__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U3687 ( .A1(n2989), .A2(n2975), .ZN(n3038) );
  OAI22_X1 U3688 ( .A1(n3285), .A2(n3038), .B1(n3282), .B2(n4465), .ZN(n2979)
         );
  NAND2_X1 U3689 ( .A1(n3196), .A2(REG2_REG_12__SCAN_IN), .ZN(n2977) );
  NAND2_X1 U3690 ( .A1(n3434), .A2(REG0_REG_12__SCAN_IN), .ZN(n2976) );
  NAND2_X1 U3691 ( .A1(n2977), .A2(n2976), .ZN(n2978) );
  INV_X1 U3692 ( .A(n4005), .ZN(n3365) );
  OAI22_X1 U3693 ( .A1(n3365), .A2(n3407), .B1(n3408), .B2(n3017), .ZN(n2980)
         );
  AOI211_X1 U3694 ( .C1(n3014), .C2(n3410), .A(n4226), .B(n2980), .ZN(n2981)
         );
  OAI211_X1 U3695 ( .C1(n3413), .C2(n3025), .A(n2982), .B(n2981), .ZN(U3233)
         );
  INV_X1 U3696 ( .A(n3415), .ZN(n2985) );
  NAND2_X1 U3697 ( .A1(n3008), .A2(n3014), .ZN(n3417) );
  INV_X1 U3698 ( .A(n3008), .ZN(n3569) );
  NAND2_X1 U3699 ( .A1(n3569), .A2(n3023), .ZN(n3007) );
  INV_X1 U3700 ( .A(n3007), .ZN(n3414) );
  AOI21_X1 U3701 ( .B1(n2985), .B2(n3417), .A(n3414), .ZN(n3996) );
  MUX2_X1 U3702 ( .A(n2986), .B(DATAI_12_), .S(n3436), .Z(n3673) );
  NAND2_X1 U3703 ( .A1(n3365), .A2(n3673), .ZN(n3993) );
  NAND2_X1 U3704 ( .A1(n4005), .A2(n3040), .ZN(n3994) );
  NAND2_X1 U3705 ( .A1(n3993), .A2(n3994), .ZN(n3461) );
  INV_X1 U3706 ( .A(n3461), .ZN(n2987) );
  XNOR2_X1 U3707 ( .A(n3996), .B(n2987), .ZN(n2998) );
  NAND2_X1 U3708 ( .A1(n3196), .A2(REG2_REG_13__SCAN_IN), .ZN(n2994) );
  NAND2_X1 U3709 ( .A1(n3434), .A2(REG0_REG_13__SCAN_IN), .ZN(n2993) );
  NAND2_X1 U3710 ( .A1(n2989), .A2(n2988), .ZN(n2990) );
  NAND2_X1 U3711 ( .A1(n3046), .A2(n2990), .ZN(n4016) );
  OR2_X1 U3712 ( .A1(n3285), .A2(n4016), .ZN(n2992) );
  OR2_X1 U3713 ( .A1(n3282), .A2(n4099), .ZN(n2991) );
  OAI22_X1 U3714 ( .A1(n3677), .A2(n4002), .B1(n3040), .B2(n4001), .ZN(n2996)
         );
  NOR2_X1 U3715 ( .A1(n3008), .A2(n3954), .ZN(n2995) );
  OR2_X1 U3716 ( .A1(n2996), .A2(n2995), .ZN(n2997) );
  AOI21_X1 U3717 ( .B1(n2998), .B2(n3945), .A(n2997), .ZN(n4103) );
  NOR2_X1 U3718 ( .A1(n3021), .A2(n3040), .ZN(n2999) );
  OR2_X1 U3719 ( .A1(n4012), .A2(n2999), .ZN(n4162) );
  INV_X1 U3720 ( .A(n4162), .ZN(n3002) );
  INV_X1 U3721 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3000) );
  OAI22_X1 U3722 ( .A1(n4284), .A2(n3000), .B1(n3038), .B2(n4304), .ZN(n3001)
         );
  AOI21_X1 U3723 ( .B1(n3002), .B2(n4294), .A(n3001), .ZN(n3010) );
  NOR2_X1 U3724 ( .A1(n3570), .A2(n3003), .ZN(n3005) );
  XNOR2_X1 U3725 ( .A(n3676), .B(n3461), .ZN(n4101) );
  NAND2_X1 U3726 ( .A1(n4101), .A2(n3972), .ZN(n3009) );
  OAI211_X1 U3727 ( .C1(n4103), .C2(n2000), .A(n3010), .B(n3009), .ZN(U3278)
         );
  XNOR2_X1 U3728 ( .A(n3415), .B(n3469), .ZN(n3019) );
  NAND2_X1 U3729 ( .A1(n3011), .A2(n3469), .ZN(n3012) );
  NAND2_X1 U3730 ( .A1(n3013), .A2(n3012), .ZN(n4107) );
  NAND2_X1 U3731 ( .A1(n4107), .A2(n4000), .ZN(n3016) );
  AOI22_X1 U3732 ( .A1(n4005), .A2(n3912), .B1(n3014), .B2(n4031), .ZN(n3015)
         );
  OAI211_X1 U3733 ( .C1(n3017), .C2(n3954), .A(n3016), .B(n3015), .ZN(n3018)
         );
  AOI21_X1 U3734 ( .B1(n3019), .B2(n3945), .A(n3018), .ZN(n4105) );
  INV_X1 U3735 ( .A(n3020), .ZN(n3024) );
  INV_X1 U3736 ( .A(n3021), .ZN(n3022) );
  OAI21_X1 U3737 ( .B1(n3024), .B2(n3023), .A(n3022), .ZN(n4167) );
  NOR2_X1 U3738 ( .A1(n4167), .A2(n4015), .ZN(n3027) );
  OAI22_X1 U3739 ( .A1(n4284), .A2(n2865), .B1(n3025), .B2(n4304), .ZN(n3026)
         );
  AOI211_X1 U3740 ( .C1(n4107), .C2(n4307), .A(n3027), .B(n3026), .ZN(n3028)
         );
  OAI21_X1 U3741 ( .B1(n4105), .B2(n2000), .A(n3028), .ZN(U3279) );
  NAND2_X1 U3742 ( .A1(n4005), .A2(n3258), .ZN(n3033) );
  NAND2_X1 U3743 ( .A1(n3673), .A2(n3120), .ZN(n3032) );
  NAND2_X1 U3744 ( .A1(n3033), .A2(n3032), .ZN(n3034) );
  XNOR2_X1 U3745 ( .A(n3034), .B(n3191), .ZN(n3358) );
  NAND2_X1 U3746 ( .A1(n4005), .A2(n3263), .ZN(n3036) );
  NAND2_X1 U3747 ( .A1(n3673), .A2(n3258), .ZN(n3035) );
  NAND2_X1 U3748 ( .A1(n3036), .A2(n3035), .ZN(n3356) );
  XNOR2_X1 U3749 ( .A(n3358), .B(n3356), .ZN(n3037) );
  XNOR2_X1 U3750 ( .A(n3355), .B(n3037), .ZN(n3044) );
  INV_X1 U3751 ( .A(n3038), .ZN(n3042) );
  AOI22_X1 U3752 ( .A1(n3318), .A2(n3569), .B1(n3319), .B2(n3981), .ZN(n3039)
         );
  NAND2_X1 U3753 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4235) );
  OAI211_X1 U3754 ( .C1(n3394), .C2(n3040), .A(n3039), .B(n4235), .ZN(n3041)
         );
  AOI21_X1 U3755 ( .B1(n3042), .B2(n3397), .A(n3041), .ZN(n3043) );
  OAI21_X1 U3756 ( .B1(n3044), .B2(n3399), .A(n3043), .ZN(U3221) );
  NAND2_X1 U3757 ( .A1(n3196), .A2(REG2_REG_14__SCAN_IN), .ZN(n3052) );
  NAND2_X1 U3758 ( .A1(n3434), .A2(REG0_REG_14__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U3759 ( .A1(n3046), .A2(n3045), .ZN(n3047) );
  NAND2_X1 U3760 ( .A1(n3048), .A2(n3047), .ZN(n3234) );
  OR2_X1 U3761 ( .A1(n3285), .A2(n3234), .ZN(n3050) );
  INV_X1 U3762 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4244) );
  OR2_X1 U3763 ( .A1(n3282), .A2(n4244), .ZN(n3049) );
  NOR2_X1 U3764 ( .A1(n2855), .A2(n2091), .ZN(n3053) );
  MUX2_X1 U3765 ( .A(n2091), .B(n3053), .S(IR_REG_14__SCAN_IN), .Z(n3056) );
  INV_X1 U3766 ( .A(n3054), .ZN(n3055) );
  INV_X1 U3767 ( .A(n4317), .ZN(n4251) );
  MUX2_X1 U3768 ( .A(n4251), .B(DATAI_14_), .S(n3436), .Z(n3984) );
  OAI22_X1 U3769 ( .A1(n4003), .A2(n3081), .B1(n3681), .B2(n2423), .ZN(n3057)
         );
  XNOR2_X1 U3770 ( .A(n3057), .B(n3191), .ZN(n3065) );
  INV_X1 U3771 ( .A(n3065), .ZN(n3232) );
  INV_X1 U3772 ( .A(DATAI_13_), .ZN(n3058) );
  MUX2_X1 U3773 ( .A(n3059), .B(n3058), .S(n3436), .Z(n4011) );
  OAI22_X1 U3774 ( .A1(n3677), .A2(n3081), .B1(n4011), .B2(n2423), .ZN(n3060)
         );
  XNOR2_X1 U3775 ( .A(n3060), .B(n3191), .ZN(n3062) );
  OAI22_X1 U3776 ( .A1(n3677), .A2(n3218), .B1(n4011), .B2(n3216), .ZN(n3061)
         );
  AOI21_X1 U3777 ( .B1(n3356), .B2(n3358), .A(n3360), .ZN(n3064) );
  NOR2_X1 U3778 ( .A1(n3062), .A2(n3061), .ZN(n3361) );
  NOR3_X1 U3779 ( .A1(n3360), .A2(n3356), .A3(n3358), .ZN(n3063) );
  OAI22_X1 U3780 ( .A1(n4003), .A2(n3218), .B1(n3681), .B2(n3216), .ZN(n3231)
         );
  NAND2_X1 U3781 ( .A1(n3054), .A2(IR_REG_31__SCAN_IN), .ZN(n3078) );
  XNOR2_X1 U3782 ( .A(n3078), .B(IR_REG_15__SCAN_IN), .ZN(n4315) );
  MUX2_X1 U3783 ( .A(n4315), .B(DATAI_15_), .S(n3436), .Z(n3713) );
  OAI22_X1 U3784 ( .A1(n3979), .A2(n3216), .B1(n3965), .B2(n2423), .ZN(n3068)
         );
  XNOR2_X1 U3785 ( .A(n3068), .B(n3191), .ZN(n3083) );
  NAND2_X1 U3786 ( .A1(n3683), .A2(n3263), .ZN(n3070) );
  NAND2_X1 U3787 ( .A1(n3713), .A2(n3258), .ZN(n3069) );
  NAND2_X1 U3788 ( .A1(n3196), .A2(REG2_REG_16__SCAN_IN), .ZN(n3076) );
  NAND2_X1 U3789 ( .A1(n3434), .A2(REG0_REG_16__SCAN_IN), .ZN(n3075) );
  OR2_X1 U3790 ( .A1(n3071), .A2(REG3_REG_16__SCAN_IN), .ZN(n3072) );
  NAND2_X1 U3791 ( .A1(n3091), .A2(n3072), .ZN(n3943) );
  OR2_X1 U3792 ( .A1(n3285), .A2(n3943), .ZN(n3074) );
  INV_X1 U3793 ( .A(REG1_REG_16__SCAN_IN), .ZN(n3603) );
  OR2_X1 U3794 ( .A1(n3282), .A2(n3603), .ZN(n3073) );
  INV_X1 U3795 ( .A(IR_REG_15__SCAN_IN), .ZN(n3077) );
  NAND2_X1 U3796 ( .A1(n3078), .A2(n3077), .ZN(n3079) );
  NAND2_X1 U3797 ( .A1(n3079), .A2(IR_REG_31__SCAN_IN), .ZN(n3080) );
  XNOR2_X1 U3798 ( .A(n3080), .B(IR_REG_16__SCAN_IN), .ZN(n4173) );
  MUX2_X1 U3799 ( .A(n4173), .B(DATAI_16_), .S(n3436), .Z(n3942) );
  OAI22_X1 U3800 ( .A1(n3957), .A2(n3218), .B1(n3204), .B2(n3949), .ZN(n3085)
         );
  OAI22_X1 U3801 ( .A1(n3957), .A2(n3081), .B1(n3949), .B2(n2423), .ZN(n3082)
         );
  XNOR2_X1 U3802 ( .A(n3082), .B(n3191), .ZN(n3084) );
  XOR2_X1 U3803 ( .A(n3085), .B(n3084), .Z(n3316) );
  INV_X1 U3804 ( .A(n3084), .ZN(n3087) );
  INV_X1 U3805 ( .A(n3085), .ZN(n3086) );
  NAND2_X1 U3806 ( .A1(n3089), .A2(n3088), .ZN(n3325) );
  NAND2_X1 U3807 ( .A1(n3196), .A2(REG2_REG_17__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U3808 ( .A1(n3434), .A2(REG0_REG_17__SCAN_IN), .ZN(n3095) );
  NAND2_X1 U3809 ( .A1(n3091), .A2(n3090), .ZN(n3092) );
  NAND2_X1 U3810 ( .A1(n3106), .A2(n3092), .ZN(n3933) );
  OR2_X1 U3811 ( .A1(n3285), .A2(n3933), .ZN(n3094) );
  INV_X1 U3812 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4083) );
  OR2_X1 U3813 ( .A1(n3282), .A2(n4083), .ZN(n3093) );
  NAND2_X1 U3814 ( .A1(n3097), .A2(IR_REG_31__SCAN_IN), .ZN(n3098) );
  MUX2_X1 U3815 ( .A(IR_REG_31__SCAN_IN), .B(n3098), .S(IR_REG_17__SCAN_IN), 
        .Z(n3101) );
  INV_X1 U3816 ( .A(n3099), .ZN(n3100) );
  NAND2_X1 U3817 ( .A1(n3101), .A2(n3100), .ZN(n4282) );
  INV_X1 U3818 ( .A(DATAI_17_), .ZN(n3102) );
  MUX2_X1 U3819 ( .A(n4282), .B(n3102), .S(n3436), .Z(n3930) );
  OAI22_X1 U3820 ( .A1(n3950), .A2(n3216), .B1(n2423), .B2(n3930), .ZN(n3103)
         );
  XNOR2_X1 U3821 ( .A(n3103), .B(n3191), .ZN(n3326) );
  OAI22_X1 U3822 ( .A1(n3950), .A2(n3218), .B1(n3204), .B2(n3930), .ZN(n3327)
         );
  NOR2_X1 U3823 ( .A1(n3326), .A2(n3327), .ZN(n3105) );
  NAND2_X1 U3824 ( .A1(n3326), .A2(n3327), .ZN(n3104) );
  NAND2_X1 U3825 ( .A1(n3196), .A2(REG2_REG_18__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U3826 ( .A1(n3434), .A2(REG0_REG_18__SCAN_IN), .ZN(n3112) );
  AND2_X1 U3827 ( .A1(n3106), .A2(n4511), .ZN(n3108) );
  OR2_X1 U3828 ( .A1(n3108), .A2(n3107), .ZN(n3907) );
  OR2_X1 U3829 ( .A1(n3285), .A2(n3907), .ZN(n3111) );
  INV_X1 U3830 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3109) );
  OR2_X1 U3831 ( .A1(n3282), .A2(n3109), .ZN(n3110) );
  OR2_X1 U3832 ( .A1(n3099), .A2(n2091), .ZN(n3114) );
  XNOR2_X1 U3833 ( .A(n3114), .B(IR_REG_18__SCAN_IN), .ZN(n4172) );
  MUX2_X1 U3834 ( .A(n4172), .B(DATAI_18_), .S(n3436), .Z(n3911) );
  INV_X1 U3835 ( .A(n3911), .ZN(n3905) );
  OAI22_X1 U3836 ( .A1(n3925), .A2(n3216), .B1(n3905), .B2(n2423), .ZN(n3115)
         );
  XNOR2_X1 U3837 ( .A(n3115), .B(n3191), .ZN(n3116) );
  OAI22_X1 U3838 ( .A1(n3925), .A2(n3218), .B1(n3905), .B2(n3204), .ZN(n3117)
         );
  INV_X1 U3839 ( .A(n3116), .ZN(n3119) );
  INV_X1 U3840 ( .A(n3117), .ZN(n3118) );
  NAND2_X1 U3841 ( .A1(n3119), .A2(n3118), .ZN(n3379) );
  NAND2_X1 U3842 ( .A1(n3913), .A2(n3258), .ZN(n3122) );
  MUX2_X1 U3843 ( .A(n4171), .B(DATAI_19_), .S(n3436), .Z(n3714) );
  NAND2_X1 U3844 ( .A1(n3714), .A2(n3120), .ZN(n3121) );
  NAND2_X1 U3845 ( .A1(n3122), .A2(n3121), .ZN(n3123) );
  XNOR2_X1 U3846 ( .A(n3123), .B(n3191), .ZN(n3126) );
  AOI22_X1 U3847 ( .A1(n3913), .A2(n3263), .B1(n3714), .B2(n3258), .ZN(n3124)
         );
  XNOR2_X1 U3848 ( .A(n3126), .B(n3124), .ZN(n3250) );
  INV_X1 U3849 ( .A(n3124), .ZN(n3125) );
  NAND2_X1 U3850 ( .A1(n3196), .A2(REG2_REG_20__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U3851 ( .A1(n3434), .A2(REG0_REG_20__SCAN_IN), .ZN(n3131) );
  OR2_X1 U3852 ( .A1(n3127), .A2(REG3_REG_20__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U3853 ( .A1(n3138), .A2(n3128), .ZN(n3875) );
  OR2_X1 U3854 ( .A1(n3285), .A2(n3875), .ZN(n3130) );
  INV_X1 U3855 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4072) );
  OR2_X1 U3856 ( .A1(n3282), .A2(n4072), .ZN(n3129) );
  NAND2_X1 U3857 ( .A1(n3436), .A2(DATAI_20_), .ZN(n3874) );
  OAI22_X1 U3858 ( .A1(n3888), .A2(n3216), .B1(n2423), .B2(n3874), .ZN(n3133)
         );
  XNOR2_X1 U3859 ( .A(n3133), .B(n3191), .ZN(n3134) );
  OAI22_X1 U3860 ( .A1(n3888), .A2(n3218), .B1(n3204), .B2(n3874), .ZN(n3135)
         );
  NAND2_X1 U3861 ( .A1(n3134), .A2(n3135), .ZN(n3344) );
  NAND2_X1 U3862 ( .A1(n3343), .A2(n3344), .ZN(n3342) );
  INV_X1 U3863 ( .A(n3134), .ZN(n3137) );
  INV_X1 U3864 ( .A(n3135), .ZN(n3136) );
  NAND2_X1 U3865 ( .A1(n3137), .A2(n3136), .ZN(n3346) );
  NAND2_X1 U3866 ( .A1(n3196), .A2(REG2_REG_21__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U3867 ( .A1(n3434), .A2(REG0_REG_21__SCAN_IN), .ZN(n3142) );
  INV_X1 U3868 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3297) );
  NAND2_X1 U3869 ( .A1(n3138), .A2(n3297), .ZN(n3139) );
  NAND2_X1 U3870 ( .A1(n3148), .A2(n3139), .ZN(n3853) );
  OR2_X1 U3871 ( .A1(n3285), .A2(n3853), .ZN(n3141) );
  INV_X1 U3872 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4477) );
  OR2_X1 U3873 ( .A1(n3282), .A2(n4477), .ZN(n3140) );
  OAI22_X1 U3874 ( .A1(n3859), .A2(n3216), .B1(n2423), .B2(n3852), .ZN(n3144)
         );
  XNOR2_X1 U3875 ( .A(n3144), .B(n3191), .ZN(n3294) );
  OAI22_X1 U3876 ( .A1(n3859), .A2(n3218), .B1(n3216), .B2(n3852), .ZN(n3293)
         );
  NOR2_X1 U3877 ( .A1(n3294), .A2(n3293), .ZN(n3147) );
  INV_X1 U3878 ( .A(n3294), .ZN(n3146) );
  INV_X1 U3879 ( .A(n3293), .ZN(n3145) );
  OAI22_X1 U3880 ( .A1(n3296), .A2(n3147), .B1(n3146), .B2(n3145), .ZN(n3371)
         );
  INV_X1 U3881 ( .A(n3371), .ZN(n3159) );
  INV_X1 U3882 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3374) );
  AND2_X1 U3883 ( .A1(n3148), .A2(n3374), .ZN(n3149) );
  OR2_X1 U3884 ( .A1(n3149), .A2(n3162), .ZN(n3373) );
  INV_X1 U3885 ( .A(REG1_REG_22__SCAN_IN), .ZN(n3150) );
  OR2_X1 U3886 ( .A1(n3282), .A2(n3150), .ZN(n3151) );
  OAI21_X1 U3887 ( .B1(n3373), .B2(n3285), .A(n3151), .ZN(n3152) );
  INV_X1 U3888 ( .A(n3152), .ZN(n3156) );
  NAND2_X1 U3889 ( .A1(n3196), .A2(REG2_REG_22__SCAN_IN), .ZN(n3154) );
  NAND2_X1 U3890 ( .A1(n3434), .A2(REG0_REG_22__SCAN_IN), .ZN(n3153) );
  AND2_X1 U3891 ( .A1(n3154), .A2(n3153), .ZN(n3155) );
  AND2_X1 U3892 ( .A1(n3436), .A2(DATAI_22_), .ZN(n3836) );
  OAI22_X1 U3893 ( .A1(n3699), .A2(n3216), .B1(n2423), .B2(n3698), .ZN(n3157)
         );
  XNOR2_X1 U3894 ( .A(n3157), .B(n3191), .ZN(n3161) );
  OAI22_X1 U3895 ( .A1(n3699), .A2(n3218), .B1(n3216), .B2(n3698), .ZN(n3160)
         );
  XNOR2_X1 U3896 ( .A(n3161), .B(n3160), .ZN(n3372) );
  NOR2_X1 U3897 ( .A1(n3161), .A2(n3160), .ZN(n3242) );
  OR2_X1 U3898 ( .A1(n3162), .A2(REG3_REG_23__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U3899 ( .A1(n3175), .A2(n3163), .ZN(n3820) );
  INV_X1 U3900 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4476) );
  OAI22_X1 U3901 ( .A1(n3820), .A2(n3285), .B1(n3282), .B2(n4476), .ZN(n3167)
         );
  NAND2_X1 U3902 ( .A1(n3196), .A2(REG2_REG_23__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U3903 ( .A1(n3434), .A2(REG0_REG_23__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U3904 ( .A1(n3165), .A2(n3164), .ZN(n3166) );
  NAND2_X1 U3905 ( .A1(n3831), .A2(n3258), .ZN(n3169) );
  OR2_X1 U3906 ( .A1(n3815), .A2(n2423), .ZN(n3168) );
  NAND2_X1 U3907 ( .A1(n3169), .A2(n3168), .ZN(n3170) );
  XNOR2_X1 U3908 ( .A(n3170), .B(n3261), .ZN(n3174) );
  NOR2_X1 U3909 ( .A1(n3815), .A2(n3204), .ZN(n3171) );
  AOI21_X1 U3910 ( .B1(n3831), .B2(n3263), .A(n3171), .ZN(n3173) );
  XNOR2_X1 U3911 ( .A(n3174), .B(n3173), .ZN(n3241) );
  NOR2_X1 U3912 ( .A1(n3242), .A2(n3241), .ZN(n3172) );
  NOR2_X1 U3913 ( .A1(n3174), .A2(n3173), .ZN(n3184) );
  INV_X1 U3914 ( .A(n3184), .ZN(n3181) );
  INV_X1 U3915 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U3916 ( .A1(n3175), .A2(n3337), .ZN(n3176) );
  NAND2_X1 U3917 ( .A1(n3186), .A2(n3176), .ZN(n3336) );
  OR2_X1 U3918 ( .A1(n3336), .A2(n3285), .ZN(n3179) );
  AOI22_X1 U3919 ( .A1(n3196), .A2(REG2_REG_24__SCAN_IN), .B1(n3434), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n3178) );
  INV_X1 U3920 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4055) );
  OR2_X1 U3921 ( .A1(n3282), .A2(n4055), .ZN(n3177) );
  AND2_X1 U3922 ( .A1(n3436), .A2(DATAI_24_), .ZN(n3792) );
  OAI22_X1 U3923 ( .A1(n3816), .A2(n3218), .B1(n3797), .B2(n3204), .ZN(n3185)
         );
  NAND2_X1 U3924 ( .A1(n3181), .A2(n3180), .ZN(n3182) );
  OAI22_X1 U3925 ( .A1(n3816), .A2(n3216), .B1(n3797), .B2(n2423), .ZN(n3183)
         );
  XNOR2_X1 U3926 ( .A(n3183), .B(n3191), .ZN(n3335) );
  INV_X1 U3927 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3309) );
  NAND2_X1 U3928 ( .A1(n3186), .A2(n3309), .ZN(n3187) );
  NAND2_X1 U3929 ( .A1(n3194), .A2(n3187), .ZN(n3308) );
  AOI22_X1 U3930 ( .A1(n3196), .A2(REG2_REG_25__SCAN_IN), .B1(n3434), .B2(
        REG0_REG_25__SCAN_IN), .ZN(n3189) );
  INV_X1 U3931 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4051) );
  NAND2_X1 U3932 ( .A1(n3436), .A2(DATAI_25_), .ZN(n3779) );
  OAI22_X1 U3933 ( .A1(n3704), .A2(n3216), .B1(n3779), .B2(n2423), .ZN(n3190)
         );
  XOR2_X1 U3934 ( .A(n3191), .B(n3190), .Z(n3193) );
  INV_X1 U3935 ( .A(n3779), .ZN(n3773) );
  AOI22_X1 U3936 ( .A1(n3793), .A2(n3263), .B1(n3773), .B2(n3258), .ZN(n3192)
         );
  NAND2_X1 U3937 ( .A1(n3193), .A2(n3192), .ZN(n3303) );
  NOR2_X1 U3938 ( .A1(n3193), .A2(n3192), .ZN(n3305) );
  INV_X1 U3939 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3393) );
  AND2_X1 U3940 ( .A1(n3194), .A2(n3393), .ZN(n3195) );
  INV_X1 U3941 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U3942 ( .A1(n3196), .A2(REG2_REG_26__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U3943 ( .A1(n3434), .A2(REG0_REG_26__SCAN_IN), .ZN(n3197) );
  OAI211_X1 U3944 ( .C1(n4480), .C2(n3282), .A(n3198), .B(n3197), .ZN(n3199)
         );
  INV_X1 U3945 ( .A(n3199), .ZN(n3200) );
  NAND2_X1 U3946 ( .A1(n3775), .A2(n3258), .ZN(n3202) );
  NAND2_X1 U3947 ( .A1(n3436), .A2(DATAI_26_), .ZN(n3706) );
  OR2_X1 U3948 ( .A1(n3706), .A2(n2423), .ZN(n3201) );
  NAND2_X1 U3949 ( .A1(n3202), .A2(n3201), .ZN(n3203) );
  XNOR2_X1 U3950 ( .A(n3203), .B(n3261), .ZN(n3207) );
  NOR2_X1 U3951 ( .A1(n3706), .A2(n3204), .ZN(n3205) );
  AOI21_X1 U3952 ( .B1(n3775), .B2(n3263), .A(n3205), .ZN(n3206) );
  OR2_X1 U3953 ( .A1(n3207), .A2(n3206), .ZN(n3389) );
  AND2_X1 U3954 ( .A1(n3207), .A2(n3206), .ZN(n3388) );
  AOI21_X1 U3955 ( .B1(n3387), .B2(n3389), .A(n3388), .ZN(n3257) );
  OR2_X1 U3956 ( .A1(n3208), .A2(REG3_REG_27__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U3957 ( .A1(n3208), .A2(REG3_REG_27__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U3958 ( .A1(n3746), .A2(n2009), .ZN(n3215) );
  INV_X1 U3959 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U3960 ( .A1(n3196), .A2(REG2_REG_27__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U3961 ( .A1(n3434), .A2(REG0_REG_27__SCAN_IN), .ZN(n3210) );
  OAI211_X1 U3962 ( .C1(n3212), .C2(n3282), .A(n3211), .B(n3210), .ZN(n3213)
         );
  INV_X1 U3963 ( .A(n3213), .ZN(n3214) );
  OAI22_X1 U3964 ( .A1(n3759), .A2(n3216), .B1(n2423), .B2(n3708), .ZN(n3217)
         );
  XNOR2_X1 U3965 ( .A(n3217), .B(n3261), .ZN(n3272) );
  OAI22_X1 U3966 ( .A1(n3759), .A2(n3218), .B1(n3216), .B2(n3708), .ZN(n3270)
         );
  XNOR2_X1 U3967 ( .A(n3272), .B(n3270), .ZN(n3256) );
  XNOR2_X1 U3968 ( .A(n3257), .B(n3256), .ZN(n3230) );
  INV_X1 U3969 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3219) );
  OAI22_X1 U3970 ( .A1(n3394), .A2(n3708), .B1(STATE_REG_SCAN_IN), .B2(n3219), 
        .ZN(n3228) );
  INV_X1 U3971 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3277) );
  NAND2_X1 U3972 ( .A1(n3220), .A2(n3277), .ZN(n3221) );
  NAND2_X1 U3973 ( .A1(n3732), .A2(n2009), .ZN(n3226) );
  INV_X1 U3974 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4040) );
  NAND2_X1 U3975 ( .A1(n3196), .A2(REG2_REG_28__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U3976 ( .A1(n3434), .A2(REG0_REG_28__SCAN_IN), .ZN(n3222) );
  OAI211_X1 U3977 ( .C1(n4040), .C2(n3282), .A(n3223), .B(n3222), .ZN(n3224)
         );
  INV_X1 U3978 ( .A(n3224), .ZN(n3225) );
  INV_X1 U3979 ( .A(n3669), .ZN(n3743) );
  INV_X1 U3980 ( .A(n3775), .ZN(n3310) );
  OAI22_X1 U3981 ( .A1(n3743), .A2(n3407), .B1(n3310), .B2(n3408), .ZN(n3227)
         );
  AOI211_X1 U3982 ( .C1(n3746), .C2(n3397), .A(n3228), .B(n3227), .ZN(n3229)
         );
  OAI21_X1 U3983 ( .B1(n3230), .B2(n3399), .A(n3229), .ZN(U3211) );
  XNOR2_X1 U3984 ( .A(n3232), .B(n3231), .ZN(n3233) );
  XNOR2_X1 U3985 ( .A(n3066), .B(n3233), .ZN(n3238) );
  INV_X1 U3986 ( .A(n3234), .ZN(n3987) );
  AOI22_X1 U3987 ( .A1(n3319), .A2(n3683), .B1(n3318), .B2(n3981), .ZN(n3235)
         );
  NAND2_X1 U3988 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4253) );
  OAI211_X1 U3989 ( .C1(n3394), .C2(n3681), .A(n3235), .B(n4253), .ZN(n3236)
         );
  AOI21_X1 U3990 ( .B1(n3987), .B2(n3397), .A(n3236), .ZN(n3237) );
  OAI21_X1 U3991 ( .B1(n3238), .B2(n3399), .A(n3237), .ZN(U3212) );
  INV_X1 U3992 ( .A(n3239), .ZN(n3244) );
  INV_X1 U3993 ( .A(n3240), .ZN(n3370) );
  OAI21_X1 U3994 ( .B1(n3370), .B2(n3242), .A(n3241), .ZN(n3243) );
  NAND3_X1 U3995 ( .A1(n3244), .A2(n3243), .A3(n3267), .ZN(n3248) );
  OAI22_X1 U3996 ( .A1(n3699), .A2(n3408), .B1(n3407), .B2(n3816), .ZN(n3246)
         );
  INV_X1 U3997 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4415) );
  OAI22_X1 U3998 ( .A1(n3394), .A2(n3815), .B1(STATE_REG_SCAN_IN), .B2(n4415), 
        .ZN(n3245) );
  NOR2_X1 U3999 ( .A1(n3246), .A2(n3245), .ZN(n3247) );
  OAI211_X1 U4000 ( .C1(n3413), .C2(n3820), .A(n3248), .B(n3247), .ZN(U3213)
         );
  XOR2_X1 U4001 ( .A(n3250), .B(n3249), .Z(n3255) );
  INV_X1 U4002 ( .A(n3251), .ZN(n3896) );
  INV_X1 U4003 ( .A(n3714), .ZN(n3895) );
  AOI22_X1 U4004 ( .A1(n3318), .A2(n3890), .B1(n3319), .B2(n3568), .ZN(n3252)
         );
  NAND2_X1 U4005 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3641) );
  OAI211_X1 U4006 ( .C1(n3394), .C2(n3895), .A(n3252), .B(n3641), .ZN(n3253)
         );
  AOI21_X1 U4007 ( .B1(n3896), .B2(n3397), .A(n3253), .ZN(n3254) );
  OAI21_X1 U4008 ( .B1(n3255), .B2(n3399), .A(n3254), .ZN(U3216) );
  NAND2_X1 U4009 ( .A1(n3257), .A2(n3256), .ZN(n3273) );
  INV_X1 U4010 ( .A(n3273), .ZN(n3269) );
  NAND2_X1 U4011 ( .A1(n3669), .A2(n3258), .ZN(n3260) );
  NAND2_X1 U4012 ( .A1(n3436), .A2(DATAI_28_), .ZN(n3731) );
  OR2_X1 U4013 ( .A1(n3731), .A2(n2423), .ZN(n3259) );
  NAND2_X1 U4014 ( .A1(n3260), .A2(n3259), .ZN(n3262) );
  XNOR2_X1 U4015 ( .A(n3262), .B(n3261), .ZN(n3266) );
  NAND2_X1 U4016 ( .A1(n3669), .A2(n3263), .ZN(n3264) );
  OAI21_X1 U4017 ( .B1(n3216), .B2(n3731), .A(n3264), .ZN(n3265) );
  XNOR2_X1 U4018 ( .A(n3266), .B(n3265), .ZN(n3274) );
  INV_X1 U4019 ( .A(n3274), .ZN(n3268) );
  INV_X1 U4020 ( .A(n3399), .ZN(n3267) );
  NAND2_X1 U4021 ( .A1(n3269), .A2(n2222), .ZN(n3292) );
  INV_X1 U4022 ( .A(n3270), .ZN(n3271) );
  OR2_X1 U4023 ( .A1(n3272), .A2(n3271), .ZN(n3275) );
  NAND4_X1 U4024 ( .A1(n3273), .A2(n3267), .A3(n3274), .A4(n3275), .ZN(n3291)
         );
  INV_X1 U4025 ( .A(n3275), .ZN(n3276) );
  NAND3_X1 U4026 ( .A1(n3268), .A2(n3276), .A3(n3267), .ZN(n3289) );
  OAI22_X1 U4027 ( .A1(n3394), .A2(n3731), .B1(STATE_REG_SCAN_IN), .B2(n3277), 
        .ZN(n3278) );
  INV_X1 U4028 ( .A(n3278), .ZN(n3288) );
  INV_X1 U4029 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3281) );
  NAND2_X1 U4030 ( .A1(n3196), .A2(REG2_REG_29__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4031 ( .A1(n3434), .A2(REG0_REG_29__SCAN_IN), .ZN(n3279) );
  OAI211_X1 U4032 ( .C1(n3282), .C2(n3281), .A(n3280), .B(n3279), .ZN(n3283)
         );
  INV_X1 U4033 ( .A(n3283), .ZN(n3284) );
  OAI21_X1 U4034 ( .B1(n3648), .B2(n3285), .A(n3284), .ZN(n3725) );
  AOI22_X1 U4035 ( .A1(n3726), .A2(n3318), .B1(n3319), .B2(n3725), .ZN(n3287)
         );
  NAND2_X1 U4036 ( .A1(n3397), .A2(n3732), .ZN(n3286) );
  AND4_X1 U4037 ( .A1(n3289), .A2(n3288), .A3(n3287), .A4(n3286), .ZN(n3290)
         );
  NAND3_X1 U4038 ( .A1(n3292), .A2(n3291), .A3(n3290), .ZN(U3217) );
  XNOR2_X1 U4039 ( .A(n3294), .B(n3293), .ZN(n3295) );
  XNOR2_X1 U4040 ( .A(n3296), .B(n3295), .ZN(n3302) );
  INV_X1 U4041 ( .A(n3853), .ZN(n3300) );
  OAI22_X1 U4042 ( .A1(n3394), .A2(n3852), .B1(STATE_REG_SCAN_IN), .B2(n3297), 
        .ZN(n3299) );
  OAI22_X1 U40430 ( .A1(n3888), .A2(n3408), .B1(n3407), .B2(n3699), .ZN(n3298)
         );
  AOI211_X1 U4044 ( .C1(n3300), .C2(n3397), .A(n3299), .B(n3298), .ZN(n3301)
         );
  OAI21_X1 U4045 ( .B1(n3302), .B2(n3399), .A(n3301), .ZN(U3220) );
  INV_X1 U4046 ( .A(n3303), .ZN(n3304) );
  NOR2_X1 U4047 ( .A1(n3305), .A2(n3304), .ZN(n3306) );
  XNOR2_X1 U4048 ( .A(n3307), .B(n3306), .ZN(n3314) );
  INV_X1 U4049 ( .A(n3308), .ZN(n3782) );
  OAI22_X1 U4050 ( .A1(n3394), .A2(n3779), .B1(STATE_REG_SCAN_IN), .B2(n3309), 
        .ZN(n3312) );
  OAI22_X1 U4051 ( .A1(n3310), .A2(n3407), .B1(n3816), .B2(n3408), .ZN(n3311)
         );
  AOI211_X1 U4052 ( .C1(n3782), .C2(n3397), .A(n3312), .B(n3311), .ZN(n3313)
         );
  OAI21_X1 U4053 ( .B1(n3314), .B2(n3399), .A(n3313), .ZN(U3222) );
  AOI21_X1 U4054 ( .B1(n3403), .B2(n3401), .A(n3315), .ZN(n3317) );
  XNOR2_X1 U4055 ( .A(n3317), .B(n3316), .ZN(n3324) );
  INV_X1 U4056 ( .A(n3943), .ZN(n3322) );
  AOI22_X1 U4057 ( .A1(n3319), .A2(n3688), .B1(n3318), .B2(n3683), .ZN(n3320)
         );
  NAND2_X1 U4058 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n3606) );
  OAI211_X1 U4059 ( .C1(n3394), .C2(n3949), .A(n3320), .B(n3606), .ZN(n3321)
         );
  AOI21_X1 U4060 ( .B1(n3322), .B2(n3397), .A(n3321), .ZN(n3323) );
  OAI21_X1 U4061 ( .B1(n3324), .B2(n3399), .A(n3323), .ZN(U3223) );
  XOR2_X1 U4062 ( .A(n3327), .B(n3326), .Z(n3328) );
  XNOR2_X1 U4063 ( .A(n3325), .B(n3328), .ZN(n3329) );
  NAND2_X1 U4064 ( .A1(n3329), .A2(n3267), .ZN(n3332) );
  INV_X1 U4065 ( .A(n3930), .ZN(n3687) );
  AND2_X1 U4066 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4267) );
  OAI22_X1 U4067 ( .A1(n3957), .A2(n3408), .B1(n3407), .B2(n3925), .ZN(n3330)
         );
  AOI211_X1 U4068 ( .C1(n3687), .C2(n3410), .A(n4267), .B(n3330), .ZN(n3331)
         );
  OAI211_X1 U4069 ( .C1(n3413), .C2(n3933), .A(n3332), .B(n3331), .ZN(U3225)
         );
  NAND2_X1 U4070 ( .A1(n3333), .A2(n2224), .ZN(n3334) );
  XOR2_X1 U4071 ( .A(n3335), .B(n3334), .Z(n3341) );
  INV_X1 U4072 ( .A(n3336), .ZN(n3800) );
  OAI22_X1 U4073 ( .A1(n3394), .A2(n3797), .B1(STATE_REG_SCAN_IN), .B2(n3337), 
        .ZN(n3339) );
  OAI22_X1 U4074 ( .A1(n3704), .A2(n3407), .B1(n3408), .B2(n3700), .ZN(n3338)
         );
  AOI211_X1 U4075 ( .C1(n3800), .C2(n3397), .A(n3339), .B(n3338), .ZN(n3340)
         );
  OAI21_X1 U4076 ( .B1(n3341), .B2(n3399), .A(n3340), .ZN(U3226) );
  INV_X1 U4077 ( .A(n3342), .ZN(n3347) );
  AOI21_X1 U4078 ( .B1(n3346), .B2(n3344), .A(n3343), .ZN(n3345) );
  AOI21_X1 U4079 ( .B1(n3347), .B2(n3346), .A(n3345), .ZN(n3353) );
  INV_X1 U4080 ( .A(n3875), .ZN(n3351) );
  INV_X1 U4081 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3348) );
  OAI22_X1 U4082 ( .A1(n3394), .A2(n3874), .B1(STATE_REG_SCAN_IN), .B2(n3348), 
        .ZN(n3350) );
  INV_X1 U4083 ( .A(n3913), .ZN(n3383) );
  OAI22_X1 U4084 ( .A1(n3859), .A2(n3407), .B1(n3408), .B2(n3383), .ZN(n3349)
         );
  AOI211_X1 U4085 ( .C1(n3351), .C2(n3397), .A(n3350), .B(n3349), .ZN(n3352)
         );
  OAI21_X1 U4086 ( .B1(n3353), .B2(n3399), .A(n3352), .ZN(U3230) );
  INV_X1 U4087 ( .A(n3355), .ZN(n3359) );
  INV_X1 U4088 ( .A(n3358), .ZN(n3354) );
  NAND2_X1 U4089 ( .A1(n3355), .A2(n3354), .ZN(n3357) );
  AOI22_X1 U4090 ( .A1(n3359), .A2(n3358), .B1(n3357), .B2(n3356), .ZN(n3363)
         );
  NOR2_X1 U4091 ( .A1(n3361), .A2(n3360), .ZN(n3362) );
  XNOR2_X1 U4092 ( .A(n3363), .B(n3362), .ZN(n3364) );
  NAND2_X1 U4093 ( .A1(n3364), .A2(n3267), .ZN(n3369) );
  INV_X1 U4094 ( .A(n4011), .ZN(n3678) );
  OAI22_X1 U4095 ( .A1(n3365), .A2(n3408), .B1(n3407), .B2(n4003), .ZN(n3366)
         );
  AOI211_X1 U4096 ( .C1(n3678), .C2(n3410), .A(n3367), .B(n3366), .ZN(n3368)
         );
  OAI211_X1 U4097 ( .C1(n3413), .C2(n4016), .A(n3369), .B(n3368), .ZN(U3231)
         );
  AOI21_X1 U4098 ( .B1(n3372), .B2(n3371), .A(n3370), .ZN(n3378) );
  INV_X1 U4099 ( .A(n3373), .ZN(n3837) );
  OAI22_X1 U4100 ( .A1(n3394), .A2(n3698), .B1(STATE_REG_SCAN_IN), .B2(n3374), 
        .ZN(n3376) );
  OAI22_X1 U4101 ( .A1(n3700), .A2(n3407), .B1(n3408), .B2(n3859), .ZN(n3375)
         );
  AOI211_X1 U4102 ( .C1(n3837), .C2(n3397), .A(n3376), .B(n3375), .ZN(n3377)
         );
  OAI21_X1 U4103 ( .B1(n3378), .B2(n3399), .A(n3377), .ZN(U3232) );
  NAND2_X1 U4104 ( .A1(n2032), .A2(n3379), .ZN(n3380) );
  XNOR2_X1 U4105 ( .A(n3381), .B(n3380), .ZN(n3382) );
  NAND2_X1 U4106 ( .A1(n3382), .A2(n3267), .ZN(n3386) );
  NOR2_X1 U4107 ( .A1(n4511), .A2(STATE_REG_SCAN_IN), .ZN(n3631) );
  OAI22_X1 U4108 ( .A1(n3950), .A2(n3408), .B1(n3407), .B2(n3383), .ZN(n3384)
         );
  AOI211_X1 U4109 ( .C1(n3911), .C2(n3410), .A(n3631), .B(n3384), .ZN(n3385)
         );
  OAI211_X1 U4110 ( .C1(n3413), .C2(n3907), .A(n3386), .B(n3385), .ZN(U3235)
         );
  INV_X1 U4111 ( .A(n3388), .ZN(n3390) );
  NAND2_X1 U4112 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  XNOR2_X1 U4113 ( .A(n3387), .B(n3391), .ZN(n3400) );
  INV_X1 U4114 ( .A(n3392), .ZN(n3763) );
  OAI22_X1 U4115 ( .A1(n3394), .A2(n3706), .B1(STATE_REG_SCAN_IN), .B2(n3393), 
        .ZN(n3396) );
  OAI22_X1 U4116 ( .A1(n3759), .A2(n3407), .B1(n3704), .B2(n3408), .ZN(n3395)
         );
  AOI211_X1 U4117 ( .C1(n3763), .C2(n3397), .A(n3396), .B(n3395), .ZN(n3398)
         );
  OAI21_X1 U4118 ( .B1(n3400), .B2(n3399), .A(n3398), .ZN(U3237) );
  INV_X1 U4119 ( .A(n3401), .ZN(n3402) );
  NOR2_X1 U4120 ( .A1(n3315), .A2(n3402), .ZN(n3404) );
  XNOR2_X1 U4121 ( .A(n3404), .B(n3403), .ZN(n3405) );
  NAND2_X1 U4122 ( .A1(n3405), .A2(n3267), .ZN(n3412) );
  NOR2_X1 U4123 ( .A1(STATE_REG_SCAN_IN), .A2(n3406), .ZN(n4260) );
  OAI22_X1 U4124 ( .A1(n4003), .A2(n3408), .B1(n3407), .B2(n3957), .ZN(n3409)
         );
  AOI211_X1 U4125 ( .C1(n3713), .C2(n3410), .A(n4260), .B(n3409), .ZN(n3411)
         );
  OAI211_X1 U4126 ( .C1(n3413), .C2(n3967), .A(n3412), .B(n3411), .ZN(U3238)
         );
  NAND2_X1 U4127 ( .A1(n3436), .A2(DATAI_30_), .ZN(n4028) );
  INV_X1 U4128 ( .A(n4028), .ZN(n4032) );
  NAND2_X1 U4129 ( .A1(n3436), .A2(DATAI_31_), .ZN(n4021) );
  NAND2_X1 U4130 ( .A1(n3981), .A2(n4011), .ZN(n3458) );
  NAND2_X1 U4131 ( .A1(n3994), .A2(n3458), .ZN(n3416) );
  NOR2_X1 U4132 ( .A1(n3416), .A2(n3414), .ZN(n3513) );
  NAND2_X1 U4133 ( .A1(n3415), .A2(n3513), .ZN(n3421) );
  INV_X1 U4134 ( .A(n3416), .ZN(n3419) );
  NAND2_X1 U4135 ( .A1(n3417), .A2(n3993), .ZN(n3418) );
  NAND2_X1 U4136 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  NAND2_X1 U4137 ( .A1(n3677), .A2(n3678), .ZN(n3459) );
  NAND2_X1 U4138 ( .A1(n4003), .A2(n3984), .ZN(n3650) );
  NAND2_X1 U4139 ( .A1(n3979), .A2(n3713), .ZN(n3482) );
  NAND2_X1 U4140 ( .A1(n3650), .A2(n3482), .ZN(n3523) );
  NAND2_X1 U4141 ( .A1(n3683), .A2(n3965), .ZN(n3651) );
  NAND2_X1 U4142 ( .A1(n3963), .A2(n3681), .ZN(n3467) );
  NAND2_X1 U4143 ( .A1(n3651), .A2(n3467), .ZN(n3514) );
  NAND2_X1 U4144 ( .A1(n3514), .A2(n3482), .ZN(n3529) );
  OAI21_X1 U4145 ( .B1(n3978), .B2(n3523), .A(n3529), .ZN(n3424) );
  NAND2_X1 U4146 ( .A1(n3957), .A2(n3942), .ZN(n3532) );
  INV_X1 U4147 ( .A(n3957), .ZN(n3927) );
  NAND2_X1 U4148 ( .A1(n3927), .A2(n3949), .ZN(n3652) );
  INV_X1 U4149 ( .A(n3652), .ZN(n3533) );
  NAND2_X1 U4150 ( .A1(n3890), .A2(n3905), .ZN(n3884) );
  NAND2_X1 U4151 ( .A1(n3913), .A2(n3895), .ZN(n3422) );
  NAND2_X1 U4152 ( .A1(n3884), .A2(n3422), .ZN(n3863) );
  NAND2_X1 U4153 ( .A1(n3688), .A2(n3930), .ZN(n3860) );
  NAND2_X1 U4154 ( .A1(n3568), .A2(n3874), .ZN(n3426) );
  NAND2_X1 U4155 ( .A1(n3860), .A2(n3426), .ZN(n3423) );
  AOI211_X1 U4156 ( .C1(n3424), .C2(n3532), .A(n3533), .B(n3653), .ZN(n3432)
         );
  NAND2_X1 U4157 ( .A1(n3925), .A2(n3911), .ZN(n3883) );
  OAI22_X1 U4158 ( .A1(n3863), .A2(n3883), .B1(n3895), .B2(n3913), .ZN(n3864)
         );
  NAND2_X1 U4159 ( .A1(n3950), .A2(n3687), .ZN(n3861) );
  OAI22_X1 U4160 ( .A1(n3863), .A2(n3861), .B1(n3568), .B2(n3874), .ZN(n3425)
         );
  OR2_X1 U4161 ( .A1(n3864), .A2(n3425), .ZN(n3427) );
  NAND2_X1 U4162 ( .A1(n3427), .A2(n3426), .ZN(n3809) );
  NAND2_X1 U4163 ( .A1(n3699), .A2(n3836), .ZN(n3812) );
  NAND2_X1 U4164 ( .A1(n3859), .A2(n3845), .ZN(n3811) );
  AND2_X1 U4165 ( .A1(n3812), .A2(n3811), .ZN(n3541) );
  INV_X1 U4166 ( .A(n3654), .ZN(n3431) );
  NOR2_X1 U4167 ( .A1(n3859), .A2(n3845), .ZN(n3537) );
  NAND2_X1 U4168 ( .A1(n3537), .A2(n3812), .ZN(n3430) );
  NAND2_X1 U4169 ( .A1(n3846), .A2(n3698), .ZN(n3478) );
  NAND2_X1 U4170 ( .A1(n3831), .A2(n3815), .ZN(n3428) );
  NAND2_X1 U4171 ( .A1(n3478), .A2(n3428), .ZN(n3539) );
  INV_X1 U4172 ( .A(n3539), .ZN(n3429) );
  OAI21_X1 U4173 ( .B1(n3432), .B2(n3431), .A(n3655), .ZN(n3433) );
  NAND2_X1 U4174 ( .A1(n3816), .A2(n3792), .ZN(n3454) );
  NAND2_X1 U4175 ( .A1(n3700), .A2(n3715), .ZN(n3788) );
  NAND2_X1 U4176 ( .A1(n3433), .A2(n3656), .ZN(n3438) );
  NAND2_X1 U4177 ( .A1(n3774), .A2(n3797), .ZN(n3769) );
  NAND2_X1 U4178 ( .A1(n3793), .A2(n3779), .ZN(n3451) );
  AND2_X1 U4179 ( .A1(n3769), .A2(n3451), .ZN(n3657) );
  AOI222_X1 U4180 ( .A1(n3435), .A2(REG1_REG_30__SCAN_IN), .B1(n3196), .B2(
        REG2_REG_30__SCAN_IN), .C1(n3434), .C2(REG0_REG_30__SCAN_IN), .ZN(
        n3667) );
  AOI222_X1 U4181 ( .A1(n3435), .A2(REG1_REG_31__SCAN_IN), .B1(n3196), .B2(
        REG2_REG_31__SCAN_IN), .C1(n3434), .C2(REG0_REG_31__SCAN_IN), .ZN(
        n4023) );
  INV_X1 U4182 ( .A(n4021), .ZN(n4024) );
  NOR2_X1 U4183 ( .A1(n4023), .A2(n4024), .ZN(n3549) );
  AOI21_X1 U4184 ( .B1(n3667), .B2(n4032), .A(n3549), .ZN(n3477) );
  OR2_X1 U4185 ( .A1(n3775), .A2(n3706), .ZN(n3449) );
  OR2_X1 U4186 ( .A1(n3793), .A2(n3779), .ZN(n3752) );
  NOR2_X1 U4187 ( .A1(n3669), .A2(n3731), .ZN(n3661) );
  AND2_X1 U4188 ( .A1(n3759), .A2(n3745), .ZN(n3660) );
  NOR2_X1 U4189 ( .A1(n3661), .A2(n3660), .ZN(n3440) );
  NAND2_X1 U4190 ( .A1(n3436), .A2(DATAI_29_), .ZN(n3712) );
  OR2_X1 U4191 ( .A1(n3725), .A2(n3712), .ZN(n3448) );
  NAND4_X1 U4192 ( .A1(n3477), .A2(n3659), .A3(n3440), .A4(n3448), .ZN(n3437)
         );
  AOI21_X1 U4193 ( .B1(n3438), .B2(n3657), .A(n3437), .ZN(n3443) );
  XNOR2_X1 U4194 ( .A(n3759), .B(n3708), .ZN(n3738) );
  AND2_X1 U4195 ( .A1(n3775), .A2(n3706), .ZN(n3658) );
  NAND2_X1 U4196 ( .A1(n3725), .A2(n3712), .ZN(n3447) );
  NAND2_X1 U4197 ( .A1(n3669), .A2(n3731), .ZN(n3662) );
  NAND2_X1 U4198 ( .A1(n3447), .A2(n3662), .ZN(n3439) );
  NOR2_X1 U4199 ( .A1(n3658), .A2(n3439), .ZN(n3544) );
  OAI211_X1 U4200 ( .C1(n3440), .C2(n3439), .A(n3477), .B(n3448), .ZN(n3550)
         );
  AOI21_X1 U4201 ( .B1(n3738), .B2(n3544), .A(n3550), .ZN(n3442) );
  INV_X1 U4202 ( .A(n3667), .ZN(n3567) );
  NAND2_X1 U4203 ( .A1(n3567), .A2(n4028), .ZN(n3445) );
  INV_X1 U4204 ( .A(n4023), .ZN(n3566) );
  AOI21_X1 U4205 ( .B1(n3445), .B2(n3566), .A(n4021), .ZN(n3441) );
  NOR3_X1 U4206 ( .A1(n3443), .A2(n3442), .A3(n3441), .ZN(n3444) );
  AOI21_X1 U4207 ( .B1(n4032), .B2(n4021), .A(n3444), .ZN(n3557) );
  INV_X1 U4208 ( .A(n3445), .ZN(n3446) );
  AOI21_X1 U4209 ( .B1(n4024), .B2(n4023), .A(n3446), .ZN(n3548) );
  INV_X1 U4210 ( .A(n3548), .ZN(n3457) );
  INV_X1 U4211 ( .A(n3449), .ZN(n3450) );
  NOR2_X1 U4212 ( .A1(n3450), .A2(n3658), .ZN(n3754) );
  AND2_X1 U4213 ( .A1(n3752), .A2(n3451), .ZN(n3771) );
  NAND4_X1 U4214 ( .A1(n3710), .A2(n3738), .A3(n3754), .A4(n3771), .ZN(n3456)
         );
  INV_X1 U4215 ( .A(n3874), .ZN(n3452) );
  INV_X1 U4216 ( .A(n3695), .ZN(n3453) );
  NAND2_X1 U4217 ( .A1(n3888), .A2(n3874), .ZN(n3694) );
  AND2_X1 U4218 ( .A1(n3453), .A2(n3694), .ZN(n3871) );
  NAND2_X1 U4219 ( .A1(n3913), .A2(n3714), .ZN(n3692) );
  NOR2_X1 U4220 ( .A1(n3913), .A2(n3714), .ZN(n3693) );
  OR2_X1 U4221 ( .A1(n2147), .A2(n3693), .ZN(n3886) );
  INV_X1 U4222 ( .A(n3886), .ZN(n3881) );
  XNOR2_X1 U4223 ( .A(n3831), .B(n3815), .ZN(n3814) );
  NAND2_X1 U4224 ( .A1(n3769), .A2(n3454), .ZN(n3790) );
  OR4_X1 U4225 ( .A1(n3871), .A2(n3881), .A3(n3814), .A4(n3790), .ZN(n3455) );
  NOR4_X1 U4226 ( .A1(n3457), .A2(n3491), .A3(n3456), .A4(n3455), .ZN(n3466)
         );
  NAND2_X1 U4227 ( .A1(n3861), .A2(n3860), .ZN(n3923) );
  INV_X1 U4228 ( .A(n3923), .ZN(n3465) );
  AND2_X1 U4229 ( .A1(n3459), .A2(n3458), .ZN(n3998) );
  NOR4_X1 U4230 ( .A1(n3463), .A2(n3462), .A3(n3461), .A4(n3460), .ZN(n3464)
         );
  NAND4_X1 U4231 ( .A1(n3466), .A2(n3465), .A3(n3998), .A4(n3464), .ZN(n3476)
         );
  NAND2_X1 U4232 ( .A1(n3883), .A2(n3884), .ZN(n3910) );
  INV_X1 U4233 ( .A(n3910), .ZN(n3470) );
  NAND2_X1 U4234 ( .A1(n3650), .A2(n3467), .ZN(n3977) );
  INV_X1 U4235 ( .A(n3977), .ZN(n3649) );
  NAND4_X1 U4236 ( .A1(n3470), .A2(n3649), .A3(n3469), .A4(n3468), .ZN(n3475)
         );
  NAND4_X1 U4237 ( .A1(n3473), .A2(n2179), .A3(n3472), .A4(n3471), .ZN(n3474)
         );
  NOR3_X1 U4238 ( .A1(n3476), .A2(n3475), .A3(n3474), .ZN(n3487) );
  INV_X1 U4239 ( .A(n3477), .ZN(n3480) );
  INV_X1 U4240 ( .A(n3811), .ZN(n3479) );
  OR2_X1 U4241 ( .A1(n3479), .A2(n3537), .ZN(n3850) );
  NOR4_X1 U4242 ( .A1(n3480), .A2(n3826), .A3(n3850), .A4(n4306), .ZN(n3486)
         );
  INV_X1 U4243 ( .A(n3662), .ZN(n3481) );
  NAND2_X1 U4244 ( .A1(n3532), .A2(n3652), .ZN(n3939) );
  NAND2_X1 U4245 ( .A1(n3482), .A2(n3651), .ZN(n3970) );
  NOR4_X1 U4246 ( .A1(n3939), .A2(n3484), .A3(n3970), .A4(n3483), .ZN(n3485)
         );
  NAND4_X1 U4247 ( .A1(n3487), .A2(n3486), .A3(n3722), .A4(n3485), .ZN(n3554)
         );
  INV_X1 U4248 ( .A(n3488), .ZN(n3492) );
  OAI211_X1 U4249 ( .C1(n3492), .C2(n3491), .A(n3490), .B(n3489), .ZN(n3494)
         );
  NAND3_X1 U4250 ( .A1(n3494), .A2(n3493), .A3(n2589), .ZN(n3497) );
  NAND3_X1 U4251 ( .A1(n3497), .A2(n3496), .A3(n3495), .ZN(n3500) );
  NAND3_X1 U4252 ( .A1(n3500), .A2(n3499), .A3(n3498), .ZN(n3503) );
  NAND4_X1 U4253 ( .A1(n3503), .A2(n3502), .A3(n3501), .A4(n3515), .ZN(n3506)
         );
  AND3_X1 U4254 ( .A1(n3506), .A2(n3505), .A3(n3504), .ZN(n3511) );
  NAND2_X1 U4255 ( .A1(n3508), .A2(n3507), .ZN(n3518) );
  OAI211_X1 U4256 ( .C1(n3511), .C2(n3518), .A(n3510), .B(n3509), .ZN(n3531)
         );
  NAND2_X1 U4257 ( .A1(n3513), .A2(n3512), .ZN(n3526) );
  NOR3_X1 U4258 ( .A1(n3526), .A2(n3517), .A3(n3514), .ZN(n3530) );
  INV_X1 U4259 ( .A(n3515), .ZN(n3519) );
  NOR4_X1 U4260 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3522)
         );
  INV_X1 U4261 ( .A(n3520), .ZN(n3521) );
  NOR2_X1 U4262 ( .A1(n3522), .A2(n3521), .ZN(n3527) );
  INV_X1 U4263 ( .A(n3523), .ZN(n3525) );
  OAI211_X1 U4264 ( .C1(n3527), .C2(n3526), .A(n3525), .B(n3524), .ZN(n3528)
         );
  AOI22_X1 U4265 ( .A1(n3531), .A2(n3530), .B1(n3529), .B2(n3528), .ZN(n3534)
         );
  OAI21_X1 U4266 ( .B1(n3534), .B2(n3533), .A(n3532), .ZN(n3536) );
  INV_X1 U4267 ( .A(n3809), .ZN(n3535) );
  AOI21_X1 U4268 ( .B1(n3536), .B2(n2065), .A(n3535), .ZN(n3538) );
  OR2_X1 U4269 ( .A1(n3538), .A2(n3537), .ZN(n3540) );
  AOI21_X1 U4270 ( .B1(n3541), .B2(n3540), .A(n3539), .ZN(n3543) );
  INV_X1 U4271 ( .A(n3656), .ZN(n3542) );
  OAI21_X1 U4272 ( .B1(n3543), .B2(n3542), .A(n3657), .ZN(n3547) );
  NOR2_X1 U4273 ( .A1(n3759), .A2(n3745), .ZN(n3546) );
  INV_X1 U4274 ( .A(n3544), .ZN(n3545) );
  AOI211_X1 U4275 ( .C1(n3659), .C2(n3547), .A(n3546), .B(n3545), .ZN(n3551)
         );
  OAI22_X1 U4276 ( .A1(n3551), .A2(n3550), .B1(n3549), .B2(n3548), .ZN(n3553)
         );
  MUX2_X1 U4277 ( .A(n3554), .B(n3553), .S(n3552), .Z(n3555) );
  OAI21_X1 U4278 ( .B1(n3557), .B2(n3556), .A(n3555), .ZN(n3558) );
  XNOR2_X1 U4279 ( .A(n3558), .B(n4171), .ZN(n3565) );
  INV_X1 U4280 ( .A(n3559), .ZN(n3582) );
  NAND2_X1 U4281 ( .A1(n3560), .A2(n3582), .ZN(n3561) );
  OAI211_X1 U4282 ( .C1(n3562), .C2(n3564), .A(n3561), .B(B_REG_SCAN_IN), .ZN(
        n3563) );
  OAI21_X1 U4283 ( .B1(n3565), .B2(n3564), .A(n3563), .ZN(U3239) );
  MUX2_X1 U4284 ( .A(DATAO_REG_31__SCAN_IN), .B(n3566), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4285 ( .A(DATAO_REG_30__SCAN_IN), .B(n3567), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4286 ( .A(n3725), .B(DATAO_REG_29__SCAN_IN), .S(n3573), .Z(U3579)
         );
  MUX2_X1 U4287 ( .A(n3669), .B(DATAO_REG_28__SCAN_IN), .S(n3573), .Z(U3578)
         );
  MUX2_X1 U4288 ( .A(n3726), .B(DATAO_REG_27__SCAN_IN), .S(n3573), .Z(U3577)
         );
  MUX2_X1 U4289 ( .A(n3775), .B(DATAO_REG_26__SCAN_IN), .S(n3573), .Z(U3576)
         );
  MUX2_X1 U4290 ( .A(n3793), .B(DATAO_REG_25__SCAN_IN), .S(n3573), .Z(U3575)
         );
  MUX2_X1 U4291 ( .A(n3774), .B(DATAO_REG_24__SCAN_IN), .S(n3573), .Z(U3574)
         );
  MUX2_X1 U4292 ( .A(n3831), .B(DATAO_REG_23__SCAN_IN), .S(n3573), .Z(U3573)
         );
  MUX2_X1 U4293 ( .A(n3846), .B(DATAO_REG_22__SCAN_IN), .S(n3573), .Z(U3572)
         );
  INV_X1 U4294 ( .A(n3859), .ZN(n3696) );
  MUX2_X1 U4295 ( .A(n3696), .B(DATAO_REG_21__SCAN_IN), .S(n3573), .Z(U3571)
         );
  MUX2_X1 U4296 ( .A(n3568), .B(DATAO_REG_20__SCAN_IN), .S(n3573), .Z(U3570)
         );
  MUX2_X1 U4297 ( .A(n3890), .B(DATAO_REG_18__SCAN_IN), .S(n3573), .Z(U3568)
         );
  MUX2_X1 U4298 ( .A(n3688), .B(DATAO_REG_17__SCAN_IN), .S(n3573), .Z(U3567)
         );
  MUX2_X1 U4299 ( .A(n3927), .B(DATAO_REG_16__SCAN_IN), .S(n3573), .Z(U3566)
         );
  MUX2_X1 U4300 ( .A(n3963), .B(DATAO_REG_14__SCAN_IN), .S(n3573), .Z(U3564)
         );
  MUX2_X1 U4301 ( .A(n3981), .B(DATAO_REG_13__SCAN_IN), .S(n3573), .Z(U3563)
         );
  MUX2_X1 U4302 ( .A(n4005), .B(DATAO_REG_12__SCAN_IN), .S(n3573), .Z(U3562)
         );
  MUX2_X1 U4303 ( .A(n3569), .B(DATAO_REG_11__SCAN_IN), .S(n3573), .Z(U3561)
         );
  MUX2_X1 U4304 ( .A(n3570), .B(DATAO_REG_10__SCAN_IN), .S(n3573), .Z(U3560)
         );
  MUX2_X1 U4305 ( .A(n3571), .B(DATAO_REG_9__SCAN_IN), .S(n3573), .Z(U3559) );
  MUX2_X1 U4306 ( .A(n3572), .B(DATAO_REG_8__SCAN_IN), .S(n3573), .Z(U3558) );
  MUX2_X1 U4307 ( .A(n3574), .B(DATAO_REG_6__SCAN_IN), .S(n3573), .Z(U3556) );
  MUX2_X1 U4308 ( .A(n3575), .B(DATAO_REG_5__SCAN_IN), .S(n3573), .Z(U3555) );
  MUX2_X1 U4309 ( .A(n3576), .B(DATAO_REG_4__SCAN_IN), .S(n3573), .Z(U3554) );
  MUX2_X1 U4310 ( .A(n3577), .B(DATAO_REG_2__SCAN_IN), .S(n3573), .Z(U3552) );
  MUX2_X1 U4311 ( .A(n2572), .B(DATAO_REG_1__SCAN_IN), .S(n3573), .Z(U3551) );
  MUX2_X1 U4312 ( .A(n3578), .B(DATAO_REG_0__SCAN_IN), .S(n3573), .Z(U3550) );
  AOI21_X1 U4313 ( .B1(n4186), .B2(n2347), .A(n3579), .ZN(n4187) );
  NAND3_X1 U4314 ( .A1(n3580), .A2(n4168), .A3(n3665), .ZN(n3584) );
  AOI21_X1 U4315 ( .B1(n3582), .B2(n3581), .A(n3573), .ZN(n3583) );
  OAI211_X1 U4316 ( .C1(IR_REG_0__SCAN_IN), .C2(n4187), .A(n3584), .B(n3583), 
        .ZN(n4202) );
  AOI22_X1 U4317 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4268), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3598) );
  XNOR2_X1 U4318 ( .A(n3586), .B(n3585), .ZN(n3588) );
  OAI22_X1 U4319 ( .A1(n3588), .A2(n4256), .B1(n4281), .B2(n3587), .ZN(n3589)
         );
  INV_X1 U4320 ( .A(n3589), .ZN(n3597) );
  MUX2_X1 U4321 ( .A(n2349), .B(REG2_REG_2__SCAN_IN), .S(n4176), .Z(n3592) );
  INV_X1 U4322 ( .A(n3590), .ZN(n3591) );
  NAND2_X1 U4323 ( .A1(n3592), .A2(n3591), .ZN(n3594) );
  OAI211_X1 U4324 ( .C1(n3595), .C2(n3594), .A(n4278), .B(n3593), .ZN(n3596)
         );
  NAND4_X1 U4325 ( .A1(n4202), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(U3242)
         );
  INV_X1 U4326 ( .A(n4315), .ZN(n4266) );
  AOI22_X1 U4327 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4266), .B1(n4315), .B2(
        n3602), .ZN(n4258) );
  XNOR2_X1 U4328 ( .A(n3627), .B(n4173), .ZN(n3604) );
  NAND2_X1 U4329 ( .A1(n3604), .A2(n3603), .ZN(n3628) );
  OAI21_X1 U4330 ( .B1(n3604), .B2(n3603), .A(n3628), .ZN(n3605) );
  NAND2_X1 U4331 ( .A1(n3605), .A2(n4276), .ZN(n3618) );
  INV_X1 U4332 ( .A(n3606), .ZN(n3607) );
  AOI21_X1 U4333 ( .B1(n4268), .B2(ADDR_REG_16__SCAN_IN), .A(n3607), .ZN(n3617) );
  AND2_X1 U4334 ( .A1(n3608), .A2(REG2_REG_13__SCAN_IN), .ZN(n3609) );
  OAI22_X1 U4335 ( .A1(n3609), .A2(n4174), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3608), .ZN(n3610) );
  NOR2_X1 U4336 ( .A1(n4317), .A2(n3610), .ZN(n3611) );
  INV_X1 U4337 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4248) );
  INV_X1 U4338 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4490) );
  AOI22_X1 U4339 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4266), .B1(n4315), .B2(
        n4490), .ZN(n4262) );
  AND2_X1 U4340 ( .A1(n4315), .A2(REG2_REG_15__SCAN_IN), .ZN(n3612) );
  XNOR2_X1 U4341 ( .A(n3620), .B(n4173), .ZN(n3613) );
  INV_X1 U4342 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4491) );
  NAND2_X1 U4343 ( .A1(n3613), .A2(n4491), .ZN(n3621) );
  OAI21_X1 U4344 ( .B1(n3613), .B2(n4491), .A(n3621), .ZN(n3614) );
  NAND2_X1 U4345 ( .A1(n3614), .A2(n4278), .ZN(n3616) );
  NAND2_X1 U4346 ( .A1(n4252), .A2(n4173), .ZN(n3615) );
  NAND4_X1 U4347 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(U3256)
         );
  INV_X1 U4348 ( .A(n4172), .ZN(n3634) );
  XNOR2_X1 U4349 ( .A(n4172), .B(REG2_REG_18__SCAN_IN), .ZN(n3624) );
  INV_X1 U4350 ( .A(n4282), .ZN(n4313) );
  NOR2_X1 U4351 ( .A1(n4313), .A2(REG2_REG_17__SCAN_IN), .ZN(n3619) );
  AOI21_X1 U4352 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4313), .A(n3619), .ZN(n4271) );
  INV_X1 U4353 ( .A(n4173), .ZN(n3626) );
  NAND2_X1 U4354 ( .A1(n3620), .A2(n3626), .ZN(n3622) );
  AOI21_X1 U4355 ( .B1(n3624), .B2(n3623), .A(n3638), .ZN(n3625) );
  NAND2_X1 U4356 ( .A1(n4278), .A2(n3625), .ZN(n3633) );
  XNOR2_X1 U4357 ( .A(n4172), .B(REG1_REG_18__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4358 ( .A1(n4313), .A2(REG1_REG_17__SCAN_IN), .B1(n4083), .B2(
        n4282), .ZN(n4274) );
  NAND2_X1 U4359 ( .A1(n3627), .A2(n3626), .ZN(n3629) );
  NAND2_X1 U4360 ( .A1(n3629), .A2(n3628), .ZN(n4273) );
  OAI211_X1 U4361 ( .C1(n3634), .C2(n4281), .A(n3633), .B(n3632), .ZN(U3258)
         );
  XNOR2_X1 U4362 ( .A(n4171), .B(REG1_REG_19__SCAN_IN), .ZN(n3636) );
  XNOR2_X1 U4363 ( .A(n3637), .B(n3636), .ZN(n3647) );
  INV_X1 U4364 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4493) );
  MUX2_X1 U4365 ( .A(REG2_REG_19__SCAN_IN), .B(n4493), .S(n4171), .Z(n3639) );
  XNOR2_X1 U4366 ( .A(n3640), .B(n3639), .ZN(n3645) );
  NAND2_X1 U4367 ( .A1(n4268), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3642) );
  OAI211_X1 U4368 ( .C1(n4281), .C2(n3643), .A(n3642), .B(n3641), .ZN(n3644)
         );
  AOI21_X1 U4369 ( .B1(n3645), .B2(n4278), .A(n3644), .ZN(n3646) );
  OAI21_X1 U4370 ( .B1(n3647), .B2(n4256), .A(n3646), .ZN(U3259) );
  INV_X1 U4371 ( .A(n3648), .ZN(n3672) );
  INV_X1 U4372 ( .A(n3939), .ZN(n3947) );
  NAND2_X1 U4373 ( .A1(n3948), .A2(n3947), .ZN(n3946) );
  NAND2_X1 U4374 ( .A1(n3789), .A2(n3656), .ZN(n3770) );
  AOI21_X1 U4375 ( .B1(n3663), .B2(n3662), .A(n3661), .ZN(n3664) );
  XNOR2_X1 U4376 ( .A(n3664), .B(n3710), .ZN(n3671) );
  INV_X1 U4377 ( .A(B_REG_SCAN_IN), .ZN(n3666) );
  OAI21_X1 U4378 ( .B1(n3666), .B2(n3665), .A(n3912), .ZN(n4022) );
  OAI22_X1 U4379 ( .A1(n3667), .A2(n4022), .B1(n3712), .B2(n4001), .ZN(n3668)
         );
  AOI21_X1 U4380 ( .B1(n3669), .B2(n4006), .A(n3668), .ZN(n3670) );
  OAI21_X1 U4381 ( .B1(n3671), .B2(n4010), .A(n3670), .ZN(n4035) );
  AOI21_X1 U4382 ( .B1(n3672), .B2(n4292), .A(n4035), .ZN(n3719) );
  NAND2_X1 U4383 ( .A1(n4005), .A2(n3673), .ZN(n3675) );
  NOR2_X1 U4384 ( .A1(n4005), .A2(n3673), .ZN(n3674) );
  NAND2_X1 U4385 ( .A1(n3677), .A2(n4011), .ZN(n3680) );
  NAND2_X1 U4386 ( .A1(n3683), .A2(n3713), .ZN(n3685) );
  NAND2_X1 U4387 ( .A1(n3938), .A2(n3686), .ZN(n3922) );
  NAND2_X1 U4388 ( .A1(n3950), .A2(n3930), .ZN(n3690) );
  AOI21_X1 U4389 ( .B1(n3922), .B2(n3690), .A(n3689), .ZN(n3901) );
  NAND2_X1 U4390 ( .A1(n3901), .A2(n3910), .ZN(n3902) );
  NAND2_X1 U4391 ( .A1(n3696), .A2(n3845), .ZN(n3697) );
  NAND2_X1 U4392 ( .A1(n3827), .A2(n3826), .ZN(n3825) );
  NAND2_X1 U4393 ( .A1(n3825), .A2(n2220), .ZN(n3808) );
  NAND2_X1 U4394 ( .A1(n3700), .A2(n3815), .ZN(n3701) );
  NAND2_X1 U4395 ( .A1(n3774), .A2(n3792), .ZN(n3703) );
  NAND2_X1 U4396 ( .A1(n3704), .A2(n3779), .ZN(n3705) );
  NAND2_X1 U4397 ( .A1(n3775), .A2(n3760), .ZN(n3707) );
  NAND2_X1 U4398 ( .A1(n3759), .A2(n3708), .ZN(n3709) );
  XNOR2_X1 U4399 ( .A(n3711), .B(n3710), .ZN(n4034) );
  NAND2_X1 U4400 ( .A1(n4034), .A2(n3972), .ZN(n3718) );
  INV_X1 U4401 ( .A(n3712), .ZN(n3716) );
  AOI22_X1 U4402 ( .A1(n4036), .A2(n4294), .B1(REG2_REG_29__SCAN_IN), .B2(
        n2000), .ZN(n3717) );
  OAI211_X1 U4403 ( .C1(n2000), .C2(n3719), .A(n3718), .B(n3717), .ZN(U3354)
         );
  XNOR2_X1 U4404 ( .A(n3721), .B(n3720), .ZN(n4039) );
  INV_X1 U4405 ( .A(n4039), .ZN(n3736) );
  XNOR2_X1 U4406 ( .A(n3723), .B(n3722), .ZN(n3729) );
  INV_X1 U4407 ( .A(n3731), .ZN(n3724) );
  AOI22_X1 U4408 ( .A1(n3725), .A2(n3912), .B1(n4031), .B2(n3724), .ZN(n3728)
         );
  NAND2_X1 U4409 ( .A1(n3726), .A2(n4006), .ZN(n3727) );
  OAI211_X1 U4410 ( .C1(n3729), .C2(n4010), .A(n3728), .B(n3727), .ZN(n4038)
         );
  OAI21_X1 U4411 ( .B1(n3744), .B2(n3731), .A(n3730), .ZN(n4120) );
  AOI22_X1 U4412 ( .A1(n3732), .A2(n4292), .B1(REG2_REG_28__SCAN_IN), .B2(
        n2000), .ZN(n3733) );
  OAI21_X1 U4413 ( .B1(n4120), .B2(n4015), .A(n3733), .ZN(n3734) );
  AOI21_X1 U4414 ( .B1(n4038), .B2(n4284), .A(n3734), .ZN(n3735) );
  OAI21_X1 U4415 ( .B1(n3736), .B2(n3991), .A(n3735), .ZN(U3262) );
  XOR2_X1 U4416 ( .A(n3738), .B(n3737), .Z(n4045) );
  XNOR2_X1 U4417 ( .A(n3739), .B(n3738), .ZN(n3740) );
  NAND2_X1 U4418 ( .A1(n3740), .A2(n3945), .ZN(n3742) );
  AOI22_X1 U4419 ( .A1(n3775), .A2(n4006), .B1(n3745), .B2(n4031), .ZN(n3741)
         );
  OAI211_X1 U4420 ( .C1(n3743), .C2(n4002), .A(n3742), .B(n3741), .ZN(n4042)
         );
  AOI21_X1 U4421 ( .B1(n3745), .B2(n3762), .A(n3744), .ZN(n4043) );
  INV_X1 U4422 ( .A(n4043), .ZN(n3748) );
  AOI22_X1 U4423 ( .A1(n3746), .A2(n4292), .B1(n2000), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n3747) );
  OAI21_X1 U4424 ( .B1(n3748), .B2(n4015), .A(n3747), .ZN(n3749) );
  AOI21_X1 U4425 ( .B1(n4042), .B2(n4284), .A(n3749), .ZN(n3750) );
  OAI21_X1 U4426 ( .B1(n4045), .B2(n3991), .A(n3750), .ZN(U3263) );
  XOR2_X1 U4427 ( .A(n3754), .B(n3751), .Z(n4047) );
  INV_X1 U4428 ( .A(n4047), .ZN(n3767) );
  NAND2_X1 U4429 ( .A1(n3753), .A2(n3752), .ZN(n3755) );
  XNOR2_X1 U4430 ( .A(n3755), .B(n3754), .ZN(n3756) );
  NAND2_X1 U4431 ( .A1(n3756), .A2(n3945), .ZN(n3758) );
  AOI22_X1 U4432 ( .A1(n3793), .A2(n4006), .B1(n3760), .B2(n4031), .ZN(n3757)
         );
  OAI211_X1 U4433 ( .C1(n3759), .C2(n4002), .A(n3758), .B(n3757), .ZN(n4046)
         );
  NAND2_X1 U4434 ( .A1(n3781), .A2(n3760), .ZN(n3761) );
  NAND2_X1 U4435 ( .A1(n3762), .A2(n3761), .ZN(n4125) );
  AOI22_X1 U4436 ( .A1(REG2_REG_26__SCAN_IN), .A2(n2000), .B1(n3763), .B2(
        n4292), .ZN(n3764) );
  OAI21_X1 U4437 ( .B1(n4125), .B2(n4015), .A(n3764), .ZN(n3765) );
  AOI21_X1 U4438 ( .B1(n4284), .B2(n4046), .A(n3765), .ZN(n3766) );
  OAI21_X1 U4439 ( .B1(n3767), .B2(n3991), .A(n3766), .ZN(U3264) );
  XNOR2_X1 U4440 ( .A(n3768), .B(n3771), .ZN(n4050) );
  INV_X1 U4441 ( .A(n4050), .ZN(n3786) );
  NAND2_X1 U4442 ( .A1(n3770), .A2(n3769), .ZN(n3772) );
  XNOR2_X1 U4443 ( .A(n3772), .B(n3771), .ZN(n3778) );
  AOI22_X1 U4444 ( .A1(n3774), .A2(n4006), .B1(n3773), .B2(n4031), .ZN(n3777)
         );
  NAND2_X1 U4445 ( .A1(n3775), .A2(n3912), .ZN(n3776) );
  OAI211_X1 U4446 ( .C1(n3778), .C2(n4010), .A(n3777), .B(n3776), .ZN(n4049)
         );
  OR2_X1 U4447 ( .A1(n3799), .A2(n3779), .ZN(n3780) );
  NAND2_X1 U4448 ( .A1(n3781), .A2(n3780), .ZN(n4128) );
  AOI22_X1 U4449 ( .A1(n2000), .A2(REG2_REG_25__SCAN_IN), .B1(n3782), .B2(
        n4292), .ZN(n3783) );
  OAI21_X1 U4450 ( .B1(n4128), .B2(n4015), .A(n3783), .ZN(n3784) );
  AOI21_X1 U4451 ( .B1(n4049), .B2(n4284), .A(n3784), .ZN(n3785) );
  OAI21_X1 U4452 ( .B1(n3786), .B2(n3991), .A(n3785), .ZN(U3265) );
  XNOR2_X1 U4453 ( .A(n3787), .B(n3790), .ZN(n4054) );
  INV_X1 U4454 ( .A(n4054), .ZN(n3804) );
  NAND2_X1 U4455 ( .A1(n3789), .A2(n3788), .ZN(n3791) );
  XNOR2_X1 U4456 ( .A(n3791), .B(n3790), .ZN(n3796) );
  AOI22_X1 U4457 ( .A1(n3831), .A2(n4006), .B1(n3792), .B2(n4031), .ZN(n3795)
         );
  NAND2_X1 U4458 ( .A1(n3793), .A2(n3912), .ZN(n3794) );
  OAI211_X1 U4459 ( .C1(n3796), .C2(n4010), .A(n3795), .B(n3794), .ZN(n4053)
         );
  NOR2_X1 U4460 ( .A1(n3805), .A2(n3797), .ZN(n3798) );
  OR2_X1 U4461 ( .A1(n3799), .A2(n3798), .ZN(n4131) );
  AOI22_X1 U4462 ( .A1(n2000), .A2(REG2_REG_24__SCAN_IN), .B1(n3800), .B2(
        n4292), .ZN(n3801) );
  OAI21_X1 U4463 ( .B1(n4131), .B2(n4015), .A(n3801), .ZN(n3802) );
  AOI21_X1 U4464 ( .B1(n4053), .B2(n4284), .A(n3802), .ZN(n3803) );
  OAI21_X1 U4465 ( .B1(n3804), .B2(n3991), .A(n3803), .ZN(U3266) );
  INV_X1 U4466 ( .A(n4061), .ZN(n3807) );
  INV_X1 U4467 ( .A(n3805), .ZN(n3806) );
  OAI21_X1 U4468 ( .B1(n3807), .B2(n3815), .A(n3806), .ZN(n4134) );
  XOR2_X1 U4469 ( .A(n3814), .B(n3808), .Z(n4058) );
  NAND2_X1 U4470 ( .A1(n4058), .A2(n3972), .ZN(n3824) );
  NAND2_X1 U4471 ( .A1(n3810), .A2(n3809), .ZN(n3843) );
  INV_X1 U4472 ( .A(n3850), .ZN(n3844) );
  NAND2_X1 U4473 ( .A1(n3843), .A2(n3844), .ZN(n3842) );
  NAND2_X1 U4474 ( .A1(n3811), .A2(n3842), .ZN(n3829) );
  NAND2_X1 U4475 ( .A1(n3830), .A2(n3829), .ZN(n3828) );
  NAND2_X1 U4476 ( .A1(n3812), .A2(n3828), .ZN(n3813) );
  XNOR2_X1 U4477 ( .A(n3814), .B(n3813), .ZN(n3819) );
  OAI22_X1 U4478 ( .A1(n3816), .A2(n4002), .B1(n4001), .B2(n3815), .ZN(n3817)
         );
  AOI21_X1 U4479 ( .B1(n4006), .B2(n3846), .A(n3817), .ZN(n3818) );
  OAI21_X1 U4480 ( .B1(n3819), .B2(n4010), .A(n3818), .ZN(n4057) );
  INV_X1 U4481 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3821) );
  OAI22_X1 U4482 ( .A1(n4284), .A2(n3821), .B1(n3820), .B2(n4304), .ZN(n3822)
         );
  AOI21_X1 U4483 ( .B1(n4057), .B2(n4284), .A(n3822), .ZN(n3823) );
  OAI211_X1 U4484 ( .C1(n4134), .C2(n4015), .A(n3824), .B(n3823), .ZN(U3267)
         );
  OAI21_X1 U4485 ( .B1(n3827), .B2(n3826), .A(n3825), .ZN(n4064) );
  OAI21_X1 U4486 ( .B1(n3830), .B2(n3829), .A(n3828), .ZN(n3835) );
  NAND2_X1 U4487 ( .A1(n3831), .A2(n3912), .ZN(n3833) );
  NAND2_X1 U4488 ( .A1(n3836), .A2(n4031), .ZN(n3832) );
  OAI211_X1 U4489 ( .C1(n3859), .C2(n3954), .A(n3833), .B(n3832), .ZN(n3834)
         );
  AOI21_X1 U4490 ( .B1(n3835), .B2(n3945), .A(n3834), .ZN(n4063) );
  NAND2_X1 U4491 ( .A1(n2001), .A2(n3836), .ZN(n4060) );
  NAND3_X1 U4492 ( .A1(n4061), .A2(n4294), .A3(n4060), .ZN(n3839) );
  AOI22_X1 U4493 ( .A1(n2000), .A2(REG2_REG_22__SCAN_IN), .B1(n3837), .B2(
        n4292), .ZN(n3838) );
  OAI211_X1 U4494 ( .C1(n2000), .C2(n4063), .A(n3839), .B(n3838), .ZN(n3840)
         );
  INV_X1 U4495 ( .A(n3840), .ZN(n3841) );
  OAI21_X1 U4496 ( .B1(n4064), .B2(n3991), .A(n3841), .ZN(U3268) );
  OAI21_X1 U4497 ( .B1(n3844), .B2(n3843), .A(n3842), .ZN(n3849) );
  AOI22_X1 U4498 ( .A1(n3846), .A2(n3912), .B1(n4031), .B2(n3845), .ZN(n3847)
         );
  OAI21_X1 U4499 ( .B1(n3888), .B2(n3954), .A(n3847), .ZN(n3848) );
  AOI21_X1 U4500 ( .B1(n3849), .B2(n3945), .A(n3848), .ZN(n4066) );
  XNOR2_X1 U4501 ( .A(n3851), .B(n3850), .ZN(n4065) );
  NAND2_X1 U4502 ( .A1(n4065), .A2(n3972), .ZN(n3858) );
  OAI21_X1 U4503 ( .B1(n3872), .B2(n3852), .A(n2001), .ZN(n4068) );
  INV_X1 U4504 ( .A(n4068), .ZN(n3856) );
  INV_X1 U4505 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3854) );
  OAI22_X1 U4506 ( .A1(n4284), .A2(n3854), .B1(n3853), .B2(n4304), .ZN(n3855)
         );
  AOI21_X1 U4507 ( .B1(n3856), .B2(n4294), .A(n3855), .ZN(n3857) );
  OAI211_X1 U4508 ( .C1(n2000), .C2(n4066), .A(n3858), .B(n3857), .ZN(U3269)
         );
  OAI22_X1 U4509 ( .A1(n3859), .A2(n4002), .B1(n3874), .B2(n4001), .ZN(n3869)
         );
  INV_X1 U4510 ( .A(n3860), .ZN(n3862) );
  OAI21_X1 U4511 ( .B1(n3924), .B2(n3862), .A(n3861), .ZN(n3909) );
  INV_X1 U4512 ( .A(n3863), .ZN(n3865) );
  AOI21_X1 U4513 ( .B1(n3909), .B2(n3865), .A(n3864), .ZN(n3866) );
  XOR2_X1 U4514 ( .A(n3871), .B(n3866), .Z(n3867) );
  NOR2_X1 U4515 ( .A1(n3867), .A2(n4010), .ZN(n3868) );
  AOI211_X1 U4516 ( .C1(n4006), .C2(n3913), .A(n3869), .B(n3868), .ZN(n4069)
         );
  XOR2_X1 U4517 ( .A(n3871), .B(n3870), .Z(n4071) );
  NAND2_X1 U4518 ( .A1(n4071), .A2(n3972), .ZN(n3880) );
  INV_X1 U4519 ( .A(n3872), .ZN(n3873) );
  OAI21_X1 U4520 ( .B1(n3893), .B2(n3874), .A(n3873), .ZN(n4139) );
  INV_X1 U4521 ( .A(n4139), .ZN(n3878) );
  INV_X1 U4522 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3876) );
  OAI22_X1 U4523 ( .A1(n4284), .A2(n3876), .B1(n3875), .B2(n4304), .ZN(n3877)
         );
  AOI21_X1 U4524 ( .B1(n3878), .B2(n4294), .A(n3877), .ZN(n3879) );
  OAI211_X1 U4525 ( .C1(n2000), .C2(n4069), .A(n3880), .B(n3879), .ZN(U3270)
         );
  XNOR2_X1 U4526 ( .A(n3882), .B(n3881), .ZN(n4075) );
  INV_X1 U4527 ( .A(n4075), .ZN(n3900) );
  INV_X1 U4528 ( .A(n3883), .ZN(n3885) );
  OAI21_X1 U4529 ( .B1(n3909), .B2(n3885), .A(n3884), .ZN(n3887) );
  XNOR2_X1 U4530 ( .A(n3887), .B(n3886), .ZN(n3892) );
  OAI22_X1 U4531 ( .A1(n3888), .A2(n4002), .B1(n3895), .B2(n4001), .ZN(n3889)
         );
  AOI21_X1 U4532 ( .B1(n4006), .B2(n3890), .A(n3889), .ZN(n3891) );
  OAI21_X1 U4533 ( .B1(n3892), .B2(n4010), .A(n3891), .ZN(n4074) );
  INV_X1 U4534 ( .A(n3893), .ZN(n3894) );
  OAI21_X1 U4535 ( .B1(n2099), .B2(n3895), .A(n3894), .ZN(n4143) );
  AOI22_X1 U4536 ( .A1(n2000), .A2(REG2_REG_19__SCAN_IN), .B1(n3896), .B2(
        n4292), .ZN(n3897) );
  OAI21_X1 U4537 ( .B1(n4143), .B2(n4015), .A(n3897), .ZN(n3898) );
  AOI21_X1 U4538 ( .B1(n4074), .B2(n4284), .A(n3898), .ZN(n3899) );
  OAI21_X1 U4539 ( .B1(n3900), .B2(n3991), .A(n3899), .ZN(U3271) );
  OAI21_X1 U4540 ( .B1(n3901), .B2(n3910), .A(n3902), .ZN(n3903) );
  INV_X1 U4541 ( .A(n3903), .ZN(n4080) );
  INV_X1 U4542 ( .A(n3932), .ZN(n3906) );
  OAI211_X1 U4543 ( .C1(n3906), .C2(n3905), .A(n4356), .B(n3904), .ZN(n4078)
         );
  INV_X1 U4544 ( .A(n4078), .ZN(n3920) );
  INV_X1 U4545 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3908) );
  OAI22_X1 U4546 ( .A1(n4284), .A2(n3908), .B1(n3907), .B2(n4304), .ZN(n3918)
         );
  XOR2_X1 U4547 ( .A(n3910), .B(n3909), .Z(n3916) );
  AOI22_X1 U4548 ( .A1(n3913), .A2(n3912), .B1(n4031), .B2(n3911), .ZN(n3914)
         );
  OAI21_X1 U4549 ( .B1(n3950), .B2(n3954), .A(n3914), .ZN(n3915) );
  AOI21_X1 U4550 ( .B1(n3916), .B2(n3945), .A(n3915), .ZN(n4079) );
  NOR2_X1 U4551 ( .A1(n4079), .A2(n2000), .ZN(n3917) );
  AOI211_X1 U4552 ( .C1(n3920), .C2(n3919), .A(n3918), .B(n3917), .ZN(n3921)
         );
  OAI21_X1 U4553 ( .B1(n4080), .B2(n3991), .A(n3921), .ZN(U3272) );
  XOR2_X1 U4554 ( .A(n3923), .B(n3922), .Z(n4082) );
  INV_X1 U4555 ( .A(n4082), .ZN(n3937) );
  XOR2_X1 U4556 ( .A(n3924), .B(n3923), .Z(n3929) );
  OAI22_X1 U4557 ( .A1(n3925), .A2(n4002), .B1(n4001), .B2(n3930), .ZN(n3926)
         );
  AOI21_X1 U4558 ( .B1(n4006), .B2(n3927), .A(n3926), .ZN(n3928) );
  OAI21_X1 U4559 ( .B1(n3929), .B2(n4010), .A(n3928), .ZN(n4081) );
  OR2_X1 U4560 ( .A1(n3941), .A2(n3930), .ZN(n3931) );
  NAND2_X1 U4561 ( .A1(n3932), .A2(n3931), .ZN(n4148) );
  NOR2_X1 U4562 ( .A1(n4148), .A2(n4015), .ZN(n3935) );
  OAI22_X1 U4563 ( .A1(n4284), .A2(n2103), .B1(n3933), .B2(n4304), .ZN(n3934)
         );
  AOI211_X1 U4564 ( .C1(n4081), .C2(n4284), .A(n3935), .B(n3934), .ZN(n3936)
         );
  OAI21_X1 U4565 ( .B1(n3937), .B2(n3991), .A(n3936), .ZN(U3273) );
  OAI21_X1 U4566 ( .B1(n3940), .B2(n3939), .A(n3938), .ZN(n4088) );
  AOI21_X1 U4567 ( .B1(n3942), .B2(n3964), .A(n3941), .ZN(n4086) );
  OAI22_X1 U4568 ( .A1(n4284), .A2(n4491), .B1(n3943), .B2(n4304), .ZN(n3944)
         );
  AOI21_X1 U4569 ( .B1(n4086), .B2(n4294), .A(n3944), .ZN(n3956) );
  OAI211_X1 U4570 ( .C1(n3948), .C2(n3947), .A(n3946), .B(n3945), .ZN(n3953)
         );
  OAI22_X1 U4571 ( .A1(n3950), .A2(n4002), .B1(n3949), .B2(n4001), .ZN(n3951)
         );
  INV_X1 U4572 ( .A(n3951), .ZN(n3952) );
  OAI211_X1 U4573 ( .C1(n3979), .C2(n3954), .A(n3953), .B(n3952), .ZN(n4085)
         );
  NAND2_X1 U4574 ( .A1(n4085), .A2(n4284), .ZN(n3955) );
  OAI211_X1 U4575 ( .C1(n4088), .C2(n3991), .A(n3956), .B(n3955), .ZN(U3274)
         );
  OAI22_X1 U4576 ( .A1(n3957), .A2(n4002), .B1(n3965), .B2(n4001), .ZN(n3962)
         );
  INV_X1 U4577 ( .A(n3958), .ZN(n3959) );
  AOI211_X1 U4578 ( .C1(n3960), .C2(n3970), .A(n4010), .B(n3959), .ZN(n3961)
         );
  AOI211_X1 U4579 ( .C1(n4006), .C2(n3963), .A(n3962), .B(n3961), .ZN(n4091)
         );
  INV_X1 U4580 ( .A(n3986), .ZN(n3966) );
  OAI21_X1 U4581 ( .B1(n3966), .B2(n3965), .A(n3964), .ZN(n4092) );
  INV_X1 U4582 ( .A(n4092), .ZN(n3969) );
  OAI22_X1 U4583 ( .A1(n4284), .A2(n4490), .B1(n3967), .B2(n4304), .ZN(n3968)
         );
  AOI21_X1 U4584 ( .B1(n3969), .B2(n4294), .A(n3968), .ZN(n3974) );
  XNOR2_X1 U4585 ( .A(n3971), .B(n3970), .ZN(n4089) );
  NAND2_X1 U4586 ( .A1(n4089), .A2(n3972), .ZN(n3973) );
  OAI211_X1 U4587 ( .C1(n4091), .C2(n2000), .A(n3974), .B(n3973), .ZN(U3275)
         );
  OAI21_X1 U4588 ( .B1(n3976), .B2(n3977), .A(n3975), .ZN(n4095) );
  INV_X1 U4589 ( .A(n4095), .ZN(n3992) );
  XNOR2_X1 U4590 ( .A(n3978), .B(n3977), .ZN(n3983) );
  OAI22_X1 U4591 ( .A1(n3979), .A2(n4002), .B1(n3681), .B2(n4001), .ZN(n3980)
         );
  AOI21_X1 U4592 ( .B1(n4006), .B2(n3981), .A(n3980), .ZN(n3982) );
  OAI21_X1 U4593 ( .B1(n3983), .B2(n4010), .A(n3982), .ZN(n4094) );
  NAND2_X1 U4594 ( .A1(n4014), .A2(n3984), .ZN(n3985) );
  NAND2_X1 U4595 ( .A1(n3986), .A2(n3985), .ZN(n4154) );
  AOI22_X1 U4596 ( .A1(n2000), .A2(REG2_REG_14__SCAN_IN), .B1(n3987), .B2(
        n4292), .ZN(n3988) );
  OAI21_X1 U4597 ( .B1(n4154), .B2(n4015), .A(n3988), .ZN(n3989) );
  AOI21_X1 U4598 ( .B1(n4094), .B2(n4284), .A(n3989), .ZN(n3990) );
  OAI21_X1 U4599 ( .B1(n3992), .B2(n3991), .A(n3990), .ZN(U3276) );
  INV_X1 U4600 ( .A(n3993), .ZN(n3995) );
  OAI21_X1 U4601 ( .B1(n3996), .B2(n3995), .A(n3994), .ZN(n3997) );
  XNOR2_X1 U4602 ( .A(n3997), .B(n3998), .ZN(n4009) );
  XNOR2_X1 U4603 ( .A(n3999), .B(n3998), .ZN(n4098) );
  NAND2_X1 U4604 ( .A1(n4098), .A2(n4000), .ZN(n4008) );
  OAI22_X1 U4605 ( .A1(n4003), .A2(n4002), .B1(n4001), .B2(n4011), .ZN(n4004)
         );
  AOI21_X1 U4606 ( .B1(n4006), .B2(n4005), .A(n4004), .ZN(n4007) );
  OAI211_X1 U4607 ( .C1(n4010), .C2(n4009), .A(n4008), .B(n4007), .ZN(n4097)
         );
  INV_X1 U4608 ( .A(n4097), .ZN(n4020) );
  OR2_X1 U4609 ( .A1(n4012), .A2(n4011), .ZN(n4013) );
  NAND2_X1 U4610 ( .A1(n4014), .A2(n4013), .ZN(n4158) );
  NOR2_X1 U4611 ( .A1(n4158), .A2(n4015), .ZN(n4018) );
  OAI22_X1 U4612 ( .A1(n4284), .A2(n2876), .B1(n4016), .B2(n4304), .ZN(n4017)
         );
  AOI211_X1 U4613 ( .C1(n4098), .C2(n4307), .A(n4018), .B(n4017), .ZN(n4019)
         );
  OAI21_X1 U4614 ( .B1(n4020), .B2(n2000), .A(n4019), .ZN(U3277) );
  NAND2_X1 U4615 ( .A1(n4029), .A2(n4028), .ZN(n4027) );
  XNOR2_X1 U4616 ( .A(n4027), .B(n4021), .ZN(n4178) );
  INV_X1 U4617 ( .A(n4178), .ZN(n4113) );
  INV_X1 U4618 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4025) );
  NOR2_X1 U4619 ( .A1(n4023), .A2(n4022), .ZN(n4030) );
  AOI21_X1 U4620 ( .B1(n4024), .B2(n4031), .A(n4030), .ZN(n4180) );
  MUX2_X1 U4621 ( .A(n4025), .B(n4180), .S(n4369), .Z(n4026) );
  OAI21_X1 U4622 ( .B1(n4113), .B2(n4110), .A(n4026), .ZN(U3549) );
  OAI21_X1 U4623 ( .B1(n4029), .B2(n4028), .A(n4027), .ZN(n4181) );
  INV_X1 U4624 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4479) );
  AOI21_X1 U4625 ( .B1(n4032), .B2(n4031), .A(n4030), .ZN(n4184) );
  MUX2_X1 U4626 ( .A(n4479), .B(n4184), .S(n4369), .Z(n4033) );
  OAI21_X1 U4627 ( .B1(n4181), .B2(n4110), .A(n4033), .ZN(U3548) );
  NAND2_X1 U4628 ( .A1(n4034), .A2(n4354), .ZN(n4037) );
  MUX2_X1 U4629 ( .A(REG1_REG_29__SCAN_IN), .B(n4116), .S(n4369), .Z(U3547) );
  AOI21_X1 U4630 ( .B1(n4039), .B2(n4354), .A(n4038), .ZN(n4117) );
  MUX2_X1 U4631 ( .A(n4040), .B(n4117), .S(n4369), .Z(n4041) );
  OAI21_X1 U4632 ( .B1(n4120), .B2(n4110), .A(n4041), .ZN(U3546) );
  AOI21_X1 U4633 ( .B1(n4043), .B2(n4356), .A(n4042), .ZN(n4044) );
  OAI21_X1 U4634 ( .B1(n4045), .B2(n4342), .A(n4044), .ZN(n4121) );
  MUX2_X1 U4635 ( .A(REG1_REG_27__SCAN_IN), .B(n4121), .S(n4369), .Z(U3545) );
  AOI21_X1 U4636 ( .B1(n4047), .B2(n4354), .A(n4046), .ZN(n4122) );
  MUX2_X1 U4637 ( .A(n4480), .B(n4122), .S(n4369), .Z(n4048) );
  OAI21_X1 U4638 ( .B1(n4110), .B2(n4125), .A(n4048), .ZN(U3544) );
  AOI21_X1 U4639 ( .B1(n4050), .B2(n4354), .A(n4049), .ZN(n4126) );
  MUX2_X1 U4640 ( .A(n4051), .B(n4126), .S(n4369), .Z(n4052) );
  OAI21_X1 U4641 ( .B1(n4110), .B2(n4128), .A(n4052), .ZN(U3543) );
  AOI21_X1 U4642 ( .B1(n4054), .B2(n4354), .A(n4053), .ZN(n4129) );
  MUX2_X1 U4643 ( .A(n4055), .B(n4129), .S(n4369), .Z(n4056) );
  OAI21_X1 U4644 ( .B1(n4110), .B2(n4131), .A(n4056), .ZN(U3542) );
  AOI21_X1 U4645 ( .B1(n4058), .B2(n4354), .A(n4057), .ZN(n4132) );
  MUX2_X1 U4646 ( .A(n4476), .B(n4132), .S(n4369), .Z(n4059) );
  OAI21_X1 U4647 ( .B1(n4110), .B2(n4134), .A(n4059), .ZN(U3541) );
  NAND3_X1 U4648 ( .A1(n4061), .A2(n4356), .A3(n4060), .ZN(n4062) );
  OAI211_X1 U4649 ( .C1(n4064), .C2(n4342), .A(n4063), .B(n4062), .ZN(n4135)
         );
  MUX2_X1 U4650 ( .A(REG1_REG_22__SCAN_IN), .B(n4135), .S(n4369), .Z(U3540) );
  NAND2_X1 U4651 ( .A1(n4065), .A2(n4354), .ZN(n4067) );
  OAI211_X1 U4652 ( .C1(n4093), .C2(n4068), .A(n4067), .B(n4066), .ZN(n4136)
         );
  MUX2_X1 U4653 ( .A(REG1_REG_21__SCAN_IN), .B(n4136), .S(n4369), .Z(U3539) );
  INV_X1 U4654 ( .A(n4069), .ZN(n4070) );
  AOI21_X1 U4655 ( .B1(n4071), .B2(n4354), .A(n4070), .ZN(n4137) );
  MUX2_X1 U4656 ( .A(n4072), .B(n4137), .S(n4369), .Z(n4073) );
  OAI21_X1 U4657 ( .B1(n4110), .B2(n4139), .A(n4073), .ZN(U3538) );
  AOI21_X1 U4658 ( .B1(n4075), .B2(n4354), .A(n4074), .ZN(n4140) );
  MUX2_X1 U4659 ( .A(n4076), .B(n4140), .S(n4369), .Z(n4077) );
  OAI21_X1 U4660 ( .B1(n4110), .B2(n4143), .A(n4077), .ZN(U3537) );
  OAI211_X1 U4661 ( .C1(n4080), .C2(n4342), .A(n4079), .B(n4078), .ZN(n4144)
         );
  MUX2_X1 U4662 ( .A(REG1_REG_18__SCAN_IN), .B(n4144), .S(n4369), .Z(U3536) );
  AOI21_X1 U4663 ( .B1(n4082), .B2(n4354), .A(n4081), .ZN(n4145) );
  MUX2_X1 U4664 ( .A(n4083), .B(n4145), .S(n4369), .Z(n4084) );
  OAI21_X1 U4665 ( .B1(n4110), .B2(n4148), .A(n4084), .ZN(U3535) );
  AOI21_X1 U4666 ( .B1(n4356), .B2(n4086), .A(n4085), .ZN(n4087) );
  OAI21_X1 U4667 ( .B1(n4088), .B2(n4342), .A(n4087), .ZN(n4149) );
  MUX2_X1 U4668 ( .A(REG1_REG_16__SCAN_IN), .B(n4149), .S(n4369), .Z(U3534) );
  NAND2_X1 U4669 ( .A1(n4089), .A2(n4354), .ZN(n4090) );
  OAI211_X1 U4670 ( .C1(n4093), .C2(n4092), .A(n4091), .B(n4090), .ZN(n4150)
         );
  MUX2_X1 U4671 ( .A(REG1_REG_15__SCAN_IN), .B(n4150), .S(n4369), .Z(U3533) );
  AOI21_X1 U4672 ( .B1(n4095), .B2(n4354), .A(n4094), .ZN(n4151) );
  MUX2_X1 U4673 ( .A(n4244), .B(n4151), .S(n4369), .Z(n4096) );
  OAI21_X1 U4674 ( .B1(n4110), .B2(n4154), .A(n4096), .ZN(U3532) );
  AOI21_X1 U4675 ( .B1(n4339), .B2(n4098), .A(n4097), .ZN(n4155) );
  MUX2_X1 U4676 ( .A(n4099), .B(n4155), .S(n4369), .Z(n4100) );
  OAI21_X1 U4677 ( .B1(n4110), .B2(n4158), .A(n4100), .ZN(U3531) );
  NAND2_X1 U4678 ( .A1(n4101), .A2(n4354), .ZN(n4102) );
  AND2_X1 U4679 ( .A1(n4103), .A2(n4102), .ZN(n4159) );
  MUX2_X1 U4680 ( .A(n4465), .B(n4159), .S(n4369), .Z(n4104) );
  OAI21_X1 U4681 ( .B1(n4110), .B2(n4162), .A(n4104), .ZN(U3530) );
  INV_X1 U4682 ( .A(n4105), .ZN(n4106) );
  AOI21_X1 U4683 ( .B1(n4339), .B2(n4107), .A(n4106), .ZN(n4163) );
  MUX2_X1 U4684 ( .A(n4108), .B(n4163), .S(n4369), .Z(n4109) );
  OAI21_X1 U4685 ( .B1(n4110), .B2(n4167), .A(n4109), .ZN(U3529) );
  INV_X1 U4686 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4111) );
  MUX2_X1 U4687 ( .A(n4111), .B(n4180), .S(n4362), .Z(n4112) );
  OAI21_X1 U4688 ( .B1(n4113), .B2(n4166), .A(n4112), .ZN(U3517) );
  INV_X1 U4689 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4114) );
  MUX2_X1 U4690 ( .A(n4114), .B(n4184), .S(n4362), .Z(n4115) );
  OAI21_X1 U4691 ( .B1(n4181), .B2(n4166), .A(n4115), .ZN(U3516) );
  MUX2_X1 U4692 ( .A(REG0_REG_29__SCAN_IN), .B(n4116), .S(n4362), .Z(U3515) );
  INV_X1 U4693 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4118) );
  MUX2_X1 U4694 ( .A(n4118), .B(n4117), .S(n4362), .Z(n4119) );
  OAI21_X1 U4695 ( .B1(n4120), .B2(n4166), .A(n4119), .ZN(U3514) );
  MUX2_X1 U4696 ( .A(REG0_REG_27__SCAN_IN), .B(n4121), .S(n4362), .Z(U3513) );
  INV_X1 U4697 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4123) );
  MUX2_X1 U4698 ( .A(n4123), .B(n4122), .S(n4362), .Z(n4124) );
  OAI21_X1 U4699 ( .B1(n4125), .B2(n4166), .A(n4124), .ZN(U3512) );
  INV_X1 U4700 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4467) );
  MUX2_X1 U4701 ( .A(n4467), .B(n4126), .S(n4362), .Z(n4127) );
  OAI21_X1 U4702 ( .B1(n4128), .B2(n4166), .A(n4127), .ZN(U3511) );
  INV_X1 U4703 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4468) );
  MUX2_X1 U4704 ( .A(n4468), .B(n4129), .S(n4362), .Z(n4130) );
  OAI21_X1 U4705 ( .B1(n4131), .B2(n4166), .A(n4130), .ZN(U3510) );
  INV_X1 U4706 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4450) );
  MUX2_X1 U4707 ( .A(n4450), .B(n4132), .S(n4362), .Z(n4133) );
  OAI21_X1 U4708 ( .B1(n4134), .B2(n4166), .A(n4133), .ZN(U3509) );
  MUX2_X1 U4709 ( .A(REG0_REG_22__SCAN_IN), .B(n4135), .S(n4362), .Z(U3508) );
  MUX2_X1 U4710 ( .A(REG0_REG_21__SCAN_IN), .B(n4136), .S(n4362), .Z(U3507) );
  INV_X1 U4711 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4448) );
  MUX2_X1 U4712 ( .A(n4448), .B(n4137), .S(n4362), .Z(n4138) );
  OAI21_X1 U4713 ( .B1(n4139), .B2(n4166), .A(n4138), .ZN(U3506) );
  INV_X1 U4714 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4141) );
  MUX2_X1 U4715 ( .A(n4141), .B(n4140), .S(n4362), .Z(n4142) );
  OAI21_X1 U4716 ( .B1(n4143), .B2(n4166), .A(n4142), .ZN(U3505) );
  MUX2_X1 U4717 ( .A(REG0_REG_18__SCAN_IN), .B(n4144), .S(n4362), .Z(U3503) );
  INV_X1 U4718 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4146) );
  MUX2_X1 U4719 ( .A(n4146), .B(n4145), .S(n4362), .Z(n4147) );
  OAI21_X1 U4720 ( .B1(n4148), .B2(n4166), .A(n4147), .ZN(U3501) );
  MUX2_X1 U4721 ( .A(REG0_REG_16__SCAN_IN), .B(n4149), .S(n4362), .Z(U3499) );
  MUX2_X1 U4722 ( .A(REG0_REG_15__SCAN_IN), .B(n4150), .S(n4362), .Z(U3497) );
  INV_X1 U4723 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4152) );
  MUX2_X1 U4724 ( .A(n4152), .B(n4151), .S(n4362), .Z(n4153) );
  OAI21_X1 U4725 ( .B1(n4154), .B2(n4166), .A(n4153), .ZN(U3495) );
  INV_X1 U4726 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4156) );
  MUX2_X1 U4727 ( .A(n4156), .B(n4155), .S(n4362), .Z(n4157) );
  OAI21_X1 U4728 ( .B1(n4158), .B2(n4166), .A(n4157), .ZN(U3493) );
  INV_X1 U4729 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4160) );
  MUX2_X1 U4730 ( .A(n4160), .B(n4159), .S(n4362), .Z(n4161) );
  OAI21_X1 U4731 ( .B1(n4162), .B2(n4166), .A(n4161), .ZN(U3491) );
  INV_X1 U4732 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4164) );
  MUX2_X1 U4733 ( .A(n4164), .B(n4163), .S(n4362), .Z(n4165) );
  OAI21_X1 U4734 ( .B1(n4167), .B2(n4166), .A(n4165), .ZN(U3489) );
  MUX2_X1 U4735 ( .A(DATAI_28_), .B(n4168), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4736 ( .A(DATAI_27_), .B(n4186), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U4737 ( .A(n4169), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4738 ( .A(DATAI_25_), .B(n4170), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4739 ( .A(DATAI_19_), .B(n4171), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4740 ( .A(n4172), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U4741 ( .A(DATAI_16_), .B(n4173), .S(STATE_REG_SCAN_IN), .Z(U3336)
         );
  MUX2_X1 U4742 ( .A(n4174), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U4743 ( .A(DATAI_7_), .B(n4175), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4744 ( .A(DATAI_4_), .B(n4201), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4745 ( .A(n4176), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4746 ( .A(n4177), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4747 ( .A1(n4178), .A2(n4294), .B1(n2000), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4179) );
  OAI21_X1 U4748 ( .B1(n2000), .B2(n4180), .A(n4179), .ZN(U3260) );
  INV_X1 U4749 ( .A(n4181), .ZN(n4182) );
  AOI22_X1 U4750 ( .A1(n4182), .A2(n4294), .B1(REG2_REG_30__SCAN_IN), .B2(
        n2000), .ZN(n4183) );
  OAI21_X1 U4751 ( .B1(n2000), .B2(n4184), .A(n4183), .ZN(U3261) );
  INV_X1 U4752 ( .A(n4188), .ZN(n4185) );
  OAI211_X1 U4753 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4186), .A(n4185), .B(n4187), 
        .ZN(n4192) );
  OAI22_X1 U4754 ( .A1(n4188), .A2(n4187), .B1(n4256), .B2(REG1_REG_0__SCAN_IN), .ZN(n4189) );
  INV_X1 U4755 ( .A(n4189), .ZN(n4191) );
  AOI22_X1 U4756 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4268), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4190) );
  OAI221_X1 U4757 ( .B1(IR_REG_0__SCAN_IN), .B2(n4192), .C1(n2038), .C2(n4191), 
        .A(n4190), .ZN(U3240) );
  AOI21_X1 U4758 ( .B1(n4268), .B2(ADDR_REG_4__SCAN_IN), .A(n4193), .ZN(n4194)
         );
  INV_X1 U4759 ( .A(n4194), .ZN(n4200) );
  XOR2_X1 U4760 ( .A(REG1_REG_4__SCAN_IN), .B(n4195), .Z(n4198) );
  XNOR2_X1 U4761 ( .A(n4196), .B(REG2_REG_4__SCAN_IN), .ZN(n4197) );
  OAI22_X1 U4762 ( .A1(n4198), .A2(n4256), .B1(n4245), .B2(n4197), .ZN(n4199)
         );
  AOI211_X1 U4763 ( .C1(n4201), .C2(n4252), .A(n4200), .B(n4199), .ZN(n4203)
         );
  NAND2_X1 U4764 ( .A1(n4203), .A2(n4202), .ZN(U3244) );
  AOI211_X1 U4765 ( .C1(n4206), .C2(n4205), .A(n4204), .B(n4256), .ZN(n4208)
         );
  AOI211_X1 U4766 ( .C1(n4268), .C2(ADDR_REG_9__SCAN_IN), .A(n4208), .B(n4207), 
        .ZN(n4213) );
  OAI211_X1 U4767 ( .C1(n4211), .C2(n4210), .A(n4278), .B(n4209), .ZN(n4212)
         );
  OAI211_X1 U4768 ( .C1(n4281), .C2(n4323), .A(n4213), .B(n4212), .ZN(U3249)
         );
  AOI211_X1 U4769 ( .C1(n4464), .C2(n4215), .A(n4214), .B(n4256), .ZN(n4217)
         );
  AOI211_X1 U4770 ( .C1(n4268), .C2(ADDR_REG_10__SCAN_IN), .A(n4217), .B(n4216), .ZN(n4221) );
  OAI211_X1 U4771 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4219), .A(n4278), .B(n4218), .ZN(n4220) );
  OAI211_X1 U4772 ( .C1(n4281), .C2(n4222), .A(n4221), .B(n4220), .ZN(U3250)
         );
  AOI211_X1 U4773 ( .C1(n4225), .C2(n4224), .A(n4223), .B(n4256), .ZN(n4227)
         );
  AOI211_X1 U4774 ( .C1(n4268), .C2(ADDR_REG_11__SCAN_IN), .A(n4227), .B(n4226), .ZN(n4232) );
  OAI211_X1 U4775 ( .C1(n4230), .C2(n4229), .A(n4278), .B(n4228), .ZN(n4231)
         );
  OAI211_X1 U4776 ( .C1(n4281), .C2(n4319), .A(n4232), .B(n4231), .ZN(U3251)
         );
  AOI211_X1 U4777 ( .C1(n4465), .C2(n4234), .A(n4233), .B(n4256), .ZN(n4237)
         );
  INV_X1 U4778 ( .A(n4235), .ZN(n4236) );
  AOI211_X1 U4779 ( .C1(n4268), .C2(ADDR_REG_12__SCAN_IN), .A(n4237), .B(n4236), .ZN(n4241) );
  OAI211_X1 U4780 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4239), .A(n4278), .B(n4238), .ZN(n4240) );
  OAI211_X1 U4781 ( .C1(n4281), .C2(n4318), .A(n4241), .B(n4240), .ZN(U3252)
         );
  NAND2_X1 U4782 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4268), .ZN(n4255) );
  AOI211_X1 U4783 ( .C1(n4244), .C2(n4243), .A(n4242), .B(n4256), .ZN(n4250)
         );
  AOI211_X1 U4784 ( .C1(n4248), .C2(n4247), .A(n4246), .B(n4245), .ZN(n4249)
         );
  AOI211_X1 U4785 ( .C1(n4252), .C2(n4251), .A(n4250), .B(n4249), .ZN(n4254)
         );
  NAND3_X1 U4786 ( .A1(n4255), .A2(n4254), .A3(n4253), .ZN(U3254) );
  AOI211_X1 U4787 ( .C1(n2021), .C2(n4258), .A(n4257), .B(n4256), .ZN(n4259)
         );
  AOI211_X1 U4788 ( .C1(n4268), .C2(ADDR_REG_15__SCAN_IN), .A(n4260), .B(n4259), .ZN(n4265) );
  AOI21_X1 U4789 ( .B1(n4262), .B2(n2015), .A(n4261), .ZN(n4263) );
  NAND2_X1 U4790 ( .A1(n4278), .A2(n4263), .ZN(n4264) );
  OAI211_X1 U4791 ( .C1(n4281), .C2(n4266), .A(n4265), .B(n4264), .ZN(U3255)
         );
  AOI21_X1 U4792 ( .B1(n4268), .B2(ADDR_REG_17__SCAN_IN), .A(n4267), .ZN(n4280) );
  OAI21_X1 U4793 ( .B1(n4271), .B2(n4270), .A(n4269), .ZN(n4277) );
  OAI21_X1 U4794 ( .B1(n4274), .B2(n4273), .A(n4272), .ZN(n4275) );
  AOI22_X1 U4795 ( .A1(n4278), .A2(n4277), .B1(n4276), .B2(n4275), .ZN(n4279)
         );
  OAI211_X1 U4796 ( .C1(n4282), .C2(n4281), .A(n4280), .B(n4279), .ZN(U3257)
         );
  OAI22_X1 U4797 ( .A1(n4284), .A2(n2106), .B1(n4283), .B2(n4304), .ZN(n4285)
         );
  INV_X1 U4798 ( .A(n4285), .ZN(n4290) );
  INV_X1 U4799 ( .A(n4286), .ZN(n4287) );
  AOI22_X1 U4800 ( .A1(n4288), .A2(n4307), .B1(n4294), .B2(n4287), .ZN(n4289)
         );
  OAI211_X1 U4801 ( .C1(n2000), .C2(n4291), .A(n4290), .B(n4289), .ZN(U3284)
         );
  AOI22_X1 U4802 ( .A1(REG2_REG_2__SCAN_IN), .A2(n2000), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4292), .ZN(n4297) );
  AOI22_X1 U4803 ( .A1(n4295), .A2(n4307), .B1(n4294), .B2(n4293), .ZN(n4296)
         );
  OAI211_X1 U4804 ( .C1(n2000), .C2(n4298), .A(n4297), .B(n4296), .ZN(U3288)
         );
  INV_X1 U4805 ( .A(n4299), .ZN(n4301) );
  AOI21_X1 U4806 ( .B1(n4302), .B2(n4301), .A(n4300), .ZN(n4309) );
  NOR2_X1 U4807 ( .A1(n4304), .A2(n4303), .ZN(n4305) );
  AOI21_X1 U4808 ( .B1(n4307), .B2(n4306), .A(n4305), .ZN(n4308) );
  OAI221_X1 U4809 ( .B1(n2000), .B2(n4309), .C1(n4284), .C2(n2347), .A(n4308), 
        .ZN(U3290) );
  AND2_X1 U4810 ( .A1(D_REG_31__SCAN_IN), .A2(n4311), .ZN(U3291) );
  AND2_X1 U4811 ( .A1(D_REG_30__SCAN_IN), .A2(n4311), .ZN(U3292) );
  INV_X1 U4812 ( .A(D_REG_29__SCAN_IN), .ZN(n4441) );
  NOR2_X1 U4813 ( .A1(n4310), .A2(n4441), .ZN(U3293) );
  AND2_X1 U4814 ( .A1(D_REG_28__SCAN_IN), .A2(n4311), .ZN(U3294) );
  INV_X1 U4815 ( .A(D_REG_27__SCAN_IN), .ZN(n4442) );
  NOR2_X1 U4816 ( .A1(n4310), .A2(n4442), .ZN(U3295) );
  AND2_X1 U4817 ( .A1(D_REG_26__SCAN_IN), .A2(n4311), .ZN(U3296) );
  AND2_X1 U4818 ( .A1(D_REG_25__SCAN_IN), .A2(n4311), .ZN(U3297) );
  AND2_X1 U4819 ( .A1(D_REG_24__SCAN_IN), .A2(n4311), .ZN(U3298) );
  AND2_X1 U4820 ( .A1(D_REG_23__SCAN_IN), .A2(n4311), .ZN(U3299) );
  AND2_X1 U4821 ( .A1(D_REG_22__SCAN_IN), .A2(n4311), .ZN(U3300) );
  AND2_X1 U4822 ( .A1(D_REG_21__SCAN_IN), .A2(n4311), .ZN(U3301) );
  AND2_X1 U4823 ( .A1(D_REG_20__SCAN_IN), .A2(n4311), .ZN(U3302) );
  AND2_X1 U4824 ( .A1(D_REG_19__SCAN_IN), .A2(n4311), .ZN(U3303) );
  AND2_X1 U4825 ( .A1(D_REG_18__SCAN_IN), .A2(n4311), .ZN(U3304) );
  INV_X1 U4826 ( .A(D_REG_17__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U4827 ( .A1(n4310), .A2(n4427), .ZN(U3305) );
  INV_X1 U4828 ( .A(D_REG_16__SCAN_IN), .ZN(n4426) );
  NOR2_X1 U4829 ( .A1(n4310), .A2(n4426), .ZN(U3306) );
  AND2_X1 U4830 ( .A1(D_REG_15__SCAN_IN), .A2(n4311), .ZN(U3307) );
  AND2_X1 U4831 ( .A1(D_REG_14__SCAN_IN), .A2(n4311), .ZN(U3308) );
  AND2_X1 U4832 ( .A1(D_REG_13__SCAN_IN), .A2(n4311), .ZN(U3309) );
  AND2_X1 U4833 ( .A1(D_REG_12__SCAN_IN), .A2(n4311), .ZN(U3310) );
  INV_X1 U4834 ( .A(D_REG_11__SCAN_IN), .ZN(n4430) );
  NOR2_X1 U4835 ( .A1(n4310), .A2(n4430), .ZN(U3311) );
  AND2_X1 U4836 ( .A1(D_REG_10__SCAN_IN), .A2(n4311), .ZN(U3312) );
  AND2_X1 U4837 ( .A1(D_REG_9__SCAN_IN), .A2(n4311), .ZN(U3313) );
  AND2_X1 U4838 ( .A1(D_REG_8__SCAN_IN), .A2(n4311), .ZN(U3314) );
  AND2_X1 U4839 ( .A1(D_REG_7__SCAN_IN), .A2(n4311), .ZN(U3315) );
  INV_X1 U4840 ( .A(D_REG_6__SCAN_IN), .ZN(n4429) );
  NOR2_X1 U4841 ( .A1(n4310), .A2(n4429), .ZN(U3316) );
  INV_X1 U4842 ( .A(D_REG_5__SCAN_IN), .ZN(n4433) );
  NOR2_X1 U4843 ( .A1(n4310), .A2(n4433), .ZN(U3317) );
  AND2_X1 U4844 ( .A1(D_REG_4__SCAN_IN), .A2(n4311), .ZN(U3318) );
  INV_X1 U4845 ( .A(D_REG_3__SCAN_IN), .ZN(n4432) );
  NOR2_X1 U4846 ( .A1(n4310), .A2(n4432), .ZN(U3319) );
  AND2_X1 U4847 ( .A1(D_REG_2__SCAN_IN), .A2(n4311), .ZN(U3320) );
  INV_X1 U4848 ( .A(DATAI_23_), .ZN(n4403) );
  AOI21_X1 U4849 ( .B1(U3149), .B2(n4403), .A(n4312), .ZN(U3329) );
  OAI22_X1 U4850 ( .A1(U3149), .A2(n4313), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4314) );
  INV_X1 U4851 ( .A(n4314), .ZN(U3335) );
  OAI22_X1 U4852 ( .A1(U3149), .A2(n4315), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4316) );
  INV_X1 U4853 ( .A(n4316), .ZN(U3337) );
  INV_X1 U4854 ( .A(DATAI_14_), .ZN(n4405) );
  AOI22_X1 U4855 ( .A1(STATE_REG_SCAN_IN), .A2(n4317), .B1(n4405), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U4856 ( .A(DATAI_12_), .ZN(n4406) );
  AOI22_X1 U4857 ( .A1(STATE_REG_SCAN_IN), .A2(n4318), .B1(n4406), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U4858 ( .A(DATAI_11_), .ZN(n4408) );
  AOI22_X1 U4859 ( .A1(STATE_REG_SCAN_IN), .A2(n4319), .B1(n4408), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U4860 ( .A1(U3149), .A2(n4320), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4321) );
  INV_X1 U4861 ( .A(n4321), .ZN(U3342) );
  INV_X1 U4862 ( .A(DATAI_9_), .ZN(n4322) );
  AOI22_X1 U4863 ( .A1(STATE_REG_SCAN_IN), .A2(n4323), .B1(n4322), .B2(U3149), 
        .ZN(U3343) );
  OAI22_X1 U4864 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4324) );
  INV_X1 U4865 ( .A(n4324), .ZN(U3352) );
  INV_X1 U4866 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U4867 ( .A1(n4362), .A2(n4326), .B1(n4325), .B2(n4361), .ZN(U3467)
         );
  INV_X1 U4868 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U4869 ( .A1(n4362), .A2(n4328), .B1(n4327), .B2(n4361), .ZN(U3469)
         );
  NOR2_X1 U4870 ( .A1(n4330), .A2(n4329), .ZN(n4332) );
  AOI211_X1 U4871 ( .C1(n4356), .C2(n4333), .A(n4332), .B(n4331), .ZN(n4363)
         );
  INV_X1 U4872 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4334) );
  AOI22_X1 U4873 ( .A1(n4362), .A2(n4363), .B1(n4334), .B2(n4361), .ZN(U3473)
         );
  INV_X1 U4874 ( .A(n4335), .ZN(n4340) );
  INV_X1 U4875 ( .A(n4336), .ZN(n4338) );
  AOI211_X1 U4876 ( .C1(n4340), .C2(n4339), .A(n4338), .B(n4337), .ZN(n4364)
         );
  INV_X1 U4877 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U4878 ( .A1(n4362), .A2(n4364), .B1(n4341), .B2(n4361), .ZN(U3475)
         );
  NOR2_X1 U4879 ( .A1(n4343), .A2(n4342), .ZN(n4346) );
  INV_X1 U4880 ( .A(n4344), .ZN(n4345) );
  AOI211_X1 U4881 ( .C1(n4356), .C2(n4347), .A(n4346), .B(n4345), .ZN(n4365)
         );
  INV_X1 U4882 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4883 ( .A1(n4362), .A2(n4365), .B1(n4348), .B2(n4361), .ZN(U3477)
         );
  NAND3_X1 U4884 ( .A1(n2804), .A2(n4349), .A3(n4354), .ZN(n4350) );
  AND3_X1 U4885 ( .A1(n4352), .A2(n4351), .A3(n4350), .ZN(n4366) );
  INV_X1 U4886 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4353) );
  AOI22_X1 U4887 ( .A1(n4362), .A2(n4366), .B1(n4353), .B2(n4361), .ZN(U3481)
         );
  NAND2_X1 U4888 ( .A1(n4355), .A2(n4354), .ZN(n4359) );
  NAND2_X1 U4889 ( .A1(n4357), .A2(n4356), .ZN(n4358) );
  AND3_X1 U4890 ( .A1(n4360), .A2(n4359), .A3(n4358), .ZN(n4368) );
  INV_X1 U4891 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U4892 ( .A1(n4362), .A2(n4368), .B1(n4445), .B2(n4361), .ZN(U3485)
         );
  AOI22_X1 U4893 ( .A1(n4369), .A2(n4363), .B1(n2305), .B2(n4367), .ZN(U3521)
         );
  AOI22_X1 U4894 ( .A1(n4369), .A2(n4364), .B1(n2546), .B2(n4367), .ZN(U3522)
         );
  AOI22_X1 U4895 ( .A1(n4369), .A2(n4365), .B1(n4461), .B2(n4367), .ZN(U3523)
         );
  AOI22_X1 U4896 ( .A1(n4369), .A2(n4366), .B1(n4462), .B2(n4367), .ZN(U3525)
         );
  AOI22_X1 U4897 ( .A1(n4369), .A2(n4368), .B1(n2785), .B2(n4367), .ZN(U3527)
         );
  MUX2_X1 U4898 ( .A(DATAO_REG_7__SCAN_IN), .B(n4370), .S(U4043), .Z(n4397) );
  INV_X1 U4899 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4447) );
  NOR4_X1 U4900 ( .A1(n4450), .A2(n4447), .A3(n4468), .A4(n4479), .ZN(n4380)
         );
  NAND3_X1 U4901 ( .A1(REG3_REG_23__SCAN_IN), .A2(DATAO_REG_29__SCAN_IN), .A3(
        n4493), .ZN(n4373) );
  NAND4_X1 U4902 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG1_REG_26__SCAN_IN), .A3(
        ADDR_REG_13__SCAN_IN), .A4(DATAO_REG_19__SCAN_IN), .ZN(n4372) );
  NAND4_X1 U4903 ( .A1(D_REG_5__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .A3(
        REG1_REG_23__SCAN_IN), .A4(REG0_REG_16__SCAN_IN), .ZN(n4371) );
  NOR4_X1 U4904 ( .A1(REG2_REG_4__SCAN_IN), .A2(n4373), .A3(n4372), .A4(n4371), 
        .ZN(n4379) );
  NAND4_X1 U4905 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n4377) );
  NAND4_X1 U4906 ( .A1(D_REG_16__SCAN_IN), .A2(DATAI_14_), .A3(DATAI_12_), 
        .A4(REG1_REG_10__SCAN_IN), .ZN(n4376) );
  NAND4_X1 U4907 ( .A1(REG0_REG_9__SCAN_IN), .A2(REG2_REG_9__SCAN_IN), .A3(
        REG1_REG_5__SCAN_IN), .A4(ADDR_REG_9__SCAN_IN), .ZN(n4375) );
  NAND4_X1 U4908 ( .A1(REG2_REG_25__SCAN_IN), .A2(DATAI_23_), .A3(
        REG2_REG_3__SCAN_IN), .A4(REG3_REG_2__SCAN_IN), .ZN(n4374) );
  NOR4_X1 U4909 ( .A1(n4377), .A2(n4376), .A3(n4375), .A4(n4374), .ZN(n4378)
         );
  AND3_X1 U4910 ( .A1(n4380), .A2(n4379), .A3(n4378), .ZN(n4395) );
  NOR4_X1 U4911 ( .A1(IR_REG_28__SCAN_IN), .A2(DATAO_REG_3__SCAN_IN), .A3(
        DATAO_REG_15__SCAN_IN), .A4(n4462), .ZN(n4394) );
  NOR4_X1 U4912 ( .A1(D_REG_3__SCAN_IN), .A2(REG0_REG_22__SCAN_IN), .A3(
        REG1_REG_21__SCAN_IN), .A4(REG0_REG_20__SCAN_IN), .ZN(n4384) );
  NOR4_X1 U4913 ( .A1(D_REG_17__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .A3(
        DATAI_11_), .A4(DATAI_8_), .ZN(n4383) );
  NOR4_X1 U4914 ( .A1(REG2_REG_15__SCAN_IN), .A2(REG1_REG_12__SCAN_IN), .A3(
        REG2_REG_8__SCAN_IN), .A4(REG1_REG_2__SCAN_IN), .ZN(n4382) );
  NOR4_X1 U4915 ( .A1(REG2_REG_27__SCAN_IN), .A2(REG2_REG_16__SCAN_IN), .A3(
        REG2_REG_18__SCAN_IN), .A4(DATAI_31_), .ZN(n4381) );
  NAND4_X1 U4916 ( .A1(n4384), .A2(n4383), .A3(n4382), .A4(n4381), .ZN(n4392)
         );
  INV_X1 U4917 ( .A(IR_REG_16__SCAN_IN), .ZN(n4385) );
  AND4_X1 U4918 ( .A1(n4386), .A2(n4385), .A3(n2083), .A4(IR_REG_25__SCAN_IN), 
        .ZN(n4390) );
  NOR4_X1 U4919 ( .A1(REG0_REG_27__SCAN_IN), .A2(REG0_REG_25__SCAN_IN), .A3(
        DATAI_20_), .A4(DATAI_30_), .ZN(n4387) );
  AND3_X1 U4920 ( .A1(n4416), .A2(n4388), .A3(n4387), .ZN(n4389) );
  NAND4_X1 U4921 ( .A1(n4390), .A2(n4389), .A3(IR_REG_13__SCAN_IN), .A4(
        IR_REG_31__SCAN_IN), .ZN(n4391) );
  NOR2_X1 U4922 ( .A1(n4392), .A2(n4391), .ZN(n4393) );
  NAND3_X1 U4923 ( .A1(n4395), .A2(n4394), .A3(n4393), .ZN(n4396) );
  XNOR2_X1 U4924 ( .A(n4397), .B(n4396), .ZN(n4525) );
  AOI22_X1 U4925 ( .A1(n4400), .A2(keyinput19), .B1(keyinput2), .B2(n4399), 
        .ZN(n4398) );
  OAI221_X1 U4926 ( .B1(n4400), .B2(keyinput19), .C1(n4399), .C2(keyinput2), 
        .A(n4398), .ZN(n4413) );
  AOI22_X1 U4927 ( .A1(n4403), .A2(keyinput15), .B1(keyinput40), .B2(n4402), 
        .ZN(n4401) );
  OAI221_X1 U4928 ( .B1(n4403), .B2(keyinput15), .C1(n4402), .C2(keyinput40), 
        .A(n4401), .ZN(n4412) );
  AOI22_X1 U4929 ( .A1(n4406), .A2(keyinput54), .B1(n4405), .B2(keyinput31), 
        .ZN(n4404) );
  OAI221_X1 U4930 ( .B1(n4406), .B2(keyinput54), .C1(n4405), .C2(keyinput31), 
        .A(n4404), .ZN(n4411) );
  AOI22_X1 U4931 ( .A1(n4409), .A2(keyinput33), .B1(n4408), .B2(keyinput1), 
        .ZN(n4407) );
  OAI221_X1 U4932 ( .B1(n4409), .B2(keyinput33), .C1(n4408), .C2(keyinput1), 
        .A(n4407), .ZN(n4410) );
  NOR4_X1 U4933 ( .A1(n4413), .A2(n4412), .A3(n4411), .A4(n4410), .ZN(n4459)
         );
  AOI22_X1 U4934 ( .A1(n4416), .A2(keyinput58), .B1(n4415), .B2(keyinput55), 
        .ZN(n4414) );
  OAI221_X1 U4935 ( .B1(n4416), .B2(keyinput58), .C1(n4415), .C2(keyinput55), 
        .A(n4414), .ZN(n4424) );
  XOR2_X1 U4936 ( .A(IR_REG_25__SCAN_IN), .B(keyinput6), .Z(n4423) );
  XNOR2_X1 U4937 ( .A(n2083), .B(keyinput48), .ZN(n4422) );
  XNOR2_X1 U4938 ( .A(IR_REG_13__SCAN_IN), .B(keyinput32), .ZN(n4420) );
  XNOR2_X1 U4939 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput10), .ZN(n4419) );
  XNOR2_X1 U4940 ( .A(IR_REG_18__SCAN_IN), .B(keyinput30), .ZN(n4418) );
  XNOR2_X1 U4941 ( .A(IR_REG_16__SCAN_IN), .B(keyinput34), .ZN(n4417) );
  NAND4_X1 U4942 ( .A1(n4420), .A2(n4419), .A3(n4418), .A4(n4417), .ZN(n4421)
         );
  NOR4_X1 U4943 ( .A1(n4424), .A2(n4423), .A3(n4422), .A4(n4421), .ZN(n4458)
         );
  AOI22_X1 U4944 ( .A1(n4427), .A2(keyinput12), .B1(keyinput36), .B2(n4426), 
        .ZN(n4425) );
  OAI221_X1 U4945 ( .B1(n4427), .B2(keyinput12), .C1(n4426), .C2(keyinput36), 
        .A(n4425), .ZN(n4439) );
  AOI22_X1 U4946 ( .A1(n4430), .A2(keyinput22), .B1(keyinput7), .B2(n4429), 
        .ZN(n4428) );
  OAI221_X1 U4947 ( .B1(n4430), .B2(keyinput22), .C1(n4429), .C2(keyinput7), 
        .A(n4428), .ZN(n4438) );
  AOI22_X1 U4948 ( .A1(n4433), .A2(keyinput39), .B1(n4432), .B2(keyinput28), 
        .ZN(n4431) );
  OAI221_X1 U4949 ( .B1(n4433), .B2(keyinput39), .C1(n4432), .C2(keyinput28), 
        .A(n4431), .ZN(n4437) );
  XNOR2_X1 U4950 ( .A(IR_REG_31__SCAN_IN), .B(keyinput9), .ZN(n4435) );
  XNOR2_X1 U4951 ( .A(IR_REG_28__SCAN_IN), .B(keyinput0), .ZN(n4434) );
  NAND2_X1 U4952 ( .A1(n4435), .A2(n4434), .ZN(n4436) );
  NOR4_X1 U4953 ( .A1(n4439), .A2(n4438), .A3(n4437), .A4(n4436), .ZN(n4457)
         );
  AOI22_X1 U4954 ( .A1(n4442), .A2(keyinput63), .B1(n4441), .B2(keyinput46), 
        .ZN(n4440) );
  OAI221_X1 U4955 ( .B1(n4442), .B2(keyinput63), .C1(n4441), .C2(keyinput46), 
        .A(n4440), .ZN(n4455) );
  INV_X1 U4956 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4444) );
  AOI22_X1 U4957 ( .A1(n4445), .A2(keyinput20), .B1(n4444), .B2(keyinput29), 
        .ZN(n4443) );
  OAI221_X1 U4958 ( .B1(n4445), .B2(keyinput20), .C1(n4444), .C2(keyinput29), 
        .A(n4443), .ZN(n4454) );
  AOI22_X1 U4959 ( .A1(n4448), .A2(keyinput45), .B1(n4447), .B2(keyinput35), 
        .ZN(n4446) );
  OAI221_X1 U4960 ( .B1(n4448), .B2(keyinput45), .C1(n4447), .C2(keyinput35), 
        .A(n4446), .ZN(n4453) );
  INV_X1 U4961 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4451) );
  AOI22_X1 U4962 ( .A1(n4451), .A2(keyinput43), .B1(n4450), .B2(keyinput3), 
        .ZN(n4449) );
  OAI221_X1 U4963 ( .B1(n4451), .B2(keyinput43), .C1(n4450), .C2(keyinput3), 
        .A(n4449), .ZN(n4452) );
  NOR4_X1 U4964 ( .A1(n4455), .A2(n4454), .A3(n4453), .A4(n4452), .ZN(n4456)
         );
  NAND4_X1 U4965 ( .A1(n4459), .A2(n4458), .A3(n4457), .A4(n4456), .ZN(n4523)
         );
  AOI22_X1 U4966 ( .A1(n4462), .A2(keyinput8), .B1(keyinput42), .B2(n4461), 
        .ZN(n4460) );
  OAI221_X1 U4967 ( .B1(n4462), .B2(keyinput8), .C1(n4461), .C2(keyinput42), 
        .A(n4460), .ZN(n4474) );
  AOI22_X1 U4968 ( .A1(n4465), .A2(keyinput26), .B1(keyinput37), .B2(n4464), 
        .ZN(n4463) );
  OAI221_X1 U4969 ( .B1(n4465), .B2(keyinput26), .C1(n4464), .C2(keyinput37), 
        .A(n4463), .ZN(n4473) );
  AOI22_X1 U4970 ( .A1(n4468), .A2(keyinput17), .B1(n4467), .B2(keyinput47), 
        .ZN(n4466) );
  OAI221_X1 U4971 ( .B1(n4468), .B2(keyinput17), .C1(n4467), .C2(keyinput47), 
        .A(n4466), .ZN(n4472) );
  XNOR2_X1 U4972 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput50), .ZN(n4470) );
  XNOR2_X1 U4973 ( .A(REG0_REG_27__SCAN_IN), .B(keyinput53), .ZN(n4469) );
  NAND2_X1 U4974 ( .A1(n4470), .A2(n4469), .ZN(n4471) );
  NOR4_X1 U4975 ( .A1(n4474), .A2(n4473), .A3(n4472), .A4(n4471), .ZN(n4521)
         );
  AOI22_X1 U4976 ( .A1(n4477), .A2(keyinput51), .B1(n4476), .B2(keyinput18), 
        .ZN(n4475) );
  OAI221_X1 U4977 ( .B1(n4477), .B2(keyinput51), .C1(n4476), .C2(keyinput18), 
        .A(n4475), .ZN(n4488) );
  AOI22_X1 U4978 ( .A1(n4480), .A2(keyinput24), .B1(keyinput56), .B2(n4479), 
        .ZN(n4478) );
  OAI221_X1 U4979 ( .B1(n4480), .B2(keyinput24), .C1(n4479), .C2(keyinput56), 
        .A(n4478), .ZN(n4487) );
  INV_X1 U4980 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4482) );
  AOI22_X1 U4981 ( .A1(n4482), .A2(keyinput27), .B1(n2597), .B2(keyinput21), 
        .ZN(n4481) );
  OAI221_X1 U4982 ( .B1(n4482), .B2(keyinput27), .C1(n2597), .C2(keyinput21), 
        .A(n4481), .ZN(n4486) );
  AOI22_X1 U4983 ( .A1(n2869), .A2(keyinput5), .B1(n4484), .B2(keyinput11), 
        .ZN(n4483) );
  OAI221_X1 U4984 ( .B1(n2869), .B2(keyinput5), .C1(n4484), .C2(keyinput11), 
        .A(n4483), .ZN(n4485) );
  NOR4_X1 U4985 ( .A1(n4488), .A2(n4487), .A3(n4486), .A4(n4485), .ZN(n4520)
         );
  AOI22_X1 U4986 ( .A1(n4491), .A2(keyinput4), .B1(keyinput41), .B2(n4490), 
        .ZN(n4489) );
  OAI221_X1 U4987 ( .B1(n4491), .B2(keyinput4), .C1(n4490), .C2(keyinput41), 
        .A(n4489), .ZN(n4503) );
  AOI22_X1 U4988 ( .A1(n4493), .A2(keyinput44), .B1(keyinput59), .B2(n3908), 
        .ZN(n4492) );
  OAI221_X1 U4989 ( .B1(n4493), .B2(keyinput44), .C1(n3908), .C2(keyinput59), 
        .A(n4492), .ZN(n4502) );
  INV_X1 U4990 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4496) );
  INV_X1 U4991 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U4992 ( .A1(n4496), .A2(keyinput61), .B1(n4495), .B2(keyinput49), 
        .ZN(n4494) );
  OAI221_X1 U4993 ( .B1(n4496), .B2(keyinput61), .C1(n4495), .C2(keyinput49), 
        .A(n4494), .ZN(n4501) );
  INV_X1 U4994 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4499) );
  INV_X1 U4995 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4498) );
  AOI22_X1 U4996 ( .A1(n4499), .A2(keyinput16), .B1(n4498), .B2(keyinput60), 
        .ZN(n4497) );
  OAI221_X1 U4997 ( .B1(n4499), .B2(keyinput16), .C1(n4498), .C2(keyinput60), 
        .A(n4497), .ZN(n4500) );
  NOR4_X1 U4998 ( .A1(n4503), .A2(n4502), .A3(n4501), .A4(n4500), .ZN(n4519)
         );
  INV_X1 U4999 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4505) );
  AOI22_X1 U5000 ( .A1(n4506), .A2(keyinput14), .B1(n4505), .B2(keyinput13), 
        .ZN(n4504) );
  OAI221_X1 U5001 ( .B1(n4506), .B2(keyinput14), .C1(n4505), .C2(keyinput13), 
        .A(n4504), .ZN(n4517) );
  AOI22_X1 U5002 ( .A1(n4509), .A2(keyinput25), .B1(keyinput52), .B2(n4508), 
        .ZN(n4507) );
  OAI221_X1 U5003 ( .B1(n4509), .B2(keyinput25), .C1(n4508), .C2(keyinput52), 
        .A(n4507), .ZN(n4516) );
  AOI22_X1 U5004 ( .A1(n2523), .A2(keyinput23), .B1(n4511), .B2(keyinput57), 
        .ZN(n4510) );
  OAI221_X1 U5005 ( .B1(n2523), .B2(keyinput23), .C1(n4511), .C2(keyinput57), 
        .A(n4510), .ZN(n4515) );
  XOR2_X1 U5006 ( .A(n2782), .B(keyinput62), .Z(n4513) );
  XNOR2_X1 U5007 ( .A(IR_REG_29__SCAN_IN), .B(keyinput38), .ZN(n4512) );
  NAND2_X1 U5008 ( .A1(n4513), .A2(n4512), .ZN(n4514) );
  NOR4_X1 U5009 ( .A1(n4517), .A2(n4516), .A3(n4515), .A4(n4514), .ZN(n4518)
         );
  NAND4_X1 U5010 ( .A1(n4521), .A2(n4520), .A3(n4519), .A4(n4518), .ZN(n4522)
         );
  NOR2_X1 U5011 ( .A1(n4523), .A2(n4522), .ZN(n4524) );
  XOR2_X1 U5012 ( .A(n4525), .B(n4524), .Z(U3557) );
endmodule

